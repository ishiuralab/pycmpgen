module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [24:0] src26;
    reg [23:0] src27;
    reg [22:0] src28;
    reg [21:0] src29;
    reg [20:0] src30;
    reg [19:0] src31;
    reg [18:0] src32;
    reg [17:0] src33;
    reg [16:0] src34;
    reg [15:0] src35;
    reg [14:0] src36;
    reg [13:0] src37;
    reg [12:0] src38;
    reg [11:0] src39;
    reg [10:0] src40;
    reg [9:0] src41;
    reg [8:0] src42;
    reg [7:0] src43;
    reg [6:0] src44;
    reg [5:0] src45;
    reg [4:0] src46;
    reg [3:0] src47;
    reg [2:0] src48;
    reg [1:0] src49;
    reg [0:0] src50;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [51:0] srcsum;
    wire [51:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3])<<47) + ((src48[0] + src48[1] + src48[2])<<48) + ((src49[0] + src49[1])<<49) + ((src50[0])<<50);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd86cf4e2bcd312285ef7eef69ee0012a09b6b3e744674e3097da79fa4a4934d4c35d32afb9f99de20c270ce81ee860509b34a9ceb42d32a8d67a76dd137299f011b28dbbe7d70b58b482cf4d5339389ee79aa27f3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f8e634e254f488a7a805c50c514e57cdcd183adf8aab2a2f3d8a3a97950e14dc697ad90e16ce73f3df4e1bbb2ec19b2cb6e41728b9b369c813ce58fee0859541e65f3b9eb75eb8c99e7035a207b46ed5e83285fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28f46cbde47922211a84fd8ec5b3e0b2828d9f98078e5ebfacbb337bac81dd8a4d6b6741c9457b26bded5eb8b32a44b2ab5db2d69732a8772e3fd7fb051e67c8e84bc9bd36840fada6978e594471121aac274c2fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60d177d03e730e2cc60af77aa9bb367880a0431d555ae9b21c4166e0d0be88ce16ca4eb77002c379bd569c1b0e8ccdef58e05be1cfa9bbbb18ffb0415cd6c8d5ebad038c6026adaa6ef609520d53669aa909551d6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h260bb61da7e35caff9a5097739a336fa777567d41707dfbe0b3f2f7180174b470346ee00d892852d914bf4f262b87f21b4081a7e5fcebf7c2bb6dd78d8ba35e70b47d075b0dd62da550bca9febd34155b211886c0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcec9ed0b4f4e62842867cfef0c8751a607daf4a2aacfb1941ca7d2b49390c2aeb39f4172437bccbc70c0d3697cbf65605a230c0529d61b00b6131f6d4789651b1e394279bc1b4eed7dc48e99e194bb737bdc1ca06;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d7e98d24db11c2c08b22c8fe801feec671ece4c864eab2a63e4ae27dd6727d83cf629351e68187c8f98fe11495b7079dcb09148783fafd91fec9288e8002f8e0d429f5b7dc414e02923de6f6d1dc5e3f197596ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc48a8fbb4773c11ed8a5a10cf6ad37147ee71d5bdeae32f928d46a383b321b480a014565fae26e4b4b20122cd63be685e8327e9d5c854996e2703130d319ff94b8310dd3bfa64137390b0385c546a7e8f41bfa16c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37a635a74bed208224e020f61c2f3b050b8c3dba2b9fd57b64cd7e20276725442b82f157100348463ceaceb56bd3a1ee99c59c14c0c5039bb51a12c900d1938cdbd54fc4ad47dec6c924268d986f1ffcde5b18bda;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97d655182fb3df0b70dce87d2de88ba83731dd0667355aedd09473d279e85f0266ac2a8fb7343f5f357e5d3c4ae11cf85dc2d3cd2ae092cb9a1e0bb55f45910cfed00a4e147ae3eec9955b03b776468bf417eb327;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9ddbea93fb7934f07639ed847d68650fec09816b458f01ca5132a341325ea676874e1d7c82d1299f7723a8c3abf1ce15027de3c9789947197e8e71ee7070b7b0ad543d96fadcdc26bb908e0858d8337152374db;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd06b1b2422d93550878d5d870a3f484b4bd7587d56090ee23a4d3e5ede2352a5be1eba8021c1864b99a0184ad232c277c78d64726a3b54dbca399c9a369394c7dc94e02c5541a78dae8d8327028b3406fc55930c9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7486ce5e0adc22bee7830fe0f552b6cc161ac5cee55a51ff6abe7503ef8391ef2354eb6a6ca8728a897f8279f58ebb579878c43735c0d7adc6f51d2cb299ad181b05d6e927822b1ae9f569d075701943680b1c842;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf88d8da388086c87121a926d3ad3b822de41b2cc6b9b921a79e90164129ee099c92baedd1b6cf18b8dc47a7eb7d5cfe9481aad0b603720672aa4adab46f76f2759d0dfe0afaa20ef98744f2384004beee1159058d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f6580c94419b710f18fb5f1b7690d0cb853a399a5266e9a51d477ca551078192ccdd2ef592b1723cb0f8118ffcccc7841a8e5cb6f0e65c0a7e20d3cf603576f74455e36c3c1f4f37a140cd92add7408d2ae8dad4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42f35befabbf1bc865ad349b92decb35977c8fce27b0614f4e1d0c742d3396bd6270a6fa467ba26d2f74e9ff4a69efc2747d19738243f0ff1a5b207888d00ea0eb47a32c29c40a9cad40c2f4587fd2a32b6579b68;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc87c735249413ff0389448e33965e2bbef1f19bd1a721d09d482039517d05167f20458205db1d9d2ff4d377f521b99c673abc5103662c6420df4fd62b762a43cb8f674f210ba1a7d40570cb1e32453d2d7d2c9ba6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e7e5c6b2a552ad6748ca1479b1dedd44aa5f81c3561f4bfbc96aa3065133ea757f894ccd3493ac4fedc456d212f5b23d11678b75ddb54641c94e442e46e7a4d274239bc01ea78637856904ca8cacfb3d5aa7bce4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha082e25ed179f4ee1079dea92c46afa5390582a47fc9f732c1b5fbb0fbf0b78deab037ae292c4a60f4f32299164dba2cfa37d9918148841832e51b90a06b08f51feb2b3b59725d02178bff8490e497b51a81ff813;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc493ab0320ab82426e5751d65d493e6a219970df0dfa9691cb5e9815b7ee88ea2f104df1d10d8265cc379b2937ea602655399936b59dd5d54e6998a50f0cfb69b763b82d652c4fb5570cccc44ef96759727cc69f1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb252a77c757dcb1c2579687e5b26c1818ac3c43362bef6da2a9b00a7074e6aaefbcfacf1e1ead7c3c44a7498d0d7159c098e23fb25d5286446d8bc3dcda2cb31bf9a379afbe8efd379651f753ac5d4e9914ed7f8e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h261866209928d9dbc91fdb31e6d0ed4c633b4581928f5df337c406f8ea08660f2bb55ead8035ae80cf56b6e4761b70dce1e0ffbfd3ef3ed920b7b0febdbfa810a6670acc124c6e9141c485a045c083771575a1285;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60370fca1d59f79dab7f8b90ded0772b3e4818a431b7e8f5f59e7e002448c9411a8e013b5a9f4c9aaa38ab9df235d966312be0bbf16b72fde5a4b2a7e70d9dfdb16eb7a8b2a3ba11741dcc32dcef7e870b66a9661;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8197ec079add3e0071ad5b3304eb2eff48de350be9895b0ad67ffdf1493ec19b5e8b7f6c574c2f36628a56a285c758a31c11c76b4737da0197715c29e9e2ae338ba0479bbe655bb5ca14d71c575b20dea18a6824;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf70a11a847dab22c1d90d2533e2f76f26529670995a89bb5d6b88d8bbbd08f881b5984369762ad2912122310ca16114bd2dbe537fe04a2e55dd27259d2efdfcfbb1f78f59e428a270e63dd685fe2de58dc36535b3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41d9a4ab7bf9aff27a856fe4c8d34f81d07823042c1d1ee65d0d4b77a792ebd2ecf73c7848fe8df206ba42a97cf6f0ecf548feb03a8705aee50f06cfd30f53edbf6ea8c7898f26e09b310da18aeeed1ed39c2ca08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67e31f75c78d6e6513e959e36bd26a2231badde265e9f72b2a5cea89890d7bfff3144996edb774b72a30ffc00871e9427f9cbb2c6e438b1da3400dfde5a0a5cb265821e9c52732c6512b12a14f0a48ab7c0e7ec56;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f8b17101ef21740a29fb48212dd1eeeb72f6e0a189e6a88ba9b24f1d1af2d1648a7fccb7afba40f6fd2f50c7ce38857e8d2dfcbe1720b25e88a0f5feca4d65abc74552d28d03de03de836409c327d1d1140cffe9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c2a2180ac47d23d759a4d04c2ca6384b132b6eb71e9ac268268b4b1d1d352353af7d699e2d18e8f9dabcd65d48372c6224e8c78dcb698319236f31d081b5ad7a6b5d573a2b5a2759e48d75cfd21e9f2222b22c3a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74c7207a7363b4bc6710e28bc275f1551d5fc7502ffaeddb25d157266b19692c716b7b4fa37a81aed272be28bb36a5053618daecfe1f95a25de1b799a9e2dc77f45e67f1da2395ca806efdcda52f4e9e5fdbc9d7e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb65a4ec249f3001005304d0125837696daed90ed49a83a54795570765374a4dc37dc602cb2f4549b1adb35ae4de8976a4837ab8192e25b0f4d29614c2f7c8cde5eca245a01812cca15fd932c459530c69a46b252d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e8558bee3360621b7ef9b24a548af8af18b76560a92fa7f3c3076d586f55e390e2e6443ccc63982fd1fbee9ed2ec93190cea179bfbbec00e461c6a1733faf8803824b632f0da99a782ec1bf1ad13d11a62d4310c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hedcb50693fd659a4358d24158d4b42767ab2309d31b538261c3069f4df048fccfb6ad1ec7f263d299aef264a228e4cfdfe4b61f503a0ad1023f7fb80519b584abb7999affce36516574991974366ec6265bc6e4bf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4de0e32e8f43adb76f2441f274b485a8e87c8ca832ded52ec5c0cf3118b1d6f3bf901816297ea8f56f2d3029660ecfc11371e03e5d95887916f5a5500a1b024489c5892efaecfd60e1a38c4ad52f76a918968c889;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb07414b79863dfe999ba943b8971726ed8599d241dfd42e33298d770ce8c090a55000062e6b022143a7a3ab38de573db2e9568bfae520a0e94d8fab239dcac11bc74916bcabd8036c711898bec54904cb7c116e72;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he82cfa901d068ac4706c047e2f1f3bfbdd21368a2e88cae5ae0351796ea19fb5bdcc1bdc267a1fc5075aeb19110cf178d71e9098aea77070916e42d15e5011b596693cf779ece2c27c53bac6d28e08a45265f4d50;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26d3107f3db6015e011915202d0ffe5d68c049a443dd85b3be964bf81e49ae9523e23b54e366d097fad6683b880e70660e1b198bcdf1b60ae7a26cc045051ca19968184fc4684a85b2647b2aa3f60dbb474c35b93;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56954351674fef78471c9b9dce4869ffe1af2a4e91c481f15aaa3b83bacda196eaad2936d0e7417d98f8fd0d2758a2d7c88cbae1881b9a8834497d71f1766a9dcea613ecb68f0af4432e8e411459e60830fbb2483;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h146f444edfcf394b3936fa7f5563671c506e683ed53935200404b66168608e7de7f23c416c5e9e545dfbc89d0554c59c2052f2faca026cdd7efc5935a57895c0773892a501f7f188dd68ad245fc88bb90aadd394f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hffecbdacfc7089b8a84ead4a570099c5c82d60cdcb5ab39acee9e08a7178f9db852530119611756ba8ed52b61bb457fb9917d74d47bd048f768df50838f7038a6b40e2920ae792a9ce86e633a4cbf7dad4ae0bf85;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h744da2e88d6911c9b2d3639f956144ff310b1733c395668c0dc8eff817a0714b6b213b79cd1cf51317f7d4c3db7f5b3bd013ef4b933982cbc38bb4c3a47775113743362da62b7de3a53fff3d92fd176765430c338;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbd71d254018dd38cf716e0e8c617bda25b18ebf3fc07ebb95ef096fab435cecd420021d4b2f78360645dd599a8ce25a75586163a431bf4115b180089c4014ad13856a12731cf2d5300b5e1fa5671fececf67f3d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3bf4765fdc6d39f5c8d5eab02f43e9adc4fcd29d39d1a6ec35f0fd9614c3221cf77f67d7f1dfd4a933b6bb53be4bd496f22eaf44a34cb2f7eb1cdb619f61ec110f4736483d9ab947b0d45df04ba0191abcda4bb4b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7879004eae37df8df6844c79f2c603b2664bae5c3717e3dcb5d212db2a6b3d16298eda461d17f2208cc85bc8bc1bc3a19d4bfa611fd22a86e60a32986add786c3252ae219a5fe67e437b6c7a53d3e30c21e8b9cf9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd73794bc54bcf6395aadd63dc6702abf7ca671dad5521568aad063abc1934d56d3d8d60233897c7f20fcd86ab81100b3ed258a6ad92ef73fbcf6528ee82f7ee2d5cfb194fb83805c0e0708a0862601e5f0efc416;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f07d22c9c2385999d0cb8805cc948f8c29e8477f9f2395196e1660eeba02dd989b7de251bf5f3978b4b314a4d0b83b12e66a7f25dd83b014946cb7345673f629ec884f43f0054d3455303cd5e62c8a231bfd45f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1af40f8f2986fc7027fbd9c07ba4c2ef62f7adc1ba01331c6c20720bb0d78741805f50dd75442fcaea7f95c40f827bcf4a04e97325638b38e6cd571a6c5352368d93a080fe7477c84d0072b2c7502bec88b04613a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h406d8d919096d27902974330e889a497728cb42968259d7ce518ba720d6572f5e019cd8d880d1f98198c496b714610f8caca07da64ad09de9b8f3522f27943ebc58f02d2a63be63320810ac805bcf4d1c9cc5d5d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1dd4afb171a49ea46183867f3b57a15ec2db435a324a5bf2402f56f47c5137d3e292de660958f67ba2f3c3232eb96ad30e2937c2d6de4bd71bd1ce4e860fc493ab72eb089d09d34c9d85b19c5590f3f57d93bfea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h768b46cac8df432301ba792b6b911fe7e04f7364b6a1bd8f3287e0f49cd54acc22bfa5e18bd76281e0f3f1685b60d7d32c3e20c03e80f6d24557ae28c5972fe4810795a0fda5a60d7b996199c952dad1c64c91be6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc666ffcd2c27460e74027ba7e6dddc2eef11320c44b3c6646994cdd005ba090dff4285fc7d7687396c78545438494564d48f32d259f0e787b6a6e09d527544379c686f52e08333d5eca5178f0be8f80c5fbd036;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd559517ea06af1804d2b6a42b99c2abfb26f74e8dcf66dd416459a421ef6f1163d3a42c0650ea45bd88bedc0697a9d2eb8fc68185bd9252b53e4dbc3c7e8208691142b04ce81e827a22b1cc1935974876d1d888e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hecd655423dfe57dd0fe9d5712fcf54e54f9284b0661b3595bd7a7690f8d2d898ae4848008f1399dc7c1b1736591bc820fb99831f00719ed85d7eae24375f68cecbb587f6dd2bc3f0e4db527605a4224024f83c04e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f90e3339b389946f545c6f405dc553525e24ab84271e5361ff097b8ecf3885df3378331c8d38786efe32f72111e11b1ecd53194092f51f33a75c8bdbdedcd2da68b0920b914d85aff310c6cbd910d8553e466060;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6838d555a5e292576744438c9933229d9168da25b648053b7d28e8718ee9319b3ecfaece522499d43c25f4f0e5e052dc034e6e42b621475ff25d167cf6fef1f8364ad482a16fcca6b64a61818a4465ccbba4c9ce6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2208b0234a07ab29099f4542a1f8f730697eac27a51ca28a8be677402bead611f5b1f33f27cd4c2076cf65f17ef4b50a781f6b1ee8f40d844bfd44687cc9a5d199fade360f407d81a6af85b287c805871ce05561;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5639dfbd6f8340e7e7aecf681ef3e96d2d96adef3900f7e7380783da883db97d98fd1a0d176be8fd38d5ac33650c241d1a167f2d8fd6160c8174ce94b45e56cb8216f953ba2457190a9a81b50127b2282868b2ab6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6aff100480c7e880b7e4fe5293d01be2e667173f922fdfd25b735f1e40874ef91139d5b2ffd87ef4dfdba2375aa0ba6cf4b0408e79fe37cf1a9edc88cffc07a57382cf81aafd640136e56ab06ba399d74b3f232e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fb4d92b31b86b4a456bb308e1b5455089d15910e9a2e4888547118c1cfbe8087684451219b9dac8dbc452031af3436e433518b8d5d8f05ad20ab9a2be83952e3efc89413ce2ff4fca8062fcaa175cc4bbf910fa7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4447d05b994a591b329cf39c612c60b5121e5e7153dcd6393e002c66b0b9b372ae57cc2669a76a1503255c261710b12b3c1e6748e65baa83a0bbdb41d4037a99ecd5874f9cf03f3901a0b7af2d31aed79b47237;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h159f75dc1c47f6468795b73ca77758912f124ef6a94ac9645435108e8d426e50ebb7ddcefc3033d79050f693a33b2d7fa5d570d5b0b508e0bdf42c187154af20347c86727e4990e76e44a6dfc1319239db0ae48a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cb6f05a8fae3c36eeb3bc022c434c29bf29eeae9762794ad872af908815b118ac1d5e2412871f657c5dc5bf82d1029c5aa1cab27c8d911cc5cd297f2dbb54821d97fe290eb743e191ff4f85e537365b08da54689;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9671da32f000ae9348ae03ec07e1cc52109126c0e45ad1800dcf6ddde54223dafb316242938ec6ea22d2cb032bcdd5924f3d514ba09e19abdae70b29daa315ee0210898f834a8443446a20e6079fa4afc2e8bacd7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb44f34b085bc877684738379b3c59127991a0df873b20ae51b336bdb40e4c1a14e9e08605fe245be48ec08c109ed86240da822748b288e9de96c48a381cf84eabe19e4cd439d16913afbd5a5bae9265b7b93836dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h456648e44438c78ffa768654886c9f36258a3e29ad73a2464544f1fe7abc22f7914fa70046e5ca28b05cfa849781fbd63e0dd1a13263807d6219b72b1f877c99fbbe947b4ef6eea130095f4bdb3105eb57fd920ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6004b19c2e0bc04c8d562f350a416ec46b7cffc35b0f322af8e57f47ba13bc1e206d3b0de6205956909b34bcbf860382ecb4c60676fd0eadbb018f92cd23f6d9dd8ac112004e6cce6f3fe11358df9242ecb6e0704;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha633905282f70037be242484f882969c86128d35a0639903d2a2b81a06c9da3f69449dfea29b730b92b881efd629efe416fbe808aa180c81417f37b49a22ebb51e7a4a7a245b636dde712aec36d570ee49032439b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3450a6c4d83922a109de3224b2423e49349eef281cabfbc2c781ea1d7ef337308838853b8b83c0e3346673f79625002044bd1c7ba1652509d6de54b47a74bf2ae5a9225a3db9e34ccea52671b8f0dfe43395bbd9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27305f216fd76b2e295c2f59a88972e03eb7b1de731247e902757a0447bf19681a2cd0938978d2efad49137ca7abf866d4d4631c1f14be018ec1fda534861f849a11b6aef53063846671373d25878e9a1126c0a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h540355caa91332ce95c7ecda82862a1a75016bc74f209ea8eb1cc281a7aa3069a70d303f35a6b40ca1f93c13efce32c3e8519672bb7aab890aec805b3ba2f51cde90430fd3adb798e805b3adad1e1ae865cabbc60;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2864cd1f3416a7db442e49013dcc8c8463a14cea7f8bec1cf5dc2ba25ca7540ccf717a048244c3def0f974cc80e55d61a1cf2a36f6a609fdc045a9e4aa54465646a8fe97c65dd1eebb7fa990c71d319d7c2914b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfbdcc94bd40f1053bcc2d8a51e44cbbd30589b452e6a0ec1edf1d1e98c1361f787e7b3c8d81b9ef103ba6c84a5d208b7f7aa803a05c987962eda57c663dd1e1a4fbe71027c98eed58f900d107fa1266d6391eb2b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87b1d801025ac7769631e8530cd206a829651d5634bc1a4c0f0e9861387d46808f637a23d73ffe789fcef4e799fb8be8ff6722c6cc1498f22bbc19442cec955b4e54e01075f31933a1ed07b940fb8fee4d578d482;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf483cfba1c43876424f20ca7815fecfb899e1fc0cb0fced5c7027f6ed54202be15db5c1ad44898102a192459d83c461fcda0edc59273dcf7c972adb18ce69970dbb7b431f3fc74c40547e1fce4fda1d885d1ce154;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a655c9620410e10815674f6a953b509d093c88e94b88f966cfd584ce6a942c3e0ed67edb2a3db55150c75b5bb55aa4eec9a884fe8ccebdb9146a0680e6a92275762093ff237e9a90fc0bc97ad6acf02c1f0f11eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h964affc424364f792a5b5c27014dc099eed03fbccca5d9927580c42baec7194ea9a77ba5ed0e88afe4db37ec655d10cc45338a7ca0a43d9c1949cd451ac02e187e19f4731636c287eff1844429b2681d3070197de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a24f9dd9fe688d9c34cf6cc6fb67badc21044e41c51682bf1e08997ac2211f2510d0efb1db8266d947fb1533c8def79e80c203c120dfd017baaca75ef3538d40ddfe19869e42c6e8d941a7905b01d214103507fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcc269e32a56b99c77f461272116021d16211f1bea8cf6b8e00e523f6a7db74300ff91673d8fd195e68afc56ae4fdd859d50ed2327f290f3d38f885fda77fd13e84d98900c2cad062854ea254ff3daaefea42e38b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0a5be579f84320757b6430e24c06f45e8c0a20fca8864785d36b87bcf7388348bdd0629240a08f6299124d3960e3889bd60f6710f279fbd85deff92b358ad94d52a33035cc26a407a9680038a6f23a16a78dfaa5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe0913cda2e67221e24732c552a02915b2eb1cdb61814b24867389900dda19a5e31820becdc7539d0259047e1debc4b1c8f3fdd0c24153519a9ad371d76b8ce8da61148f83caa9f382c5c84ffcecc3163997babcc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58882e5f6e9c8950881b9e6c65ec1e82c9de873f3fa9fe5b23ea8873204f4fb357e44555e3eaa47fbb3dd0c87b90e505b4c60d8c0d7119d2d71004d595afb2873f12416063a00605453c86f06804521988d5dc16b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4459483b9f3f32f99b8fbcfa27811ae804e285ff3f47ebef5e49929a02fbbf725e80aa7de7b574a759de48006199110dccf8924a18221ecfb63fb84edec93e6c839c8dbe0a1f7aea2a61563d5c0f7bf432aa9142a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5541060f8fdbb2e72e56a55df7bff7bd78fc2f8fa5ac8e6855e0bb582106da656894d30ba543a9db92a4f0f1ba51216d74dcf0b182d0a0266c2030e6e8d5d3e6d4360b6644c996d8f58d04c28b1d6e48a6fdc3097;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75349c7f80f0d483cbe02c26998758e04bdb81a9c78141def12d532545315bdcff5659036895244dfaf702b9577e218f36f8006e79d3c9d2bcd88e9cf25c46ca089b883a0b9a8052e4122523899c14832abb2ffde;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d9d19473a715f729bcb61458fe49454dfd6956887d235b32d57e59457c5b603458eb14ac8346a987b6d661261aff752e96f153c39324593d4bd55e521f5fcd9920e1c4a7aef2b3cadd72172b6a248014b711c3e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcabbb83f57f885c1d6669275be3769d06ebb6311f2e9353d83018d648d51a4b5c7bc0f876dc75cad1ef919fee501c377898c78cf91c8949ce2f06e04b562be06a7440cb8e51c9549447ef72864045a76177958226;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcde7ca69088f8765dff7ba5c8b5d6488468a58004a54bee1b34355f95e0d085a0abf10c00ca350d0ba7a050493eb22913b6a5e58d00a12c9b766e9e079962ce5e125e4fa9c213b18300efa8a0e6951da41c4b6efe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a998489ec64c81f8e8a0aa406d2a132bcfb9227c29d5ef40968521ca4101c443e9e18d1851c706b60e37cfda3b55af277b1f9e16d577e08b836d0248697bd52f4a954ddd91bb7ae8ff8e03262bff317c2457a67c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hadc69ef8d8eacc40b9406c2c0b44443088cf57f75ae4ea8b4aac2d0ff3a072761ba242592c3fbe1e45db86a9a553b49312f962efa594bab41a651e272872be3bd77e8a6b33e24e6ced0e9333f8f2435439d0af30c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb380eee5b9320701b0bb3d43c2b155a70834b8bd5d0ebf2b23e6daa34da1d06d9e994dbbf0eecc692800bc23450c0d833de8063d1fa8956f0983f15abb40d529838e7050a7de5feb0bd6eeec4238db6b23c60802c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1468e173fd16e95151e462efc93e65502ba1169e5837c225846aeefe767fc71c80cf5aeb944c1d485a7a09b2c9b0830a5eb154b1428a8e1e9fb91bbf81452ae2e63ea4627fbcfb6ee95d70fd44d47bb2efeb254b8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e4200820d6e8d5c4eabc6b5ec2899f47d89be753aff7adcbe3c1195083c735238e7562086d958e173740c02b92b72bd173f74864922e983df6e6dd9b6c14eece3a0d939a0f29551f7cbe6c3d7b4bd426753ef1ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f4b648e88ebbf1aa1caf2bf2795afc33fa7ce23dc695039cca549869b6c80acb831768ef5d11cae6c1cb8961415fcbca1957b3067865a8e8c7310f64f73fc8b020bc2e8935607496f47e86ec7852288cd3a590f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbbe3ae60da81d7b4103852017221ee5bdc682e677717b9e6416775070f4a553b0a9a15d17a2e1dbc8cd7b817c49276b9ae86494716392e06426dc13c8f4e3cb4fe642f7a5b5242b7b8b7c64466a24327b005ba85e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ed4bff0e0f461dc42c60bc558845567da94687ae005e401e9423774cc38c59c176b5f9c397ffdea80c79de324b60fe5aaa5b1d5cb21818515fe88ae1602a2699581a1fb0e750ac8da358bb20f9af69810aed8de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5c7bd2eeea4ab5b13113907a595abe5482f043ee2974f65ede0244c7374e99aaaa773ef0c82276b8e3bc67d2e669278c65c6cc853ca37ef7478c9fd32f5045f48aa3e2c452d2bfbb10c60103d3f9f288f7c5c3f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h86e93df642787e9021a85a85aa895a08660967c013b071534dc2705c69afb2218ad5908952ecf1b709146db3c50e7a730c4167de88a744de17bb74f6d952449632abe7ee27de7d4f040b6adb2ba358e6177d0a15c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b665d45d46739f148064dd88d39c2636bfa312e4bd5e3cc8b0c547e6bfc191d45f3618d805a0674831b36eacfbb4bdbe91e7b66f564917d97b4941809ca5a6dc7a2f24fea9372dd07205847fd3d7b8c8536f0d4b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62aa284571db0346e61ac77c93aec5e5dd8dfc1a4afc6e425ee035bdb1326b841470b25a84ee7a3d2a3c54c9e270367576f184a8bc7b7d415e386ea33fba91e052497ea52cd6da4d75a476844d41aaccf80c62aa8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88e2c5575db0867bd70587c396af2303604f97ffde3daeea6fd2ddc5ddd385ae215eeaba2013cd22bcca0a834bdc79c69b6bbdffe2437e4ada9c4c61d0d885856f14da09bee832c5409e6c09ea799d3341072d3fd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b06f977b34940fac9b139e0c2613b94503637e428a69c16343568424b1f62752f99aefccee52ae682dacb525c3388818abe6d7b8be9998f02e276e1eaa4562173a75810a7a02650e71d7f79c2bd94109c340526d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbad9e683e850e18700fb1582d7695c2b4e08e5b1aa5d68d78594a4beeb70923ffa9159859ea7b17329c2cc1af5027f05dbc577d69e7b875a51ca88f3b5733ebb66408a597fb89672dec7894407926eba774e6f5b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61c41203b2b2976effdb4bb0a022c7e77578bed990a37f973a50545b49f72a3210d4ef7df7306eccd59ee646b5b4c3a5a8ec312dff23d157b75e45947cb1fcb3712e74d7d593924f6efce0d68e61a67ab2609b6ab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5beb3e888b3e9cb375f5de2c2d9d76e0be070ac9403b94a5feca804fa1b40c679c416b0d1f497d8a454e9d23484053af40b41a73336986bf3b6428989f775c9b5c84f4598f66ef2a9c1c1b9e00d8e2685c8816c93;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f937af7b1e073c1380d0d08b5f88ef40f8e42dd8d3b06847b60b9a4b6083be5cc52ebf559570c1f7f38a02e4d7158dbc32d62818711098b1c34a91687d08f4b3fb9460e04bb497aacdb516225250e9272cb8b2a5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b3b68d41257150b0d8351dc76847ab3a474a3ef8b5ec6b45813fbd6f4d040cd33929c10edee42b396009915ca3fe6a6aeaca6b8e88694137d69adc3e9107fb9e4fd899f165ed35fad9a83149c19db6049d37e62c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c413f63df9b5d89b85ad8c36857f4f0003e65ccc850f2bef4ee533d61b3b9e97ee3cbfbe35f7b5b4c045967f3fac891f510291904b51ee12f581b4c2a378b86e040018d680b3a230155da077f185c891efff1d00;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5db1f4543a85b55d7c8b7fc585d94b442e68afc0461140be5c8f6fc32553a83c1801e327a787782984e46221549e59304ad9951405a3c7fe7183bbe6450aae6ae9f220d2b801c7a26ccca1d1d317d2cef9ad8eeff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12b3d060490f9baf517087ac3cf188c86eedc175d7e355240feb0d404a7a8f312fe11d456f732f775557f6844fe30a51f33784e58bf69e3a164a3c59f55aa8024285c646763bbed1f45cb4cf5ae79e4eb5004ed0a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf336d764f83dee4b8eea05d9d3e1847ab8107033fd91b7c6ce3fd62d0bff8c6181b45d50468dff93f9498a9b42e454003fea76cb7185cf7cfdfdf69d4623c002e547fe12ffe33b5519f8171aee1ae16b4e75344cb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63738a29b6cd8e33e3f5d6c07356da755973d96b4721e170d333178e88de830374298b6f83bff96eee42a6e165b389e67381b14ac91f158c807bb252f0751766bbdbfebbc61d6e8aa28f42f3af9f486b5f2b6dc81;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2f78cbe718249b21dcaba370b548178ce9e7bf6091ce4fea4b53ca6177ec59f7859c0c6d778ddcf59462afc622a0dfa2f33ce985fe3f4220aefc6b206751b552600d17ccfe339dfca5db397a759b1a7650783eba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a30196cf493a0927531b28ff005466135c1e234a61c4911bf963c010e561fe1a7a179a669b7b1db5d5599ec6e69ab9d10548dff413179ef171c224906f58fd2ebbf03f4e7c7fe82361441828c7b1454bfeb419ea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e9ddc395d8ada355e9de8f83eecb93d67f61747f7600e0ecec70a900540bdb302b48661250fd2f29898d4ac2d7321070238f666b334f4d2769ad5944b4b33e057174b4e371198552f62d401b603bdd3c77e3da31;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59c28c92fa7961ea2ebd5592d449cf5979bd72a8a9c64b53330f51dd42ef61c4eb3c293509ae8c65aafb648ff966d1beba89bf5245e66cfe58c8852766a9dc6f871f7ec6839754f2d0bd5489e18837caa3ee9a664;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c501a04d36bef128daf3d1466315d8e8186a0b5da5292ee8866e3ce05f0537515281dc71a4948c4c13a3363fddb80a174a4b81a94a55217ac5049354d0a26de983fd3c11a55492de323836501a5deac2e140b974;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e3b2dbad94c700ad3d0eabee0f0ea765cb15d309ac2f248a21df7d5fe3bda2e74a9a00d7d74a5f854ab2d5634198c6a40bfa27cbd95c74021bfd66619e49533ff848a9622a24da08e50382bf0d50fde03ca7197a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8aa2031f415b9e54d9b307fbaaab7a30bcb222265bb2873acae2b821e8c804593df1d17e8dea8a8c05d5a398dd6f86a8a829513e1cf2a4539e32ba3d46f8bd7f76923191e62025b7217566940ed3ee540775116ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a8c3eec7c63cbaa9b6acd43bb092c5d9d637357bfbcca3003a2eadef14e139057223c925fc7bd682d9939ddaee53819823f2ecdf0840a096d5ed2a32dc7178d33cb4cb04041fca0cb35707f804cbee6b023dacb5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11d3d158f3d2e3188bd1d52e1dd98b1dd5c383de75135eb65d6c911c8eb1d2c46d499eeed5a8d0474603bc6332a809d00e2f9820c94b1b80c96512fc804393a73ed59c48dfb86600761549039087015a2d541a30d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee867a0c3102dc5a564bf54b3ee8013bf2903d69e37097b164caddb4e874cddefb4af62ce11034ea5645e54faf9fcd7e788d2cfa04da9b4b34a4fefcfc5604cc81cef9ab0a012d15a9148503828fcf17baf374657;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4bf49813f96584f2ac254e78b069cf95be4ae6eb0e55d3dfce74f6f84b066aa46914ba887ce8a41bcaa973792c4a4d6f673189e73fce37fb1187b7415be41c33afdc354089f9993944e0355c08b11ab6eecb15d08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a9ff465eeb5efc9fc98cbdaeb625b1a20527f91b00e85a5287f1f371ec63d70d1c655ba2e142e853ee97a1e05fdcef1391d47f46c647a9f18188b08936bd663aa9f41c3eb4c6a28d051d2dd7f8177cfe94d3cfeb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2047c2e8be5db7b688759ac1c56810244cd45c53c7259e16e1c9c8589825851209a3b62d422b414068970e7ceb7a1b6a7161fc1b4caee1d6b634f13b565d5946b77c8c87c7f3b1feaff9f17729d95a8b2818843a9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83d64a7d486f29655f1d70cc3d3c3d1e13e44b0d96bc0e7ebafaf0222e95a9d15888612c5c6ea3cae103ea1d7af42716bfb48d2c4e3d8fac05b080554ca5a7b45c0bd625cb98d15042c321e15383d8587905a57c6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40d438b7acc3baa6a0b6d2f495db7d773dadde8661b1147367b9475911d3056e9dbb9c28bf5d2fac5b63855b74fbe04130b7b69f9db042c283dc8e0d56f63c7d1f98c3cdfe5f79f30a17b1e5ac6e1c877daee7d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85bb84be2ffe92bf9e1af12243541c9059c873b683249b03c58b58fb2c085b0ecad1f5f7bc65a4fb20f45bb122aab277fd078e71528e494008c865ec3053e8f3bfebf5343a3c6510cec7f6cbc2ed31dc8fa953b6c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a48ac84aa0d0079a9c129b2d07ab233d6127ef5115b6a6cd9414b5a4dd94833778c11b2980ea2c4785f7e55d85ebd171cfbd22ee8f90cf65d3ccf814f00f7456be260af8def4e9f5a477f800a1d3d48e060152fe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha33b1b185c42becd864d275625579801f4b1d76e3da096d7229029d94ca99949ff5894dd07bc4038a658f3067d60bf611fe9b32eec3b3c676be27a8f885f88218b7c7a8ed7aa813ce39b81b8809b58bec1e70b7ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd608d7617ff7d3aa0abdeaeca326d998d1f6b50f9ce0ed6d8c8461481566de332ab84cfbe93d1431ac9faf54fb4c3be3625724835ff8856d2f868a0edb9724ccbaadd3b4e9293627d59860cd3ed03011234918800;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbae2a7a869b9d954f88518a0baa472aef896a53e4faa6e89a4dabf302e69cdaf78e3e48d671474d4c8630d7d395c16c266274549d8fc2b93b257d4f2c79311bf397cdab252e1316bb38f56a3b525fb792d8702914;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h335846a133b786f293ea53feea24edf9177d448389bc70fd9a8035afdc0106fc776567b29a41489779642002322a987b607c785fe7d3a105a37dbde318e057385d59d8f761019547e99818d6e7ea796940e0373df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h803e1bee51506a254546bb335bd26fed3c218b7c40a1546cacee6707ab2864c5d0460bbf1f1c5fc0b82f20582bd47a23a683aa26b826b43be27eacf17db2fe08e66ccfdd141ad58ee623fa74429a425ab2e311ba6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha99c3020ddb7d8b638b5aec16d47ddafe777d595296095b45fa40820513dd334a5e4572fa7c3482732f3ef682fc4893779ead292e120d7494dc51d739a78b25d6bbd2adc870dd1182d78f3c849844c64b03e54ea8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e92b06c5c4f68830fe9f4741143802bebae24b12fe8485d4723ace64de33c91e8090334720270e05050355b5ed2158f00d2534936e95667b80301bec9bacbb0c4dc3961400af337f9a9f186f28565f270dc59ec9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfac158d7a13e1896117d30fc4a711472e16dc8f3e079a88dc7107bb06e66bc697ff6f37a7534d08b18705e215f0062082ad0479debb09b564ac2c915cc575ad560fd3223a6dc1ef7b5b816b5f0090c8904234831;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5a54a28189289357bb7af3249812ce5d420480b264208ecea69cb248f82b8d68b9e2aa03ab87c36fb6db587e6efa6ec30e3a6f4e9ed21b8461b2656293f80885b8380e2f8aa4febdf5ea37721c42894985c9ab34;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1eb5a4510b2dc393661e87f594a01cd04a509b48778b97d595b2271d76314c08b5528c3c3b18b33bfe1b5ddfe32d7faa06daf5cfdcb84d58f9b7fba35c26a1c88e12daf376f6afb6e0012f9c830423a7eec4387ff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce21115f2a8276f0eef46de6d7754ec25cdbd446518ab7b83ab92eb62b1bb21e8ffbf2d19a7b8d2c7658b723ce9200b60a45f66362a7e89dc102f6c10efd6e7dd8336097a39b2ee425eb7ff078e5aba4ce9114c8c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e0b6ecee8adf2c67d63f095636f0ea51bd6e56de017aa0c16cd747f822fc4b566c0eabf95567046525314fc73608fbba19e2e91a3d9681543410f2ba6daaf875aeb85ccf2de36e9649702fcf86ad5d1cef9794ed;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7c1f0ce54c1382164c68ba1b0d6e59d302284864694b64b415b3e1e4657a741dbe26764d4d71793b9bc4921213544ce29de12418964ce7f42ce45691dcbd3c74cf9a88f90a48e5865bc6ae6ef375b16db4f866cb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a77a82175051b1dada88e372f7f76f41988af9fd6b51369e55cbde0d0d54e486de292962c766bffabfbb95a8c3684a51e24c2ac32a71f601f0555bab3557931f65889f776b5d2af842abbef427dba6e1910aa52a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8a7c0fc85dfc87ae10e4870394c90cd343a72ac67d9890332a17e096d64514514e3a02f58dedd1b008f6c4fc8f58db9cac678c06290794d1dbabcc673dbd94630d51cb9f29f611b77dde3f7c986981c64939ff8e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2c3b8f9fd09b2c9a27c687bdda6c9d031a5f52c29a03182266b601c5afac494c94843cc8a37042701c41d42378aa9e74db0da38cfea23b7905860e087935139a2e5d83b47cbdfb140d9b40452bb69747ddb2c998;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76303a1db14ca0f7cc1acff3a546f1c114b211dbfaa9bfa4ceea094b50d1ae85ef3bb40f345c7903ba63e65c499d8b142d0b8f786c9d6abcf191b38a2970393db958c872626399e0cd34a36b8d65dc5507685e4d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h262a6d1a38081afc37479be3e145bbccd52d2b497eb2a8c8554a27c5823582a88773c8074451619a5a343a71f64b96152c8c07a909f5bcae66baf41d7468277a4e060b4726f0334a3cb421b1b0ac519d6291753ce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18ed4005f3152b35c290c8e13201883bc9c41b7e2a1b01685220169ae9d59054dbc3db53e8b82224e2e0093b029583f070fcd99f7cca58ce339ca22fdafa144549f3ef8bb8b936d8421c88af71f6e64d7ff1a8259;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd09509787c4cf4e0bef3d3dc616d75ea819dc9f5fa9b055538a3cc50840aecea890f2ec38964b9b9f7458a9217c1977cde3dde16a9cbd152d5dcffc6b9fea1cac889f182b0ad3dde1da5ee8b40e0ff4e1629f8ad8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9be7fe36bac0fa5ceb2869efa78acda16e5b460525d0e501a48a0ec6480e17890e6634a8a7380ba2de5a88eb4e061b24ad91512db1938cafdd89f6f95808053cc2b51dd48e894c94a89d9b0bad6bf10998d2b995;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h136daee53f24ae8d0fcc60af43be51397f70302d2f6d72fbd2e7e10a45e5ba0f3d22d392e5c1fc4a45fe6bbd9b65e456143eb12d3dbd28a1f4bc145acfa0ff39059e4cf3189c30ed58c68a6d594f9f7e5825c8fa6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19f401e05702d69d776425654ea7dab01d47a251115efbbc13423791aad88280c1664a970a8ccb9daf03872687eb202895b9de5271587a04cb5d783b5cc65c77bc698501fba1ce8b4f3a661fe8d306c533096cdf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac73483c5daf84e772211c0cd3b3dab1cccbaeb92895ae9d08fd1fb8d42ade4105001940046749deadd2d30b73d83cb9482d7327b01fc492a82fb5ec78eb7ceba99d25a55030eaa09ed1dd829670f18c98e238fba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12bd8c9910ba87cb567851c7be112b1b6f55346e9bd28d93bade544436043bd71699caa0c49844047a1b85d9917e4cda902196b1414c117e150b4bcda9746533dc841511e30be66ddeeb5698c4c10e850f003016;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a6792cd4427d7ca346d92dbdb86c2d169d3a4710efacd8524a98ebcb2ce585d1d6e0cc94ae485f65690909bd42a361efc76f75e97dfcfa9536b222f704f569f7265ebaa3b314f43cdc8b181da39c6caea2bc8c21;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4c122b7adb4c9f1f0b86a287d6e584d4b2e1d71bd48d0b49943bbe4954424955e249681f80a4d939be8e9e9de68747e4dda519e9e60ea245f67ba6f913648907463c3a552c80f4a8d000bd7545a605f9a3803821;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h225dd93dc4edd6d0522316d79e9f302a6d7462a48fb2aa3425f397dbb214c548358db985e0347b458461b045e133d3fe4b57f74382bfe7be4004f123be9ec9601c1bd5eac6d37ccdab3938dcf123c27361522ed13;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa33d9e906c4cd3613855a69a0fd14caf2c13cc33f01482bda212e56bac8b1ebca3065d2dced38e5856b1d13b2372291cea542f47c080d63bd5296de2936f8da67fcfc3b54560e29ece7c0590d51516d2c3520ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c5947a385fe64abe4599913f797e294a6bf556f9cef517cdd13e458ab5019ac6d65ba9014b3be272f09841f23f4d12d95e10261f74932ee2401984f6fec07d8e211ab8cac0b765ea37d0158b519e2c5dff5ed4bd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6f69482c6216b53167efb8dd29ba3d5070f1f85747749bc2aebad121cc1cc3e089f7f4a783c50723a4d202a8446029f7d6a64cc1c4f38ba183b2aca58719d5f4d24c9f31a8d4f8232d4769924b63337003ca6e53;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fa2be544f137f1becd04547db63b5fa1dcfae0807e15b5e3917f13216eec39be230c6aff80fa4ee56344f76d18aeef45e6002085e1b1143772b5eb42f90da5548a98d5d492b989b1e2205fee90a0ffb58b95fb76;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h956ebb5a12e14c713747a1a606f29b35cc347c883d114d4f37ed95fed0c429b054ef01304010fa3736648c0468046f64a08e08135c651f4ed5cc10fac711c74f97635c7b2707c653a82ace8898927a3bbde43b2d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3dcfbdaf780b5342a994721e9e9ee59c1ce20cf72cda42fe791b4a10fe2eccc4b7191ed25ae07adb18ed65a83bdf75cfe538d1a65b70d96bcefe71fa92e94cec0f72001db8db7897828730102a907b6a50be45870;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac39dfdc1a9dfb843c2e76d2ee79a74e40a17931da49d09048755a6588c1364ab1fcd778b5ecf03b4261610065dcbdddc17833408c388951823b91c73ac1831fe3858c278b908dd046a4de93ff7a156eef2e0977d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8385559217e3fc00330bba053046ef36a26822aae8603a2b7bd6ab66e70f950ffd28416a22e0ea354a33affe04e02b6be3a1dd2e9463cd421678fbbd5d3b66ae112f2054a413518920a86fa7a46212f81dc18ba83;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1a959c36381e138a9e9fe9f49d16eadb53f495f3e5cc94c04eaad7fa196c6b0f02d4ed4fe225a40043098350dd403276e53b6d3dc25236ee2f9a3cab074f645dab83a0e6815fc89365b9cc5c0d4ab08c581bd874;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a250ad35c66d09e48595d69c934a79d1c94788b336af818b12fa8795512423cd05012ebf466aea50bfe22700eb3312adac024f4e08a72700dcce93d598af24b10d979f91381771290a2dd7e1955d3b86b7d9fa8e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd6acd826a23e7f508a02f7e803a9f344400cfc37dfbfb06ffeedab8e95812d778000465b8ef3050dc6ad9c5f4ab2f849456073650ee477f78d4e51c3c9a95e58258a449b5065ba2789fcbdf16be84234ac5fc419;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a6057956a038fc9a24557d929f8bcdb18cebe1be7843b9f0f460a21bbcda45c0c7dce282d0660e614211ac2444d9f152acb880689b594b21c934587874d184bb51991b07a9c84167e0526d73d57efbcb9e083790;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93a0af2e57b9e31d269fed10925cd20fdd728cafa837d0f09c188d032d081efb04c1eabfb2b7f11fefd37cd0d73a75bf0da3427c47d160adafc55dcdd13a9e97787f59119895149ff051e106a289f19f47904271;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c50f0660e5ad39c65428a6bb302f92aa146012cea68a1d50e73fec9efdf053413d2a69a4fffc9481b135bb890af06955a72cdd556954603ad8f86ec67a0552cbae63b410e35cd18c3dc19921a3ff1dc477aa80e8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17c80ab34224c429425d0b25d70197d51467da497f0217ef340e8fa889d8e29f43a407b7d09f78f5b78c73094e6471fc728303bf27f86428e4ee47bee110b3de35fe50781ef6b814db3f0b82d44efa7051f1ea6d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cdd514cbbf4404e836d325c8047356dc9935b719b7b498b874b7a968403173e653fcc6381d05eca2b818bf2a0a0eaf6eebb48066974beec3578dd947e02d214b777309c8b16d7245696a183f65591dcbc4ef3e29;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0b8ab371811ef55206ee8c1d651a453acec14389fafe3a5d934cfd1552484bcae948a577b1116dbd1e8a80691cba74fc274bdd9333bbeb75ee1f228d8c9284391663def131a05c1e088b61237266d34164770d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca2c1781cae9c3f5f7f3a530f793f5555aa2ca3d1d115ffed1e89161acf3a65f43421bec95042ab70c177cadb85a5ea2c9885340bbc8c55a3989eb706a5e5cc19a047284738e62ea3a586382087f9c8f1b4b15bbd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57ac8a60564cd885634a014ec5aa31a1aecab026350d20734464e92e2f2ce887fd1dcf699be61429baa01d4f14df23a492de50203b88e5dfab901ed72c4fc77a46ca6d3df0652989e07d52f5394463707d6672985;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fdc4b5bfd9b941bcad8b4d378ea3caf6b97f540e0382fdbe657de890ad318de1afa38a382b58c317eb429ce81f6978d3eae294fcd8fcbcc345c4e4d2ee4e00edec7f8ae9e17ac3cba93f7ec07e395a946f14b489;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc260ef032bc5983a1f922590428af1d98b3ae4bde1b5537586cd84e2b3728f71887d1b410781bed2a63e91bbfdae895ce477163fb3cfe1b5ba7f45ea5ca1c019bd7a2e878e4096930b0637077507d96d5fd98382d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d9764ec75baef88a8d5a5ea0b19e2ddddd57d23418531f584174e14bc7e32e3eeb11c16b9458e5b70d7c01dc5763a4295771accd7ed55e5ed1d997a62b7e85aa226a68d4dfe4dc846fcfcbe1b0ca95d0f077ecec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98f6b581036c1d0d47e5bae94166498eddc5845438a8201de568e54974ae485812444bc243ee9608c090068311034b13aa577cd63bc21d6591a86df2d4ab131e08d35d03a294fd59278a6e7bdf4d3b9604c310288;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12d727dff753fb07a69da60686c5e140c3a66b826f73c7e2e8d2ddd020ba3dc6614528b9b574e22e1b79e3a470c77d75a359f9a3dbb512b4da07d761952ca1123a66236c83c4cf8168d11e97afc7a70ea2469be43;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h605db68089b1ff0d341dc7c48d21b3ca711381100624dc083425d88750194db0d58dfddabad701c5a01261cc0db3d4b1a90e9a12f5f2f075e5772794459eea31525b0ae027e9318fe84b046977529d9b37f5602f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91b4082e8d70f18e7568a45fa23b859ca2e07e82bff8742e2320e9c6f0dcab9df3edb0c24eb0f9a8182b3035e14522bb1ee7e95ba1a72579ee1ad9fdc894f9cfef639ade5f511a48a9d81917274006668ee91f38d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60f8bd2338efa07afd8c1feaed0605930a421f54d703d2f9871a38c3d5f147120b5b1c1f5295e1094f5bb0337ad13043e5de958c594d72e8cb33272cc5069e57d09b9a21174f58ec344c6047a0e90ab5b8f1e32ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h356d6139257950151f62b588150ad2dd8e3c7a37de9205518c9e58d1f7ef673e69327854ac7056f5fc56dcd2f36fc65deda31c46d2890f743bef23eb16eb6452ff9515923db425ebe05941286ff12a4ce617df2a3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hadea239c7e1518aff1d66006e0d498d1f90340ea1823e4074933205c182713b54b59744ed8334df577cdc28edb50b59d0ac02f730f9f8d985c1b7655385497b093a54224779a8b02cd54f3660241071beb92e17f0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6bf83b2d056c39f82f6849a53425c3aefaea391efa274072d0c1e4f45f0cd6e1d861ae0d20740d159239ea5e4de4d2c28a70812a47cf5681ce7d039d2e766216d2abe9f9010360b78bb53fb5dc45c2d278b809a89;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hecc125c9518d3f4be3bdd8087e9d773336ad1f4c61b7dabb40f3d4f3fe6816b1bf4732bc4b58a06bfad5d756795f8da4c5b42719675c335691830ffb96ef6ec43cdec8f5cd33c878021d43f849b8516fe43fe62c9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd02f75f18aa28758a753f8cd1994d4ce6b58904c801b5f55309d0f26bc4dddd49e8dcea0fde7add03b7db90bd770b66715d3bf2542b3b67ff73eedc8fb6d696e05c1aa07d608b765c696c3fd823339620a5e481a9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3681701c269e368de44f471222c7356fd3f8bcdaac8f9998b4794a0bf6aa1a06ba8656e23a4e1b6cf7666b6759136b37ae23ad55ba08b3667fe9af585a7ac8292bf5db2520b04de0943ab47abd9b03f6bdb0b6dd4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdacb24386408ac7ee1cc9e3948ab47e882780d68a2b86c9dd2c2a1e820257b1129f19859acf6647f2efa4e91eb26c81e76e026decf50f1bb2dddcf5a7e2abb9953b778205d4cd83ca78e44d414ebec187c051ff49;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54fae4606f2cd0e3ca8c880f7d9004d316f37e7c8055fe47fee81500984f703c13071b3ea570e14ef8120bcac01280661569c5dff7f86d39ac29bd8b9765269885324a5f54ae31ab91f6c19f7a1f50ad7bf777608;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61df5a8ebe93d41c7888f8a5065dafea47a1d453ffb9454468ce3bc5c9988035eeaeed4480774e161ce235b1dd457b8633d04fc926cbf4424ef1409ed8e8b94dad94bf0ddb8f497fbf8c478113e181b96872adab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb60fb257e3701230796f23b72c0da831579496aa4e2b5a6d71343fe1e351f420eb93c86afa2aee1769a3cbd35d4fac2cdc8738d71b44e324ec805885072d5be1dd635099ae245f975e86fe3f2818dd8a75c942072;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he88bb9a46934d11a2a815003978e19b43f6815801cc207d09ba45fee8387d50707dfa723d56e1877fa050fb0debc8c0f8d7b61bfc008664a5bfedeeaa599cdfea5bf04d67bf2f5e75e0a146d7524eb8cf3a474ea9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha781cad4c7b7dc5e3f92d72c5a1686df92fd33e2ea7a33a8f67c56e0b4fc6d0b3a6df4d9cfdefc28b5604616419a126eec4ba25975d1200006654cfc7a4e4edc953b3413741e6bdcbfa88358536dd6801c4bc1a50;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h738080834b8c1e4b1d31a662ff065cca30d3b011943ff7d5bdf98622ced9b43f89ddfd91c1aae8e21ff7020c5ccced1a0988f1a532d53b25b05feb2cac5092253065535ee3869c618edc246d0510b8c44b627df1d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7447d773cab4a188f298bf486892d1386978751a4c702a69c942c0489753cb659131a8a38679a5b457fb784a3474e139aad4221349d7ff535ed62cca99e7f8bfd5fd4fd9403f5d497b148062fc71e52b04165616d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed80dacfd59c7145ae8a34f6e84f87cda73bb1bb988f8d65213fc037b9cf793006e9dd874085f61df5aa7fadf66f79c864b8f877f779c2f0478e227140ccdb2b85efaa027f07a3985b35f75b3a465bf9dcc8cc5b3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7cd53484864279793cce20b95f6df283258032771deeb81097fc92ab60db05bd120f391dd0c59dbc1fab0caeb4072c33e06e965fffb51ba19ed85dd9908789462eeca6a97d4fefe62e31f170c7c1f82ad5face7e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9fea919189883343994abab404e3a5a72c1ed9f0f8de32f570ed94e6a23f1d1fc402d0fcc3ff7cc275bdc5bd40fb8b73001d04725fb6af80e9895def9ca43dd29e9c2c6981c94d7298ec1aff7262380ca4bbbf27e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he105f553f5c2f501a9c10a03ba550ee2e7a588e3401b337082ade117d01c763bcb44b94f213be92193300b53de84e5507aa40ccae3aeab5b6b672a4c9bcd761fadc4eec17fbe32b19fa8b9ffafc92eb8654651c1f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55acb9ff03afd8a2970fa7b133a84849b744df6520fbd3c0db519c9aaeb4a5db416224cad7300588a7bfd85f44460c2fa6a3cff3e102b0ea2bfc894774dfe4ce2863eadf57e086f33c637c600b0b503b82cbbfcbe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h278561b763cfe4975e9fa01c83d94fd9ea5fedb5f4e7b4b39666383b6f4770aa320678c82954907c277c7b3204dfbe72b4e42bf09f53ffb0dc6a7db72be5f8b181934573ebf7a95e42023cb7db196d23f3a00e1d7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba13cd4e95e62bd38f247aabdae10a52d0df464ba4b7143f670ab8ee45efec329ada8b5aa6b2a86b6fc6fd8bda103ffbedaa1d20003568c3a3401de5788a200f3ae5ae3ac90f11e7934e61ed161f5d24e92950354;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2e90feb8cd4d4300061b84fe5c6ef072ecb70c34af1aadad0184eed011283b22ecb15a322ac51336e5374da8ab7da826b95fbef3cb335e759870283910e4def27d1c6f1d1cf7142118fa4874e344b3377151de9e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdde8ec178dcde824a4d8fd4c484e67a3d893ea9b92a58e492296e418cfc58efc554bb4af46a49899bd8be04d8f807b40c95a54147006d65512d0a2dc6f9b1cae496dd9df0e440747d21ab58398a5a7d0f43fde68;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99dddf596fe26e0893032444bd97b41ff2b80a9494c2240b2118281da7f3ed419f788f33b26da26a40cb9be256d6059449f7b49161ac31970260aca3b1b3c412d0e81d4dccbefbe78e411826f5c847b9bcf160ad3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7f9984676154e45cdaefe582ce9e980b31b24f32bb4f0545e95726fe1548d19de2e2990e67f36f835edc66b0c4372a2ace7cf0e114c99157a5d0a9d261f027f7584be2bcfc739731fe221de112997c8edb86952;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h460f5194fe42c177b03e8a4a72f7387816fa166b5b15234e04b3e05b6bf7eeb90a98756467a2f27e009d9884d1d05789a252ee2519cbe1fc4300476ccefe91bc415e83a30d7a3fb3e64fa66184826825fb47623a0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6bb91f3dc57004caa7b393785678a97e96afabae3de72793a118b4a0d5b2276bf584d5f02199cd13124aa842f50646547fbd36714c5117820aa01735e71c71b4faae98d28ad38b1ede03ebdaa831dc57dc2a4cda;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h282f08bc0914986ef6b45d370804e6ebb361cae989d7a701f9bbfbc03b37e113971706538e0c999b982da4aa11d522766b8ae72dabab09c8676ca6a4ca3b1574bda72439b1550a9d0e1177e46b05b32bfae6d4af5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15da5d614cbf7025f8fb2f37c0363270577a249d80fcbc28bc3b5668d3d54b0859ce01d2c8d387701b7d3dc8031dca4af0e42ada302cc298fcad68f50d410a8b3b659390b76722e6e8a260718111e55d6982bea81;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7158b709033c42c598df557b438c36e3b869f8f573a2b4f77b5964b35f206df42f6dc254ed36f7b85caf35b9e41cec72217cb2d5867358ef716b3c7b330d435c0217ad5ebf73e63cdd0f54194c47439a22f78df89;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddc57accd78e0af61c2f45a6a0629c727c301f7286ed1fcf639b25fdbb83dc93e121bcee94d4631f200fe17552428281a604ee12a460ac34e827bf2e9367298cf7c0fd6b8d61ccb0c4dc803fb8d320eb8c4fecefa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6535d7ec64f640b28db72ee0736c186c549dc041fedbb02d8fc694c634a3628ba3b488276cc18e03cd3e15d0175fb650ad963a18d3b98cf0091b4e2be8b8df2b8051c0d5082a4901eb5c74381d061bfd919d39a70;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57ce50759e4ed2c630168fdeb275531555ea12892125f162936fd7a94ba045708654ca433ef2bb28980da574c2086e15f935f5b7245652a7e0a4f37c50fc66693ba7b232d5a60bba8ff06b057fc000d4d02c90f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h273b20204b23e4f42f4db8a01b06a9145672ec9e59d3cc371984272f89523e548c8abd3c9ffb63b4add5e85bcf1195749a46acb479f5c6a892844eef5b3d0d207aa1596ce631b56ea09fc2e56d7f24b496b21750d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf975e191549dde0ac23a467d33964dbc8dfa3e2b06188dc6a5bc28b4c4799484f7d230a8781708e99094933ac3b6137abeed1cab1d7132123b86293a248e70e93cce4a579bd95decbb60ef9fe83d3e59c7cf5214;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c9b3b15c55eb1ceee7008bafaf64557660a6451cc03a1e691f4bc9379eb7065edcf93d0de996f24472be5b71e1f21b6bbcaf4b5cc693cd03a917903b7f4c30f3cb9404daad6cb1de9ec7e947c2b6f4ef8e6c3983;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd80b9d05a8494398b4ccfa7e73828d792914f51b119e7628999b8b30e0faa42799a2e19264c139de5fc2124b7190195e3872a5b36d3967b808f9a9f3d3736b26c0fde486787265efdaeb3cbd869c9c40e11b3733a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e7914d19782e1f318a0f1f8da677277e7a7a1201f728a23dc97cadcea03b19a6b656b4da1477d1f933996a4701d538267bc7105602c69dafc595f0fa161cdd84602193b1e6717b32a52ba5c824fea4d77a7a8399;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc690708879e41b32f18f8462c4474862e856a740213579a6582954562d72b4a3ac9ba2053e3c4ae4489ffe1ee15c716a7e08056333cff679dfd14c72d5b890b89fd42b9fad18abf0fcada42af7566fcb8e79b883d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2647d1b7e2650b7be500c21b5430d9fe85dbefa596cb7dd4bd170e010f45555fcf7aea6e6a63c10ec216266d5898ce252a1412817d1e662945965083db83d2e53e2f806d23ab67ce70d19ac9fab58d6824214ffa3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h361e89be82bf5f600b1ccbddb45acb2486d27eaca95b1ccbad6fef9348b1da5275428ee5363d9c80c5f5df7723effd5b53e792562f38a9d9b0379ac7d625281aa12f7d52c8aad972e3449382ed8233aafd231f0ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51e945bf60edebbf3d1f19eaba94d4f45c0768d99503f9631f2567a7264aab7b8288f5b65d19c5eaa95d1aa48d37c61ba353f2c00ff5c9630ab7ff668eabbecd024079c7e8b334e7bfd8ffa336cb6bcaeec4f2c6c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9860721dcc79062590983f565fc9c32b469ef97cc2d7fdb68dbaf8b896519c20be911d2913954665dca3889df195cbc64fd0b8203317d5aae53e637fd036e267ce27967ab7ec9cc058b9dfdb7729e4bc80b560a89;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h239d044c8cd46041b84fc7f4209eeaa27732c529b7252e8a09d81e4f021e1b19585860af5d0ce41ff47d8724a26c43829c2bc4becf65369a5e963dd5868a71e141a668f801655a4d330701ba3eca23248588d39;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h750f6c8b0b08305e4df9bc7c1485cc67eb87c53f9d97c0215fae9f928b3fd50514c3cc91b42b0784e13839b122cd52ac351a962bdcac24ca7ecc25107e596da9a5d5f4f4a782bbb597db3a873c3aa9a1ba24165eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf011e09a96149ecb2745ab3b596a8c0f326c08a3385ab8d7a9cbbba3168aaed4a5b164bc98e9e588a635652181ff4cdefff6b8a31c3f78743d51f727b513a3550a683e1f05f0443df8ad150a31dc4a88c6b4368ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3087ba5a5ed603a9dd026832a815ebb6312c9e0969b56fd7046639f069859e630e1c4e1404fa032e951fe335e40c2f966de032f3897e7c2b6eece6212e936201845443b2613cca8e9701e466bbe243510de37b68;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8fe754f2e585825fb6b63fb17b740bc76a73d85663b2284e733730a16184ad5506b9ec92403b2b69d9f3495eb824eca0ba5e00e139fecdd9fc9d6b73088e7689324a6686af0009a6bd58dd515e0be813c0407ce24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3dc6b02797eb0ef94ec8e803587ff92c4bcbcf6ffaa75bb7f6c00a3f39e5d533a6003c0a20263bc1785587b05352bf87b0167b0de240f9c61973380e4a162c8728a788d2bfd7d0abb8a4243c2bd0f28793828189;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc96a49c978325cfa7d85b1280901454988643649ef84e3a96a2c5e12a5b0985b8c6456a6ab8046bb69620438fdc11b9fbc1b3f29fb196134b73fac768113916382791b8c692c1bac9d12d4746bc2ccf3acde296c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafc506c7a538d3e4cb9f588cca207378ad72ea49f09a330afd815679938b8d6990d7c961e2116f470fa4188aa1a6983d2a757c17d7adc8b61cb1a2e86df481a95a753b719f18cc164bb8def44d9723a43225a4388;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c62c01817da029f3c26fcabd51d363043681694b70433a648521f5e053b2c1a24efa575b18748cec521422496b911f80d439a07a941f6290b499fd0220205d7e262fba7b055a4e40a3607f0f0e6303c90bcf1f81;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6b75f5ed5ca76b2c1f2a76535cb116b2251774fdd82862dd25094581bb578c9e968ac1a5f2b5e5b6b528174e063551e56fa2ee1b717ac2cb323a3dae7987cee5c885d17c79d707604895ceab1388a9853a1f587;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb456134a6fd6324bc9b9a598c6af8a1e3f258264c18d71ab89349d31b83d25ba626c8a47892e764c15791bd2b5bef61e367882f2d0ddcaa160576155fe74f0279072e4d1c90454234fc6d76efa5edd4843f458a04;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d5bd63522ed024164cadeb327cdb2248706bb8e2b16347a652dfaef9ff420e428572d80d484caa0c0844010636a123b3354e6a981fd655f698cb4f204731ee2cabf00512cf215b6336cd9be04428746948630222;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b719c4233f43e07f2b88cbdfd4886611e973989e7b6699c240f05d4dff1c6360d925af5c4ce933d4d521d6d0ba8923e9d6aee1f14e67348c5e59ded963089cbcbc8e2560cfed0bcecf7c76655f59149dc14a174b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heacf90d8f748025b7579a1f0f0069975ee91c909edcc3c75eb9900bd963a89561e2e3522eaf5864deb8cea856dfebc8e4ed3dfc0abea9f5945eb5890bd49ae997ed8d665c8ff8016c6d1e77cf086e25e6594002fa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26533144b8241d84b765bc25dd30743dd8824effe4f16d3301880271e9fc1d2d095c4bf998556e8878c895a7874a6a94dc416e2fb5f753ec68cb6a6e3ae358c8eb9b28e148fc912a6b40dc11b04f934abd5fa359f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93b2407387b45f4ad8fe67eb251b6e19506ec0ba51de74bfbc3f3903f34a42ea8891aab85fd3d04feae261888e76453ba2fc4f803bf693dab108dda914c1c9ea3baba313593193263befe92e47ad6125c910d383f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50bd1244171da4f9a853515d81341c1a2dbb81d12909eb3e79cd619b03ea7c0cfaa107a98beb2d4d83d948124c68ef86f910ca1aecfbf94593675bed7807c4f40fce1eb23c177ff8bb462135c58119a9820315b12;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52e6eb6e042a19a6591810805ce1dd89c5e701796839e43055c491cfe506298cd6880b47fab3e6b47e8b6ac876fe01d480d19670e30e1f7d1402732c2487450f53ceebedd72d4fde138e858f8726c16cc40c95545;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61e4ac8845bd20e06989f40b97e44058de1efa350706c7ab1131a50f8cb8644212a91c8694144740538c2aaac3d7b948ca5d0e2b5c37784289667b71f1339df9ffe3a0a66c448565fa5d6d65ff885c5421b4f82dc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb29ca112f52899313db36832e84e08f2f3bc826d861a5d12702a543f596ad47b3b8259fd451544b80eca5ee4f9be423f1c15fa84c01b3d3e0189f163f7edefed7a2f28cec76233e5f684dd0c9bed6d56741008e40;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0510f20fe860b6ee640cf900e64e73582a6310db034d69285c3f6dec7b4ea1676f8978f47fc1945dd9c7c08dee96e43b517f9349df7cda20f7540a0a618f89a72440821ea365467864dda734447c3e845b751e5d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h580b8960473ac7fbd08c7dfa2fe31a13148c0738e544125df9a9dc650939b94b158421d6debe4f601bda74d8350c14eba11f4af1af1feb3aa35623b78a05c77dc68f8d599ecfcfc5fbdbc3fb2a25be2994171b403;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h516586951ae58279fe8b8794bc58db0f9e8fe6271aa523a42600b30926934b41a9a930056c294584afb2386afccd5506f856d60cd8e72530674f365dee1d514ebbf625c3c5f4f12deab0fa1a18ccaa34093184409;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h427453a8ff9efae74d7bc6c3aac2d6efbb36b61afd97b509e2c74a03264b7c7d940eba09d99d9a6244e4801babd8568dc9ae8456b92220b5a0918f64af52df939ccca704d2e79c09f850adcd439d9c51dd1f9fef1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc5fb3ae276f17f5c83035266f08a4c137564cbc6ff4c19a0391a2228881d432ba95a2305f7128cbc7f2324d9e377ff56064a942e690da74bbb55c4f7d041834cebcf30b3dfe9d162528dccd77f174dfd059cb973;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf808d791c397651fb556013b5ed09110b002ddeb1c7663e78aa491f1594e2d432109b927d3ee6db58d559748a3f1f6e7fa77b6764bc2963336404b19136a82bfefec3ad2abbee5a4a13b62f3afd062b64c90145a7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1010d8eb7d8af21d8f759db133630abd73743440324236a0fe7f4ad4f7bc5c706153eb14d90bb516219f824e8ab3424bf622a1b1ff536b6a16e84ef0869c227fb13db47330f24d4c700a80e463f89a6137969fd8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2818167b0d509bd3273a5150094955b4ae7cde7de53bfefedf3c5094cfba3504c624cba4f79d141e42c7e2e853e422c679687552a0a5443c24558382a0805db5c6a3352d882b17e58b2b79dcb942431c159c0ba7b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2a56561856369ab52199c97e4428e9e8bbc3bbcf34ce3208d2dcb2e7cf2b0b061b3c75ee2fff4dfada315792feddfa885c3e66188a21358b0ba35e46c96b130ef67a7896dff6a8686f1fd32b1de7d4e92d56f80a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc1faa2b55cf6b6fa01adb6e7ef73583a2e268a23db690624bf5f4c4af9b17538da5c0b8dd94085d8ae72b0c4646ae7f89d6975f5ec5690009c716fafd25020a8cb2a80d434ce96c1611209ce5c9fae88211d3fdc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a454b3b041e670c317cbf2b3c56ad96695330f978a79399fab44785b9d76ab65a11cabcb65cd964e8b12a35f2bb78b516a81a0c65a8a936cb0530d96f40abc3170d2294141916f324961da30c5cc5ce93ad92a07;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h494c6152e24833b0821248fcca3830e40c5d4892a568c8ce33cf3eefa9ee0af2bd481192aa0112e7ceb57f9b766147a47d539a9e58c80f76ad669d2d71f4d7d5d9921d30d8993cdb8a9c0aee06e4a09693ad7faa8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c55fd4d5cc92e0d15de32d961ca3ac210f525cd09b3638c47251a2cb6973dd4b5ccf052596020e1539ea2cbf01bb705939388b7ee59d982f767c9fb3399b5d3ac71acea787a60c0bf4504c08a2de48cdd545d5a5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h538e85e4d5e6c1d6a8ff0ee8271dd886068dc42f4aad6abf11d8c1d4ac19c59a295c215189a44a63bf999dd38ef54f356b6e37cfa2e04ad7047f884f06b235c418616ef8d843a53c7adbff6f6214f4a2038a9fd16;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1c8054bb1005dade456aba9b213cbb571157647715be87904142b79a373aab532803d94ce7a668dca69965d8806fac81dca6a42e6ac90f0b4e8999169af70e8329ea19f94f6f864f6fae9959d826fac71f09b59c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b70127630c68aa3c165677c45bf432e224dd2aab336fe9e7a64d61610bee1e56a7e752ab4ed4cee37ef6b042ed818bd4b001dd2bc4b0af73ae1881641d5939f8acd90e7574aafc7059db73b3930e3eea70adfca3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d9911b1726101fb1eef0c8b527514d1ac0d77d186e86e6e1f3d476905ba458b6a5d50a7736999d584688f4149d560381be85da4c2f6c096bc60f5d0140513858c967ce7e9f24d5776028a254d42006f55bad4803;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he726536c2a1e110caee7eb773ae6bdcb1ce0f4a2106fcda1b2d8f20775e60e5fca2c27dc6fda72dc5fd72f1efb1f3c802a353beb591b426aa856d998c7b50fcf56c5fdb6a4d9287656191bd2d3a24b03f53f95d0f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc2a8ff416f4d8aa296b18074db641bcbda4a7dc1b33b70054582c3079fc4dd7be0cee0db90e222822e2ddaaa6b05c1d49a57fbdc93bb80eb1495fbba345629c8de55777a82edd52a683d1462ca02ae595a2f4712;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2460e3c630932b885f01e02b37b7bfde2d8fe6d7fa87851f3f1bbf1c21f298e2483090037a1a29963773f40712acc8147669cd1ac54bc0f5f9a34fb42e1cf5dc52a42175dae0f287c24eb1d33aa5e5b59e28d8fa7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heda04b1db6e7da0305669d58d59d137937daf3846258ea2edacd01f66555deae0ead4559c0e25edbcc4c9f289e332297f65a2ab2c8607bec283c2b24935795919ec68a78606319b47cb3f1513dccd50d30a93c7d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h644b1156ff9dde8fac9d7dd1c74cdfc88c6876de23431e91b8367c44732d690762237d9d147938a393024c1d50aaa44c0f53789b4f2722925cffd959fb122349e16199f5ab6f5af95b7ded55a54794f466c5f4cdc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h628785950371e0fdbd63d638f44943303788a4bbbb06c9bc5b72c2b8d676793c09e9c9360ab6c31ba44d5ca2712d7026a26c7732864d760822e5bef2b4bb07b8d9a0f2c6b05bd79864f532e04a6373044243fccc6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd17fabffdb85bb5320dee9afdcae18fe147f05ec1d81ef8920a83dc00dc884b5b9c0c4a505e7b09da64ab6e55fec957974a5c4eba0be18c2f5b2882e7c0a24eb46196ddff0222ba8b10b14c86b19754bbf52085ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe10d1a7b8baab3398a104fe308004e91523713ccccbdd17b9df3d6ce5a9608be5a5532cf972f7e9a0c4dd9670596b75345461b25013c75e6af9b22aa9016d621f0843c44f7229a92aa8a69a99340d3258ac0b792;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc09e19ef3743d20e79423495045e76b4516c58f8fdc120a7363cb32730527cb2bf218e8d140af0f21fb56a9e71dea7ad52b590ea39564db09c8a62781414645e0461823a03dbffcb50a6e573ce64782619e5b968f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ca97be56f57781a9896cb10c6a2682ca84709905fd03ce1f550b37cbd0e2cca67807ab344aeafa20ce512b9b803bb8c34a61fd8110cc3e5f65d7f322117fd6f8c7eb47eaf69216174a302cfaf749bc4c0c209872;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f8020135b2591accf8199f433da1050b189f838cc1d67838738d3c42ec0ac74dc289e7b1f130e43d943b2e39e89e139a068f706588096ef05b5ad1ef65dd5f09b961168fe06ca500356dca087fe6482176895672;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7bfd24210d9632a4a2ac01e03903c8f807795d372fe0143f9550508ad7df0411fca7d5f62295d375cf9f2849904aa99a9beeac44455bf325f6a3dd98a252068ee0aeb9c92d0f73b0e2171b1893c7b37fff5cec834;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc09c47ac001c396a988977dc12951362b96df2aadb685569ab4397e6bb64b85e5f530a8fcdf4d6870aae3f5b188ffe0282c32f6d39a25ea02e727a2ecc575e33f443bc50b29f042ff8f00ec2f98a5d97280ce7b93;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a9ee635b59c848fbc245938f30dc98f9c167b5e50f9a33366e4cc8e74251f09174ce5be206ff7691d9164fedd5616951fdc29dbdc86b2b007ec75bf1f84978a7d60e2ea73db262532b07c72c109e6d1fe6394abb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb21fee6e874e2650c091d6f93ff44616f5af6324c3930aa884ea6355eabc16e544ff7c194e23a734bad18a5e030b6311b7704643cb1a81e5428cc0f6efddc603425a205e5f80dfd8f60aad1b63f1d19f2d95e916a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74e104b186a1f386a364a7f47a37a0df10df5ef74a90ba33018aebd1d99bbe1957f446730343c6512624ed8dd6b23ce52536a9a1d9482835965cad09ae70722037cd62cff81ed08b306783c4dcd320e038d04932f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d87c16e4e04a2c9f92c854ccb04aa68289526889742cab7967d6f3755eada348e76c39decfff8b04e9051903f2054d18dbb546d3cf6d84f7b343758bef212288387a779ceaf384302ce933e03a70145a71e3b19a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab646eac6ca22ce5504a424602d378177e9bc0461d23b901c13a8733f6a5a105a5b827e5cf31f923514ea04c82ea07ee3bd8cba2775e635e2bca8c28ffa55ac58cb5110f50e442fd07aa570df68a39112997d3688;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7b08e400a6b67418edb0710917989e0498787becd877a26b924a02556090f698bdd1dcf151955a24da8406f8dd7322af06e9822d14b5ae04c8a4d183b2b94b48afa347d2580d937b6a21e751489fefb62821aa7e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a128bded6eaf0f551e531835553c6f4f3a6d3c63f7d4724f488088ee98bedf3a2690ab36dcdd0d7b628191f820c6846e910be2739449053cb91cfc502f1860c0f8060099fc0118484bdc75e8db51cb3a8c5f9e1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha345633be08a7717c2752ea3b48050b32f707b05fb5ebde4c2f90f700b1e750fa594ce255f591943bca6da332b44f1409ddded212fd423c063c5305f91a8f3997b87733bfcb9c1a8f59d75a0ef07c4ef753e19f08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd40e796ef2abd19e3168e5b6de0885b72dce427873ae9919fb0d2aeab07d4378b88ceae1fe81a55f05f59fbd67a08a0950d673a0b5c4ed700bb43992a8cc4797af13bdcbab6e74783109e795cd3a82c4d255849ee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6409067619ae5cf2ebfbb705e2542f69eec7366d7946157a47ec6e62fe8c868cce3ddf032232dd07206b50570b65529f2b88ddf878d8bfad2f5baf08c52081e9d382d036ba9bd0928e651ec3147ce9483a7d02990;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58450a1d9dfd17e0e76a200e2fd55ae6b50673555d106707b1955d4e75bb3a6fb0c49d5255239f70749644a6bca3af69b4e2aa9d728d1d6c5abb7c5e63f75dd987f5d7dfe75a16f853c3a8b4224455f61b5e438c2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h513a9f9d079a3361c4915bb41e054d01afd93577daecb5586fe2071b5d2686872d434765b9de8d8565b2d709d162bfed1190fd072c63b42b5a2d0ef5754c6bc732510c66ef90dcd4bed3b9e584d073f63df79ae78;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha467b1c96f9d370ff9e298ec678831504e9f92c40b8a9026a8f56dc953f835728ecc794971ba12ddaed03225ea34791cfa2407c52d8e0e82484ee521b108ade2de1fa5516589171bbc43d7a9cfed3a9e868e14138;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4fab49c79f8873bcc7c179687e3714fa77ac6c387d62599a0b6bc374faa80ff697cdf8fa628a74dce8f18391666d1fc48bcfb8695825272d0e709a6e5f8031e4b3509102d90a89318eb4331d95aa6192061ffe677;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24c04aa4880856476d8b1b84e5db1e291b50b77cb1d9f0f0ddfe414cb1abffc56e79621472625d1506180c8e85c4e98e73cf13155d3b356b4b38fd8313680dd2cb0b8b526a0ea39db84578fbe62e79b0670b19591;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h324af9269f30bbfc8219ab539cb88e13646cfe030070600ed8397247391f7bd5ef02d402070acbd8c684438497a8ad092dcd09e969b5c52f1aa6729ec1dd5b634ada1449547f6f8f48c220788db512eabd49f0993;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d361891f355a575e32b9187bfba424c688ac465c2ae0c72b77267e7f6f0836fadd7a9373dea041d254aa150bbaa1f44c672f69bda23df9cb3e94411d4f0321179b69292d82bffcecdc40ed099d809b405e3b2a32;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f346ffe6f7dc20b524e5e7e5ae31cbc7132421ef5d880e99362465200cceaf328d1f1ea0e0510f0ece5918e23a290a9c1c363d16017ee8ec59b594c856fe8cc990f67867b71d658ee641eeb238f6802b5c7fb714;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcad7756625992643a74a92826ac7e1c64ad717ab43328ecc9c62d9df8b5bf92de1fd73f829e4d8065931e18069d785417c6fb0dbafa05408c7433275f3eb8393242da62921365b11b4453e70db20ffd1f41e1b076;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57c9f9e64b87695036acb8888a9a9fcdc895e2ccc6a502a42446922063a6c46bd5d28c9b08c837a1981c330ac81d73ac8e287525c9c3f4f5834fbb936f896d8a08f8dd5be0a4ced1e27dd64e2d7df867251620217;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5235b9a2a2be1c3b307b8483d5cd0d15a061d404c91ba972f850dfd3d5b642cf36b0c60b320c84ce445b6aa7a02ada021423e2df33d336ab236695f72e10c93b9420df85b07e87221a38ca797f6ad0bfc8e3ed9f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9765790036d5266da69445c91cb480df05aca025eb5714b33b74e65227eca38295cde339c10ecde7435cca701a7b1d50f1034434e21ce2b319c0b4a8ea5826311d6c00207dade73d71c40831cc68f441f320e228;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34eaf8d7ca25dba96407dfad4e0e2e7984b5a10280b884f4571e0e8b460c0fc25a609afc8ca42f8adc244ac7edd9dceee98627a9ab804fa91f9413ba4d4412bf88f5b29c394b874ccb35c214fc19dc0d9bf4d8b5b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd42433b92d3a40e559d9753769fdfb9ab325235cc0c06ec19953299cf646eda50eed8031d7c3a7bdd09527e951ef1a5fa722a5a916285e4400a05740581716dc5aed019fae1a328390473011999b19baa88837852;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc907226db5bf4b0cfa311ec9c1cf77ee4f5f5d7a51b694a7df846062cd6391ad71928c9f4f3ee1f2671236808bfbe2255e1e6fc991705514ffb4947889c00f8944d8c5a2f497ac0d73d5d5a0dcf6c94804444f06c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c94f3fdb635d100d0e00f9b6d9d3bf8da8720c7416d0f1822d1575f2fa66538f549e6f857d078758096300d1002d627e9ee239867d05c2777ef0e24df34c7dbb3132fa457b020eef691ca870b68236fd6a2f15d6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c98bab0c79784d992431f3f7f6421824fe1a6f0aca6039678753000e39da9c4faee9be355b3b6dd3132b27559101cededa51ab94933bc83e55a946f626ba682ce71b8755a1555ae5515749562bd2129ec20c1b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba71d88430774efdcfeaba7ea44de0791fc5e90d5434c1d6a3bd9bc7844449deb996c6c576ea5a4a307d5cc27034ccc829db0f0caab77d1bc724f7f1a0a94adbf69e1829fbddde9400db8461035dff7f0f95785bf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c38d47be553c4a9f2ab028df3c566c0253fe76658a3bcd59c464e71bd82410cd9de1c81cea3baa43fecd929f73e2fe9192674ae9f17dc32531b0627a35c2a9dcac700c9b2b300d7358c3aa4d293678fbd731e528;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ec1f9d359382a36af59a1614dddc3f0f7f5ebfbf14594a28f079d29bea6ba49e36cc71a6ffdac47175476e54cc446a21ea8128526271b7d3bfa455d59c700ce7b3900c135eabecaf56a5e87b02eb984836b86204;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e70b7947b24405cecdc06bb5443faee80369e2b19081476923d55428c3b2c250029633cf1e46eabf813706e46862aeac8a73740a9d4712eb00fd79b59399203766e09325b44432cf7e140121de6d0db7620ad1ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee7ca8b9ac9937ae086b80cacba527bc9f2a60881f1faac3db4328400b36e5c927e26a93655d97b5177c23cd1527e31a8de3b8dd03347fb5d5d75e3cba49e666ab6f30726bc98f5b191dc6ac09d584074635076c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15c54ab020682a5988e6204ec92d6122f795309fa9f7ea4d10f66d333a09045511ff582e9009b56362efd424b63e483359b050458fa13970a6ac2c40ca251c6c87368283c3a7fb89c91ad472ad3d9d5702bacfa59;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb06703d059bb8a131e5cf4be2a31cbb9319df3772a11674da2513aa09e8a017dfd9521d6051a3fcdaaa421aba1632ee3ed7efaba290fe97aeeb672e4ed70ca96adce9c54dcf7c468014e638db71953b640deafed9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b47ee839b9f9ee9c14eebec729b44ace7341b34a7476743606a9fe2f2cf27d8d96dbe9b862275f78f560fce91109d238f85cc53530bcaed25e9cf9922d5a37ff86e10069e98a24058f67a27b769dfd88ac759efb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b9ed60f23c971aa3d442cfecb2c26e8a373390565bfa341b42e190510d0117a621d60b37920ad162e67a1aa22769d8171535280c16989bf9ac8490f092c7b9477986e4410fa82b2ccd1733927974aa26cde29433;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93348ca2b4483d1fc9989c9a53b6a5aae78f3cdf00407b8a5b574079344ba935dfeea35276e247e5f0eb56c77b5d2009abf2f0ab83233271518604a65b187d6c8b48730dbf30e9e790dae56bca3d6cbb9f3e1d102;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3887c994bb3017405ecf82186716da9b507654857e3d370b90e78b0a530e27d3858f8182e32978b8e26998d6470bdf3a91fdf8f1c747ec9e6c86381626d2f43dc33d25de4464cc87466b26fd5095784c051596ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31370bf9c341888e70ce92bf698869bfdfc7eef7151c433e2f2244968425adc5ac97e1a8caae3fda3b1d30432083764d0a6feb119a97246a67e9ace81ae45740a95153cc61393ad64ccc8c43bf7cb2fdc08b94cf2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a22bb55f877659f06e12bd0875385cce115ae08243c6056c4025c1212e74cff1f6405dc6fdb0f23e6c1108c0279eb2dd491ff9fff1d7025609d22ba64b3ee33969bfd14f32aedb0795ee17f42820106f3ae575f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha47db77adff6f74efe1e6debee7c26327ff8633c0a7be6bd288b753c6913127248aa1bcff683058893ee90a0844bff984b116a77b97f94b6c5fd9fcf3f83fc77c11b10963ab7bae635cd96ccecab4178d39d1fd78;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe896b8306f0c443e9d441d6a4c45a1314390a3e72c90a7c6615fc1fae183d67ce734bcf6fec893b8114cc8aed1076c858eb1234038e7aca4f5360dd5c13506bca3765b52073074fc49b60707ac6a2caf1134853c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e5f446fa5320d884d8637fbe510a318293802cfeccbaed341c9062fb6e7247dce060d126359e13245fb51228c180a29ea9a22cf3be0b668bfe55a10c3a24ae6ef0a8e223237ad8a2ed60d2cf8d6de6f8cf996317;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c850c3a2988a69321bd7e459ba8e99cebc89b8939188ed1eb76345b1fc310a8fd13607a49a801953a4f1e0918cad5235f8ccfe87c67bf964ba26737465aac18b81edd3141a23c8dd7068036ac7538e7ef88b297b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5fab301af22f4aa0ce07eaa64d28792ba1bb177e0c23dc5b3aeb424985ac41faddf442c64ce543262b13337f7e06052ba899f94f83fc05465b5d31c41e4dfeffef05718a9fbfc78813105922fcfbdb358768745;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41c7f854be4310b4c9ba4aeb1708b37a33e5249a3b504e79e93eadfe37fa25e6462b951416fb2f95c74429fe4bcb5eaa9065d0b7f45c134bbd14da0deda187566ff37aa58689e10c10a9ceab16d9325ac05bea756;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e129bc264b44b5385bd87945223af83257b347cec58e4aa62fbd62fb933dffd33c4a66e367ec1ef799f35f4a666f5db0f265e43ed4e3483bf6763ce0dab6dd8b66b763067a154b09a1d9b208bc1877b7f68018df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f0c17030f42954042c5f64bdca212d7edb949712850f24a5a7217b4c94e17e742fff11538561fe3de17a834b6cf22f0128d30099ea87b586738ee0e1ba40b53a3481802f0ed871ee5e7fbc4a9d026c0ccb92c27b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haab89c9b379e938510b52f5c5a706f3d48b005068ced5e7abbb5222b512d57316d49fe02d9f0509dfa7ac5da5a2e6055b9e57d49b3d04e619c9705a7637b00a1515e75f1a15e146408028059f003b54b89d8c5e64;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74791ba1580104b777b97f9cf528f18d2ee7253dbb61ac317db1f36fc34ef0a04a7b962522ffc3c6bdfd0b6cee0769455ec1ea224c1a4112177de088d1e0cfdc22af619c90116cc8c77c34492646486d2e49bc08b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb79a1026cf1febda0c0726e15ecc0adab51b60a95e57f2939b31643207444208e33eb719e032aaede8174f4bd1b780cbb96db950a79712e5a39f42be34a62d2e8c48c41c3343f0a4eeb92c54bfd1982241382dc81;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6120c5db09c134e5cd771bd9dd4d9c9a3e4c1db35d95e5e6a2e2ba93dc545e436fce23f13a0c84bd10e4ee2df2e958a1feaa337c7bef398ad3beda1a5a1a104a6c79a7e60ac94f421bdfd30d180c5624ad0214b95;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h924469e960f49299989e5dbc7c08f607e494b33acfa05c3f90a924ff2d0e5f1700c383d2c6bbbb754a1152217f3cd4be42082ef7081054ef0ded46f855bbb9f22ed48860b250816dedfe6ecab9de2d1a4fc9fc6a2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h158a71bbda507c9426cba014d88cc0035ce66c5de3f11e0ddd09edf7a0ed2f58d19a961700944f37cf8ec0c622df396c1b08b45757390cafa9929398f3756115051f79eddf0610e9cdd33f0796edd9f73d78a810d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4bce0b8930ef8b27c853a12c2f21e10854a1328cddc4ca21326434ffec75e46a4d3cb7d0a339127cf515753377d6d80f7b3e270a47cb3189f6395ce43f75095498042be933970280a9437439aac17d4d2a0bf1332;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b229fbdf175d86daa4ab95edb1b32e66bfa4034cbcacf3d36240c67b32cc4e475e07a750809126697b193f2397a00bc0d844d47bb467e788c174f3ae40533e0be82ae0661be18527e34b51b6de1d8c9a7eaa3a4f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6846e178d47f322239a69c3273e6c509b2cffa1263bff832ac828155e0f8ab0255e8d5050136f2500797be0e1209eedbd093bda0136f4966ddde644e56140885b9e269193942f906841527311650b805450a8530;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5e17a43aefca4af2dc926efbc32231911b87254a00bf7717290de51d12158a2f8aed9a78dd3307ce92cd29002da1e5efb67acd0054e01336d4eb2562cc7e2b5407d983b2ca0ea8c602dfffffc5bca2e70395fb2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93ad47ed0eeb98635c7bb3e498d8f6aa310a9262415f7af515e3deb0fdc5c54a9a20b341fe394bbe43ec267c58684123aad48342175f33e096715196912bd795cdfd3ae5166809f0f24e8bbf3542676b393fdccd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcaecb945f03233ae36246b6b9fc2e4b29e0c30eb9deaabbe8cbcfe391a8f64981e69f245d5c9df0e95d5097e51b803e48f78524bf308321bc99e2fedc1721c8d2e1534fc179dcbfcd56a689b7565f6ccf279a159;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a87bb6c590e7739cbfd01dd74303a17844a8078297fb2ff955e1594f48a97951013d3e00d900fe35a6eb2479f5a5591be7638d513f3bdb1c9861af1b65ec2ad30637c6c9a5552e23ea9d4b20362faf0bb4cad6b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8554ce41bb7c8f0f80f4255d48ad4fa5148397c90d4fabbdc14cdb422250796e4c5d1ba426e3b62b48d73168c12706a433d4b793a08c9b03247d094cfe1b24f910a42a755b7a57a73946bbabb7366f16366b166c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfea870203df6aaea852c0e2c5d414861925d01396ff720ba9f329b6dc6af7e739d03fd987dffba8cc890cfe56693b57555e32a0986114bd5419e138e6c404f8f92716cd7e7bf1569249febe197d16079118ba3dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd9f9ceb14dca1e6345f9105fd055557e62327bc518ad63109d5eb3dd6ace79c44b62c1303cb306c2ff801e46d958b91deafe8c513676e4f08cd6d3e12c29b8c1014a6dd207fc4be39b0f2cb6809195ab56fcabe8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h723448b0ebb5e69c99dfd396a84d6dd57ed359fcfe986f0f584647211a0a14563e5d3290fde7333266b8f0c1f445d6304375758a16d4d2f8cc1784a74d3c7db9d1feb9d5db4a9ec33cff1d6a90d425db1cd53836e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdeea23c7457cd2b48809e687b52054d4970ec466f37c9b18811b1d1cb60d77ea5c43b6160804341a738f2b295adb69d3f4663cc3a2a341ce7fb404af348eaa8d1ce574e597643517e13cd5d927757b91007aadd74;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a13497de83c188585191731686eaedbfd991612e64a51543332df1e61e2e39979fa995e3f914bf26b1610a074f836c04cb0f6583b9a331b0973540861ff4f516d6c98ed5f5a4fd4497455d8482305bbead32be7e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c3da1b150d94aaeb9068c5cad6af7781fa6b0fdd69e80457a9430558d9eba8eb0b36b32e355683291d548e848c0057d504340408c68310d40910297104887497883dc0b6b2c851c63070f62bdba0ac56e1a915bd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f66205de2f6257e8b456ce473723c3298d5e05130e9e494447518f664f80d7242e02ae5dbefbe23c7188b4bebb6d14ee17d5c5da176c163b495241b2315d229992c5955ec0b348145a0ce1f1e29afab20338203e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b4509a06066cf63da1d31c8f8ccb37b8102641fbaeb4cac524029e126eeccbfc31baf1dc744435334d0a84efdc8ba92f822fc5f0665e94f9d564057b42151db221aed6158befdda47bb58fcf204a0ed18c81ba39;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8718587466651aed4a1b0fcfc2034603660c3122bd4c7d4223765f4b62750d768a364501a93a57f37cb275ebd0f0e75e0c4406292f1502c55ece0a5a46fef32c17cfe05c600630268d7a71a16734364b74302047d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac6ae174fabdf1a574977b9c217af40cdc94785afd8b28298b2c528a12febd910062e99d3c414885b2ae64e4cb6c45b98c22db44edffeb4addba07e62883d4e71ffbd8bdaf83288f4f85d2a8eadfc24e41bad7b35;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h412771a1553051aa274ed38c08c68bb18adf8504b75deea9285494553be769923a851c6b798e3689bf57011e00212dcea2df945dfe0999ed62be4f4fe33dbdaf836028a0b6bcf04687559df47d618960ef0d088a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb0b067a1aeed4dae89d11f2c14fd924e9320d0c9c0bc1f468472541a2624f50102c2d44fa2a1163fbb623ba279bc6a557c4850e7704427554dde66a649f7beb82a706cd0bc8bb09007734e32932c3c5b30fd2d5b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5be2645b4b85e492b267cb49e53982d298525af4fca969ecae92e5a5fe6b9eaa1b367cdc5e0ba3e3846d8eba8ef8ccce30600aed52926ea2b25969544dba41d7213d7377459a8f8b4ea95c345e50b12423a35472a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb12851a1676ef54fcb98c95dd328e4cc4544b69d2167d03542b96ae726f37198c139a433a9ad297e0af74847a66bc993e23441044cb72b687c5164f15846e9a7834d76bb02ebf44b26a07ddac5fb8f8eae3a7d65;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haaa023f1643e579154a83a458d40fbb1f912a0da898327104106ca21abb81b94480ca9612ee96fe6486cbd667786ece76991878903e961ff5f76218072f3d0545e88816ca7d8d81ed7fc87877278add26d60e2634;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff658d0a10aa96209bfb7798fb755f4109c79630ba56026125049ed3b7845cb8b8fd4d55b7f98937f4c78512c2cdfab358bfe3c52201782809a2ca331b81a553752c1207a73ffaa29df3ad6c08dc3c295c9e9f11b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf89d0f569e48ae5a137aa627a9d261ce06b93c34457a54c37c85ff23141073287a02a0763f07c5ad5cf6b6f7e7ed32d2760a77799274c558b0ace8f1acca3ec962d765336933b30d92df4d5e57694e719cb9bd52;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53d22e74bf7969b1a55e450d912e3904b7efad630bc00147cb34f3bed943b8be4576bd390a912a5bd052799552fc76d54051b6328caf48eb5fb1b078042bfd2f4f10cf474222d71856b06d5ab1ef5b8835bed7fc8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h939dd2de05dd8f43663ac2b85df50724072165100087ad026c2883629fd7cf733a876d0796c8b3c7f4f7de5bd43a3fb460048f9c92fff8d1e4245e937a76b9a711603c009570c014129614855d6d4695c62e08b28;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf133e1a5dbf87d97ebc9cf9806cdc49ad6eea9492526abcbca3d36fcb73bbe18ed66339331ccbcee4cf84e68db6fa4922b644acab32cdd9b09c01bf5d8a91c0890543b6cb595ef0ef5b33d11367d22f88243b11d6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d3cbb0e7918a139641577d528ddba349ac81b2978f72f4c0724f1e82b4401b390df78e28b2d469630762aef7bcab14c8fc3297b617d99f9b05cc27f4d1c905b6b489b2722ad70299c6ad6436ffe58d40c22c9a7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4b5a782bf1e0a86dce3dfda31841335b9314827e5f266bfd15448bfbe79ce54fe54646d388e0fcf86624a8f725ba2fdfa3e23d00fcedf53851b740d78dca99f2bcbbd2863f45fcfaceda443115f3162b170c8b60;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6453a13298e5f551427c870759d844fe9e25a5cdf3f65dc31a91231d4752849123c086db03077d99f380cd490b604e9da9757a15ae318aef64d472e87113d6b5f5ca12ddd9281528f1a4d06efd5e46024ec0ca03;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef14125c95a5861971179ff65b92c325a10c1fccafe57156cc773775dabffd79c0eb5cef05e7ff005861687326df40235214c17b7cc596be9408ff55f33fd52b2693066ffd004ebed2dc687e336498d6a7e118d19;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6307dabcb6bc97f1cf18efb1c48f3fda120ea9bb5b50dee2cd28d2939b9b2a84eec2ef7982675d98926473305e28d29718c2b6ccdf775b309e10967bdf1a4e0c5438743f128d0a955a15686d2f460d6e240216023;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h808ee4f32c724d956e85c49202924b3da45ab783ce310c9412a735810385e29a650dc8bff5bf1401d318ed564b652988c7b1e573cb3ea5aecf2e17ebcb8f2068ba1e93e19aca035523870835a550af89e3331c156;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha335c59f170fce21cf98d15fc2c94aea3df40aef38ed05385eb54f7d15b98436fa96c6e6501fe76e50d36d8961baffc8cf45e56745bcac0a6f04099afccc231bebd1e93847a3f68381fd0339a947acbf9c8cb48ee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2eb4efea17572cfa74acaf850711c6f21d118580852b1ed0695ba0aabc4de79d80982e731fac8ec63930001e554720d933c6e7b94858f011e6b9176b42cb8e4792e5d745358e96edb73131e207d57847c2ec75d1c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h846b6957a2dbb8a325e465181ad14c0cc00f86912061f8faae382832993bb725fb5b718b4fe87301d4af4b48da09907bb1464faf87f76fee40ca6c94b28d87f0d2562df0483307cc3d3431817b478dc6b8e63c5c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c52004c1d81f3152277aca7ca6be7875f84cdf029f75e72ccb8961ac97fd5d72ff1b0f2c135c3ed8fb3c8b58d90dae8101e6e55cb8313aaa348ce7b137d0aca86d69de9d41c2a4529ec3e199e5315d514de415a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd87fd9a7dbbe13e8c87f5e14cbea8877858292eedcd45628eb54899d63f8769265c5d53b3eb99a1e7297299a6e8bbeab6d280228e1d733b44c8dea1134f3f9d94984afeca598d59c218ab126571e7870ea75f25b8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc91f1c74c3d431aec16e7c4d17cf1e1036318d2886668c5607a1ad484fdd0735f0b6e042adfd2037e94a8df5a5d2901c57df0c5dbd8aa29cf24b03ca211a13017abd791f0a7e4c976c1d16060c2463572a3504a84;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e0bdbf1768d2e85c7b50f88470ce9c0398a7d4690c43adf86968a6caeb06ea4f33dda30368335506ad31ff6df990189d15eceeacb5d310fdf185a245668bbc2cbf9d0364566f49c47318297b9838cbe258d3cbe2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had06d1a16c016eb15d96c0a308892c5b92f32eaf389c4df2142fe9e0f23ded3415c26bb25df0442d2fd13484f06949609c2442f1efe823619830f873fa83f441e65346dc480d7cf488364814f1e1aef43e2fcc136;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e7e93e40c33881ff734a101bb1a3bb1b2d8434ce2e81f26d97901d22c6d4234d28787937bf88796fc5b4f8125db911f976a7c47e609f3feb875976abbf43b361664a07462989f6f5c1b5159f315aab8199f5c902;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17e015d4e2d3d931c74b8961511ef719d3e11d20aaec4ddb9b91cb8f4d16c3b2205c3282a21d999f4e9cc74096c2e089c71ad599c2429808a3ca638c3a8d26feebdcef1b86a5a10c8e61f7536ec3b2c0e7a108f40;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c818c339e015bccd0cd8c09ce23bedfc419f827d55719ca9cd903f7daf99679ba5e0e788d43f765cb5e3657500b2fda3e6a0e2c66ccd656413beae78690a960551fad7ad4836571898f1123d62de52e158953b64;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd092d91dfb27429c75dcfa1cf03746b7d14a1f2c29bd0f760b16477b69c4f33405b0a689e60f0eab6d21e3276ebf4329adb6b61ca19e82eec0704218188ff565685dba9ec2ae53c0c6c8d54e3a274b87b98a7253;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4eaf9609a54737d32950ee93286ce485e63be1d394a218540b10a73a72ea113a313c1998e45a3ef2992b9570cd45390fed445930dffc6a8b4cd0195130fb228998d7f7971f07e1cdf870c67497d20b6327a656ea6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h135e75813f11521da1e71415c45cf50340154a740d0c6e114650094f805a15ca4f5bbf60d2f5f068103283f755606bbe5fce5b61a29dc4e7395eca6fe1656e1f66c44418c4a4ec27c170cb2ab0e8eabafc108d32f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb7d1d04439455dfd49808d8d2b0e5d1ecc517998d66b2abbebbe2832be3e3e000bdce1096b4e1a0c5a1e42a31c1aa8ade520ad927484215cf78f303cc33a112243235316acfc98eca83ed929797e2bd3581a2b8a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc60f75c2cd716091f71a67a517d77f4842d21bdf3d4900b52b07027114b8ba6e9eba8877542224c537b89284b56ecd235c42cfd5201d5609fca0f5ba6318d7502d06ba7ddc460cebfa61e6347dbcec8896972363;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb33f6471b7ebf331876f98756964ce88127f1487f41b78f8bf3a10c6d2d29ac95f6e63d1244613cb4b4cd7481bddba524c2b41091496124d79852b221190b91c33cfd8d32edd0c0b432818bf90a750fbb215f21b9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdabd1c6ed5d99297fff06b466bb8d70f055482e4369aa8a746e0386d38e32a30e96331a056fcd4587a8d03962e78fc0f6781ee6d966c78c17c40466bfc5a1b459024d3cb51da5d9537a3504ded4a24eac4df53e02;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e1a3f8170f63df2ca6e712addd2ad771156c7574734c12e6c56ee0aec03185d6cd0dabc21d97529304681077eb9f1b66435c35e75e2c06c155f906b1bc506c6b91d94456b986023fd255c65e1caccbc97687a3df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h86b5fe279557cff60029cb38363866f1fab4eb057a44a5f2f5917851c74a567fed2d2d1f074bd4b5e14da38e9ec59cc3d932492862cb0405ccaabd92fe276ba970ecce4b1bbbc2378e55694128f32dd6e2d6a0150;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fb5c96399f2479e5f8d657dee5bd4be589ae7319277ecbda23223f54210a84e4253bbbcd510b80e4d3d7bc6e60852587b3bee50a163b46c928c73f662efd8af018cd12c01b2ad942c030de688ce030586a31e453;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb7364ceff6797bb9c101853a0799f3025ddbe96bbd951453bf73ec73f1567b2ed842f460a7839a0c2480b5b44acf6063c4948e8ab231bd661e903ab60be07d0f2c714fac05b49643ef88bb652ffda68ef51cfa5c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95abbfd7d3e59d6a8519dbe253e51f16e7ae8016725215f9ee59e8453a6b9d73d0fce514bdbe80dde598f7d71c0e67998aaac9fe3fc475ed572ca8a035e691f6643bd687bc7bd4b6793595bdb1e6ae7ec6c7456b9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d58d60f3c91c8791c39ce593170e1899ea4b3418fe57894c93b72c9e4d893f6bcd382537faef389946f6903054d23a2ce2abf3458591309ffcb4e594163e89bb80297fa12c7aafcda978ef7b5f5ed3cd88a770ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfcbce3f56155dac999ebb4b35e987c9d03c43b36fd99d59bda9b9d3e200df818019623dbeef60c5013a45b3a846cf9032943628dacc499f853a7edf96263978e37bbcf36ba7d568450517c8905a3f26fcd7689eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e906212e392a56e62923f7ffffd81526ae6d461154ffcf343b22bb4281c5858293dd31e5d2e42b3c546c29eadd73bac60e3904ec8b0170150a8baf1a094feabd0eb80458cf0da98443e9cd1b0fa29710dd6aa280;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h886f1b498233ff72c531a73da216c6aefce19eeeb5b51ec91a8cdfb747364079ced70a08457674ec2470f4ad6478db7ea29f0e35060d0edd3089222824fb27d930202c37a1f1c2e3364e798b4cacce1e345fcd930;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f96a643bf19e51652a14046d63e524deb40afe4b722f604caf9c65d1b08494f2d276d9077cd545279bc2396e1719b1df6ac55b377fe4c5dd4e27a453ea7f38c51a51ed7572a72f2805523f7d270d77ceff9c8a78;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcdf00a010e89bf2e43e046ff9867b58fdfd73c04ff8f1b36b83eb315d4e2ec3d23256db41ecc07acdeab431bf1fe9c803023f4ef9bc5fea545577399a5216534a56da0532b85653a93991e90d47902d49ec62f3ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4a9452743cb300d95d38e7ff0ccac06b973ad01e664ca254d1451825bff01d40f9e37df18b6f75fe3691e14678a15de9148842ab8b9e6b9612699915f3492b56246a6e5bac9f3c3d141e74133715659eeef5d447;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ff33c859b2ec89baa0e7c115e0b78a0b641180e971137f9226f2014cfc8375db29264d492173c748f16f04650ce431334d3f220baa9315378a42c38f321d191e5c3d9345c13bf0b4b26f2fa345edf06791ff11b3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h614c70c0760529e39e797e9000dcf3b9a948a02cdc4a9350f8b5b4ae110e09b20ab09aad64fd4b0943082b607fc98344befc3727cea1d3a82df8191cefe7c1bbba6375134a4551747d0e72e487ae6e0aa69debf62;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e826b9f05d7c5e727ff2548df9b2e5d80b2071d757d1c06288e8dc09747cf2f2e596f645b0962036fba4885e0f9a231a9a5c59b0bfb3522b69fa0501df6188a51dc8e2497d02b88f090445275cd8d89eb06098be;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d6fd887d1d6d3d90e36d8bd5289e35036cd6a0d49eed5c5d6eb932189123554dba2368704085bdc7cbc97f44128ca9a024bea721ef2313998e0ddffc2872e4b73b49afd71f55c38a9237122a464e34220f13318;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ce6d26e4f49af448d2a0b83951e9d85c2331ae69fb62c51210da5cab81308de48f7e944ab5328ddf4aa552c8a55a01f8afbfc74c8ecc8d7f0bfbad3d45b752911ecae50995361a0a1c59fd623e0477fb158dadb1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d42b7c9275f847bed0de61208fbcbefb72ce8ff2f0b5f0750cc812666b6b8a3b00244bf29a012c98890ce3bf15f34884b5011bea28c6f23d8cb2f67c86a457f40da208a8a0504a5bb845a37b9f5baaf433890f23;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb8391917da69877138be830a1de57468d1a895357c4b91f83f4a9cb0fa1bbe52ad51aa01ceb451af961d733fcea8c2b88bb694205588252bfdc1f028dd3f7f28de1a3e40f6c4158a472c5b0657cdf1f43362480c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce67069ea9bb564d7895adda44d1afcc66bad7b60f0da404be6b7fd583d5006507ca9965f116cb9f03500c1539fa3856d1436f1b5434733e90346a633902732e82e7e46e158d21c8779c5a8e41d7490c692788d67;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2517d49946f6ec723e8acfd7cbc575d7bf945a4da463c38a4ffa98d7d4cc56bb07455051940bd61fe773bc1c8fb2e449408fbe8d44d772157d223f378bb3211f4e27635375d8c3decd46e4b1109c20496b17696c5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92d766e007d50d647c86a964a6da59a3c67bbf0b2859fd87d6c232a06bb22018764e66846b971f7fbe4afbf76a881ad966671da1bbf6617b62cf386576bdf4b3d716d8a7413a702c9980ae5247e0c436b9235713a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31c5a85d4ddf0df458772171d19eda66a05268b6e9a177e520393aafa009ea000761c02fb204ce1fbdd15db7aa4661ebf8ab0b5a837e2d9f50eee289ea1adedb789203aa96c5c93b0c5f7b813f8d1ad148decfec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23052c785c41961bd155841cc2714ca01a70b133e9a55cb0e617b5c7877697256295f64b40e14a377cbadac47e6a30272bd81017732e031149675ea807f7d504d523d19afa942aaac80ebb54140b8faa8f92ef8f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h961a9c638535ebfe59684ca47cb07a7c1488fdb4a88513657d7d9c8ca389f00a5fc02348624d962f773b68db2f23637e4e8f3acc65e0a9f6a7e8b81138d7b1eb16bc64567910f1706cbf15bc9a40db94ee1b7ecb9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1cb09f3c4cea0a1f4c4d421bcc499c6f548f9456f5952f8d2f9fed01a50be698c1073f4dcf9e8634af3f712fc946492e556184789103bdf8387221ef186e495de1392b508bacc060d8af565ebce60640b4de65315;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6df24f614184a97be51455dd0007c86cd81d8e617bff0c6aa64c116c95ead53717563128ed339122a4e7518a932518852fc434f7ffe1b3d13b8955dbf87e897594e92d2327bae28566377adb1085d0aabfa460e0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30bf67931427ea4eb0d7b75c081993d328dde826f58d40c2e5c1adc59908c7f824276d849febcd758baec9a3cb8485b2ec775f5ce33a14a16019aa6d50de171635891498aa3442f5eaf6e996f45ca693269669ec7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cb3756cd7cfeb4d6dacebfb19e17cdfa34fc4a13c4540f8dfa68773d72d4093f67d5983cb00f44766f2e109e8899d36c4fba77e8347cfc681d38d6ac22c912146b9936a563b79217a824149bd4c6356c0d525ffb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha315d6bd5acde76e3f813b2d8dfffbb8612d059223566450460b2a692fb87e20d86a4fbddc1f984fbd12b3d15a05a0a8c00ceff0f05ec7948fbe90e3ed36f8a3627c2b323a6c6dcc9059b1cccac572de57f48ef5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12c62262e604b4eabc43379ca120e3d572a2c960f99e93b206a5848b2128b471318d3cc8149c9c6ba0f0f36b37953c55a2243d93764180c3286a1a4eb95f4c6381a8ff6c553215ed585436e407f77316ae1374a6f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29579f3186392bfe01a03f1f8e14db0b3a8dd642446f4efb6b2998b4397f9b21dfa53acfe2b9045d4d0fa1ca57ffd9469c7ecce2d478dcad73335c2a498eaf859941c31db00736ae8ccd8ffa98855ef64429f1225;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ef359b10d526afb11d373e0df520f3d376390edfeb876a070a5c2990bfbf775a4cefddd0454ac916284af61145c676372e8be67ed14c5ebe1f9cd6772bb2f6dcbb8100eefcdbcfce2fa53bc48edea0c8a9ae7d8b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb552e4b93d18550c18f2d9f79aef8578e348877abfe1a9d092c7930e67b7f86c42029a136a7f203b2362d0ae34c2e3f8afb8dc8b2ca82679ecd0ea9e7711306cf208713210856fb0c4f159c40681e33e21ecee6b3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a52dea952dad945062eee61176b6aa86045b5d5c1c8338f375d3d664378eb767bde627f6072a99002c0b96887c2ab79de6c6b88f3123949f52d01ab5c54d8a53db3f4a92c6d10861defff4288d09bbba01273d37;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hced32e6a16abcafa3228285ebf94bc9029713ff82ffcccf202d6e9953838d53a4184d07f0b830c68d4ab8890b61237252fb75c23a2938596caec5f14be5bebd1c5689e2a9fdee50bdbf5711417bdd696773ddca99;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7801310484d01d31d3be3b7a530fcd263c955547e3e04536717eef6ad0dcddb8eb8857eff5a945e3793e34e361b219851dea4ad82b8c6bd85ad16cac10cb9774ae06a865349e8ebcbb70a53015060f22f63d6ec62;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96adbe507b5f26acf0ea33bc8dffe3845970bf623086bcb0166fc4047bda3e09ad874538d36d946cc581b9dd5a2a6583cf567291d8e85fd86f3f393d360ef06b183437c90b47dcfe284f0ee3bfa8bd37e652ba3f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce5923ef1815c5ee5e81869718abc9faf9160d84d3ee34899e9d875c603e5a95a14b84e21f00d19b6052260cfac62e6067236a27782b4cc77ababa29dfdaeec7870e5cdb577979601b26360b255cc447253a575e6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h286fd1f6d58519d80e8a9477d2837d5299f4c3b87977dbd49a5b3b33fcd8889ce62b53cf8d546f9883288774a17511deafaf2abb707c1b10b7c8bda680cb9d8a78f00dbef908ccde8b38a8c8e4b427ffa8b53ef7f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0ad9b6e56b1b5645d70b64bc9a11fc1f420382bfbd76d3343f24c108f50fc006c7ffe26bf0af8f825c45ab0a837dcec3eb11aab9f6e820bac98cb0e81b03e1f33277436593318eedd2589aae4bcc7545a82917a8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h445309ce9932e9df60113fb21a7d6e3d73bed0d20adab72fa9cd46788bee5757df46aa4875d54dbdec299ab6351cfc2ac0794a1c5f27c1a782f53265ea8b7450bdce70ad7ae059a83389f587a8dfbd7f4908c2753;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h444778a89607c1e928f3bb030c0e0d1064b89d70eee127f1e8556d6f49f8ceac0805c2c9c97042518556a913d369c345f87015ce6a0c4a72fb40fbf041a520c398f960a6aea2d168cbda3fa88c1ed8debe086612d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57fb7cff2c2fcf93c65da936f154efcff49045ea53faf2e82bf21052503caa9d437bdea6f104607a511608708afef360dd606f851e528035bd499c096f018d1387aec9899cbefc222b095118eddbef7d1c2fbb58c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb04894f863005c37d8b177132b7b8503b10812d3e72d7804e064c2e8d45b1ea5a1f99b9c6e84f4844c52ee4d68477983ed1748064bc84273c5fd5dc92fecf435d04c9e810bc5f7f113d53572d596b13f4f0314f55;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7540d921dfda9e5f6c2ff39caf00c06ddc0bd24f2f97375d9b7e258b7d82a42cf973aef1e7f061eebe3b6be6b86bda98fb708bdaefc554ea06ece1d4053f8e42529f76a7e63b856271e8562266483b8602af96e6c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d71a4eb0860eb7398ff9f1962f0406ecb9dccd666a0a8b44495d2946db0ab203b6e9264fa91716b174c5c5a7ad1c73452eb9e6ea87ee2a2abd0f49e312ee0c60726faf6d15b44456951c4531c592dd8b3a2610eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h525ec44e782d477023739029536ed3f6a08db4efd8fc7754598c27086978df8f114bf7fd17e54963a986d1b744c7ac97cacbb60b85e4f4dfe90e1ba06f85dde7660fbb79543eb1bc8a3a7c2466956a23ab6f835f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e6e7a9a35eb4dab6c1e87649f5202c4e16478296696e6aade3f43de3e2c96656f91a60d30d819222426b4d7827e86f9959156417642a75013efa63c6b8740789fb8935dbd4b6a2d21e0c2e428b7158efbb91847b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20fe034f0207b9a8da374798460f9052d304237fbe0c9139225dd0e673befe3cd12dd24b79b6c2526f794895717e5863fb29575ec1e2b8f3ce59ec076a86b2a4597074462d84c2ffd9bbc14e81b21aacde54c6829;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4301227d0964cc75a14f97a8432586c22783f4c2d8267947113b00286876c39aaaf058dfc75bbbf2c8b921d428be0c273610e375a2d938ec5bab9abdeb7f2f60af0b96ebe0edfe2f4808063dd584733d806d66cd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1dc91a10535d795ad8a3aafd5e25d10212bbea5c624722d7431071c4eed13d2479b9b4289df69fa786971b0a5607eabdf101f7a9345960d07effbfb36ec5f93e3a0c1e02e7842b0d9322f1f6caa0268dd2bfccbf6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha035be040501b222ff96eb353ab73cc078a583bbd78ce4f840cdb3e44a4fdd353a8a992872cadbc4914f1c38b8ab99bcad36d144f2cb0f6ac1215cbd1a77ab918792a5a779dc394e46b7f7ea243e90c423a81fa47;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce45c7302690b6c0d169d2b806ae81e9b611f92aa58fa797354180a8c7f50f919a7c3e51e9e51bc5e638855a7b7342c42ff8b4daab9339acb801acbce04253655caebdc1b1cf19337d3ddf631f741d54befe6b74a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a01e340f3c6567bf34400e249411c018b0ecb1b818b53ab125dda51b240b3498bc268c64091fd9c9c5ae181dff54f73a7b74ec0337e5f641d0bb4e00da789fe35ee2bbc83838aa866cd853c34162e3ca3e05004b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd87ce646556e7239dc07065a2a2d14a4d9870031bdcddba3be0cd6a84858154cc98dbeb8921703cb365b5638bd7eb8f509e6229042b6948022a451e43e2b39d9a96fdc9d5edefc23155b3b85dfb309a589057b172;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a86ab316009f3d6602f1f529efc94f46ae4e186db5e453937be5b4cd4725985ea6d66c88c62b936400bd282c16b641b64097a603a47eea01c576c87d6ef0c3f3fd13192587c9b38c1cd4f56d4ffcb634e53e1021;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8caf3593be3ddd8a5454868e1f3b993282b7f11b2fd1a81c0c6dd870d2a78477de4f270a87d91d47fd4179b58ae3994ed78346d23b1587e63d6c44daaf735af5195dae5ba1991148a23753a10c095b011d36a057;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h130c7958860f9aef6f2745a769fe51a1746875f4ba781cef72f201ffc1af1f46ae9e090bf1efac574b2f5b2c7d8b6b8b436da6767c4d3d311e6c9c5eb0481aa12f2ad0a247eb8d0a8b5e28fd262542969d7cf18c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cb3ec928f1b9ab3c8a566f440b23c9c4e70b2af7917d8882821318b36c2d3925f7f2046a4741196a692fe04adf5aa8b2c86b211e8faca41e9ca11d5a7ef3e1b23cb9997c5b186cd0608e0b281e1cc3b1d6874c34;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b4809850e028a1ccc2312716d2f733346d5f6ba542b2936d0acfa4b5a7662e676052be2012a145cf6d9c73c4999e3ba7fa84fd2be669e140edb6ab91b60aaf24fdbca37c613d08e9c24e90e39613976a448611a7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h210d1a2652ec82b1ca9f6db027fa0ab134415334d455ba0a113a7ebeed23318f1aa6d7b5fef80452ffe7b18a711b40bc89306744370c447791c33cf4d894f5efeb069dc19956f260ae5979f3b8e4732b0b85621de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2a242aed53a0e26732efe3a44bb7d98f599a0c1fb104ecb4cf81597cf412760de019c05903ad7d2581da8db67a614ea8cd2e16fdc6d2fb3c4deaccc515f71ba5b7851f2663b79f21b4037d245a18b36569e8f197;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3e1c420d0673594c09d35277630f8461c567b8faa386bed91cb39e02095ef808d78610b7a0e9e4dc85e665ebc56633e3a1b6cd81c0e18cabbdd2358446d1b682193f00719f332210d9f22d54914492ab1bfb9c3a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31b149dff117eaeb100c10e1f26752c7b03d1349ea08e5ed50ebcd50dccef34e46ca3de05753f769d5e813bccb0e890ee91b84d9539f690ce0676fd00685ae28cf081c10613911fb63e40a2f2f048b0458a497d5c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfed91e05338d340e1e80b6a155550ee0dbfe1c2430c82aec843803bf5cdd09c711f66245d505962eb655059d7ac7c122c8a591d81e7495b02831edc7060d7d03aaefeff66d1dc542a7e39a6fe16f57a45d2e9231d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28c389dfbfe0cf7e30b24caefd8fcb8a1e64990b48bc7bbdb8cfd87a28c9b52f1b4c51f7eb168d5eb9f7c02f22c48da69504c1f169fd02d8ca4558df83823b69309a8db60717ee370077f2daa15e99026f09df0b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f9c45ee3cb90cc01f2b949d17c72da87cec209be08d6d222b4b5587139b3cce85d0c9b6a7f2faf6ee5c0ac73c45a55f018873c0a632d5745fc4a9d0428ec3ddd9b5e270a8c8f68afd882edc89d3cbb4521e1e9af;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c0e1c716e611d1938f5248e251dc50ad388de371b5fed5734f5527eda7cff6c541eff020cf35a839ff8796fbfa50e8b65c2329684b5141a9c48edf83b65c5c98621cef3db0965d7d3242e2809ae05975ef21ef91;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd5a68855017e76b3e1dd90239960d0c8e90a7d7c1e972d88f718efec2b88b12aa99adeade89779a803c60c94d65e603706f6f11f9e3bc40f704176a86f5be5a45974378079363d22ff9fa355d3d615bc55cba761;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4f64806963671b69a039dae078815245e445437cac0e79124bad4f11a531bb37938cd46673def225c60655f45c1a4690189c0c609f14119875f067c773dd229e0f6820dedaf1006688ea9e9a4ae8246998f5fc15;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0d43708dbbff5fb75a331db302a88da0e8bc374287e53c22047fc328e28e76669b9b7b60093c11efc50658bbd80eec69540f6e9b14d24eb539703c63b93a281a34a97a1474c704af5e61228d110ad883fc4f0431;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f9f1288c8158ec07ce2b4cf6fede17e2f4e54560c45d1bb57197ce1b621ed9aa34ac9687626da962fea378dd6f408dbb598b501b1a4c00a7a1b6fd2afea8fcb868faed8c8cbb23baa8650e0a4e582494d1025397;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f5b3e0c4de6286e0a51cef42c72743fa8c62d2b1ca7df91671bb455cd57b2fb1687addb323fe1bce8064f292762bb994f13617efbe4e2efcfeb142c4aa402012082a5e6facd26c12acdf85fd526ae0328f4973d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde61ee25b7f27109b1f8a89a2b85771d87e7db635407695c6345d43552b3d770a154c77e42f7d42e25eb0897b6a000a15a32d7f614b357475f336468bbe53ed24dbdb7cd0f9226ac8efc6519cd1149ccb179df47a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf835a0270d6aedec5a1ebeaf462ecaa06bfbf1c94596f7f20f9c4bd2d1679760b75bfcef35f8e4b3464581cec88c853d0cc9b1291e08048ade4c7c9c15938b1c70c04cbf7f69f4d06f6eb5bc3428b4a33a8d0e45d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h957b3555b044ea2585631660f541682515e4918d7a2c69f8c6fb4e6c86ce07c7295a09c3d57cd5ef6fc1a10a3a0f23f18b4ad2dacc9560cf4d0379fcf58375cd687c939f30c627dc75499d093c6255d33fe747001;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6752adb61c0b33bf318d99030d0c7d19b4cce029e9445a6d536096de24423531305402d1c7e1b5dc98006b1737cf31a0f8d3e27267edc2ef8132ffd4862b2fc09b302f08f6bea9ae1d51a81988aade03fdd705be9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h182b796d63db12239f05216cb64f6923097d25a51b5d44eaa9a9b70470e5f9bc84f40c581b28c08d282f2b99629b96cb2ced1423bfe968c59ad892df31188b8e05740cb49f5fccb2448dd5b1768dac4fc5332ec11;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48b93651ad57ff508407bcdbb300bf994528d9b8532b038c8b856eb93b0b9b67188541af304e39cf2646ec829e5e95fd65faaa1b0f73c9747bb31b0f3ca20039b365760a9e695db26e377cec8ca33ecf05544332e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h997e468a59aa1b2bb3ec7a7a069d69120281472f3ffe81533c4d2de001e355fdc86f5fc55a8dc788997591e4a2ded0e6a35a1e6321827aa87b20b2526ac74792e88f093ef6e20ae21878460f3763c2c6ff3c4c88c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h517315c51a774523296e4a88216bc5f1fef9127e19da2bd8db0b61af07849c3b71b5c0b2d3c4cd7452f19554a2bf0772ebd09174c77bb9445c8239778948a811177447f24c018b30580cfa525fe471c4a6f60d169;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c6463a22e455c3bba33a88a14960c5fe4bdcccbe2fefd84ec59d9f002264d2713bee80d451bb1a83ee27c17942c91967a812c398a58986eceead919cf75fbf9bb7867093cf2e56962fa8daf0f03e6b713291eca6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h405f5ea52935ffd246ae12f949c2b775d4898fbb91e59307c95206b9a11002bf3000f0ce9c5ec0b0fc773e38736426e0d40118c6861cfbb42467a16e777b6ba8a6b45b1fb3e1ae9a2fa93f7640ae9861b327e8e8a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2011baf9987366fc4bacad5864d69ae78f1f18b4d0860a703049db5ed1738dda833206d414fe4bbb1adcba7e3adc383eae9970d6de3b21e2c4048a1ca3ab2570f34c85f4887bf9d5c8edf39ef70828fce5cca7c7a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3075aec59be63b1cf51882481e0cb199d57982fcf82f8c60f73b370186c0fc9cadca8ab3274045442496360c801a6d75452fb68acfb9d0d28685c76f3991c662b05087d9c349cb1a23acc522f3baacaae5a7f31e3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61582fb38cde37366db777bf13e03e5374db1f64287403d6f049463a9bdd0f21c7fac486d98df80bc81e041e15517f67eaacda5897285a443fdc2de773b80c95e2adb7980495e369b3813f1f69859be1190146b98;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7730391e109f708a12617947d80fe6a8a25559ade0991d557388ceeef53f1d8c4ab4af5f37426201be419dec8c7080e72008b32fa58efe790dd4dc3803efaaf0e4307f9290f99c27ce2e5487fb07f5935d38faff3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h237470ec46b8349622129c90ff2e8eaf4d92c06f1e69f8985168e5725c492b155e220e12e14fbc518c688986bbee70ae99cd9293b25ef3709b10f5b177433696b96a2fa4f5aa6ac1d793fe146d5a042b95c2f31c0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3337b4e18a62799f03e100d2200587fa5041d5e5d447b7ab84afbf9657a9b99aee2d07b1ac5e6be7338e27dc406fe27dccd8081f7d8a3ec8990acf3fa78cdc7a8ea9000bd142f30882174a9857ac281bd4859949a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90f08d9884be5fceab6e98e3f47f43d2302d7ee127d924a84daa1add3aea7d7349855de724f84760d48acb21c4157090352c82f465762daa3f879be3ebe97e2684633657e7966a633c030a7762dca48dea26085fa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf344f50029d63c1c3c9f06ca4401634d6082348930d8d9b6c2d17474c0b2526a670e10cc4c05f99f8ad478d15e4b8bbb873d63e9262260d238d70e2dddcab0c0523620f73acda12b1f59222a5fbf5b457bedbc94;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9cb399c9cb6c02f39d612a21be1009cd1e73e1a069945ab129c9d678e1ad1ea0fe90aa014565ef1791ce2cd431d16225f9711b14ecc3760c8a6cc18c44abb8b90d5baaeb86f433b959cc4f3ef6b94a0d9fdea7c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35d5f936928ad8c63a56c27bcccc66b7371595aa734924804b6f5dddd4a77dd17482dc052881f23f6a731602a0b05782a500ff64b8da0a27f3f2c6eb61b1c7e655523850f21dca388d31681a48cd1a4759488770;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a7e7d2f64160f53ed5dec20c76f12db1c355ad92e9328f17012a1543310acb6f1feb9d46763f9f6deccd9e0a11361c9553bfdf21d15b55b292bad482aea64aff641292113ff734f597c2a718649389ca9d760093;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3aba760211a8fda2c0b4ce5a4c63fee52a6a41c23c6ac8a2cc753848323491a9235f25d94923e971de538c39e45357e313dd2348a0e445acbf8255b52fb7888f7309752f4ec22247cac5d0cf9e3c3338cc5e50890;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b1048acfae806d3c032f62e3f899fc742fe4747768529a539c9a39968ac0dd2d71b35603185ac21952d367b178df54efe9da7036aa0f02bf56111225d32d22abe1c596dc2af34a47ecd29fff7e6ff0c951b6acb7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5cc43a0017734df99e7d2a3d0717f3d24f8c78e37ad9ad5db96b2ae2d1d7ffb9ff4722df26130e6563e072f4b5d9267dace39c8a6880612fd32150da78d9209d52c3d5ebc94acaf2b2e5c8ea5c3f443d87979a10;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb197a1716c10e38ca6597f96937fb4633d5b5b31195242782a255d75ef7f30b65cb922c74c0bf2d7e106a74483c3fe2c5fe2b92097faa8d4a2722a5d39d45baaf4b3bd6d39434bd72431111b0d28c241a509ce09;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b4438d1238d7261fb8292637881f2fc1121a2d86868c7ff00b8f5f7917666e5fb038cee7f94f0e80e3abba5b02dd238ddc3274835296a042723b44a4c7419b7b27a76e5d58cd82aebc257d8e6ab593f80c3c7ed1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5de6dcfd5c06c93586e8271a7fe449ddbf533386652375ae69a2b87ee8dccc50c784d51b4a6d52c07ddac5d394db53ec6ce3949cfa9269c7ba3aabbb32ec038bbfc398d6674793c9cae59b798b0102d16518e1c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9bf70d378ced7395e146094bec77902ac0cbddf3492d14004caa2b64920a770675ed67fd5f6c9127f7a41eeb8ca0d4c1e31d7719cc863c9d78a4b214f41be492ba2d8b4f4fe8dd2dcc01589461b68de375f1d4b8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b59518e42c610c4683e030edaea4dbe534770f0f3dd46cc98650e53d238b720c502e6e1e383be8acc71695c50a5e5a288132794b541da1f8835d00ee9c2364fb990d384a479102afa4a3d549c43228c2185264d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5926a144951a508fc4530cb70ff7e275e7c8322ad19502face987aede13d2073adb508dc5a04b8ede8daa9ee36b527afb1c1accac74db1ed637de9177d3dceb2f1363916e2018e937dbc710e0c7f15ceca4f11b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdbe78cf704d5f5bbc63999d5484081dd3dc9465faa62100a54e63a77cefba5af5068687e15a1dc2f00460dfab8b26d9b026ff83426c835880f2213efce1cae1a8533f1b96e0c2b99a97c5ab08e6e3b9af906b4af;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc17745c2b04d711a09baae8090ec13b83a8aaf93ff3937909e91bf9b3720d8cd3506fac85425490dc60ed182d5f7fdab15c397837cef96c19aba0a75a41974e85ae05cf7b642311d389fb1bbd28eeb965c0a99586;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf1cb83ace957c9710d2ffb6c25c9d1d625889b3fd214fe24ff9e60f8e12ac2d006bb391a7d7d32353f4024e4113743b32c81593fdf40bd5b54f02f7492a2d7735cd5b274b7bb2739251adff6443c9a51d7c62e6d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5c488dc653fed8006f6382ef1fde7faabcd88fc1574db2237fa9409107a9e03df90a49d41eec4e537ba9af2fd5bdf16872f2b5720ee66ee4e7af2274ebe51a9ff339d05b2867b7e78b072a2c7283a7d854526407;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfec72ddfbd15d00eaa83d0ec5cddb0a9e68dbc13eac3051b6c7ca8856c2b89d3c622dd545efff5e5cf0ba185c6d1bd3571911d1c09fa5368ad6254447af8fcbce4f7a0a6ff2337adc290ffc3d7dd25f76fab9860;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h349728a90b34eb077b7385a5e8a899d7b79cc0b70871ac328e7e6e831dcddf16314c50ab7d1a1963a79971dfceb59934194496c6b59d3ff3e7d31d26a92ed2957c8e8165e05fc2876e2c0fb410063bafeeefcf367;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23a41b03cc91c8c9713397823967e06b65b4b5a4211974aefd9d7045aec24ef47501c23fc8d45d68d7ccb19623e3bd6aa4105dd4ca275f45f2ec0533189be6103840d5eb06d788e92c35056e01343b973afee54ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13fc21eaa4d6bc2f00780d84903b4cde35ecad28853d11bcaf27b208a3af8f2d0e875b9682ae4e5d0f4d72fa954988466338b0e56e1d0d6b7d7ad9f41db14da087cdfb7fd2b92dcf6816256cba9adf0b59fcde33e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72eb14f6258d37ee1abd24db08dcef157858e42af3fced70ce8ec9cb2fcbc3f1af6bcf4f2256be6c44986f7dc89d858ef305c2548429454ad30042e6e2f2257f6837eacdf45a176d5b435e25d70b24ef0ae9b75a2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85c138259476df5a162544e188fe328677404a183f955c3eaacb9c3d1e994be83099a9e7a8248c91b1cb19cd103f1f2ffc0451cd327bb3043565dfcd565d2ff973113118a847827cabe0a2170b8f638c0d7db6fd9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5228ed276726a2297a6107255fb9f57ff17089f7d1164d93506769d4a209ae51b9e8840969e9032b4cdc850083e414d7ee7c88a5bbef1a3a5eeb3155bc8d5259b53526d903275f640abbd9a25775a7daec6c04ba3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8e7d8dbfc2f323a77d94c957d68d8f38895d08d9e57d02808b32cf7abd7fa287ddad3ad5c8c743668172972577fb6a28a86e86c9f7b48484bbe51ae77eee16ff0db55da5e2c69c8cf19ae8afbb95a7460b8b98b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6cec3ea46af057b3761cef8a36fab6528ace96cbba250ceb606a604006e6013987b3041cb47162862c91c5558b9541158b5e841126bf106398f159104466fd59c97f0625d13689ad90d44db5e325ad1ee5b4ccaa0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb176700081e7c766ce6909bea596dc7d97bccce9de4381b7589ab7e1ba52536943cefa9d4953c3dd7d3d2934a77a4632fde485ad2820b5e21ebba93cecb7b66c2fdfa368e4fe99555900a1a1cac494e757a5574;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha825d85c081579f33f71728f0f273ef0f6c9e972ce46bf7d3bd12672c9a64c67b98967936eafed7c2e663087c184cd289464b9d184af1c80788f5890ae8d7b4b5590b294525c1fcd9622d56b048b4f81d05ce2955;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3222e4942a7641c5d21464b230d80ed1377a9d6b739f7ba75664cc96abae5a43c80325a7cc1b25df8e58e627881bfa8a043ae121c3e7b64cf544318fc9fb19daea5ee8aea8226f0c478da01429780602f585daf7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7eba1fbf7b029a966c0afc13b29ae55b9329f756f31f5d461df0f96e8de7766787373a17b88f9ca9f2771665b9f1e6fee01c539dcf136908d14ce492dd70c56cb1b7da9d3774c193ec57996725695d5862a53aa3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ba2de3df3669e1af0193a650ee83cd492cd282175fbf593326d0463cb261c7bc50ee622cffac16ff79719aeaaaee1b6c621b9aa7f27575a1fc287765fdf170a1948fc23f77b96629ce805119036cec991b92a785;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb75b8b213ced489ed32fd6345c787f5afc5c88ada1e0456b108fdd152345790953fea017446341a74ceffd4effa32d4e181aa6a324d6b2c29484eb99fbff460798b41e7f7592a4c333b8ff75f41470558b5dbbfb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha53ee2e392827328f1c9b43dce6151f09d4575f4ba55750ab568600b54943c9cba1648b428d9b1f28f4b802de1b65c4ed4eac7c81a293301988541b46505c0013ee006fe6cb1cd6bd6e248f17b3aea58be3e0cc62;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3dc42e338e2474b10fe0c7640d6b80273fb18befc65faaecabbfed429af93b37c2a0659f63a29529f0508daa5ac5b3f38aa572e8bfc9e8dcb717e47d1c30b11b0afa2d8d116dc6d0dbad4826741c15183c2e98285;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe5f6436f4ed668495b69d1f7b57c92a2109eb9ef564c0fb83d6075235999a9aba6464c6819a76e00f6eab25eb906a32e2d4a805141b9e5c3c18d56a141814da416540d205b565cfd4d0a081030869223f020219c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1063fac0ba99d7eae5907307c9fbbcff5ea71241015fe39ec5b5828210b6a748ac068bf7679e3444c1820fe7e99a689ed29095b570b1f915d145c8cbfdd7cc24c595eabae9fbc2b06aa50290835e8a29096f69efe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25023627517b92d3ed23343af3c18e072e51260cd3ea169874300ee292630a317c3aae8653b55265ef40f50c09fb46d6eda1c533f3642aabf0b572c942b1fa725839ee4daab79438672e3a8108dbfc84bee1c8bd2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc384d6c1bf68efb92ebfb5a450630e64006a3d8b043cf6167f56a01c2e8131b2b11ad21b28b7548ea422ef48fb2b2a7aeba35937b26c2ffe2c0fd3aabaa0f82bddea901e7e32d555b7b4789c95e9fae7acbcccecc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71b8f7b95ca2b674bc0d9632399bda212be5899748333f4b86317926588dd0991918619c948e389eeedf334c21b148d5645e72e9a2cb987cfde02cd5184ea90bc0469dfaebb15de4affd5c64631eee2ab8893f453;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1e45404fe0374c1a4d4a3c3d3eb4bfd7e7d48d967ea4208c70e3cb91e549a22efe50948681416ee550b3a09a13b1795fbfed78de4c6175c72999dba940f84d727332ef18a34190cedc8ef2b08916592bb85553be;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ccda827332f3aaa9541973054b20c77f9ff5f589bc6f8e7ec193a04e937e556c2f0c447649acbbf4a35ca9a14dfa9a7a4f190197baa5527c3e5575c0596f8da460af0d5063df31d8f813127037c6bac7167ca754;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b36ac3531bd3778fff38b1dda0f3adf178f27350182e84373307e25ff7e8d356c0b7c588b60516313ec11bbc01c57eb423bbf84c36fcf75dd4d4d41e52a9eacbd018737adb360a52a982f0396eda82829e1f9630;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1980e8cae988e23600c71c134061f6d98664294685388bde1aa77364e02901a93953d1c690f3cd3eb79344b1c367d95ea8f3d8ff492c9c5deae7e76814285897daaa6013eae791b486957a30f7fc871c358b8e27;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h872f0a1e3c4631cd9c6f7e8f4bd13b101584dea8d1b954da68a095e6cb1111d4d8ba1ec22d22cfc109e42cee50e9b12df4d45038620f92f6370c5e4fdefb7871ffe8a6f4b5a477cda4b7cd8169d5ecdfebe57c8e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72dbc55b43445f277c964d3b0f20b51d8cea3c80df81682e483e7f851c211f305c9156c69bf9d9c0bcd288b3f7551b5e48d837d984c462f09ff54a1924d47c5517188f8ae37ad092edb4ab1a1012743c15ec56511;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd308c58c4ff2929000e5ec70bfb7ea21d322ca2a329042c9678fe1ae6bc6571e7d6af09804ff5916e0dbeba5eeeafd3c0375143416ec3f9376207d2ab4796988470333a7a477cb0139d9d58fda7f1f52606b59e6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf02f8b1d5fed496aeed6c17cae10c3ba8c1eafa3d9c101fa296acef48399d899bfd470f46804f9c34a094f04a8e6f083b6a5021a67247ebb208421ee8a4f74a11caf6366f05bd0d954f86a8ebd02f1748ef3a4db6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fc90a9ee7a0625b9df0c8d47722b2b042a77c4c843cbe6c267398be1fcfdb8fd93352a968e542f9d806cf4e0bd542cdf88c2a15a2756fce8f1bf0f4f7fd0bb9e5b06a4cb04b04e990b3784cf224c0cddb080ff19;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ac2d49778c6ba1aecf72fcd2d2094560bc787ec1580b1e71a26d2922efa4cbf26a2b0286ce6e730efff03169d11bb6e1325a718fe2f6937a548a6a5ad76363e585ba84e4b970f0caee946faa6f43f0f94ea7ed05;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8098f60f0c5c423e56790c44038fff2cb7f87c8ef792e1b34305d2e479688ebfeaa0fa4a4ff673935c94f4a9fb0e2b4ea30e0acded768c20fc918a344c09aed5e6b7f02b30adb06076290a3e5716435d72c40d754;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdc5f67249407481d1172d6576d21fa03e281a9ec61a125f595dcee189a923f9b2bf314d528c9d19466c415faa3849572aaa13006a9238f99a4cee0ef12651aa6a37033221643e184fd67936d25ef1a725216cec2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h427e889d6155131a74e74861350c85f12f7ea873681325633dc00ba6afaa588156ce65cff8269e492cc7aafa45c972cea8850a81642f56c41cb4a3752e5891686e0e47fc43355fd5d5fbc77da34c1bc49fe58202a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf170ead2794be385172b4fc2c17abdac9b3bd48277a836a87287147a549fc837368099c7afebbb975e38614e64cb193ff9cf2042e328f404fc6f35958f26d9e42d723883f3fa1153c3c87aa9fa836afda39da15b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48638e51a98cd203eb0d83f54d312b409e968c63d04b782b2bb1d3d668308607c0bb45e21da014abe9ddb1f40609838bc595f9e73e5b7b49a6f9898e57468774c457e878fb1d474f0ef772b909bcd52c67d95358f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h503ab7627cf845a22e28bd77b65013274ab5557d484958591867903ac0278be6ce1272ba44e3eb51611eedd7843f541c3e31364509928d67f347be29b3e1f9332c65fe5a3d5d6a17cedc539e7b271f514cca6e337;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3227fffa221df922c6714964dcf7bf07449e1ad1992cbc0d13da4a881778049f953f55bbeaa08d78b9f6bdb00450ceb8e7867881910a964c1ddb6a55ab7e0ef7405bb93a23d8f3280323cb219703b1c4f4a2af070;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb22d09b2b33c1c50f98718f526375b3662fca5db429b4c3ccaee7f95998b5fc4724f9b4bfa4098d5e6bc516ee134f9b3b2bd3a153d6fbb249011871c4f086762eaaed9173cae9d683a464e97dbd428529e80f109;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd67672992b705421755ab23f1ca3f5016d09e4409b5252dadbdc156efdd8ae0ca75e3292b8bf41c48a796a701189b55d38df31d015777d6827f0c08b822c06b24a7db7bac9ca2f0bdbf7358484e35e90eb788fd86;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44868d3df16c7c4747554ead12dc0aa3366410a6d14161eec095ce7763b9c2cfa3446166f9d908eea33c7b9bf8937916738ed1215c3363d2d828d20b5ecfd43cd658bfc093365911566cabeca963827a35092a328;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7df4b41a197a1a5be1ef9a649609ca1e090b8bf1ebc49547f5202dbc1e7e5f65f98efcff5596cfbb4f209a7dd1b23fe40c82d043564563897ea185f805b56493fe94b9f6e9d44dba5e8c457aa070e3b3303deba35;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he45f9b9870a9f23fc763a14cc7677c19c7ec4adef7cf4df7e5f5b0e17621a064395a677b27104783a80672588d8e65207e01faff3bef6d62b0f9975ebf4a2bb02fc511016f9d3feb8ac1cd73d968fd9c40be75d12;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29f86e896bb798f9ce8d8e78027ea0c3e242868b735d661bcc6cb4f4f512b7c66a62ef077cd8cd1ab0379a271e09413e3f210ff797d662892eafc6a3b3ae81e43d98c2640d36bd5b608c316785011386c07e68444;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa3147bf4a90ef1219b1773e7401ddf6e6b6601c867e286bd0204a882a72ad7dfa32d43206cd2d2cb55e51ac91db7434f7a9eb3e3af7ff638475d71a108a98553ec81c2789f9dac1e34d922f3fc1b887ce6c81e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h694a08b02c0aaa5b4721732810a96661672934210bd0eb806af66bc84006abfa099f59e32614e1a32b0d11d8af406fecf37edd6263594d2e961bf8ebe5dceb693f83f285776d672e4db503143789d3ae5f0fb6e63;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4eb7771705a08ec462500009c91bac5d7266a45ecd9a1a072509c1cfed180a270cc3bb1a58a5f4cc7629ddb70af8e1cfd5005575ae2a1db5eb1dbe5eec6e3105a887baad49effbf95566d27336a1c7d8559a3caad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5be35c33c1375bf70e5ffe3dd2e752756b814cfe3dd6744e6289c7d922d0d0c855ca9a6321f93092f7ee67b896288bd2a2a529498265204c1f129267c3f70919bfe2799aa44a4221500a4293b1eeec1c291d8a549;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18401127302c0be684858a70f12ea279839eafca3a890a9ffd216ce6c4fbf0970094740172f37ebf6fe286aa6a8e73dd2f5db94484a364e15499b752f9716647fa701b56e95160434b4cd5593433228e1fd41bf91;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98163b89c94288319a2c5912ca505674c29ab4ef1475748827af6ff555644cdf2c5a7c232389f051204a18219e85a6373c4cd52d295c7418688ac78b25ddd048703f7440ca9fc6a22fb83ec05fdadd7dbfe96aeb5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63a056c28c37e1f6f5857c48aa61d15329273e9983b21204a6b18d90404b4028bb2f62d194cc7ffd142a77164ad16ebd4e8834e2093114d76b7ed00bef03933d41aeb490808d39d4d2dd7110df74229497862f38d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hffb9befe927c0da70d06d259dd12f5d43256aa2104d956f4c43461a88ee9809275e5343735e0d93c1cd8cd17d48836372157649b6c8b811f4e949d6c872334a5abda1529982fa7655cea2f8a2fe154d9bb53272f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h595825dcfa8cf7ccbd1992f843b19ecc4f4f7b4fd999ea595d78e38fb57b03d1027fa80f9d3383be82977dfb5fb8e275c699249dfacdda996f32e70ac7279ae4170945888ccb4b297570b937cf71838f1125e9ce9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3efd0c4024133bf80ca57645a83fccf28761dbb9e9edf273f733a817ac4c842199c55b046b1ab90dd8faf5bcff04771cc8fec1454b47e9274c520b3341dab20bfd7c4bdb3770a00fc75947aedb803ff466b3182e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4f27e794c5f0f3ad799e2a4cf703b7f4c82a199ddf2116a5410545c1b92dad951912e4fedf5ad2d7e8c61db73eca67b8729242c0997600b3949bdc4fc6204f87160e11cf5e1bb6b85f16f7a4d3583aee0618fed8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7756a106a541451b2d5865c360b52708cca12a3d773780dab1b8585e9ab88e5f78eeef75266ba94c8c0ccdcc699e600565424fb2af4c6cf35a6995359c8d1a5657852367dad479aa87480284a4cddcd52322e188c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h689e69c1a6d1f09dcad512a43e0c6204b89debdc45c1d4543306fe21387331785ca727ca050b0f386a8e0d2a9817d2b6a0210c47adfc0ba9a23b256adb29032e6ba5ad8291ce2f37b7b7648483f08a4140a3ecfc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83a820dd1fdc6dc31f0a1931e966ba07f5870c9f06d67ea7ed0a36d315aeefd889853ee493986d1d4d1b748a3dd4629165e537c358eb6f756214fc4ed7ae3e1eee97ab90d0237431d41832a08271a54d79f26b584;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75e6a15f29ede2a4e1668770c8b7330ef3634454716bc3113d2a2a4d11cd4a44970da0c2b5f16251ff044c2224facce710dd724c9f69060be66fcd4754842378b40a61bb935032cd499d8e3337dd21295342e92ee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h677bcf66ee782caa4010b716e1eac2df3fefb33d7268f6b797fb2a76eb0c4dc1aa8e795438707c0156888c7e3ba68819683cd75b6dbf11375e09c61f3c911e44ca7f6c37c9eb24062bc555bffc2c6970e687fb513;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0c01f115faa33f8226f7c8bebd4f47f08462e2d4b2f9c9b6599928b68dbd5d7bb45de032a840c3e2b953e0a5371cf8e2f328f00bf0eb9a89d8dab3903c03e126d0bba397c22ad2b38e47da47710b4a4b90782357;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdeb515e97b54d60e883a5ae4a2e3e3f7a87680f7be28680baf81499a4fc65f26eea56a19e8dfda1176c4a7a468e12386268eac22551aa120796f87cddda35ff2df1cd1cc4cb47b6fb32f5b4df49bd7fbdcb24e775;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf88d44b50fa625d26557a0b78550a51eea69628398474a5e2445e8376f55e9a63c789aa43e5481de298566a2a85b859bcfb570a5497046a35ba17333b49dd5a32b050c301471776fdfeecf115c2fa0b323691a9ee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ef1b23881dd7ab1a68bf56b922fef46728d4190ba3a342a13fdd8982e17f6069a57db71165d980851d9158be633cd4e6462be44bbf3afe45e146934787d41ee517b84d540029c0e1bf50af38b81af5faf7ff390e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h310a5499a938ae2a45ad700c125e5601fca9d211d1eb76dec8f597e40bc588d6d8fc3f5f9eb4eb9d37e6035509d9342e7b6e7c467bbba2947c5c784d7c50d6df486686c25907f14966c54f037fd492693eb18deb4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8567beb24833f5538eefe00f1784183b58da0f88e09d5bcd6562542df8b26f9ae9db29be3c37ddc98608b8007670b9d9e90d01c83fc19a58a8ab7e7380533d1d9ecf5b19fbf472e8c541a9da52312220dc147930b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9062dbb49cfdb23ed298358e65a8af0a922551171ae1f680d56ae91b652560aa3fd91428b263d0505ad9e1e13b1f072305db8f278e972864ebd6f9baf663c25735da385d62558fe70e3a0f407d24704e569da586;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71709d1b52719f437ed936badd2f121675a8fe16c7da3f9c2fe1589cc808d7ec411568657b6b43aebeb5d5801dfc97fdc2eeadae7b313baa4c8d33e40b312cb94355562cd46faac7ef58d7aabbaedbfa780bb33c5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68eb1ade69d184cedd3088b28f465e3d2b707c145286a5b863ef55c10db4b349f8d3b72edce2bf789eb8ea4cf3c2bfa32a5bca8f1e651cc61ce47f5b8dde20f3550a550524eea745a47ac04d3233f234b5d4e391c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39348f225ce95072b08a6cf7bab46a217a492f5ae94a75acf303331ec4a9ad5e5fa930d3dd25b7a9f74fba2a61b67558a0350226636e5d42d0f9d2887707995a5b2a1d86a46ccfae4d2fe81928ee0438d8df04fb3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a5298cc1ca8d477dc60bbe9138c2237b551606310d47e0fe659f722dcb45d626253453df09eaf014f35c6073d7611b19c13bb71c88c8d604abe2c9dcb475975de28d447721a5c7faa0778b1d01a1514f368e0573;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d1728e1da2601c834270ee1bb919c42032b4bc740a9dd96b365bbded36504cf5b860e04aab7bbb5a7baf82a9d6a6203318b027f9caab6e9625c9ca7e95dbeadfd864d4cdbe67633e8db2a53baa33c713a012e4f3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c1c64b5858a9aa89524a222028a89647e935097eb5abfcea41dab6fc067ab7276a3f5aa865f6d56b6cedddbcd53a7bb5eff657c1f4c4739ae98770fd67d9b056d7f803904d2fccfd41de7e2dd216befe24556334;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d9178411f6fb809ca7f21fe8f80c914d7df2f99b9d88739a6d5b82f089580b142a7bfd48ddb5f94064470953a1a2020ce2b8143b873cc5a843847c7ad9598362b78a97788e9c63e49b0268c5614f84ed5b409312;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78335fbab2d41d161c710a6a47c3472f9f349f48aef174d58173029fa1bc4ab3935169e33345115e83693d26d3d4f954e70c577a4c4858fd64b0ee9901e10448f3092dedc38d3aca9e24a2b45ed9bea646f74058f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79f5767eb720e7e46e2a647f71e4c0c8d69f030bddc05c55ec060e9b32a9ae517f78b3f570a7c6252942488066906c17e0b039558b918a3ecb9711045c0a6944af59ebb1a30eaac33265caa44a3e0dba8bf5cc48;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfafb60d45e67550e927794fa19625f17ab13661857ccb39ca57a2b209d366ebe9837f4c6124df778300818e929f984d3d002b4b5e6a97898fc53f2547eb09a0719c58361546480f7226e3a114ead677449cfb2de7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha265218209ff56a92b1eaed5d5c6660b275b11e70b45fd72074e446c8bfa0b50e62633c35d305a3156e40c01947f0155e590a308b2b8e50920ed498736f2a24c469e0ceae29f2dcef2ac079d893c08198201d1cc0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4cff76ac0c45806c60dc2817fe019633b9a3231bae35369254f1bcceca88a1a6084dd97ee167ccdac58495498e29062eebe45af5ecfab58788834169f00da44ca4f85c27940d227624b765acf71578a890a9e32e5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a80798bea2f00794a4583f582ba55023c4a37b4ad242fc4c659c723052c6f507e5068c79c63cb9125c48f25e43308f416cb4781e8c813b7549ee760f85e10b977627fcf45e842726e9bf4b3e26935fc46d60c556;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8fd1957c15fd239a29edc2dd5abcb12d1cb0a5b167b7090f658e5dffad59af3d5a0e85cf61e6e08606387660333d532af58af23ae72d871a12d8d43ce5270d4a55b650701ae1fc116b62c7947e2d97660c125946;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h299415d2dbf549ab01f28d2966724e699e763e25e2af511445bccf96fb78266c6e8552d8a26c56115caa21ee542269a99e879d331da0b68d3ef901aa8309162b3d74a18c5e89e09f528c7511239042c9e5560a9ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he416a3dee6bb3f88d2db1424b2d51d1f890b7050b5c9331acc991c37595b4eb8ab7cbd95d02256e65c9bd7f0ed0303de8291587e2f948902357b47b64ec5455e9080050389ac5aaa774c78c3e27375ddefdde3f75;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h978bc56f278b86a22cfbab4e6db684962b974ed88383800c02f6878f63c50784475e4ec53c0f7d8f031bbc377408a36027d724b60a976f3434adba17740c1d941decaca17e25adfff580ca466f77ddae91338ef80;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd438cb8bd8b1d937f2eff2f2064385d8fe3713fa0aa767f618c7c48992ae20ae5f32ac0dd8271143f298bf2d745e3e1aafb8901a5ffb2c92753de30b5ab14519abbc2bc4b0536abf26ab2597513b137f14d8e8e9f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h133fc2b61a1e340cc970cff53f634b64427474b35e16066b25d6b538c14bd79a2df939516d3a8ca3fe712dc61fa717c1b69e651433be3f751062a57c70768e1a79c4b28417afbc9beb6541ce4f710c80b89b40c7f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6f7e26a6ed125f2fdc1dd3d04264846dcd45f5e11eea1e8a0752e2f83a772f263f384effa666495fc05c4f6b01030e046d4a9dbf4cc0510cfd1bf5b07262cb76b7adc0ecd671eb7e4e748048971a1e9d900538dc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51871da878940c2b5d4ca640f09927e621205e0604ff7990f6878d2985992b321db58ad41ee813ad7172950f01dd1799abb74c0762f5bff660595100cd2eefeb5d10ac6b04083a60b4d5dab80ef15782efe2d2c0e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52a6e3a2b47297d2ab01839cd1b4943a03a898cee9c5ea601e64d5790a42dd648da76fa4d80a10274ddf08b0ed8ea10e222de797365b7b49e9f2d089c8e4d2d3219991e4ed78683c469d4840dd1eedaca0ff28ff8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8a0853896fbf8addc39b87ab683256fc033af7af7701a4edd6360d9523dde80442ef9dbd538521f38c385962816bdac5b5ef51fbe2644e19c9e8912a910e2401bc6602b3f87955096f611e09ec6bfa480731257b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f7d0029265c5eade3173b4c00b438aaecdc5f189838e50a9bc947abf9bbd306673d7d430c6e9cd3122d6b93dbb26cd4f1ae6cb806f149cdef783656a3fa3daaa672109b01c0b25ab9408004a840d5ce7f183820;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63ea78a84cd7ecfd7e5fdda13aaf134efaa2d9eb0d21b247e34c93d090dd9d5efc228da2dba99b6f3364dbdbdd555016bd1a85217e51fcdf2aaef41c3c260666f03cccb514e1ae17b4c0c3d35c316e7542d77f2a6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1f19d6701b57d31d80814af4d21b4c3878594a29c459dc992212ed4cd63bcdcd33274d89b9b78374fa39326507ba0dc42f4a97c4f34ab4f44b078aa95c82c444be3fa25e00e47a11422a72c7bc7cbf4b2733bf80;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8f9c63c234c65782fcbfb4f6883a70962ba8f7582446258895480c5dfff85fe9337b8f3be6a8f6d7a7b52949cd7a47ae229427af0c93c7ddeaa6055caded923a976ecf00e8de6259e5cee3298fd0039ba7a0a688;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h499c8c46794c639a544e853eb6f833851d65fca8080d4f81b47077d48ff7d46194b2ff9ec74223499f2b75c9fb4e08d3ac6e540c4913d69e32a0c1706b0eb49a6efafc531d48be2a8ac39a72028e6bb43c68ba97e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3bc4b95fad3ceaeb5c5ec9b3c0524db3028e9a89809252157c359c516bd487e5ab0d8b0e6def7c1de48cc968a9c8bfc3cbed8d1c7f61413f9daabfb3e603dcfec253b93df0813cfb2e6a864a0d890c7f1f4465b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b2cf2ce7b7814f54de913c19a47b204b39d947049d715745d98644f60855b53257c3edec0c748239bd3ebec0efc2c6ae1792498027b630550f7b7b12b2430bffad3e9cf7590b8938bc7f20a2f178997330ed47d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9d080191ebfe83b76be17faf9f0be9addf5a98d5855a58ae07e2d115309b233f958494ac576948c50646fade96be5414c3c6d236c9590e97e55c9bc02b097c5816ac72e4b0abedd806c5377dd1a0deed15711e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h786050ded078ef3e299bddf856caf3c3bdc6f20de2d4c8bcb7a10f45032c32f0d01b43912610d4166db783137570604515f94c80b0a33139f4c0f5854042e1638508c027304f485cce36ed961a9de64f9302ae4a3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c989cbca82e7f8c13e07c2dc653202f1f02b13813c0f06fea05d3e8e8498907a6abac295d41c539ea91784774d71a0fbd7417ec59f53b8b3ffbfd8f9725762fc3836adfe9bdfdd014668e9c17b70fee902a775e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc67b6cd29a8f8b745397e0087d468216258622040added18852fc1976bf8f62f661a5c8d45afd1215feab5f4a2b526e32d2a7709be1b1e2a846719e0ea5423ec4356c210e229010dfac79415a4acbb118100376b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h641eedb96c9d0974f6091592f7b61c08c1e590e94feca4ae25d966dad72d9c10e307f6a69c47afed977db8613ed5c484af3184729b41877ae4194641a25273f568a6807eb63086b065e1d8f9b3653678f24f0243f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdaeb2d99de2d3c2d4b0dfbd3efa394d3764c127781fe6ca9276fa18a7cde58db86b258e76a487f5e8d88af7eabcb8d28d463e974092ae4057aebb6879fa09d034ed287dc0192c40c1b4066e86083226aded2071dc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h719950ce6955aab9c7e55fb01172403d06dd6d5c1e7298822d3c2d466ebcd1c2942e08f80b1d6cc93548570eb2d4d537f2bca45259d3bd56eb8cd27bf8a6321c595fba32e03f930918797b22c9d6c1e51e7c4916;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94ef20cfa861a8c31065928f5e53b4b010372ab48b9a7b0f7a261c3ceb9cff3eb70d17d5f0eb44c2057b6cd985e5c64c764f082ff65058db6d895019703fe760cd3c349f1e1e5386e9ba72758a475ddfdeb4ab502;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9b195587548325d0d95a339f576a7b809480e59db13f8a4d54ef02d3403c48b451c64a3f8e0b9deda574613c4f6ca7b8bcbfeb55b039e916530ec901a48b3c94f3c1631a5dd8f8da9b43b87e305493356fe5b3da;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d4a00247ac453d87c7dff502608935b9003a14c127d6bd3eaddccf24a23c37978ceefdb22efdf554ba5455b11de46df4ab01847eea777fe0f9e2c57025924f5b042db4d7d796fa6427489428aeeba2bc3640dc20;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc442cc41d4b5723a1c0874136a5b8c89ab71a6fe81d74a726c51af60ddc4259faaeaa581e465a9776d7da979b038728f07024abb23a152eae4181700f816e39838169107259edfb8553dfe36b6a5b4b3e66aeeaac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc62ec2686239057fe1741e7675489f9a964b08de7338f0e1467d1d9e350761160355bfc2fc867c0b7473a4d23eda4900e0911996954fd277d382b04461a6bc07b2ba04492d65d89a34d2ade90967dd86afcfe9317;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54098a5a58003cca70ed4d001c6d4a414efd560cc4468424c6536adaf801a028aa875fa7fb1ad567dd3eca5c7584f77f9dd9b8b9530994e3ba7e7e85452cdd587b4a6f148b0de924f2786b7698c94c8e606e976bf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd27c719477ef0a33e411cf817b94e0ea59fb58af2cb8e2b821f20cbb68148bded86389ec675c132a7e9e9b3f9b033987bc6cce5b17e9b7977461aaf8e9172a158b874858d03e8f187405a603d8a7be76f0503163c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47418d21d52e95111baf3ef6b82f078bfab7405d43bb81eba3a7125771fe8c83b3e0bef75009c020b1440af3faaf71a3c48e4de1a1569f2acaf7324118abcc089af0555426a07bcd36da72fe71c2a81986a020a7b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5b83eac897b3370b5e23cf3fb1539e1a04b53881cc81806199eade70d17981d013de56a6bd00b26ef3805c7984a7e325c618864d7d71d324ca5494a6b123ab9c8d0b137e08ef42945f0ef57153efdf1e643a8a49;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c5582a3583c5e4438d938b728b0d0781513effe6ec7d8be60c7f4b92aba160fbe713dda77a248305ed90745878bfa4e2d3343c292102279d70c131a1468089d9713696c6acf14f949d4a300594cf4334356cbcce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b4a6d888d5129a51719f826821acbdaf7fc6f47eb285cd7215c04caa63f187e0917301d19893963576b9df9503f5ad19394a9a8393f5a2ef05f97b24d917b7af25b7d60f8d8e1beeee3b3352ea3a65ba13a74daf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb1f03295df2a2acf9c70e2d1fd2a9f43ca92ae5cc30fbbb1a86b6bac58a34e608a67764ae195eccab74a93b2859084fcfb5ca7a1479569a7e84416168b2104e61c0f361f410b114943bb8e97b716751a18f6d7e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23b9c8e1b5e9fb5bfed8fbeef8ec2904d162ac8b4bcbfd739e230625ea0fb7d9a8ee36df2714d0608c2feeea780499520e80c331878a0666e1f727273271c1327ac912696d7b51876d5ef8d208b1de58b47cc2615;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ab14b76ff7a375b906149e01a52eac2c797b3bf2ec3553f31c0a415cc42b63776c79b8c9610c3a7c989f031ec8afa5be5f75dacfbac63ad0ce1cba5c0655abffa3e185ee6544d499237a41f6f9e9ce632ca4059f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c6d10f01371257a13f5feb6e9b6a445268155122b9e0c38e446d9141465f508fbd71f591ad714c8069f0e7382213c3378682bb6fc278b0d1fab52c1d10d43730b0158af06b3771267d85ac467a6b50a667b0e36f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d04f1331bb1893bf5da37cd9f221c3b30262fe53e827dd21d94246b2da3afc86e8734d64baf7253986a8ad960ecee5183fd23b3ad678e357f6939ed89c3af23e3f9c8a3825953d14e766db62806aad7c99bcd2f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0d908642a58c85c37409ec390ad7ecdef23d7dc601771aab7494156aa0870761b58f4cbcbca858713a5534088971e61bf95e427fb356a9e29b4134c50586f11ba31cb8bae3cb422040edcb980a3a7151a431eac2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f8b2913049d12433b0b821f18c280a4c0708c6802f1817d44f40aa686eeae77e81396fcb424176b1cccddeebb517021541e9ff86fd11cde95164c32c0d350ce66c2ff77a067c51ed1c192b5e9af0d2d050967dd6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca516c7a6cc886000b131e449340ae716d6a3609cfa483cac8a2ea0f1272403bf7f8766a2a799b14a39a45f2c4b3322071e797c60a7bff323865d3ac8ab94210e60725cfb8c6b9d61022dd783966919f69aaa80b8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1abe8754d6354d9b5c720a8c96040125279353b5c4da9bcbaab42da3a5cebb332bde95d106bd8f4d3c2ce616097b26871c60c25a59bce56d24f3df4763078afbfcdaf01c0ffd68eab3b15a0d6ad4313b84650952b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4c1f8532b237ec4a082c6cb48cf43edc4970538651a860f352a00f6cc292d90dea56523b42f2a840f32c3cf0df3a08998d517b27072088c6e03f857925e82d11a10a124a19631897bf4436480f3ccbd1574bc338;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7161da6d7195f2476144349dc51a865cf946e07e014c502203a99e335aef759d75020c7a91322f20848cb8d08884d9c31dadb088738038adff3d2e2dcfa81e4eedc83bab07cf4be94a0437ed4d1057902fa5510d9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h538ab094fd033396f9cef468df13acca2be5e2e453b4635f5365395d1cf1dec593b3a857b79ce91874fabf0de517d439a97ee444462f446b5dc734a76e074610b8f9476b04c070fa496fc4b06c595e83a28412fad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h417fba55d96ed3a50481b957e794addf13a9747b072b291e9ab41ad0a171baa3b0496d459ba330e6ac5272bb55a2ae6092f7430af35bf5140b0b17c5d057214b9cb7445fa3b607729a2af6b2f406ba16321b809dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57d629791bdb96e6804401f0b893f64a748eade6ee98ea23eccdb85b711f243303f6efeb0e3057ef17691d7ab2b9086a96f5e458614457668849d2085855ea0051508bf4f5b3f3884943ce4c8dcb9f9c0bc313887;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7a804484def19b402865f87271c76d02e95f2e15016ed5cdf98a0ec4be66c627bbf3238a4ca126cacf71a1265ad90ad3b8fb494d2687895df0184b852ce7f1851734e852e52e3406c24d94946992846a22300abb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab507110e541f3795b7a87b224b87de2245e8dc646506b8d60ed7b13a01cf5efd5e47db3a203690e8033613be669fdcecb85de70919084fd4374827e013d47d55229d0f0f29f23b868e16ae6666fbefabe6e95def;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3dd4d8a477aa42efaadb491af952aa7b852fb37de18490b745de9640ee90cc678d54544096858cd06a3f40dacb083cab5e283e5f6607e5c82bc76a6a890f2cd80b6e3fab6669f7b0fb9c42fa553850236ced5f387;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56357022aa78813632fdfadc297c33f4127ff15a7080ef588d3d5899830d380da15373571d5a48f99279223faeea6c343a0145ef90915e995fe0b94a012e1995ba8402c0ff6c949bf2a0feb9a94a3024bab33209a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb89a2f4b2e155e52f43e325ffae04bea1caa39e30314f63dd0d806b9ff3edf32ff59fd599679426d6848fd07ed19da5add66d71883876bf4af8bf11ed83e1a7e89e7aa107b7800ea2abf07cd358a1afd9b23705a6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e8e3b6c4c9e3a796a02d062e086c98a00e6a5b2cf1903f920b92d345dd98c7107ff8ed2569e39e26037cc08981731f83e281f611b76def56668f682cce88a32171e9a26012261593acc8e5468021bb954cf7f2d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9caf1a5d0703c36367bf9ea08e17fc1dce0a6bc512c1e1fe5e906b5e58e0a76df41c86234258f012e1aebc19b67742fd1fe0254995ff713229d4184086b00d7c6574dd73cdd74936c33ae1a051a2196c68e799949;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf3d4125f3e159c12b8cf86b0ed814a950a048424d4cf7d64a4cf123bb618c372221aa283a205acc58f7408b90367382c95abb3f627192e643b32f05cf1345e8320f66d09a15538f615a09079a7a4b7f51eda2ef7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc691f3c2be685204ddc84ef8da204a0d85cf8d440a4cedd2379558dd96216d1317df07db826339e0391ac18c88490335d86270a492dd891fde2176aa605053c91844d383c473d20f733c64d2f2a6f7c903641f922;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7af65d6d12022206a2cb3bf00c3896a1e7828a6423819946083fefcafda1b3d352662256d4536d940a9e988d17a7f57733a95a02dc94258611fd2ad87e1601fe078075a4f26de31ce70aa0e8c980f76acd8fe0a87;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h916ed1843150a229595a6376da8c392044ef3b7abf7f0c8bec5ca854adb44ec066b9715049445a50243292280c6f1d625657582ae286a0fe04ff7fda4ae1d91308bf69d944e5f381b45fc907c15196590007ebff8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3209f3b63425f2142d72b2fd3a06bbfd99efc85e9c9d9d705ba3dcf7f7cde20b2f1135a9d619e5cb75313cdce1b98ca302f1f81bfd13c9e98378b14e32eeb741e371cbdf1e5887431427cbb8f8e437b42391a19ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d94ef38a0dd6b50c676463caaecff728d833445f2778519be3d466479dcc5a915845c916e81c7a755b03d7bccff996d37986fe4e9d76b978268b2dfc3da57b7918d474477d0a72beeea8239144b0c2afb4e5042e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3239c3977477ef9bbf62a6dca98aeea0dfb04dbb3283212d442f952268da43b591f2ea620a98c9657a224b65ec0f7781387ea527913afd10a0d7b938785e9861d6a6ff8de58c09eefa0fe5c697a39e0a9ebcdecb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30f76fbab96ef99c511d79cf94623051117f8da8699714fb2df6f6dc0a3c81399cd77d306299e23f9c0dd62d8989be3c86a3c6a68b600be6e6f4559c7d9e3023ad73432094f865b95d0ac227ced0ce21b8b7f8a19;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b80bf56b3be7e56ba63396772a426a2f567e32f019fb9b5dde3da2ab5312d75c84cab8c518b15a1e556ac99048158670af9ee9116319fea430a0c7ec50ff9cd90377cb0752db5a4961ef60b8a74f0db885ebeb4f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1022fd22989162d1b05ac1f822bc88d4364490cd8894bf5fa2d32b46866b640545ba0518cfa28033cef5cd4697de8aa67392e1dbaf205d162926e8dac223edb60f0f86f1a078e65d0215cc3cee4a764b3d9f648e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c77ddeeae6ac563d11fe4ae70adce1ab758ac9e0141cd6a80179c1f5ab2628469eff0ccd0778b9c68cc01e674c242cb97a53436dce62aa338232443c64359b81d7a79b18782935cf28e1c7928d38badacdc722;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ce31e31510785064cda43b4147c81b566b9642560cf23df48ce7e3e79e6f55aa15a16a1609b97b6d984abdf43e4e42bd676e2e1f6af5827a8b742f70cdc39254085f8d97388a0c7de3a845a38bc773d092327627;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c965ee19704eb3284363bd51d68b55194acdd19140d4cb82c402dd8da2023e3043896154c395e6126cc4e44aced339698420b185d86538535165f062f4d0c8eaff96c640b058fdec5ad3af18c1a387be8a677207;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98933dd802e0de0d99f534259b7cba287058320fafd7ea9a3f920fa6501d61f7729eb3c4862092df4d251af31106dc581348fc67dc6afec3ce52e0ab18bd186f152aef1ad5355291bd1d296d53da8f0b419cbe4b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hedd52d564b5360b1230026b35b92b2ee4acce8a4b2fdaf191586331b76b76e710752defd085a17d512592100f70bfd099c874adb10479284cb9ade5abd6d276419e8e8f2d4f3b471f1356e760d97dbac2e33f790b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9655debacb7eaf5445c4a6b7dbeb52b4264a24579a7e045158d75f75fac4472f93056b1e0afcf0ae60aa92970364da37d52127eb61c0e49ffab608c077dfc618e6778a19fb552a103e2d928e4a6d7d9370c80e4c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hada40f28e767e6bf42ee80008e708b7eefb759d5a7cd6f126da2d0e988e18ee7ac3ea235c1c1b301604dd6041d84b9e2da8bd7b1c426a2f7d18e0e09c700fb38d7172e5b117f4a4d135d7bd75b73067df4a4c2559;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ab9a207c205f6d9014e798f338961c66d8bd19c47b92b819553cf3f591b63fe57815baf346896c9f4e813070b2267181ffb13e6f30ce58aba1600c8c23c9a34d5a0261f86f9fcd6a22f03e7ea5f7ed7dce35e79f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h403c58ccbd93d5b774d5b1a99026526828ea059e4a8326dcce2305600b3ae98be08171808e70f2c358b7f54ef22d08ac87da0c9b74771d71a12d5f096fcab2bc80c5bb4ce2e680f5f14e12bebea496852865c7459;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d81a820ef9017d27fc369b03f70a7aab8c3a3cc46bc03d92b4e5ad36ac661c48666554c9a628e60f0d15fedc7529907b4d3b8ea8ab6fd76b0acc01b86ce3404dedaade695df91d2d6c83c2f9229fb14e4e0dda3f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa42c546444ce8b666004bb3c57005ef1fa9ae8b82f2f3150b38d84e6052a4cda777a7d3929139c5a57c6e8ae4e4bcd5d876ed5763e537e86d0c7d70d00ee02cafccc17563ceebf469fafb0b57a633aee0b259abd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3345296a252e26ec91736181ed198a8f5bb901aea2cd49bfd0044629dee832eef4d34355219aaf420825c75574916e08603089fddd339ba84fff19373696252a719278a35180cbd3f1d579d49833b43b230f107e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he871a099ed2ca8bbfd97161576cb44eb9916308d0e781d623d31c954274ec22467f87b3e6cd490b6275bc42fc9cb9b7db08e0b4844931a5f6fb9ba9748f83d4dfc8e4fb592afd7b81ec68ece2d9bf62214165ffa7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc19b1c0edfb29e38e8a67c73ef5a10ccb354915d3a27b96e30ffdc5318ded6c215345ac1542a9c9ec1d2e71cafff6d9f48a7ff3b8bd580709554110ee932453578d7ceeddab0f78c9966ddc9bc6d16c80d6a5a6c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb15211d527f91acb151bdd283dd3910889073e8ab1d1bb001e328f563624f99037522e7e89772d74a25d257c7be3134882208d908f0c0921e67a6d81b86674c17c1c86399cb2a50d1146cde36137c38ec34bdf17;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb809462b652b42314af51a5e70f75a0eee616bef5eca95ccab37c1190f4d4bf6fcd5bbcbaf97be9c97351d94dd84817998dbac6d89921659daa0662510adeacb74b4da38b58e220b95cf39b8d3bd15a3fcce925;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79c88b2dd80938ca67c14a02afeebc6705fc71a8a7801aac6431b227c96bf07c29d2d8ba0471894466b2336e395fcd02425fd33a2c044af3eb2eaecd774dadce5bedc082a6fe789e567c1498e4a2e9de718ac347a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h421fc2a9be60a661cfab54182ee493ace4639c7c09dbe837b7aad2b8b718af6e4e217489351182445bfd8faaba20bb38d92f6664cd8bce2d68ac4a3416116dc11a93576b4423e9ed9b0fc80b05cc9ce6a1dd5129b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h876a82a1d0e689fe67f5ec13afb5b173d2fc580aaf31130a70203bebcbf0890e7b909cdf70b6c1a1172c04b2676c47f118a22f933194a6417c583cfedd72d5dfcb6ad0d94a657b9571fe59391b97a348ae8ade66f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3992fd98a9b45cb5c9061ee6c1e03569699d14f71c450af936a9c33b0e67c99cca7f90643c7e601745cc7191b84ce87d4c8ca2459fe420c4c8bd95c8856b81e3d63105213661c21c25ff6e764685744617150912;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h74720b2186781b6b1ad6a5b10da01fbc6b11ee2a2abb5fce045ec942ada80652b9a12c46fe6c5a705102e30b5367614030685560cc672dc76b3e642998bb9a3a8c5ffb7140eb931e023dddf88e94522d06db5c60a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a26b9d5afe9cbef1cf855bd6ee199bbffda81dbb726c48040347c0f633d030bcd2d99b2c7896d1c003dc162b8fe376c8026d20d137c584dd99755681a7a296121926d101a42aebc20a46690c4c346654e287a157;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c26e17e9f9ed51467cc5f4ad1c6202053c41490dc1f892341dd19a983f3d50c89c47049aeaba8e764c1e408db534819d49f515d0bf23b2f6ce4aa6fd77649631eed68e8e2fe984a785d9737785e6c4e732aa9eca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc695c929adbac68eaa9128bc3b55f9393c7ba0927af353cf4528e3ade76fcd38ff42f55c382dbe8203caba5d004c5f81791ee1b6ee23730290518f5247f9bba1d6df6e17a381f43d4d417deafa7873de616b9963d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb366fdb11b66b60b5aa1928e2a018990f52fd4434c9150313b780c46213c0602b3866d6979c7bbb93bb0caf25290fc0259363f5e130a8df222bb739658c7a2ba6bfbc105abaeefdb5f665b10472571d6aeab6a86;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65449c5a28cceeeb8f18937927e054ab8c08e802632a07a9ce12f57f486fb2f06c256d688ff7e3b7be9d177b3b0e859bbc4169db116a0c16e2d8c68e9cc799b9a736238d3e0f16a91dd857283b4c238752a55f857;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28a7195d1a688ff6df120c9303b98c60fe93350ed97c4c27ee4399dd3e98d45709ca054f73cd80c28d65c4b4648b4a4a068ea070bf4b10278b72268b9785e620ec70bb07c91a612fc0fbe1f3f799d01d22534a215;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h721c0a3bf658404b40067bdef5a609909a08cb100aa90b1569f85b896e5ec7f9b26936d6ef0f91e78988c2670f2b2aeb218d68eecd4e75c9118fb6c0df647adccd55a9e659b0630ea6f387379f5bb356c42112d14;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac1cf562a1e7c883bb10eedcb976350257c46247b504cbf992c00502b83ef47112abc641f046537eed9c093796719a4b8d04d8bdee21fd5207c07587cc161b9da4eb306bafd5448a2db8e6d1c795e3f8bd74fb4bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f5d67109c4cae1d8cad6ecd1dfc622e50d7a9c6f1842d4fe3b8eeda73261e1d7727a095fa1192b14632832dc45155049b87b7332bb26c16b961f40e41608d1053098645997121954f4928f88dee272cad5d0144c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88539a9640b15d99e0e2d052321912eb45f299a29367a2d66174308393709f4c182f175b8502daa77427c2d01cb2a0f833e665970eec94a5d4d57dd69a1dcfe5013935645451f132c4c34bd04ecdfb1076b32692e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h275ebf24aa7c3d39149b04364eb432261d0bae04fea1fcd3e908a1710b64a442cefe14f062dddcd0fe7627dd824ece597bd535b8e23130dcb3f6bd7c7cd185c28480a3a5ac54245f7c7ed4ee1e5fd256880b6665;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c2b9c02115a5c6fba332538ce3c6eeaee710f57c3eaac604da5e0299320005f2726f99a68f51f18a91b21a5fd215771f007b8b43503f5ce03bd40c140dbfcff715d72b88d302c384fe416c56d3f44feff709c1f1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha4203ca5cd5e70101696381f533edb9158708dd58fba90a17c3597185984e5ecb0f9544ffd6cccaddbe99907ae1e773e26f786c79bf73fc82debd786ca35609813cb9132324e73c86d90d37fab8b16698f8ff059d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5115b7464940afd5286a2ea4255815b7816f88ef0c18e4ceedacb5f780e3642f1c79638633ec6cc14c7f5df3786754e575c26f22890e333c312f70eb5a0b8f5c8ba411db7a1d9040aa9f1a7971c72bbfd50dc1adc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4086b89e315b4d1d4e923c3871a53a47d9b4eb76163c7b2e8af8a7786f6107379dd69efef2a385898b56a9b2c6ea8ac576de53d30397f5f988d66c89694ae460fddfaf5fed89116e0ebb1240a25ea6b391f8c1e5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h190dda6335d572798e2d3be3cacf20a805b288bc65efb6710fecac519b81375194171014ae9b5a10aff1e9de8a78d228ee743cca267dd455c7485479dd2fb28adbc572d986f16830e0c1b0b9873f3b092af7d1262;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf513a681a9ab65a69ed0b35511d22b96b91338361d3494c93791cc05891060d5c201572ba95bd060b4eb1d2386409adddaf8d1de20bd6125629a69ceda5a4891b362e3ad6c7fcb669ceedb3bdaf90653297edf01f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65058b2404b72166f12b7942f217bc5df09e83f52b19a490a5f9d7d38837d9a6d2ef878573818c967aa35c62dc6e6ef485802958d6552b15e4bb5469126920853b726bfa96f8b125fceb9ba2db774e058936a2ef3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h152fb688bba49febb56e424d71faad4526f1a62c66e27a2b24bd5796fb17a5055d8288e287d36fbf1539a312cb38609f05bfece5ba90743e09a1102c7414d33948e045a8559884612cee5a56a0031cbe19e7babf5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h573993a9376582fbaa3169d75418017a0280a07bc52885fc81b50172db576a8b5c97dae89745d5cd0bcfa79e9ca174ac383096f6ae3443cd14f06ad0f37c56c4670cc0cae41caefa0fe7172943ef4937a75d2b34d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66744f8f9a792e3f45e03b5cffbc00945b6b4165e358444909a8d908d22cd681efd7906ed8cccf278629eb448d0fda462acc00bc996e74eb20fcdecbff28f3efaaf46103d8536286d5eec98e8d80883401f189e29;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe9d9040324262106efd4e89c5bf6b02d4b0d83f60faa2a1c75a66b4f26fffd571ca8e1f1694d151753472cdd2bd4359e428d60cc8eba7246a707a6b2a3bc8dc12619ac34bb778405752962df9183c2514d4641cd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39be5cacc958970c4e89daee18f6b345150894faba2ccc2006d15be434f41613e9c8085c5cd583e7390b5997f26ed4b9957351eba58f6921a09079d36ef25ff6a15c16e4909fe26d8db9f2e43e63c529601e9e0dd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha4b561984644bb5a6ea53573cb51bfba087070e841192003c88f9ca30338da25f56457cc401346029b4c47f8245b2c604c13d9f7d2a61bcaf96696041b28a31d6a1885ea2759d6dd0f0ad4940d24ef8bb24a5d96a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbebe324b4756c157dbcc63d66278ac6344dc52d8cbf5793d2eb73de54722d72f7fb0b0f32a2530faaee669e060d9d268a4f3d10b0afd93bbd7c92a1b9a8319586b396b13bfb0ed05c1910b9e4e1a14e38ed1b7256;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1441f162bdcdbc9878852b820dd4b7da5a265c273316f725ca3c56990cbea51fd786d5a1ee685693eeea2935f7ed86b0636dcfe991789e561a1e9e35b69b2c950ad5a0b9aabf71992fe78584f1aa05afdb4f3b394;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59f8d6f9eeffea516235ac90e3bf00923a223130ad635c9ddc1a869ea40dd4a763ef8459636f1127a897a581556edba97c0682bed498749df6cb78ef226a329ea54c90be7230751b429b1f8136436de4de7ff0af5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had6d6770b6f43ab3a701d5f9a06857c06a0f088b8f7f2506c00a15a33994a246abe7fe54b65fd0cc70f3106b06ba6d2140669e73a7b251eda17f61abecde40d58a5faacda3b819e6e8f48dd728b3f89ea723ce82d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3591c5b5bab99ff8c33214e664c268c45e34e9b634b65cf460052b7c03c0b2cc9369b2bd923335834eec072b60297f9ca4bff324c08824b17b352f742be8dd28b45214297fafb0f6ffb35179ee3dbbef3416fa3b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c0d93a64a0b594f16d895fe39f92a2546a84089d0cbf13aaf21f9dff920ba1f00c238f4c725949a6f1eae0d6109f46f8a28826f22433ca43f141c13b8f115f1b1c4e84366890460962c20defbbc345ac02f5e277;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a12d5386278d0c7babfcbcbdab49c2e4bb3e1c1e6eedb650c30a4590f5f4bfefcca6eb283c4325d6f31f88c42a738428e757be80e76c17cf54b4e5a86df762cadfc18b8b0dd1b6a67add0be908dcc6a99e337fff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97039e8be9d4c7f53f26ed8d4af656a1453cd95750528cc566eff44b28aba369854e1b59dff8a0a73e9af484bfc4b7cfd1f2c158cfbc4431d4f9a6e6b730032cd987c590d6f38692d697fde4f51e1517e97ad1795;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h828505e8e5abf00a9c7f834fce71c64edf0060f5633b8eddd3567118769fefc7d1f51ccd1640a1c32df09cf168c40d51a90e9b65910b2d6ec23a32938c30cbb396fb6353991accc91abd0fa947bd1fe53ced4afeb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0f1544ba674faa2724fae6431552649d49a2dda49745f562da379380367e87efb812d834477cd4ee0449c8b2c5ef9e6cb6c0f49dcb6e83849f0b7a703ec119b90f9acc0ece5b5feb07ea41a027142f991bc762c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdcb616f4b6468524b0f57bffb3baa58431cf905c01221efeef4ceefadb98fb39fab02aead330641f6cecda213281a1fdebc8df1d0022fd29e7e525f7364c4f920b1c5e8de24b88f521644761a12f0e49cffc668ce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcdd36a60d6d965917a8ce7e233d7c8809ede78d603f7c984bfc2c19a5ff310c55cc9afd6f9e14164a4c1b7ae55ad39b0e1918862b630a601fff35f8323a9cb47014c7344319d892a0df30e9daaef8160fab5ffb5a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc92ebccfdab728d7b6bbac001ce6acdb00e5f59790a1cb22f0c2c63e50095ac1b83d5c8b7c2a7cbbd8a2b27632b942956b347c32b683f825da9dacac72537d67d63b6aa8a9dc1389c088d2c6782599cfe89841a52;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83f3b74b847b86ae77fad57835d4b2010b3ec63a759280c29e14127a28336853101bb50b1de521dbd645a1cb5950eab6fccb4a0b4826b0fae3be850a5c19f41063e0f76003901a950f9f51d648c7e5a7c273eb136;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h639e8c7bd7b20c42209971a98fb92a7d741b2ae626d77d560ac4fa51537eae961b0c910163abce1f4ea631bd5efb9f2c44665423c18f2da19a890408bf42b6e8ab25271dfdcdfa5b32760413daa1810b5d911a4bb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34eb904fedd8f2479c7b746e10fec0c69360fbf6b67670ed0f86d0179f01275f574e67b0b37a6e07b800122f52bb01cb52f2c1a779e04d4fbd9cd59177c9c2ac62ebb67cf99d279f917a785058eff734478399fb6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e244bc8ce73801825aaaafac49de55d328af014755c8fa50aeebb81305bc3a76d23e6bc09a575409bd1a3d6843a462b663f037fad407111ddb33884eced2dc19a1a631448bf0bb42377bb0265c32d5974782ffcb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80a25c1466c26ccc62badfc06d92528b65aa0f32ba57af8ff5ba9aab47a8f0a6ec41d1e9620813c7873af2a4c2977f765839131f7b3f47322b8f217b9fd9949070587ab556c0cfd07f468d15b2b9ad236b5d3b756;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4de9c218b6808d823c3153883d32a3aa90eae127ae3bd77d707f0c110638a4d29735ed05eaf09ac07161405f017ec56d5c8cc16e9d4fe2362c27b10baa147c724a570fdb0f3b78b2c4ea58e8def6a8da4fdbad098;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h319f78ea992e9393e93048866d23a53789f10b4eabfa07784eb8a80c38b3c90a9e2776ea1a156b81b78945849cc6b539fa9ab98d37e573e5aeb68aac3ede9b51ddf69942b5aeb533c73d8f0a7186a706a77b16e1a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68c2d29347b8c32d6a6efd1195de680db1726234e2a8baf085fb908162627a6601795d6cd647662dbb78b3c85db995a1d1a0fa7ce370955670d772c6ddb6e236fa275fbbfea562193081cbe325fe0188a423676ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58fded157945017d12d94b03e97cbf01051a81dfc078543f07a1db9f372d8acefcfb6e92b95d3996061becbfab5493e92b5fa9f838c718c17633a0a85a7a905e0f45d322a88c4044e7877c121aed4df63355e8799;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he02f471556d6fff4a5eeab018f193e9cb3b99ac3efa09c75808fd9336c05a26036020e9dd65b7bdfb8a20f4bc51df88ad31b5b2b7eb42d78d8ae53cc8949a1169daebcad20455f48918e0df3691e7107e6f8fe761;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb068bc2b5d0f2d0e9738b449d1871f86ccf409ce2b43fa13aa4263b8bb8c792404c391a98fb445dd9b0406728a899573c4da5233fd20c52f48e5ae5969f682035306c61f929529fc7ffd0f9cb94bfcc29e29dafb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfedb66e3318b568aaeb52a90f1fd189cbae22dc2c4859bed709b38053605bf880f2be3ca26f17e1af18f28ab24efa5a4701829e2abab0ddf9da6b38890e1a98e5686cafcc2e6ca6fba4dfb668687239ffbfac1207;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7be30799093286d1fe7730bd07dca2211ef42a3af5a7252c86d054e64265e23966a8498ea35a00eb2d322af0e10ffa98000a1d410172ac68b5886c720ba4aca9a564004507a85cce6c8c788c8c99b5c37f220dd6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33569adb49c2c055a943a7bf7289281c18f195f6b02e880599c3302fb2f55020c01dde59c0dc9369324e36cf83f90df48c44983f53a2df7e0fb00dac39d2b075cc5c5311b00ff738e58ed7a2a8df42b8f31f90964;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdd33ca5dc2f912084d593cb5c58c8efda162a67ef6b6fc19fe6fb50d068eaca9fc5b7aae6fec9a2e31afa024c5f318880d2bd8032a54873e3803e07f2c15c1f99e52e2640233c07f14d57f3675ef1701a2596d6b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h960b9b04dea352f1f07494e3df783b72d048a0b37f4db131fee3abb24b8209811a918a82f1d471748345601fad408aa86ba74a572588a0d6b276c07929c77ed4a193a15e3b77074bd6a084d28081ae2843cc16577;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd48e9d00e168d47fc5d400a891b3cd7c20d2234643b4ecdc039172b44eca788e99d13bf1bba1d3855b59c5c44eb7570df7b21d4d7854c71ab0eb723bd9af48be27da26c1dd02601f3e586c28311e51047d72ed779;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f1de75a2a6ce6a561b91014eb361869c07dec566ca5aed5a540c7ad24b95d92c59212ab66fa789c12e3a076189ab502bc5433d5e4ad551f374d0178b96984dc2739f91a71e547132565bd9d2a197b607785fedf2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h580ef904b90cd219ba8e9d4cc9c5c863bb12ebd31fda2bf87bf4dbeaa8663b09815fb981f1abfa2923e7e8017962e9a0f95f55dbc53f1cc49a081b577455d5940fc787906d74d01a197d1f98a344f3fd4eeb613a0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7b862257ac1a960efd27524ba679ff56d5a2c6714ab933b7be59e5c5bed490da06b63ae6ef977ee761ad21cfdd488b83e63e71bbf797a531afdd950b57818a27ffc81e7cb9fc127aa762f8e4dd6541b115ddeb45;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a0a1a3e2c9fe1dab92014dab9d08665501c031d371131d4a5d421be27077b0c82c24abb98cccda378dbd1f92eb681a8a32cc43684e0089e0fa98bb894e2803404af9658383b51cd04f907a9600e77cd7d82f9e12;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65678cfeb4400cf8aca09f991271c29a2e2945ec11b931c7c185f7f52a1b6ca883f768646ee9c179da3475f4fb184d9558e3d8ce6d32aff2348a22e035d3978c96b370b8391f579659dc1aee935a16e0ca489fa03;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9883efe8a871139627e627846f87f002487c2ade2eb46c911c0527989c060ad1a0f1fbc8dedd79d2796c21a137ee1e2de1f8065f3e8a4808439b2ce7a3cd6f60698abeed330fd6abd02a61815d9215d169a8a588a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4bd25cacacd24221d3c3ebfa5fd1f55b2540548e408cfe5d0e744ac30912348c6a39bbe2c9c584c62207be177b858cf5532bd290e835a0df233ddc2fff55fc29f3e89a068eb7b8e598dbe1e5536c3b2eab3eea0a0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h457e074c27408eac2d5b4bc9261a27241fd83902d17e3ba87a40b25e2c4e58b091d42f28892d8ec555ee0818e1eb6e52defad5301526fcdbcb17576b200840900dddda2dadc340bf62e7902cd3191f8d0511843e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h552b51c404b028b33ac0db4db1d32c2d1e3d241245dfdf3d567b1dc47c70078c0e34a18255efb724fd955fe69265ddb7fa0f033c4c764a383a6a5766b12b599b8f8d73a4593d2e2754b873e77f6681be48d0bb5bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33d02ef6e1c8eed8d2e1cd218633c1ccd6e64b66f69bf163e3fd08fbfd6575aa46311f8879a37d9ead801ed3112aef47a6023de2fddfecd6ae864491e8e5bb884bda2d775a162edfc7c8c9ecfcb4fb39e2702d438;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc01d67bb11064fa7033fc74f768844d1d039a8e7b633eb4f134a0d44887127128656c9802df6bcaa856da8e3a1a1954e94be06321d4fdeab40ebbdc47f4498df2e63f65b3738b0ff92937bc489284e37952d95cf0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1dfae169424d07f26ca334d6fe5276812729ee01562f39567c40ee16701454f3e3e67bb7c6aaea5eab89ec7c7eab10c7cff95a01d4e9a752de90e1498715f0f0db0446cd8e54f82a05aef887d0b463e8a59bf70fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7cd774553c0fdbc9a7750d29cb530c75a6e53e94867a3715cb71b0e19ba5188ebfe3b4b07068d8399664abb9b4465c5569dc3cf1ab4471ff121a648ff79829de78bb63b8c1aece6e7dd1044fcbba49b4769c4c22;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3bd4d0aa7fb28265164f81f9012b78129990d83e2bcd6ede9b6c4650b1e140dfb7a5c54b8ab8edb17273151ce13500fd7c329d43c6863a5e9454a5f6fa710e139f3dbeee330cb44e09f989d80037cbb3e51c1bd28;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd51509297cbac2e5e660c625e4c43818654c4a1861cdc290343cf6646432ca71031dec11241334cde81a664b918218ebb45a50e79a47826ab8cb4df8ddccc8c4f6945b23af212379061766c7022489d447aaa5f57;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc06d9c662e90253b7a53211047252d1faf77e7bf9e147c46ef96cfe56482a0d8515e573b0e0fe566ecaf0236c23bf9ea6a76026d778ceaec5d4ce2a65b3d99d248d83f7535bc660cd57e73b0b8de0473bddacae5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d3f59a3b6719401130bee95a69d53ff485554028521bc39924d2e3e800a24f6fc3da622f1a620fd9fcb3fa3c94b04a1db5ab2f97f977cf5fd7cc21ab5d0055d7fdf080b3b1720ef8abaca158ec8ae7291f7daea8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3bbda048f972bf59506720d948c3df0e6e027405ec5e1d0c3694fb692293a76f58985a9d6ebeb0e3cd94ee5b57395ff3812d431ccc11ba0f4fb74b6a371a76aded1750fc417911d46e06d175c1d79fd45099da738;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62a1d36e083ada67eb333e677e74e497c9ba0b802a6e706d2c4bbf96c09892ac0238c1a0a966015c279f2f6e16c8545877830350325cbb8069ad2379f75ed913d5f08f8bfbc710ae2718a277d48578385e78e86e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1a81612afd8107e1111e7f986c06de3f6e3817a79bdf6161c0810c33899653c1b05ae554c4ac61f55eb339f184acd4175090b13cb4fc6e529fc1e6a59d2f8b3c10221135743afcea71584af72ae01aaa871d89a8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd299257349ed399645eb73faf315459fe4b50c45caba89bc983497b5d2b5907f82dcda3f3f8ac276c0e559de5d3d77c6389b780c28a44a6fbcffadc3179522df2b573864ad54e92db4c15119182d3115b4594fe56;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc516eb9f8f2a0b9f37bdd56809ecc6787cfd95422a0689196b058ecbe3ab5326457f70f9a230565871072cb4ab0902643b123d440c329f605eb1cf153643f05c8a88e2e5e4ae65250ef72632e79fb5df8d93b9f29;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b0a4531ceb25e623fd5ce9fa4595bee08a6fbb8f0cffb9bd2e3bc5e004b2983ae9e41f07165c49e49602cfb64d98a978f1fe9d8b3a1ab41516747085abb5f7163f17b6c59a068fd614da47fcc26124a7d5540b4b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h341e35d88f4859f4d9d6b744ea90257a3819973b68567634de2a3d8605bf2b282333a4baa0eb0eaab84f41203a0affa475ebe6ba0a5db8e23c06d86675bf908e3be0d4bd59bd0a16d1ed8c00943c2e2eba796dc1b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1feeceea234794bd76efa6c53b3c69303f0d02eba3ec33b111682f35dcaaba18056ed28d2d6cd61a35c092fc69a837f55f02e48a63a342785ba6a44fc711ffe11fa3534d9024dad62307046d7e486ae97b0856bd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd260adb437d8dcd0547b90eff061821da5af4be7d4aafe1f9bb2d980b8c6e0f72d21397282ef0b9e4e3acb72b842b8d5f5f7871812ca3eca258afea138d9763765af09c4be952dd5972c7cb956cb29e2e9c224048;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h602f6bd7216fcb104c9162a12c1a6f00c0eeeb6e2ca176db92dfe4edd7c250a292c66a7612b6be38c236cdb30443f2b44275cc1d9bcb943113d9213c3ffb6675cc8fd82d0ae90568cde1d63ef179226e2d44f3c25;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heff7dd66c6b684f596e6dadb57b9b1c603acac7a53f26afdc4773afb173d463a0b690cd2ac43c55bb0fa1df723f7aae118abb2078ce3d8ec801066ab92a07025730bcd9ba84334843444c502ca84cd8296a4a2873;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he16bf4d53c5776f61c2b347e7ed9e0c795998efd09697ed2fac2f79a9b6fe4fb31c42d1fb86c3c193730d579f16edf5440f79f06addd69c4469c518964e4b1a269e31da0894b640152b2409ce44f96f52d159ea78;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8428928f40d968914e8d08e78eaba3c38283eacf6b073d39781c0aecb1a0dcff4f5bfc79a9f022504ea2f7facb7c3850240957ac46a7de2028cc3211957ad03e0232dbe6b89ccc5fa9d8f83c71d019ee175d7bca8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1e47971945bc24cba4f1fa6a9dcf51d9966d000454f9f827950ef52d9db9e3bd66153d713665c29538ccafba0b26737cf7ba91c2fd4fd8e96c59b477fe0a40b96580fe80660b20fa2a928fa910ce43bcb69ccbe4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d3ab98170bea7bc0f2caac2ca366d0808ca168dcd54e5720478d66e375507c5f5fb01a00d029dee7481200e8ac961f011127a9d6cff64213a86ccaee91dc56f208444578d504180b1fd180d712c495300214b207;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca94dfdce9b6c714fee6935c7ed8c5ec35c6d3bf973dd3a91802fa6dd417e473eddcc04871ce99a2eabd34ffe7fbc08571c7e557cc522af2108bc3c1ac4b8e19e54de9d7c8be27aea470c00ce75ac621d291ac209;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17f5e4721cbc15e8bbbf91564438cb5eacac49dc7939ec0339d0861cec243dd1a4e3c4cbdaed38e8a305568a583fefb8279b168270cefe4fe939ceeccdddc8fa56ee1a1c6c0554c0d9f04fe1c49ae78b9c9da8e93;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5c53a5f0d49bcbdd7cc4336fc2e3f59f7f15a4ebf16156ae3e1445b5cb9e8f7f4f441bd76f4a50e4aef6d1bbf276368a7b4ad911e6a68337454f0f0b15cf592888f4188658b1e67ae8a7ef7b718164af359a3599;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d28eafaa5aa1bd02aee7633fbc2c8ed68a3682c74efdbb96c7351bddc2db2cb727c8340d34a0b4be46bfa8ecd404b036853249ca20d36b53a55b253ec779aca38977ab574823e57c52754dbc9983c40b7e238a27;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha56e82d2a076b3f13f277c28d8d861dc493ce4120e0e42552eeae5ee6fa8dc09ae89cce77363d89da63e432ca2aaf2162e06eac1291c8e920937c0af474ca44941ddfae4334628e556e3a123d429fbb6e29cfa2b3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h154f62e0d1bb78c1a8d5670cdea01aa24e85f174f58c797aa23f56e687ea2fcdea120e23cb2125a94d5c3978bc0b1792834c86491bda005f5dbdab581f1c404586bfc70e4a998b9ba67ad6558b1f14887e1ddfae8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb80abb6c6cc41005abb23e88228ade89aa0ce9d6fcfebab6d39b16e0c82a043b2850f02885c69314fbd32d027827216ecc0f2febd43aa07b83ab913e2a938dd3d8e6b5ed39669b489545e964abd9d6971e93414c8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d2adb43224daac3fed33ca4e6a73e9f2529009b03f3dcfc903c6b406659778bf1cfd318dbed2d1a418644bac406fbeb2a4bbf53fdc2a8ec8b434e3654318cbd4034b70ac67c6c17773ffd6b901b6376b759621fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10fb188992f0faa5841c7ef066d1c7236c4713f0ab8cb4661da18493986041f248c32e9f4b6ba2ec688b10f59416aa11f7c1d5c224afa3af0d9315b9f5d7f4ced4cf8a719a10ca7f45fb11a2b6876bc017b5a3919;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67ac3c287f5916ffb68de3ec872b789530e12a24ef4c41f733d029b9d4b20c9c33b05baaf07cb27d81499e65621ce669501c1a9aecb36974b39f68e1a8c890ba2099a7d0509b77694ceb52163b488a274ff4d974;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97bf952593da816a3789dc28335cbf41483bd72009a7133ecb3a58eebafa9a28c43392e47c5f3c47c77a2f3a267a010214e73eb2fd11852ec6c7514753b283f509bd2fed3f3ff8e2a847310d124f18ced6c2ee664;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcded2750dc0332475577ba2f7c2ec22ed93fc20035b6e0d859a13bcaffdb0e55e89d4fe4ad5c01e83c63ff47a3f445f645ef68ff4452458d7fbbaf31b7e0f319ce626c8f2dd3f45f8cd036b13abcc1c73786d5f37;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79ad3786712eb091b45a76aa990b61a61b5c07c2c311bda2785129232888b7428529bda859873d5ffd4b4df65df77b8a4efef6d037a3f4de8492e6e5a951513aba73d39a671661977a25ad2cfab875bec35022655;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6cc408e700cd608eb5884407ca2d9d305994f3658b51ca733e932558aa093afc279bcea2d6d3357129902ed4cec3cef4b002a499ac58c5c8f9f1a7ed90787b2e42468b06d23bb8238f056e591e807c1ed547cec78;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56b7c305b75df16f139d3bd95cf58939dcf9b50dfa9835c0efe2512881aaa302571dcc2ecd4131db75bda9944e21895dfc21b08b8a66036a753ffe4873714c083d9e5568f82fe90b3848f2ac7490f3c9abb05e1c0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81ee10668c824c16af13381b046170dac98246058cbe03350c71ff2e813ccf71926e73f8f48952a4bdaf0ede8282c54aaff10b1ebaee1e5ac56693fc6eeb33507afbc5ca6ba857fce6bd080799cfe6544730fed24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h487c043e81123f0a6083dd1f913c7469ea0f889b14fc1ae00f2b5d558b57452273e6a04f35bcaa2696e1f49233b62b1d890e3e56ac3792ad86e2399d8d8cb608b96dc48ed39f409ad8978957cd8f0732b1f068433;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c2946c63b3e738cb78c0dd41098b5920e5ca19b48ae3a9ffd7fb20a15f462d499a538b526c8a678b9b28dd76c487d5f56ea1cdd8305568db9815138d0a0e3384115fb5cf27e24c488c085cadc513560325c5778a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe011a02b783e850f9839b775d5eca8230046a6d70109011e32fbdd58a0715b0df316734247ce93ec6932e3c67e0490ffb2a444ffdf8d82085884d5b6e2a73d33239d9734201f0968a6519adfac38b98ed620ea5c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61d1d2b947665508e251b8345d3769039699a7ddac2948d3cde85cf630f2d1d2a45b820b55d65f5f9b268a73584a711da1ad80042ea86816cab6d9d6a89568894ee20c03e015912c3e25f60103e8374f8d27fe576;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h471dfb5d7d063c6e9469f03c0b49408282e7e7c02aaa1960fa8b25d1d874f0b9d0795b30972044a0da72b82f87b4dbc62ffd40ea601b02731acaff38fc64d0557562d333223923fe8a14bcf8d2999747b0a672f82;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ceaec2dca600f2ab52e9f03c111fdf7d70ce612ac076e8008a7852aa0bb582f1132f7619445087a93a7700ccf566b3a598cce725cea61f3c7146262895e08c5ebec6e2578a022ef943c9b3e83a24d5387aeaa355;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf9ff0de73670d9e1bc26344b68a9a391d2562c2d433563407ddd4bbbbcbb800598b222269f75bbe6d180ed2710677c26d11f20d9f266e59031e89aed343b8a59abbd505009d73e27f8d8b79ce710e4c313e64c98;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1cf05655ac6914a32afbba687a7d410b6f5ca8c6c2637ffe0b5fd582e265d6192d521368d98bd4d0305bc0a9939504a3c3c6037a15383c27e572823bad8be429336a8a06580389c424d62f07092d3c02edc6ff23c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70d2f4e63fb4e06dc2051363af0284c3f630a92ae947ac7f35b29160a607d63195254e11abb3da750379e36d0f6a2352a8e63b166381a3f6975bf9a284939a0e57af70507931b7ee570e1f72a8918aa4cfa6aaf4a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ee6711f958fcdd31c8dd36487d0caf021b0501337a6dcc7db0dd8b2a19ec44c64fa0ab262e738a5f71d8708ca4071491004ac229f2d8d37e46a6969564f9402b9d23a08774cebf558d8d022d046e768eff91fdef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5bbaf9c8ba8136d31281f4fbfcdac0a89e41d24e797f9f81cd43503388045137c30df46ea71a10120208fc10f7f6466c2bac55ac48287fdf86b852e4a5403b593cb4334c86e6fe3e85dbdf146714c6bf5613af1a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ce15191bcee3046e07e2116beae486067f00d511e8ea59a278cab035b6ab78b5b98412ab9309fee617a005da8fac1a039828b094ec214402acf2ea692e49a9e16d74b4f365b537fa414d8f449c4b542da4f7b784;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8fd7dd3484c965d93828b9909d5e703e3566b27a73477752e72d59df504f74da771845ba0e620066bbde82514ab1f6879fa8de9c70b6928a1a9a0495231c052a610a726ea765296151d53144190cb1a2fb009055d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef0f9cecf9c911fb05df763b64aef13ee41995e76bea045d1b11d747d206e3d61833a7632705ccbbb25a3096800d240254f14853f6331556c6825feded93ac3f5317282dcba95d535b62a82fc63132d8da42af389;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50a3c2c66f0440d41f7549d0c32ecb53713066d18552890e03732d3fac3017c71bb850d0ae3c0ff12675927284aa59cb6ed1b01cf77bb54d33516db97bb15247e86ed3e02b922ea95d64f7f5abd58cf6957125256;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h488be17391584b74d653e76ba14a9ced69ba6ccb55feb80d4cb46f2ddabf4470f6094dce6a41c196a1e7804011d7dc419102a6ddf685f55939870854a5911567c35605b7df58ebf4d218d5a06ad12c9c9cafd6ced;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd6cfe8072771056623acc8d9c31662626fe8a1c03823fe1ba39e644beea68569025eedd110cab1f598efa94ec4df34142710d6e931905f1dfeaa3a6a3a85796e3b010c2868ddd0546692f074eb860e6ac375d47d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha43204ad66021fe95e61c7736642838aa6b1b0883c5b6abf998867aa28dffd36d7fed6cf5cb303ab394fe286c8e8ef386aa0c7a959aa564e05249450c218d7183bcdd5ebb1d74ad99d717b32628a2a65e24e60cf7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f9a8ce97e3ca60002f5ac0ee1948c6d6ac52c05dd20c1a57efbb6fdba94606661b45b80ed8aea58aef2af93dcf45535b18ce34d537edfe75334ccc22fa28835d499c255b82990ebc13a097271fb30ca19657a10b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6399e89237d603a9efee7f005c9971074d69fc7c5898709ee05ab3f5798f0e812ca1e380ea4d7e29770adc2ed035db3f2288c93afb9ce353df0ced81cc31c916a95d8b5b951c3d7126b8dd4e998c5cf6f8f7c666;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bdcc8a7539d8245e554d913a10471b311c6b00fba12ffe5d8311f5a2472c4ccccce45556dadcbfeb1367491b87504866746f779cddd7c1a893bf96173d3f780fc75135b8950dacac4e38b2267a23e2b1c4f425a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd68434be7b58ce16c9cfbf50b66f551680b00f08d715e63f968ddde16b466002fe805d3da36dcebef1c0188445fcd09af89a021d6e0a63bd6647abccc93ec4b046558eef9e87a7ddc12effad1d578675750323a7f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h848ca38deaef314218e6a7ce7235fad8413684ff966a22737fd5b7f09c071b41caa4345e005e378e58865661297eedde9c02c87b058023323db6cdff0d38ff523b2a52acd3821f907747e91daf4b059c4052d5c6d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a9fbb6c3e49a7f355f6854aba6dfca0a037c497bf9c30faa3357fdc946c371ce7108aaff0278bedb466678a9c2fc9071082e0ae51906b5473631d16851bc7a51cf43b498a34cba2b49332123ba538edcfa274088;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f00f9d0bb30d6f21dd82314ad47f77c18213543a198c294c7163157e6e8ba7cd02c8a2d521b2cb471dc218f9110fa425b33b799283c2712ec2e554bd88cbe59a3f6f8c0507358102567805e841fa2c434bdf38b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc6d8554fc93631f34a7f3fcf7d4084759778b364cf1dac3c04286a5d2900b927c989e13c331d8bbbe0b40e1867a72ab86be786184f29135e68da202125963cf4a6d4229915d6e237cde25edae70a3589e8253b43;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66e5b43726d2b399e5208751b517209feb6fb893983020a1c66c5381da9afd0fe42845f121743d75607cf783f8d1934c48d4cdf5c7288be9d1d7a3f0a550ffc5771471bef71a19eb229b1fb38284af7c19cf7a0a0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39066b9fdea8f29016677b76a330d101cb04396d4555bcc1ba91b9e4e110a8a4f2493e0a87411b766e0e4fb83f913f56fae5f9032fa07dc81fcea5b82290fcfc6463ee99da0cdf18ddc2c9fcaea30a0c91d868b80;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef314ed57450dfb8fe59d8371ff22f6f0de60f214b03b2514866b6fd0834d6eabce07e2da4e49ab5c798ed7ba7fe094f39e9398ba00d1fda590e779f30b039dd3ad9e747cbdd378d09c1e27aeff08f93611d17d8e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1b6c7c6979f78406ce3147ac9eb6b45e72305b460fdfb2fb8ddb5c3d0df6dbb22cfcab62b8eb5834b6d96ff42cd31994b915134bac61e404f59c8e7c85b134a57a5cdad4a8cf779aaa7a66211262a7186cf698e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdae5054705228c915414d4e153ba8398bd5feada8cdc8a8d7393ebc25f00ad8dbf01c6f100fdfdbc475bd4f51d9051f3b42ac881742b55207ce8328e1a40d7e765720d31c5de3841100f2f724fda879791f343df3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3418b1ce2409fbad7cc2f6bf13169992fb7bef183c90b63a63f1178eeb05e984629c1f8f50925d21a32d56038641d00fee5389a360956d49495cc77315eac6cde40bcca2cdebba0e11e8dadf212b1c5f77cd7cf06;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3e62fe97c1ccbd60952c6aba3eefead946aa9711fb4e2e5683acabdaafdd55a3b755fcecdc1b2a8398f9cabc5a3981807d4b2220d674c5203aa050107150eb52758e758e3403970dc982f0d13b9c8fd4e6545624;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b2dd1ef5709cc3acdbf8a3ba0303beb8a17af2b5b3cf87f0a48029139d6b3864ce954b81cdbe0296cbaec8bb3a261757f74072f6d7b1ebf5c1fb50c2bd563965c3cb57561bc35197d8e491104bde0862d29054eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6dc551526f6fa79b6b178b05603f4f325d7e6bf0d4f120982bc4839b50d97d3827ec59a62aa7faa62e9ec33a7c80232cd11fbd71466b179cfc0dc15fa571c95ce8649706f8d562a2cda12758693c32680cf6a724;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcde6b91459d6340881116445485e3353d27bee4cb2e2d74996e3fc4017e652f26cb9093acb4bca647ee08aa8d1df2dc85346def0642f6eb89396e88416fdb3cd107a1d253d4bcbb5390124f9d76a6322ace9e605f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc7186401c1dcd193064d4dc5823dbaa67b05384d78ea5361aac6aa2f9695fc29a1d124d4b190f47e1e455c47a3ebd662334ec0253470a571ca941fe2ae18199719da59e55094062c298286d58da03d482653f57c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb40e694e9c4fc91ef7cf053f2245d8a330e30e3c244d0aabcacd9d23e537ce3b4dd697b674325e4c25c675426944a3cb0ec701bf5e9fe079b0e986ae4e8d84307acd1f725cf78c559a006802a0701fe083e74da1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23d12c4e892c8d97e9620b81db7a6d99e3dfcb22dd627373a5a8c854d94b384c08723b12a3752631e4a38819c48b47d144ae422129bd0a8a0b701bf743bdc04eff3d8f195eb2fdf8793e3c0ddb65557f043c7253b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d214220ae992b51ac9a4b228858bb99ed1bafa8db47a24c0354d4a10e410069e8639c4b91b9fda6734afb4e2ee70bc794043eadc33d8268579f7a38c2fe7a531fcddd68e43c06a3bd33e3f3713474024c94920e3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11e1d23d24e3dc6f8d1becbbd137101978a4d675fe386254c3ff0f9056b32a6fb2a164cc6e2800c7f6761fe089e87dd198a1af92dec6df3250f8d1909b1244e0680f9635a2e1ef986f57c3c23cd59585e6bf42920;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he234c38374ce55a7114f7c1dd9f28546ae4c648b90ee301546c75cd817d5aa6ce08686b787b5d96ac78a1477396ba87c275ede0f97a47615673cdf515c415953d27274752bd2cb47ef0d66fa38b8c69e9fc40148a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb7f1a838562485fe26d7fbb83cbcac8a4104f9357e0f3c95c19190f6d86c55f98f4679ab163952edf4814faf0b8ed05c7e8abdc9767c6a306ffee268568e78fe4a691dad8cb7e3c2f3c43c71c5c4893299fceebd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha827c82065877c518548fbdd87a1966d1b622f55233162639a2b448f4d893b5b437d670f20ba7a5a0c2f6f389e562a39607fe7867995f737bf5ac03f6afd3621b18a84f1ed904852e64bf2f15ac458db3cb96bf72;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19e87aa5c43efb0bc6f4c36190ef79f3e02345f02fa90dc02cf25128abbb5069e6713df64d442ba41cd9ccf44e9097660320a8a6b228df625d494b3b04d6436f86b832f57ea9b83ba9452862ece6ca56da30c30f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8444a1e593c6506029cb3b448f574233bef7bd8f5d268f47c902298129e95f68531a711bc802a4b46b5eff923a7833cee2fa7785e0473a7a11ac652017ba85a13a8c08ad2267707171b2c958214e5d1eac1e84030;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb6bbb56814b157e6bee5f71dcbb8248e5baa71698fb45f61a9c84d0f2fee53ad6e1584e9a387477b94280042d2cc9541c9cdf4ed26c211d11e0db57d1d0362b5fd8740c4a326ea287b8f049a0b67c8a83e3c86d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h449a3a41d52ecd3e03791d92b29750302fb83afad2ee0ede75a4b4399898068836aa34639876d4710df347df4516911b499ed14309272f5435673bacc7fbd44d929b639766999bc368bfdccec9505fd0cf8ae8fed;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d4a078bf9b029d7666eaf52fcba8a1392103b675536880a851193e57a64236962b98a60b620b36b037c1ef9dfaf2005de01d3660ff71498191dc7622bfec2497af858cd8b3301c7c1b8623c24672dec53b4c9e22;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2473334d62911c6a84afd123b0331bc0beff9ac1913b586e7decdc09ef8df54e0fe2bbf1223cbec9e54711b7f16d9aadd5c046576f4c6ee5180c20b42b88a926364ad082be0ba01fc5c83ebd9fb2ca5d4955ad36;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee66525e67c200e1de41e1127e8e826f6183c6ee6cb842183433bda9b2e32d00cd76c5a131d449fc9d1d9af166604d154a49b12a241d5ee4a44153342c9875d58bc2b22e6e7641a04088fe48935d89a55bc760777;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb7195261dc97c910feeb27a363d6e0f4b8a9a979ac1d3776f6cc577b1ecee04e5c400f4e1b0b59a9e88ad0339f46a464e49df820a103bf06653c38b6f434af01fc7d04ac877fab477e70ebc72ee2d9191551c8a8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e8ff461d51bac72f5cbce00db44e5cc8004b522e729dd061a865e925e8a193839c215d6194ed434e32a72038b71f44a0778f02726ae1e1bebe0ea92f4691bccd446c49a53a7d7c2af90b13cf2e3a2394d1621635;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc555300fd6aae2403a766129df261eaaf28e23186748350c7da754703ac11f2031f7ec8f47f1a15e9db4502858d0253a914565bf137363dcb6d015fd9d6e15be458cc4514ee0f18cadc08d9abe33383c331738de1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1dcdfda1a40877375a9b56f98019ea31016a402624c63a070a62672d03798b7a1b17b3615f9ca69ffe3cb9a2f5479fd69402db16f3b15d5dc8482e0ae1d5d133137bd3ad2c0221ad564d7fb5fd8ad0337b284c3d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79ff2a03ace6b5e2bc2d0e07a7b0ea46b4d81da3b263484313499ca92ada178a65b41c0497850fc7fca1a5c548c7e3cf56af3aadbc8134ae1649907d13b43624df4856e9a06fa0b2117c501b3a5dd997078e451c2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hffc9272dcbe0fe1c9de63c05c14af333834552051cb95538db6f674df815c4fb3dd39d0fce2e8cc5c3a9de93fcbebe167c1f9dbece1d914212b5727abb1f3dff132b1ee4d455cbbf5a3c0ae4dbb7a191f3dd828c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4566b6c0d019dc1afb303970031991357bd0294aee87090e3421d2bd6b7c66f30a40179600af4396bc6596053c33132c8ca8aa24daa4056c15d9fa504dd44d714aff67eb457b4f2837c1e6ac8f2f3166247d09e09;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66912283ba1de4fb37dc5c0dd1abe32106f9856e1a45484a5e48ff2c5771fd56e98cc822ec5631031b604dbc07620f2b72af175fe7a13561425ed03d8f73b8a4bb95d25fbc1969b939090e4a076bfbf4441f60469;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32a344d073834abac94f2b94514accfff22ad6eb5f2ea24326330aa5f1dda17f535cd8208c0bb0ead67c246d685eb4412ce5e4cc1b213a1435f026c80ea67cb5f143dbdbc4057c764ddaf3208f3c4b803bddf8e9a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef5de041649969138c767deae20185363362866e85daaa64d4360d0cd0a88be18d5acc28021b4cc01f5048e8529b93e6457f119ed5b758fc5649f50b5baab875dc876fd7410eafc966d501aa62fdc09ecf6304622;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h899870fe000ecadce76c99b0573b20f224bb419a37fcee54ee0f55a97c8488be3f19996a8fabb2d80f0e122f8b44106f681a2ce271f43a3882b96147ee4b39f93a3d062450f95615480ff476d980d628f1af18320;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43069996919a60af41919e996a7e8dd67ec3281531bc90ebd1e580ac8f4d38b4bd9c75eb2ea61483068401f7db468356ac0dd9e910d151acbabb690fea2c6b721468a751b88da406e2551c9701dba082e6ff1b733;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha30abb51c166e4c54bdbbc3cd2bb20a61d780ee37f13af8ab1428e378192df894257fa11cbda6ab39ef02e8ab424a2bb04b8d8c648fe8e2b0fbb64a6a5d41e2c87ef0a9ae04da8ec30077e1d8e0d9a560dbdc6ac0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd42a51979f8b301bebd7cfd73ccee8cf4b9e38c4318755dbde56eed407660519a90aea171e9afd761524a57070872cb20f6c889639ea71906ad6bcb75a15ef8f85c1523582a50e598e17a2957796a34b12a20b5cb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c9bbc1c535ad51a0a2b5d711dc0bb7463cf6ca8125d3308ad4f433e78f4ace08cacd06efff5e2d253dbf9bf5718e615f1bcf839b874ab5b7b4fe92dcf3bc92407d3369a01928c6f95d81ef6e73a5e88384ce272f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c935a9b7dac4dfb9f51b16a46fe11c48758b64aa1784328901f4bc6c7f0a90525ac0a2ebcd32df7b15e464d4941588e965785b287eca29da1cefe37918aee037c6ce80bd0c821799e083ce6aeecda25cbbe67df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf490bf6831110f8b5520a622b0ead38ccef804d903b4aad966de38ead324fa3d2792a7523e7ecee482b8c327d0723fab3f9a18b00ae0aea49518ad123e1dfe93664e2d064050bf2e37a3bbbe31531936708c29f47;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5092374aea332c73e1365547c369b4202a6ee3c566e220db71ee06e31e6971e39e90f15292419d1a82bd1701b542cdf73ea55fe48ee45c22b290c80d2b6073d9c94e701f44c521ef23f85bdcfdbb67760a43e030a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h435464c7d528dabbc92ef8044b6a96dd69f284cca134051f2458a5fb638dfa9eaa2484b334023c148adc2c4f34d4f45b2f6f5ee95eb24feb7f9f50d3c0bd4ff3fed67a4eeedebe2a6c9b4c562775910a0adba53ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2bb116d154f32a24500b53246877fdedc35dfaeaeeb7e921571d7d4768ccf467d672a72a26759c42c6cb83a1dbfd640afb4d9b7978aa1a457b9fe1422769f3cd671b442f0060cebcdcbe542f77dd5143b7d49abb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h550fe0c3578c9de0adc361af570a6ccadcb3cac7f6e30e5e63346abcbc7a7e50bf054e7e04a54de571bbafb457196de114a43c40b3e5ca467ded844d6818adc44f9bf3beec219a20c937b8ad67263f12b8e0fe106;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb6cdbbaf6d71077b32c533f6dd3191fb805cc1338f8379a994ad64a803164815e6c3727323e8f8391517de9f48ed235d3aa65137432357fcf963886cfa268b3e23d6bd44d3fe0139a45e1178f96a151902645c6f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99bf62ee70406bab08c0c155a230179e832db9b7a2fe1f4d446b16e4799355f5187c80d06c492ab163d84a59a1c590b9bd779f1fb1f2a96773a5c3b90c0c02547b65e9384e77c1ce91f1f2b3f2f073af23be9422f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7bb857ba06189143d2af2a9245cdd907389b872936c2ca8d732d97d80fba57431e60275ef65e1f708e033b5f52151c60318046241b745538360e2ff6126b53f0ebdda1d9c592f106d05dc56fb78547005cbca748e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd79f5b91808df8571dabf27f8a41facad0a8b6d7926cf9c7c89bef574c34fdd56a4400a4529b9bcc123156c011288c1cdc3e16b8143d7cfef3dda3bead30aaea64a18e974b794835bb4795c1f81b81288f10bb865;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf2fc46ec028a23038e66f1232e27105b9cf9503a7893dc79df831ac61e0b93fe5b6c37f0d908f86b60bd33494d960cff5834ce6abc3c4ef97b2e62427bb05e0934f4b99895519a798e1eced5692ef025f5301870;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbba9e6c159cdd348ce5b940f61ac3355cd27f5a1231e9ae2a6451a0fe1d2078cf4207cc59591e4ebfe4c72b9c144e2f29cdff855b5a3347f965eb3148dfdb6baec80d871c35ae0b4bf0d6edb7373c7e1d9e34a2d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1c75c28c6b16bee9053a928833c1cf545d7f6bc9ffbd8df5b6a2b563fb63163de5cb5ea2d5a439ba03418adc4f10e74800b43a7f9a85777c7c83455b46c587dbc37830a0094264190426a9bfe0cba8fbb6f4cb4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1887fb3c24f9f892274912288937b1eda1970f7025897e092742f4ca973e975e77bff73d71c6f127804cdf755f91910dfbf4ffab5830e089f0766b98964e9bc93242efe1d4cea05fd9f69aeb94cbdbe0faeab88ef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdcab3080da9b4535f5fea94acd1896b22294769e9c839268a1acbaada056732f4cd0022fa0fbfaf22fd54fd72ba5d7758ec12eb57d976613d7fb4c34bdfdfe496ce69e8ebe232432fd9e37f3e1d1e18f2adaa9958;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f7fdf9bf1834828df116b684f1cc26984dc6494d8ce6028d3834a28118e7d5dbaadf37221f6959be4465d45154867988001df72661735bf80089da74b6f83bce25ece5d124ea8ab3c0bb64a6a0754818ac4e8aea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8204760bbfbbe686950b4542e821802c80e80281348e05b17d6955cdc7aba4ef31a9b12571ff9718695a20d91e5743f19d58b8a3e18c3c601430ce8da74dc3581b6a87bc6cd82ca9acf706abfd135ab17c7c44c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5f5df39ff86744761dca0e9d810d941a66ebefcb6506d18632e203b9e705015a3ad5f5598aa77ffdc349a3cf32a42449634ab13a90a5ec59740be0bc807935166c8203e243a51d2a2025f537513efc3dfbb26f2a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d980db8c0fb14d008f92e022876a7c1b51dd185a6134460824c1c522de2a911df0de9dce8746f4c28606a263beca475c75c9e9b06a5d49246140006f4362c05e0080e02d65768e97877da0db4fce54f348945a5c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfad40c560ee8f0c71e706fbf50a228e10c4c92f100baf57a1e034a978229ed3b26de91ba24094f7817cd93043c57456bb0bd8028c55dffd736558d18e0309f4cf48a3e9e3f14b5842a043d80e9f31b4ad6332d71f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c91b94af5795d6852b51e63bfb4a0770703ef67bad5bf6ded71819139437ef9e0e995221a247f0ccab3785b3c243663f2b160d1cdc6c42131c644850e2fd3bc567b4b8758c9197ecf7de73536cbfbc1037023264;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b96abb20c1acd360d1c081016b720f37eceb0062ba56ea0b3af665ebee509b42f6e5805137555249a07c595728d92b4e6984cbdd90b96329d845783bd5d32aadd62126f3fc9208ef2dea028ae8dd4a25fab6c147;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7ab6ae452be615831e4490b95e0175af632b4dca4880b6629634d8d010f85f0183e75373f33c0e1c9c1560ff499013a975c426c6666ae1d5a5c80f52088a6fb45103ad283e0d19d8a4aa1d861f33ce978bb303b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h195409e3c407ad8578f53d2208fa8ab154381cfb8a66da23872b067174ae29b5b12f087dbe66746789882bca15a3b66d2ce3d9d3ed344600c0dcb48bd32145f2c954e5018f7bc950c0a84f3501218b7f7a2c34554;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd081c82b163d4e757fa7c4b3e3c45ea32b3df8ace69f4142dd1da630f1dadabd71c5f94fb6f1aeb7d7d4661306c98cef5a522d9ee0c721816db133449c27164576540ae9de65b182ec879f89c92f11adbc477073;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcacfa21674fe3e3aad9c4ac9de8142b7e15d3595463bc439f6703de9bbd0ba69571023230fb0a30a61cce81b4e3ec6c0fd887055b207b49f2127fd2f0395e0582e2b1c9f5a2a72bb53867c711562f8d542b69050;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h447df8d9041857135ed795322e62b80da982c72c2ce1cfd7766eb243fbf9978538708fa395ec605a577802c857f022862d84776a3b495035e3651b0f4cfd19988387973b590909f07842c251bfe73b087ef0e2d53;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcf8cc3966b62b33e161d2728104816b7dc792f4e360d316f0b61fa244cfbad87a9f9fdc4a1effb152552141f2f01372d1d5e562cee8d0c56e62dafeccd2112b05540b635e68f792772b3504c256680f38f4fa0ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcfd6515b84ca69b1c86afd798678758c86dd588bafa858bd1769649b5f28582e35bc9f68f2b41f0aaaccdbb2418626b2d6d3380975233227fec1f823a13e17945e28964ec520f3704c85033f1896890de4102d6f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a58ea407c69d4c54d388b9722702a4bb0406371844f4d9f6addbabcc5ade155053ff088b7ca45469e7bf5ee646d5897c66fbe116adb03323ac568952f4f24706958d7623b700ae1606a42592eec94be8798c6c8e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdde415593434b32ec2dcbdb169defb4c3117d996691849c065d11c8712adfd63acbe73713f9eddc2980842ca3882d05bb816ede4c2ed38b5796e571ad517a0fc208756ded4e512e7df70c2bc2d6d3a7d3813c04c6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha693c5b6cd92a9920bead7fa43d518647569c69f00639dc2aabb93fe200652c9554dd7e7036ba5a4b2526f969b383275613faae348c9430f4bf70e2fa56db437642ad7e0e65760373df08b8ef8c8b009faa76f676;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe7128850fe5f1dd4472ec1045b18cb8f34af2459feb926dfedf2fb410b8942b2cf39657b242af357941e0673281fe6ee3ca027e30fd2547e0280e52e9baaea073d4240f73c01f472d5d58c1653d58ceea44c5b2b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb057ff8fe33022b18a3e3408c60832d96df438e2ec814fe4c7b3efcfebef0968d2422dfd057d5ad0e0e56f6ed5ac327467e16bf3c9fa24e5027661fd759df44669f739fefef568b3002a0d4c6b29ee0c6d7fbcd86;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6d064e2d7783d8619ee362b165fb924f37c44d868c57115c937d0cc0b03e7ade07823219b273fbd3ab63926bcca443d99021e29b04c86ba32baad4a57f912eb83e69ecb43afb39fb91a8aed375f89b204e752418;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5c247a6f884c480fa42d87ce9b9fe218770580ed47612b4537ed78e17d5a42d275ff4533db5b62343867482f8d5020e49e451fe612383105e3627d1ab4da8414b6ef15ec217783fdd05e49ac76c7ddd2e6ddd32;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8cc7d99dc6a7d24b8a116140e6fd4fa3f31c3a8db44eea04404d9b4eb1c78298a429746119690af86d67381ece75c2c7b8dc7e0b76b6d8c7fedfe3ded54263f8b0936dc5a2645ede40c0fe62fd264065b359875b1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1d2dd20df422b2f8ced8c4428cef0a7bf1fe8130ac2553d90693ce8076f3366b720883240bf61ca7d3cca525e6ae66d722a200de78965db899d33e945f08ecfa1cf6c0ad40119f98e82e0e0f1216842be390b514;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd03f26c6ddabc1adf8ce34de770e21d356fa016a2f07cec317f40c1dd1d9f29cc5eec0adaa81c3d7b8a1c9ea9a4fd186cd89ed354fd2c0f70fc3c86b43568880528d7575ed7dd8cc29492e73bbae49b18c96c1689;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3fa8a94b7444b7325b0b326f597be187b938fc8cff703bb0d72d8d698ff27cc427c51fa0f17a4f5e4878adf521bc33c8874ab02f18ddd8b91868eb4138d45e7f712ca38a2bd21c0531004acb975ff734cb39f346;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd867f36abcd57a487d3b52ce6550d2153fd1165d81a0f18014d69bd93d8734f1dc7d77ac174de7d45ff5190a34f41ef1668956b195c9c36bfa14cec0decfb1ec68710e19340fffc9c06a7e3d41e405bbf3828d5d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60c67dc14c659788f762fd6bd2076e37ce76f426d5c2202f977e5f4ef48ed5fdc6bfe58d6ab9eca285c649df016832ba3b1fb9b5ec4254d216729f78c6e4617867206ee071499d2fa865784c11d8f5823bf1575b8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b733b28e31fca0a49a31afb4f89af1e20e2b6377c8332917030ce1924aac8e1d259c42bc43296ceb0efc086fdc6b6e36d3721a8421ac6036fda9155c7b6aff7bf8587b3ce8c7567ecf3e2f5f4d9c5343ee1a6d10;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd104445a5430abd20d123aec6bd2d9c02496d2711bedb488a3281914c2691f783c3e54d0c1d5e4a5096ac52c15f7fb3a16575f982a0aaf402c92df8e4cdefefb3eab491a0aad5ef607f526d3ae0ba5d45509c8d7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d16d7ec93012345e29092fde3466e40f53b6c5fc835f7fa5631ae2b1b62390b43532ef5e651f54d79035e9b92aef0cc3833e6f97b51906a6c856789d3d90f90417cf0e57965991db7a9f677f46e0027b3e31da6b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6f4a529cfb8180f9c14573a786642abb8d4830b0dcdb0a1aae9bfbeaa3c3328799737131154cdff746cc7d36eab8973fc8b66bbfd3bd64210ae0652a26a4e9b369d04351cc4fc6eb7e40ee5dd2896e4e4bd9d26f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h234d8aba9ef230897b558aa3c4d1e5de0db6fbeb1a9746fe758b136ecde5df7b5bccb657ed4e017663554e10568542fac3f42bafaed70ece952a6eb8df02e2aaf4b0b3bf9400570523f9d463f36c2414fe31ae0e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6fe9e49f13d888999141cfed2bed0be5a03537655fc5cce5a8f528bd8877cdbee62efbee3d203dbb45a2c0ab7a0ddc957353da39c8689f599ee6d52007dd9d408226a4c55b49309dc65524faaeaee8ccb90a870d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h685bec542a12a4bf9473d022b8aabdd8e464953866f3aa5f2296cce4b52f80f25d88593c246764362fbd2baf279e211d7d24d2cd383b1d631cbb959aa2bd648123e39e9c658b3cffd769a526cb9d70c49f9af2f37;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6060b022886d39a5f459f59707055af9c37a27b62a7937644dfb552502b63ee4e2e11d3879fdeb6456cfac18b04e78eeaf91abe8ce26ff775246454bb591a6e3566efd9234f01be1fb21a02b5fb33ec9ab58d5e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30c6f3cd672b706f0621f176ec7c14610a2eaf7173e4e2028b20bf6b32bbcddaf81cac3baa2d92dcd5dd48dcbab59bbbf4520b1c04823dc55061d54af562614240cbd04a8b44f8717123fcb65103b9386bf668785;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h874b8ff838385b429a8cb3e3ab97ce82cbf51c6cec85cffb5bef9f36bac2472392645c4fffdf3a47b95ca25f6439a9f7c428745fda79d0de62277a74e8b2f3c2f58e7219bd29fa54874a57153b9b98e3a3d5f4fd5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31bea5dc9c8029f41e692c0359f98021ebde2ba3b92c6b57149bc90d0a6bbdadbcdef73d5aafce24160531b77891780d4065636e2da7d31ce472f67a0ba9302bce44ebe48ac5948329c6eee66c3425fa9224830a0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha531342809897ecbc6af32e571037c0e5e70e957033a9a3a5dfacc09a6a2a6596fb788be13619c5e28639ba20c2641ecb85bbf0cc6c78b2b9ccbb6b20face6eaeab3c2aabaf881e88e2bbc34cde3ba51e134dc05b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48753a4bedeed4eff7905843e1d869e5fb4663ca7c8acd1abde52e6b87ce8ef18182c687c97fa2fbbd7487d69022b7c2d0dbc75f8b91209ac146e7ceabc966df7d389d8977ca742643d138ac9ab1cee4336b4bc67;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h890f3611870070458cbff24f396e65565f0eb09c2f78cb54e753243c325adc6f9d5b5b7df8852786171d9b272a597ddd93e4e9ae1a041925b2fb5fc1c55a9646bcdcb14d3379f37bd87844eb890578a079f507463;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h381087ae665da22be1833880b1a448e4cf97ae520bd32a9829e2ec603851353b4e45fb05be4ce9b9b4b327a314826883923557fc522aad89e8244c699d4ab892a2d088c2d0c0740f3bf433c673655d89ab23607e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc13f911cbebd019bc7175a699c94324090d5b01ac3cf7a6c22e63bcb07c201c6ed04de70c4fd9b62a102f7676e1150581a37ebab39df23cd5e7a2bcd1ebc17cf7595e4e5fe51e013f0d2c65a24ccfe1f1f8ea984c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79cc034cf72ff44b6b9f4d8c7df776d885710a6ff63bf87829a8df642ccad9171f677a2e047a57c7af5856921809feb69bd9811d0436642b05ab5fd00cc4b412d12dd613b1a8a258ee42d0ebd197c9f3b2b1916d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7d8b2c5b15206cb8b374884a8538d453a6fecb56fa4a7552068a20ed0197a69dd7e8ecccb940f81514f63bd594b8ee05e51e6863b541d3da80dbeb71c6e06910a12a02ead070fd18c1c294ee906dda5b92814720;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47313f635de380156fa6f4cdb433b0f0c2f388150e4e330eb42fc155d22035853ad50cf2316b758a2c2d3a0a2d7902fbf5ddd98a9694c48460f0669dd5ec83995620f75d61a86a02c636bd59ed27d2e1615aa71b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h712e70e6ab05043bcf9fdb84f0f973a1f8bfc59d7edc0d3298b6d20588293a21cc33c7096dcc54f3c99872f735b9260d5f368439eeb9b0ba2e8940a7aa50739fb6a5b3379a6866134c295620f42a95fa9fe2e01ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h852b7cca59a72b78eb3e33b276adad6214aeffb0acbf1bcd4a0eb833e055ff9a1c48b3f84979f215ce5b57305b2dc99a6b94526bd7f45e1a3c8cd402e1da51331cd6dff6492ed73b9a7b0f936b86f552f314ba605;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf42b094921e646236b6b0ee3f78ba2c8038f187144a9a4ea87bf354d7415cce721ae35ae3af6ad88a6a35f855e087f66d274485bbd1555b84f52a676c7d45d9b31cd4264a96acfddbca0db98580bec962135ac226;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf33276a74f4f4afd08884608c3b0d45b7b076d1216520bd81d37f2ca4bfaa62c9f4c8c2e157abe72de4662089c8316acb6369618aab0517484ff4bc51658df87495d0355553cad316a806e6bc810ad4e000e80e5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf625a9c56e79f56d76682d15aaeba0f7005b9314723447376535a4265e3fa488a04724c98da7434075c83d59e570e93401e6d3c61aa7e07710e1a89cc4352e60c6b885469fb5bad7e70033b34e6613242a415f3d0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92d7996066485c1f393700ce403dc8b893e2474562409fd2b0fff2f1bf1cd15a01f5a16e89415cda6d0fc2939651f22ac137f84125a95340b37d9d51643794f8292ec744cb125a388cbb67af78ae2273e10b06378;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdbf4e5f6b522e4c66c63efa3177ef5bcc495921c879e38d8bbb9e842a7544f36cc5764ea648007a2e62c5cc5199a987b3911dff2364c233b9fd3b769805eb2f03b7d172a011d2d4a90e164039aee1c28ca18e04d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4427a21404229e92f37270d90faca0181a096d0e7c76405e03adb6f04dc0be4e2472187d1fae173a2613daff12769e23b714de96aed72a844134233c04baed1b5eb64321dbd6c9e8df8a131abf56bb48b3bf277;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f98dbd6c79b3c351af47c30decbd92f88ace3e18de9c70f6dbb7b7fded7008049bb4339a7e69f1d5510c6f67004b1d88815186b8eced1ff05b8097f01ca3f14b994c9ae11b89ac6e7897beb1b33747cc8a2ec611;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e65ad7cece1153eabc003dc8ddc0dfb63a6370134a731108ca741ee137d4a4ca243120c6b2f03da2672ec886d58e5a2ae9d3889b2dfb22215c949cae121c6effbd4e14cb9efd42220db7a8e3ca15d46bbda5ddf4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb8f39d56618d02720f22083e9fb0d4df711a34d0c472b090cd2f4afa448e7f7b885a8769e27bb9a209e0b3ce467b296b808c49f5315a4b42516dd5b9af2adfe67b10cfbeea919ec8c465ba31de57f04c880ac766;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b8b86689e464a06382364c92d9385ef930d65fac20bc3712f1e0faf4da12b73dabfdef16da2735093337593902bb1c8ec607e04b5b61a0a345ccec5d48d94211848bcbc09e5f365344f284673deec0c64a72dd5c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c8ab314b39a972a4b55e040e9aa76527bb685285db95e90ac7b1efcf44b8db4f23bdc654b5c842f78605e5fd494c6f2a24c137c0bc360c6e8785ea92d056bbd2e497d77100e05a87d0b111f8850654a6d26ad150;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd72ba7959ae0403227cf79342f5b31297bef5d67adc9324e0631e4fa49d369327802594868ce8820c36e7a6f3af0854fffa6ce006d14b8edf98a3226da5a28d667fc457c988e2ac2f9512a63b68f77a713ffba02;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcb4ac42725a77ba98d5aea59f0defd3381685caec6eaa58d81de15c8a756c11a73437e6c2e0364f4bf4dddc9c96bb1dc45a26fdbe23282559a36efb5bae98b4161363655e5990b3e46012db4b022cd7484e5188d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h302bef001cd9c975185c81726105bed32c11fac1bb409bb6c8032ac258fc98cb943b5d0c65ff38c699efa7317a786b513dd6d68084dc688e1286d1668a2172afcbbd1aac429f9b57ff516d9b1b4a5d19684f8d099;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bfe30cabcb24e60ec8766772697db17ea98df95ae946fe4e7fea6d21db5800cf79ac5fdae00758e86df6b7c5ac438d6c08b1747ab314bffda29e4e501ea4facd2e09871b3503b35c136918a6bd0c546b101227b0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he687e7c98c88ae9bbcaa5d4b64c4c62d63af090347574814f194d3372a0bdf5acea6974b9e2cac1b3729eb58e172cfdbf1898cfcae9f9f77e2b94f6ece9c853ff4364f7da14b69f58287d69c39b12ecd067f3fe3f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h556d9265f21e3a670b2e337ff6331c4ba8a152e74487d935b880a0d56050681faff2bf1d6d626f26296c44e666dbb8051385674c4ff7f6b3fd4a471ceab24972d487f4148118e4b68cbafb913e4b36765e3a52401;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf97414ab2034250ade5348b0086c73a1b9c74ab93a4cc720fc46ac714121419cf69bce2b85145709373f6e1157d8c0e53952dbab7fab5a9a0594d9f2630f788a856614989f2ddad450ce1309a76330465ab33cae8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he935a068918e62bf891b447548a54b71ae4d95042dd8eaed1ea19cd72560b633ea7d9483b1e3da276f159079873c270e7edcf7761584d9ff299603656aa2c4089b390503b54763b552adafbad45ed304183bab19d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a5a759a04feb14fa9291db16ef8bf3353892f0ce30f3ffc1ba189164e8a932cf9689d8c08d774775cc181e5076007e29260484674e22e33d0e0a0cf56556465db10d4d5e6af7f05a1525e14ebb48bca3be3b49a5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b12abb8bda489ead57195d5eac4c00013f88f216866b891d852ee161311ccf8dc25f49489cc610e7406209b7cd838f4543ca2bc2aef2c31e7f6f2e5768f6a3f984fb76386bd0ed24f64fe8e12414f191c26144a4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2199e4301f671d18da102c2ef1e9c0f55cf60f4a85b213552a778b332e470c19d49ee6d4e3d0b4fd107616febf13c7f90fe0b205650b7706ac8f69ef2827ff1a7ac0e37a635698c91d2fcbea4e3e93e516e44c826;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d11671f122a45964632e386307a7966b1f05ab5d42259247656ad8599acf3a361453a12a040dd3bb43bb31d4cc5fcbc9c92a62cd95e3c838f9547aa06aa17921daed55a4602ad294f32a80608e5d0a9aa59b3506;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7cb789e2c6bef2ad1d2f1780a91644c5a5e4cf64ce6108d14d4617ebddaa4e44eab565169b1a76f7fa747b160755ba2c217e7bb32df1bcd2fe949ae22d239c29bd99d865f3fd33555bbd5d2cc646c085868a95e6b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3146d0f731a6d53640fa923d678442f2398167c5380bd14251ff39f718fbee9eaaff107b83be048a92536859fa5887a37bafaa02138d5b79bae02f27ecb2a4ec5ad0071eaf3ce178c1df1f1aca7a40cf16b9bae5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3ff1f14479d7557ebacb7fe55f7dda70c35e5e879bf7212fc52d31c30e411b3bd60c2c7d52a12ac436f384d2822b95b2afc5e0703c36956a6735393090383cd66e63a10fab3ad6884c58b68efe28fd7bf44bce7e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60c4f31c5538e4367a945a3f3c8beb2044ae70e90915920f4650442e94c7ae5fc2484bc0129dc5a06b915dea1fe13e407c1de56aaab262d453ff581a606db76184e769530b19a2f074b4589625b4ffccd5a6781bb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70c88533ac1eea302c1ced9fe3aa64fb89a7d7e1e45bf68c075fc624f987f5959cf2077b3d11f8b331b2f8b10ad632e0ea28e9eca897b884af2e2149a9a219f3f007cd01fada7e63d7d7edf1bc3df1b55fe0667d9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafafdee89ecd6fed8c9083ad616f2fc028c64de58bb9a48a97aecc564e70b8ca9a3d1613f9795726a6c87593f4639b5b1741ffba5682c14b1aad484034e2ac650d191fa11cf05bf2027a683c8a3cd3aac9de5dba0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac218ec0104dcf1e6fd3f6f487629d1f32951483eb7a6b7f0ca12217bb03bf5353c47ef6276509849ead6c91b241ccfef242d92b0e0f9a905b7ddb1afd08f21b924e9277485de98a40e336fa2b7e3f9ecf0894a35;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31a9f76474925f82049e9421095c467cc08355201d8b0a454579b2d6034328a45a4350c7795d63ddf2d1cb30f51695a44f44d2ab6db23384043686053b95967b3990776c44d80331c1d8ebfb1fff4c925bd2a0bec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd67e9bdb5f3b114a4e566dddf22ac24190e477e4dfffa18075bfa569e11ebd14aae1e7cbfbb5437ac8d323bf229ac27f97c194fa73633b0f399a3ca9e89f026d3861c5e04dbe58da2e742f41086cd00a4f13a758;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3be2d9391db0f6ed5ee397518f2a80a86e13827b7e6312cbfca8adef476b5db2fa62a554e2a90c2452978da7c049bc19338a70516f261b73bf9222e95fa6877cbc7aeb941dc828860edea02263f2ab75c02c83fc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52a043be21e9abbb7a535db961ade598fa5d5c2c0f70b12ca46d6168c0123f79003c4b9290df7aef6bcd8a62c3835cdc21899b0e1cc316363ec9789fbdc766c032e8f12b716a0a9d8feb3d89309c23220a6b4fcfd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f715b62e5d7e5e9b425565661f7217b76e3c691ed585e9d4921eadbcc919e3cf82cde60979a58c4cb7a0bc79ec57ab0181e3da4795dd9608e23222accfdaa9ee68438abeeabd850b58a83db1f04603be42433321;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h986608e850c8e5d7514409fd5bf4ecf03f7e2ba1154558ddaf4ff18b848277436f4e19c5a920740f469bcd190521bc8aa2a0240a68ab3658e41e4711dace67a7872b143c1e25fbb207aa7c08daa85cc3d75923074;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h981e050c0e6886bff0e8d0225fb51322380d6792616ee94fa65754dbf36fd9dedefe66953130abf0b6e327d80b79530b60ab34e3851856aa02998fdc123385a202b794db34df4bd7c2ce2cb4e8b2aed831ac5031f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b8e2b0039dee36ccb0b976bd843c9b7242408d5c3620c999da1a26825ef534050105cd79ef97bc49460ba01931e32c493f97df19c2607f7099fb82b591648782684a8963d673d33b8418faf5ab2adde28aed7123;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0e535688d0b483e82a69cbc0123a082804e607b1221b5739c735f641c585a67fd9f8940a96bd6d8a104c015dd79828b1054e43c4e5406f1eab2919c0d80e53501f88fae393161029691d1ca90edb303e6fdd032a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9aec033199814ced5bb127d47fe8ba9cbdc52acfb1d62794d8323495133828fb408006260ceb55a32b89c503b3de72232c4cf3379643752545199dce04c7c9ee17ec04678f1fd94e7c1978f198b057378738a373e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1bbea495ae0de55ab81079aa5d635f7f696478c9d95c9d6b9ace7390370a2bece13f34cf27d374bfbd509268b56c8c9a6b7e41bcee71e2b1216074655fa5fce574661f739c5cd1ee86e317a32f4caa0a338e086b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f2b63529b7990af8b7dbbbeced4e5f8fb5327f3b9225d8bfd0b991e305c711e9b8daa43c4a155385618b5222a83abb89b3eccb0444ad0b9e3683dee190692583012de42ceb2d52e09665a87ac53da16704f42362;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32d761c1e463f7f02fc0fb5c1dde62260b309bfa89c8931e1e440cb03abe1c3de3c2a515d1fb77c4b733720088e484fa2af00220bb74b7e8d71d7224df251e9a6e2faaabdf88366c9914717a1d9fa6eefd3607918;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22829eeb39c648e56ecf51da7cc035f8b522a1f4a4ca223e0825e0870588d8d7255bf28958cd10fc211bdda94672fe1cad88c71eb92453079e39d6509bfbf07b591072fba0a3383708db18a5814314387e38ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb157c54cec9a6a3b65b6f78b43c32736c22d3f5befd9343da8cdd3b6e08cd64a0fce8235e1eb812da70afb04cc219d5e2e01a02323e995cb5b35c636e9edb2d7455479b58595d52cc49fe186268989329150218ee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e623ca303e5bcaac252f66095c9d402b0b7e373dfdf395cfe56e308c7fafc40d9f737fa99f8c8f3151dac18e4362ba55c627ece984772945303ad75f61429107707f0e4356a414740b352d2a12b245bbb123826c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff8f713b455159119efacd64d181cbeea57e48bff9ac74d9ecd20b7e302a3e4c989877ba99f6d6173b56430563dd91469ee66d03c7b36aeec2367998a8f2a6c6c302a5c1f5762ace6ea16e4b5ffeac46ae12f3282;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2879277391dd38a6bd64e2e42067fbed047e021b38401f56aeebe984b9989c2db69b7e63375ed1a358342a8683f93006e12ef018b3fbb5148944af00e358f5beb4336d06314d08542f116b4538c7afcd29196d5b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24319143b8fb7995bf6b4a05fad5bb8f63a2f66db2a2b2370931d47c416f519d87b5f8d1cb719a5a26892690bef1031d60a2ceee8737ec8f59f4742b8df5b2b8d296f25908d4f44cedbc8bbe063abcd60268e3fc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca6c000557244c5e23530a54f6172244d16274aeff46200f2818260613c73ef299ec123d9c2d5d87f6ae15af538407234626d2b53b4fd287dd219ed7fc10eb416e9cd3fb1c97123c00bbfb7bd86307e5dfe9769ee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf39bfbd7be0c1e57b5bf43b2a50262ea3218a593722a5b0fe6211e43d3f959910695a3058d94e46e9f2fe828d3c4d15f7dd03c772fb98f55f65d6f974c0f656bafd993bb04e0baecfc03faa07bd44df9401e1949;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h867e3759e398e9c5497cbbb13705689a897fb09d75c7b7c9ad282bb1bc706924d8b8406f771ed44eee584699fe4f87e4b7b8478af4c539dbda3a00fef7f36e0b80a651932c743f87cfcba9adc1deaff340919401e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcaf8639dcfed6f6b661f31eb77641f2c22811f9ce810ce5b32cdab16772628e8137a543b98e367018d20c40ee6efa791929a332697b05c09481cd983f773a187b2f73b7e80122cdaf4b79e2a6148e2e0cb0b635e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha137b712b26accf7759e9b87288ef85763c3fa7cc48e2d1bb747c82b9ab7125936d9d1d54de11af21e3129cbbe12a35c7d8d41fdaf9dfdfc97bb408246f2857edc0c53f4d07a6b32e83701ba3aceca5ef9d983c5e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8995b4720b4b8e1c1e715138c1efd4045b952388ced33eb3a7e67c73b60826f4dcaf64b163e9745f2dcf4da503e4e0f7da5caeba4866b56e25147fe819e59efacf9d4e72ef5d564d8a0034b5227f7ae859083e10;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cb6890c034b26e18a32389601d77479f23b83476506ffd75e3e24e27c4fa6871c19ab866dabc172da0994856c06d27bcfffcb69b1c3a6a8ec534b8ab59ef9e5a61712171bea44fa968eeea430e7534a83dc9bf1b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51ecf10ea08dfe6198e944ad7eb9e6eb1d51ff7f6d2c1d382b36363eefbe664de1b74da93f996994bf63cfe1850046232c8393e4b029a0bff90ee24654e8004a7afbdda97371666c56a39e1ff2517b4598e57d3b0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a415ad66b1816c1f78498b9567990922e35cc8f3b5ce4da3ae44d74050096a5c24ff204f0851d48000f86cc2025b7c7a2cfb3fd376c8cb2dbdeb31b21a50e27a2d722593fd1b1d4ae831a9ac4026a0c2183f5a29;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h479e2742c2a26444d9c589124ef0aa67fd9d8b313fba6341eed7a74b591b23f408a3083f384a96038b610e69357892fb4a84f4f403771e333457f8e1f1485b04759cfbb543b5d7fe31c2f138a12838035cdbf6a38;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e5c8e8fadc4a52b2e02c85895ef51cdb025e64fe40eb1ad1f8ee8058088f8a1fbd93da9fc936421462b470e8b47eff84c652af0f324eab23c74c912c06aaa2db06031072827491c6ad7d1c6dc5aed72b50d5dea8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbcbf075c4cae9c86efb0f2fb46d1d4c76caf081da4e9af57544638beb7a19ff972bd262789606c434fe2351a8872bc6d42671b655f9e695388f65ff6b21ac86e721389d3d119eff59306080f045a46a25f54b6e8e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0eb8ff6f478001e4dbbd8d25db0a6e668d68177a0295d3103d5bacf3c9a7e7b5f1276371f8574be8f96fffac0b294f35d2364a157ff3cd9dadb219dd75dc97b7d083c39a525b712d29dccfb0b413524882812565;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha524a406fab98e566ec53ac8f40b3c8a80c7ed53aba3716a0b4c739e2831bef889b910fa428b59c688bb41f75c3b13191e47e8e6352a66cb259636461f27d29fc87de693725349664ae2eba3b9037f3878355c6e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h660d3a8aa2f9b258b78f71f4e8f2aea6a49f1840514b8363a88a2b7e07b8c964e68b9b5f6ef403947d1e5f3f88768b4e11bbfac76753d8c06bd3c4ce8b4ea3495ec6fb52cf5ad01d1ed9de487fdc2132134c1e6c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21ee7d6ab077bbd26a67267bcb78b765c9f450a9592c77f45a4b1c3d1ca0a9c29a4758ce342ec5dcc6967412a7c956548a114867860fff5760b42f42fb7e9671d50507660e4785d88c00763258335218c0ad87549;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h373ed50bbf21c334c50c65b33cc9bde0754c3ca7f4955daff976528a8e85d996b1513385008e9525de88de2e7f32a750a508f88904d2962c46df1dfbe1cbbd2ff06166dfc8378b6748f0b5f1bb6f0079edbe5030f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hae2b1d15bbcc5bc5ed42a00f0a177b9a0342ecc95bb3888f81e689f2d61f08f1acc28adc4d66be5bd891782da6732d910d9164f9f92878a568efdc89137b5f0e3456bfbfa6dad1819b6b9dbee10c2df0130c2f8bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2953e879d4dba4d9233baebfa464bcb0cde66bfddb898cc0d57644a15e4f96d73f2c361274e58c5bf769332ac569262c729da5168543a624692f131df031b6a79b01c1d1eaeb4d767b3378eb03d76954e860c4739;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e5334b09d8bc8d6c15aabc4bcf86d035abb4a087d55cf546ab8f48792bbf3c9c6804bf659887dff388a5747d80e180f52366f305be3e32cdb0abe9288d6497d75c0a545010eb3664ed1fb10cb8f853de5837b14b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h765e629a58a361fc1e62fe1d0c37649fb932c017a63c8cd33e6c1ee210d963869e9e6c1df15e0579cf763c22f62717b661d8168bcdd9a6d92ab29fa19e5bed763665c08c548a645922350e9c4a78f87bcbeb07910;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba14312b48a85c3757c628bc9a6eca1e4926c35bcb9acafa90d701b65b4c511c13289caa0c13f6fbeffb9960b3d5145a7c8fd4e4285c76648c4bf65ad0089b95a6009d2f0124f570e291c6ecf98fcebdb2e89ca3d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb59f027732e3d05a85d4fcd6c8c9bffccc068b10c0d9fdef4e7105bc7e29be4c889c2acd28ca3d1ed347113723f2fed60073544305368a1bd4450f6625838f7ad199784f22df63b73c2c374888b1b0825d45aaf92;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cfa5336a754123c183f9876197b54e547aa09cc95862a133108ac3ab61f546a9f2381c389e5b893e33e70043e3c1566501eddaf07d1d14c7c718314f05390d564db8e3957a90dc770e6c4e41e40f7c9bc973e7ff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda756ac0230022e309c7aeb202cd800355f4ba22142ddfccb39e908de78dccbb23c95da9013fe915a773a41cd73053f4438c5dae50886b5c9543752f23183ba51dc41a641ed8c2c33505ad0a85c5f44367aa7d6c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5be4d6c0b4df05a886230a6855200e440953583ba0d22644a1dba2c99b245949834639c3defd941898b83a4dd7a67381fe7c765c2b2f7041356680302981a53fd1acad14e10179299c5b4978b50f24e1ad07dd7d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4eaf760f03a02cc201d49b7e31e3243cfc73014cda7167cca50a00e0504e14c4e805357f0a5d8edd48318c2f86c4f41c20b16bc84b5afaf6d5878c8335a142f4e78b84ad99503c13e9da227b105cf8a11a1086864;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hedfb22616487ff97b865630fe505d294aff7c6d128be2eb2156fe0274cdd45b5e10f9595daedbfa2f8adb09b0a2f3529ab5e5d6a18334994217a7a17920490a4ac26417b6752843b8db32ab6be5828c39ee9f29ef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc77297d8a299271e8dd12110c3f9c082a8b004c1d73a5e3486e1c05b92195a8588e13b132dfe8e3695933c628a6dadbcb87f8ed90896067872784469c7067834662572c3347ff8735b5eb6917185d24e850e426b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h732e9d65c1367213b5e653df5e3ed5d770536db00c905f082f752f0b516e2ec09c791ac7ee4211bc79fb861a9a7dbc7ba79a2df4355483b772cf2433bb5539affcc8b6ab6ece8b03063062885cf2ddd48012d7620;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he217d655f84e5f9d77b564be8465f01bfc75f8c47f7783bb13891839142d58b778e6dbb76353b0c7c26878c380e6a14f129931c65944f8d64d297038d9913ca29c6f9717251f0c3cc41ddcae4f92550666e61570b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb2a1dfe51c67b171ced7a178a387012ac3e5dce783dfb32098b1f40726875f4051ac7be54ee19d126530095bbc8b8bb291502d8d596ace8628b4af1619f653722443c6a97bb6d3b5b96d23aacc08f49f22e9eb66;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ba4ed345bf20cf09f39db56ba8bc8efd2931dee19b7e8552a0c8d593acaeb3d7a4fde1f52a95b87a288c3367e62752c9ff60aea9cca082ed07185b27ba668fc3e205c19ba7360e2c1b2026134ce414d630594953;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h408d99448b2f768d928685e48b3a257ac88cd8d9d97f1eb7510312d0c8b9fc6acdde39ff294489b4ea09e9d039cf38abb77d3bb62a08219c3371beca4909facef65f9c45b77c4af7d69fc05267955b25433f1ad91;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ad77287029d49f8b0f60a4f4591f06b1283d99b8a2258ae0a6629d8fd4c104707aa2da477439b19e37a7fc8e4e093402cced2675b4b7a71013d796d53408970f076c0fbee1484e7129c79ea8844fcb03166577ed;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b0bcaeec37bf25c1db200a791b404003b19d278f6c5f28c716ad6307df4683de342baa447d59ef7bf55a6752ef8904dab2a556aec1c5bbf53ab746b3fd0e3f5a0f07a52a50cdd8884dbbf59aa9ace91bb422d3e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac6f7c25fdc5d7c214f1b0bea14442c30aaa10a01067fae45e49b872d858045e28b5f6092e10071cb3da249f22729b6cb2bd03ffc3d22b2f079b88d2174582c39cce29848061df8d5382e97c8f21383ea658e618a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha09487f0df50f3a268650ccafcb1256ec17d00a2ce0ba00932e1ec6729bdc7eba64d16203a854fdf80bf54d1b184dde7737d032f6c2d3adeecf209b7e4aba886b976b1001c128e73fd0cfb4528d2e4015bf42f989;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8fec5f00146ef1685f19c0b725c70621ec203bc33e102de9db8312fe1219bebcfb99198caa6a53da1dae9708345689247d93ed77c1c17f6c13e30e90b0527cacad9c79aa97c097b377520631bdd45e161658616;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf30f06565b6106af3602caed6ac0644bfe7b0ee7c335d95687832cd96ff9bb0d93b03951e54725be732f6604bc806921d775cae86883ea82caa9987b6cc62c60460d87449952a3dd1c232a28349710f52c5914f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cd21033b0968ef8fc84a8f4442b74f3972ddb392473c52fd1256dfaed749f0f2cdab267d289e5b6e6a26fb2fff00e774d8f4e98b1b6a49d180be247eb57e32a8d198b6db688e117a57410a2d472fb364d3df6ca1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f9bc4e354f9259416b6376f57bdda023ca85aebbf85f7ea243812fdc65edeb3331e1f99befb1bde46e0f371347bb0af9bdf215d4e3ce2364989a645e5759e3a6dd01a3ff69a00416d76c0d65ad4c7267f877663b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4c13ff61ba18294f15b0a3fef016fed277217abc9e8e3e47748ce7f714f94064412b5d1b0013c46bb1b108732f8da738f9e280223ce241d43e9bff2a8e25b8f91a55a281b330080a6be2901f3c23fc4560ac9e36;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h445864ff3866d1a81220d90ab8015a238dccea0f96ce63a67c01fead2f6f3c62f153d3e65dee7bc0446682bea41a3d61d709249d4b2810420ab09fa5c2e621ab0e078e066ffff510229348b18f8df0bfdd7bf320e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9cfa65382a408828b8427bfaf7624767f701268cd0eeace8ff06bb1af16b363ad1eed2770872459bebfca21a9a2d43f47dbca53ea939d34ceda58f3a292f4c8cce0639a1e5551bc44adac63f999e9d623413d47e8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a635b63e3a57c884e0c5d5c2a41b3a425de12be40be3ed091f55ec2e5787cfed2017e7279faa2bea00d2f805334d80f2805f3af5a52ab7e27c7e85eb62182912a953696cd2821535acb13a2bb54098bac6c7304c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34649a6cdcf040ff0bd4c7992c8c15b6d1f3ad6cca249216c8822929be5dc3b97ff1bfcf3ad45ef0daca1d6e76d5c98d26a98247f0298b6bec54f9e374941e09f3c167b1c8434e00d0cc927888dbc715f4472ab82;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf50b79da28c1554c15e3440d3513914dce2e6257bbae388d39da84d76e8810c9e13d5038048424d1ad690c14789ab01e782a64425982acdd2d3ac4efe1bdd559226c9c3447f44e9764d569a11a3a43d134caf82a9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc71c7c26ccde1eda0fb2c7e1d60054df548c0a1dfd78d90f7d5c6cc261168f75d51d7a449f8effaf74946102166cc8ba1b5d08f44c3f0b2a814310abdfaa21f5367111bbfa74a82ae929e7893eb715b326dccb62e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32aac6e49ebcd8fb4f512a813deaf9c8941e116436e3b2ca78d27d37cff5b3e87d5cc59d36e49b113dc7d7a20fafd9e0a4c5a90fb38fb7b58f8c61661c2c024f103bbe1701ea9c6aa33af606fb3a23f6a6263e09;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdc2bef26b5cd8039bbd0b4580119bdb4adb516c720b80de618dd5f28de8e8fbfceb3a07ee20be9d465e91e0e84525acb5e93d4d879cd3e96bb4eb34e1564467f0d9d247c76cbe03973c46017ffa53dfc662c11e3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf06cf4c4d7ec77cbf63d4b0ef55b63d574b6c9f244d734720b9de5943018edc809f64ce382d0bc8a141d520b1b813948bc557fecf56209b75460eef044f329878bf191adaabeb7c35fb21133b219912cf6eb1617c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f9b96dc3e2363a46d9a750dee23c04d2361b3ae98072331e493444f1569ac0ec16d8b5bee5d25c1cb4d3c20a8fc21c905b9328ac0eda524569857c4ea93fa66016a90d3b0131d6c481656a4ffa8cf3da4f17639d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfeb95157186e693a91fdd8e9057696f085c8fc0f8ca021300a2f3a1a28cff3a5b30f669e14fa9ef0fe3e0fb3322011d94a02d4af6b04459fe01a2f7fbf63646f083d59e069e67df4d5941d691657a86986c370883;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cfce93ea89106a8d0e158f3b5db8c36ecadd526653c04e9727ed8396bd4e573766c45ac5551356e652b4f278e50b4ff8839671a00b2a83e336d0864e7f13b26cd2ca905c912c0527fa2015200291cb29305824ee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e1551209cadbf83f6e333e4ccbbbbdb9610dbe8b192e1a61f1bc7b272b154a5ca2187db56f6d43ee7ebb36d69f517c9cb03c883d17f0f1a0604581d998a063f03e3942f09f989fc8a1a739684411f6c6541f6e95;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f08d9f19e5f3ea9f7b5b50986190e4bac094cbf061fd00f703c81c03f55a20f0fd62e6d700d07936363a2aad7aaee1e69ec7e58fcd89f0194195ac2b503ebc5a5e093f93251acc71f4ff253ed7cfee86991fbbee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7decbde9504e7c649932a82a61f625aae4bc0c5db734fc286ddda2e8eba5c75843c30b1522b64c5d785313032193ba8ce4c35bfee37ffd834146178ef9c9c1b690f64437df0169f345042f6e074a6fb4dd9b90f0b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3c9a5191590183dc0695ad9665603b78b6d7b5e7706ab5ac7677e8b4c1a107db3c06d01721db7e7e766c16c76509e82164ba1c1a2e9ca0c0b294289f9db2d062ea24a0d252a53b4a4bb12446d2e5f30f41daba96;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h510c37dd995a729c98965580bb4277e1fb469a39929c970251998ad36b6493ae8d5c64d478629a7f1ecb2a38228bfa5f317dbc72cc06ee60f5225711b26648ff422685caf8818c1fcaa859bc8a3055e8d445a142a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b43c8efed23f0543a5e2173e5806636ba734fc9047ddab6675af8433aa767887d3902b582b2bc553bb63b789f5d034084fcf92030d5599536d5d784a35048972a74fd1025732de65f74ba6221a6888539ce21724;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f650762f117bc3b237fb61980efe169150ea88c357cf9b7f3cfd00ba412fcd50edf1a2bb56d48bc90f937e2efd8f1e48a8e4f15e5d71a1ca684d2c29265b673e261f3f07843e997df9eb9f932e2be3519a1f2e05;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fcdcddd43b4e9420e5ea78b0560c3522d08a5ae7330b2c0b677b49acbd637d543dd504e8e2c8194dab3336d610b9684c80f96f595c957c8e4d60fdd6804a31b2153019ab4e3cf4491606b9c27c8b68433e4948ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc8247a134d391d83137e07d2b064305aaec1734945354753b1adb82df9d19bf515b9fbbc2c93c26befe21ea49a6ffc1dead7d01aeaf3f66dcfab7daf78db1a33d67d6cfddb54a8e1c74f7ff04e5b5498b108c06e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94bbfedfc19fa2cdf7a49fdab939f3cc13f2a8eb6935306ab8e1cdc6fe58477b7613a78ab8ae4eeead07392e220384bda5f4d4786955b5c54c5b319cb2c739609b34af458c41fd68b4ce1396f9375e1b918a61fe3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49fd69c019d1c9071ea2bf1a9c40a31ad57df8cbbf24e85192dccfc6fc8bc3d9b8ec669e5fe2987d5911ab5a05ca7f33954bda39a455172c921e294fa49d895082221a9b1ce4eaeb9abdea10b5740d5cde56b185b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha46cba5306c6e4f9d387431574f612214d0ea9228bc29bbd4cde66a1a8366ee81b46a83add6e9be017e8393b45cecb9221f7421ccb22ca0dfe70c1976fea35140b4853e98e1f92552d4bab577597f78582591077f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6502145227b6e8415ce6ebca7574f57ef81eb97c3aaa447de32836ccb86b50c23fcdf388af3ef8fd7acf2bac95e3f46adb51220881d4bcfc757c60614f0959ab772259d03a5165b4a9288df791420635c562f2864;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17632f756fae5cd4c03ca98b27737a6c6818a9e12cc373dc1a501ea252014490f719802d6e89eccdb3f27689b41350793ebaaa9a69847e692c33405396c21449eddcbc0814f9eb7b0811d30e5c0f3882797519739;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60a5c7b2e866f21a840dd307f816dfa6acb368acec3412504eb1a31941d8f4f2c0749687ca0b044c43673b315daf8e1cc91de0fc85f1525bddbf52cc744d231112a1bf286ccf1096e6d934b1103334d55d784e15f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he854bdbc3f8dd0650cac6c6240d84c917edfed500be91121d9de4bedf16ac4d6cad94468270d4b301dc0ac99e07ad10666b1a2c82a1c1a1647cf124ae51ef470823f36f34c43202f0f0e9c6e4b9fae15972c5e248;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4075738e5cf5295139ccfcaf6e822bad491d570127636adfc5ce4760850226bacd442e3e54667c4a6fc91bb26d7a9a1f96ac3bf6b54ca39a7ab16425768e6b736c1edd8fa940b17824c8dd2425363c4314cb06fa3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6bea4894d08a5313f0ebd2b80af85875a47a8579d7503d83105a9687da960d26f3344ff699f543ee75b8bd4d4b845c895b1b10f2857f96e4ee41f33e66f8d16297355697042a26a8e19150eeee2df2b6865b189b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf18df2362445594d89898a32786caf5c3b151a9bb03b26b9804c374a736b8dd353e19eebb7f1f74122245fbbb48677f0c38c229ae4877d95d1e7876a1cb40639811af09493cd927bd62778b9c21a1f6bf8090baa8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6bceb6c4411ac2b401a69dad219a504eca4f59c0db98368c1815a5b967bd52801a52a0caa4cf2e395924958f1caf857a1076013e5b8660623970712d6c0c47a05810451e16b0cb53e8301f7e6f8a625abe2d59824;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3dc0faf641640c16b9c38b2ee292fac49cc64a402821530161ec79fddf29b2abc97bf6f36b343d40f0e310757319d23a601df8728bf21b1871444dbd8ae92cd4a6847404032e31225cf1403c5cf46ecce50b6a2c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd294bba444fb0814de2dac9791a2d0fd0ac48ff5e2226e207c6ee92b664f62e013dab0ee85754c81cc657ada2d41a5c755a1841b2645119e5eb71ca0c376beb23c750b95686b7ade9658ecad10b5f9add0cf6e905;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7aa75f0f89e6384beb5ae6edc8d8b2ed06e4a3248ba2d27ad0e73b071c5ff41a31dd58d4ca8ebbf9a3fb502119055ce68f2f2397e9f9596cdcdd51fc92bf91fa1493c0b09a3fd70f6f8f88a6c74e3effbf89e12ef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b51b18ce5059b97f984a1150b3ca8daa20346278f8b203525a6eb7d3b8959639f77a0e7dca9f9795fafada6839109a7b0ba8db74fa62e2847c912c14b6ef4d2070fa878365aa09297bebe2d3e694414512de2267;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93a5536f85dd00a682cc54b6942720679b4caa0abc0736950be2df1369348da2282122ec904811d906b8e6a7951778fa4ad00cce7b290fa74a8b5b7ff14e24351a9bc43b147dbb506bbaafc8cfc9f2233b4bc90b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44a15d0f54a3dda80ce9cdfd2cba92f3f4ac1fe065869aceeef080c83dddd0e9292590b5da65fbd394ac87db66dc7fdd27db58f413339ea27c1e1490dbdbd068ba1e19d9687be9407a4853f85b3847a49076bc711;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb816f24781c36155ce1a96cecd691abcf5e8fb939206645706b0d018f82cbe3eb32f05a65f8a788420a1ed439659df74483f546f9a17b2e6d8437f3b583e69ee5c10aa89f0e981b7bf751b97f0569990bdfc6f07a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4ae70159d0f3692af7772898b86354ceac108485f6bb6fc8cc26c8f5da01f40c8d6d9653a8361adf50b5a56bf47995ff483a99688fb47493df2ca4ce5756ac6af2721874f519ae2b1d2cec282afb3d4e42557c92;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8401f1919f8614c81028ffb4a6dda569e1d33da4743dcca8ee6a6a896015884ca7115a9e20f89217bfb1724abfc424e059aee3092a16a25193cba3f40f70801c0dd8d6296e8efbc3792a808a21d087957bfcd0a91;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70c0ce32cc783bd3ae7079ca5136a4e8435454a5e343633f3e782dee99fd45b64bbff41b78bb6ec29942e0b4118e951f74ab5e923f02471d17ac1966ce9fb5f052d2545f5f4206eda338b68cc9d7aa7cc83049774;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5784e5e22289432bd6fcfd5dcd9063216dde852fe7ddb828397da9407870f926c6f68f718ae8cc8a5bca3f9bdbdbc4fa24edff14724da7eacba090bc773c29f6dfec5864dd6db85e39bc88662f535478ae7c13562;
        #1
        $finish();
    end
endmodule
