module testbench();
    reg [7:0] src0;
    reg [7:0] src1;
    reg [7:0] src2;
    reg [7:0] src3;
    reg [7:0] src4;
    reg [7:0] src5;
    reg [7:0] src6;
    reg [7:0] src7;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [10:0] srcsum;
    wire [10:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffffffffffffffff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16ad399df3f6dd4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e3432dea5785a67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35f0ee444e075d00;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h794988d466e6b921;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacbc283276580d45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f450bc044936682;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15d39c0bacd9ec5b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haffcb1d4f1bf9f13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7131a939eaada8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9d77c9a81ce14b5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42e8a56f883d501f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h210178f4dcbf8540;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e9beeab00f6bd20;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9c2ad73bca97d51;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9235151316f0a910;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8a53639106233f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4d61de16cfc0bcb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb210f203460f685;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7263592f34cccd33;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f0da8102b1af207;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf152544b4385d3a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9132d824a249cc8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8332cb54eb7c4ef7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3bae91f2f80a94c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8aa8949d37ab348e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e8067c965b1cd8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45bfda3a5af2505d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3d750e8e1ed9bdc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3584813dce5983f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h459f4b91535f103b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h679102fd1845b3d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf412980f4378580c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a72799bbdb1ed24;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1cf4fdbce849859a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5cd8d57808303f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99b607ad07fa6859;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32c2f09a1e970633;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8dce9000c97cef1f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f6fecf270b16ff9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8471f00767e77721;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3655e6d9187d6c12;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2b287aac9d2e6a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ca2dd0c5afc3f08;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9951d30ff95d87eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d5bcd5af690f721;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70163a195607cb0c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0baf7b571886f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2cdbaf046f24ad6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2850f52e9ef3aedd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h411847ee3d355bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h229147f516ec0bc9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he77293901d67f402;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b3e7ab0ce46cb8d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfcb62ede1425f99e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd947c6ae690ed420;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7061c430d822ed5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcea3b6c5a30655b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb807234e2d7c116b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1aa2401c149d0ef4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61bf95111253ee76;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h368318fad3cc32ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31bc2c4947893dd8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24a34f410c7bc2be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee94476d2cff3656;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48e5ce3adb3a1500;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a04e6198f835718;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c4577eb94876f77;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80218719516500e2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf1a329a72305de8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab5a607f11d7f8fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a13559a81241c05;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c50b01a32d6b97;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedfb74d4b334381;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha81898ac404e753b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h103ec8510810c32c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94adb062029e398c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e28917f15619e8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f22b135ef89d491;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35d6b1c6142c0c81;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a4eb6fbecfa6f70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hccb27fd9e25d9ea5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h566aadee7a513a2a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h458c7378d69770c7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h967d550d75bfbfcb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7219e7ff504e11f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h492a45f9209c6095;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ecdadd3fe9f373f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he933184e9b822f58;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26058206cb3ef992;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h684bf0b544e92204;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e350c505bfb4a88;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha19c0131698f13e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff9a57a3e7dc00d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5db0d47cfe9d98e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h134a788a9c4c3037;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4962024052c828c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5164fc3393c044d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b67cc8a2a60c83d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd50ecbff8b332ca9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfef55f7323d3c403;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9051d96085fa9ed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64024c9887674c64;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36d27c53e97a0dd5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c6a0cda2d2215a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he77d052dc39c6c17;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4fb04eb16b474af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7dddb498f2c23138;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c4abb61e5d00453;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he04f08ff7fd69485;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16355a29c13bab10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4d1b314b475fb72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2df5ccc9936a50d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73d9996413b46e8c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h744a2da2601abfc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha11fad334721cfcf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b6faa33b2648918;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4d7946e74b65606;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ca0a62e76ea25e7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h705ff0580318857f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0cc83f2eebe1e7a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6bef817daa765003;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6085420c49471bbf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44471f5f8d7c97d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24782ce4c12e1648;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54fa45f5b95ce564;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5ad966db6a52709;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e11f57d505d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86d9fc3123793309;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2eb4ca34bbc44fc7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe89fc861e27c7b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a661dd4ba7a2620;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b8dc0a38242a08a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b1b50c29e542c67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8919b7c25e680fca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4ac9c900c2af0a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb7924f42c2509cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ed95a898c2ce8dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e7c1aa524f2786d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadd2865e4d3afffc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c010d9a003a3400;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha439a5fa0236312d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32fe1f78e37249c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a7cc643d0487853;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h835f1b1e98231937;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf16cb1f262b2144b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea39dd88df322e57;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefdbaa1eda28dc00;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdecd9b678591bfac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf85b65c477e00d54;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h966789b49b2dd697;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0464e9cc5dddb34;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habf306083139c65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b85e3ad0db8f84b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5e352b82c24f00b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd698ffbdea543be2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3079a2af7562ccc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77c49785fbc74d65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fe8611c0b819a0a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f5cfe641435e117;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0f3949a2e8199e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf1d9ef663e83fcc4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heca7a299ae3398b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc17755ef4ec39a75;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50a1ae1ef0430d1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8fe3884132f9dbef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ff915615bab9da2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c698c4eb556a2ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h400fa4388a551bb2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h639c3ce28f2fc4b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c4000aa4ebc07dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8845408179fcfae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h899e0987fffb61d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd957bb7a99d07b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a1c28c37ef30721;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd730729e9cd42497;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3fcc2d692c1cdc90;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a22f2bf8bbabdb7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32294a2fb6224539;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb4cd9e09451a784;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hccc1baff95540296;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa60580aea2f93c7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67acb35251a68c6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefab9f76523154f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb44b30f849538b5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he11f056a131ce142;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1da42a5301e0b5b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7cc9317ad03e239d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1da90734ede3eb6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30a66ce828496236;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c2643b82501dc33;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4c776a297d77cbb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6bffbedd80bdf4cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6cb309337514a01;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h782097d6a3ea9787;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba968718af8e6b0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6334a8129e96a28a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce53fc09e047dc4a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d3c9b2fa7528a6c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b1d8ef03171c4a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d3d5c6aec81a201;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9344ee20c0e7bffd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc21cd5fb9a08338d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8464088285cc176d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1fcca9493f734e3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10e3ecd0c5fd0ea4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22999488cbda1a64;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h244c066970ba6ab2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde6c02f9a66561c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha83e0bdfb5cec276;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff15802295f4ebd6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2345ca00887a7c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2f5e1c945603204;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf80ac5296ab131b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb2dcbf0b19aaf9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c99dd6d927f9823;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h858558c53f271439;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1726efadfced860d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e0fd66c8f6f5d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc62b8dec15671859;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h409332b283fa36e3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef6d5da716369c4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha75bee6957714a48;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7a6a8ba0d98023b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5df4ec4cbb353cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33d2712139e835ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27607f6cfb595565;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79d51b8b692c54cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6631ce2ec998560;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1dcad1e86bfa564;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb3cc5d9e974667;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h766e1facf95c6e48;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a3b92c271ea5332;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h579c2528c1d791c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1cfcc6e1affd8846;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fd5a3ebeaed5ff7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc896e02c3dabd37;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h250213054154d8d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0611a19582bf20b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h387b8f2c8496e91c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52e51e45b2609439;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc45b9e49d18c11be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f49881c0736c726;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5396e642b319a3c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb72dd78726b2bbdd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b664b5dc0d8d1c7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heabe0bf88f079e11;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd030d4bd9a437c54;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7c0ecc8f89205e7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h473d129f511eda9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h789a8084a835c34a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1293f9ab5cea169;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88a6b8d1bafd30e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h286d4681746e8460;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he1e1d7975f72880c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h158c9e40c7e083ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46fa2a258db4e659;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9bea763bd39ef35;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d8e23860b3d1e2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c13f62b99a0dff2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha66c4b42544732a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14dc1ae9fc73a290;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d21cac90ecc1f2f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58975d60a539fcec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haee2f2e65f622f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc034a13a83745c67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5070b31aafc9d8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8641f47094982d14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h343771a7c67db053;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5e265b4bc86dee7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5fd48a5b8a77f77;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee1d10a45c95efb3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe212f4fc8e13578;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h491fb3136b07dac3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70adf2e30758966a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36cd1d97d0d4b147;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc406987185108be7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2385af0064b5e81;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3648982b8d8287bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h521a8bae10e9643a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h146516847c30fe6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c8316c0b20d0de2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9d8693b16ae261e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f646f83115e9243;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5cb00a425bf1a233;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba0833f7ee7ca89b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb45b5c4d9c3be560;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd026a9ce3e70099a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49113da5f349053e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7159879c62b8c5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89ceedd96ec961c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d34c241e3127b38;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefcaad0478435233;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e3cff8ea895b80;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14eb12ee914ac717;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6faa89e0de18f092;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf2470ee4366d149;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8995ef0473a042c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e2d66885eb47f9d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h726349f5a4bff7d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h392aee4ef0e72076;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb3c661c19632aff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4e8364808b76b17;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf22b53b17d622e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9424da5fe63fb621;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ff99ca6171ce765;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7c639be4d107f71;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88100c55d8a3457a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hada56942320a98c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd245f556ba63f8e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d36889b79cf8695;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8ddade4643c3110;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h338cd678ea3dbaf6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6451cf2e0c28d0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbc17e6847cd9531;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93c7abd6c8f2e595;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4135795a9ea7cc2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc18e0f68c7baecc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ac4d4b88617815c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d96212c066c4b2d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62b66d432433f420;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf604fed87a8ae0b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf00afa74eb784c2a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ff9d4aafa7565a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5ad6ca1cd49cce8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d317bf85a5c5b53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57cf94c3146412df;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6541c3764d2358fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd1930973f5db242;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84f2e34cca940de2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ffd4f4771f9d996;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a95d3b3b2d08620;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b911ae5d4bc675e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38f98a4d30596d22;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9248aa406359c9fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a93ff1b578d263;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5d3fb5ecd00013c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51311c941cd0f850;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9bc735a5410b061b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79b007f59bed3155;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9963f289baea23a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c40f2f19b5a7ad2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74b8f55c55537471;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0759932f510058c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe11b731b637a0c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc409fe1c818a1091;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71053605fc0b71f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5d4cae5dfe05ac3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94d2fe671c794cb2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc95b232618fab43c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e3c8c11a92331f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h638cc35b2bcccf74;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha42056aa9bde5699;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95f16a0d1dbb6e10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4409c1b3d23ba79;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b5ca5f28c2d527;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9dc91e706f99ec28;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62ee7fe262146df2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1eade93b0f48de5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde9fb2dbfb8bb5f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4399309c7aa7be7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d627ab17fecf5d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8472366c80ecea5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdef63b750aa6efdd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1158418bd38f586;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5adfe9e61ed1a40;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf799bd84df6585c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd354c2818232cd2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc51d65093004204b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6393a65306013ac6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb232ccf0b66f0b53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he416cfe60368e09f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51e2f23f443606e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h963704cb1a48d825;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6193da4c1bdae7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4634211ce1b66571;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77fb23bd8e03a29;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84d51315b83bcdb7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b16b88f72ea312b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91138ba8f4cdd063;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65b81f400602c350;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79b418bdb7393abf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe54db5780d87b2a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had23ad742493dd14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8aa3f81f605fcfc9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ccb874a0be26208;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he066400834f3559d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadb402bf3dd30e59;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3bf9a42b333d45ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e57008be179489d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb362ce963a65563;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93750bc404461e00;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5652d5ae7786eab9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdee95a9c80e41574;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88d4020ad5480133;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd6141c3c5e5f324;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64ce095913a3a2ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha87270ef67912d66;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14ac7603f5d2f575;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e9002b34de10c25;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b2d8a21c85147cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h496c4178864bae5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47d17bb62428fc65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd22521801b8b880;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37ad0c6f6539d7de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha95f8e3dc6d88243;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe452391c5eecec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha900817124f6912f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d1e7fe56ba39f5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24ecb65da0cb89c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he856d2bfc8a1c4b1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa7211d8bbe264d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h332a99b2a9fd9bf0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbad3efbf8c70f0ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfea76c5c9b34684d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d21137ec872982;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcd32a7aed36143f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2f90aa812927c61;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2970d0d9c3c129cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c4d100157b16908;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he921fcbf69688441;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9c00243f4eb62cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf87e227ffea21a10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b673d9fd0ad73fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5cea86fd5d280029;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12926269d2e33fe9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a3726fb8461e5cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h124ddbae641e1ba9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77e2b96be30707d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h297aae2354c0cf6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22fea2c4cc872250;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3a003bd0dd13571;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he24494f830467942;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he38cff951402f147;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd5cefb72b7176fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3886ea958a9bfbc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3976b1a7c4673d32;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3839dba1fa7e460;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1786a7b125e694c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he46e4a1123901626;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde2fccac5bb79467;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h233adb47cf7dd7a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc6ef4eaad38225f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he566cfbc6d44db82;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9cc63def298b56ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65de6f33d46160b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79d635c4e35ba47f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72e581dd1a65eee8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ae5fe228714ab7e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5edaf931e7c6e4e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0935169d0bf9c78;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90d017f7c8675eb3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0fb883f6780a663;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h369ab69b7fab426a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c4c36b39cc8d99c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hccdbf0ecebd643ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4ba02cc5d901ccc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb951aa6a0971e0fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a82245e09f5e286;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb53c7f2a006d3927;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e60f6f190e305b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2433c3a59aa6cc44;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d47063e8687be04;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habcb05d6f8a9fda5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19dddde0b24d345;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68b1dd3024e3910d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd125053125bd2a5a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h161e6fde0155961f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h205131047c99c269;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15e682a45974d37d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57ba70286fa04d65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7867b318d662a182;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc45edce72974f09a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he89c809eb2cc39d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddbcd03874b3ac8d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44e41ab9002c8af1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4acdc7bd7312ae4c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32702e9a6cc20504;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4010993c47c7e542;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf58ba2a310e1b400;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha96fe882af83cfc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d6efbbee616d2c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heccd5aa98cf710af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h337c1ac1b970f850;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf27d42007a30d4e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0687c017ad0da82;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfdf2bb0e5227e7bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h101731c5b4a76868;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4f45c6b006f9c9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44e838c93fe317e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb74a7fdfea508d01;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcac15013cd80622e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha75fce8b5c916d2a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef28f32de61adc76;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6fe527e507daf22;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hceaaf0b01f886996;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha58d746f2d437710;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had8eff19016f50a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f05da68884f9a7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d47898bd0044227;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46a732f1be43b393;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd020f1fa469e2b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89289faac670bd35;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7177c88cdf802d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h560213221109cd88;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85ad96d707461797;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63fe2a63077b8d9a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f5309cc723c4bdc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cae482321d608d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb6fa0722ac83972;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h492679c09e1fb04c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70a25fe4c455ca9b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65c318c09d9acabf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha553806a7366b3c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa955ae80c7d73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he76c8aada8e7f691;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ecd8a7a37c79ce3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b1315389f649ccc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71f89007d093b3d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf1e7ff30b71849c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66a1bcd91b415d38;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he39519f1038ce35a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd893be706d37099f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc823b20e0c208d5c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92a06a99ff96ae45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7089b35c63889c46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc18120c0a68ba5d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h205f901f791c41af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb80b233b7715f41d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7489331d805c05f1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f501653e8b328a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2e6c9f436aa0776;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f1061c13598a91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc34e9eacb81eaa25;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a4936c6d918183b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee24833268a9c29f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f109897d010b714;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a398ee1f71afb0c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb09c6d15bf2fa279;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a419f3b83ff4dbf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8b7d955092f67a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h833d9e2b547eba24;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2021dc4d0e804efc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ec3d8fd6e565e7c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7471bec08fe6783f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h681203f43352e906;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd861501f2c301055;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf5b02ee8a4003bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10f6925bc0e64e84;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51c3a9feaefd7057;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb046f8bd2bb8ce78;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd968a2ae176abed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23364a3df142846;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f59226258d553af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79403add9cb0bf12;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12dcbb21e24aa1e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4714b71f3b6e461e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d13ceda1ca7f56e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31751bd5b0e0e8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcd7c874b0b8f7f1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f784bbbc82717b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7ff2a1dcd6efb51;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfdad560b64a8519e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92fe4fdb23475b2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h194343ebb66a6cb9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c3500ac5bfc12ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf2accc12e77f525;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c8277760af6af02;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46f735a180f78981;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9bed6a6a7cf251;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d54e306d056e9bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'head11f081f36bc69;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h435e2c0d55b278f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6c041797bc6ec23;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5831807b3eedf7f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h187a5cb4eee200b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h309b929a25890c92;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55a399ddb1be8419;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5765d29977177b5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e2544f4f2659a04;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91c2af127dcc0973;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he19cf5083ce28253;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b9a1b91ae349dab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h399b7fee67c3e1d9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47611423eeee0c4c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd52778aeaf23f026;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h105529d58fa9ee22;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h192cecc9b47f92e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3eaeaeb5f931b96;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he052defd813806a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcd01050c178e9e25;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5052e377749c7733;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9865af82522dbe7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hccf499e820930953;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36689a53dc8096f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d9c0b6dbca63a26;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1999a883eb766c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ee5b1125ca0b616;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31f7b8ae1bc5fa6a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h226492a226ff4979;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae820c696a4e6fc4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha542f83d1e74d772;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h82aff65ae8246580;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8bbf3735f7a9c855;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25d366aa2d0b7eae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc00b9f24c0dd875c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1624528ed0397ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he21c05a65da104bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55345b2d48fd032b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48886464e900a184;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdf01273d9eff9aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc25d7334146370e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd6ddc66fa0729cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc7305ad6a0449e2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5d825ef4330067e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8962eb516fcce194;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d2e1514aace9ae8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94fb3368504e86da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef7f68c9096faeef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd19a1645746cee8e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb623b6921b7427a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he48fc6f1bf843d9c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86ca7750b95a851;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb1f8addd391484f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48d198846d8f392f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40f8b7409cf19e8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbbe953bff0d2f43;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc017fc7d011bbd59;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7cfcd589fd43f413;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49de2088d563e066;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he21c67f7d9451813;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cc84a3602248fdb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha98db2b77d3fe89;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he13a707d1d320549;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h910dbe06056e272;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7115125c04315ce9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e1faf044966b83f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6be2a60477ec3fef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62121bac1c527ef1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b44d5c3c5c21622;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h530ad61dd01d7e2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5efd374a652decd3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha45ad811dcadf356;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h176e8f6e39592d7e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b6fea62c81a0bc8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had6ee417541c5020;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h724dfb50919c6334;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9ab87b37040296e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ec06f7da98153f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea6a16fe1c9cae6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72de229fb209bdd2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85d6a6eafadc5a3a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b7d91cae47b6638;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd80577d2cd43478f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1284da4b6667c863;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd840cf190f57de72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc9d4bae1e7dc0e2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fdfac5095fec050;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4042c83eafb6e816;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3274c6906a6f76fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c066c47a913718e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9507f0d5fbfeaf53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b943ef4a649aa68;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24d312821c446850;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f4b62456e37ea95;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf35e8f4459307739;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8dd23114e5cc524b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2b2860704c8b07e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h987b58c57d61c535;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3bf69a4e5405c3a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a8118a0f52ba10f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h234174c3273e2da2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0df0d7841bdb61a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55b5a1d3d1ed2d06;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1a90b1a06b4a178;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62ee864add039c8c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6bc1ba008ff990d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha16df468eeea0e6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90b92b6be0fc8d29;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3b9b351c4b13277;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0f37e22bb147f3e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ff84a6fa5d0bb4c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde7c77c1c7468485;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98469ffc40611d46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcaf8dbd61ae9d303;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he1e0c4f7977502ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb40a742493eea8e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbac2abd5de86e74;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4cfef6f748933a2f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2987e62f5841e9ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6ef63f414ae46b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae5e0485bc1177ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadc908d51ca461e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69806bef63f63ac9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2dbe71527abc8fe9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f7e43eb9c18b62b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6581f71a587eaba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5e4223c4ee51e85;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65a8d1562272a04c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefa1e831485bdd40;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99612eb1e02aa112;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h962c873382133450;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd653a7730bb0d74f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdfc0bd0ea152f845;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96cbd1500f2fc853;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5a0a7cd5a4f625d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf05f363395af316;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf89b6724091e55b9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h315b752a4feb836e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66d79131b367fe05;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0a5160dd43c8766;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26bca557ef58bb32;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6701553e6a51c8c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f2dc00b71fd9272;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b6f24252370b2cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3a361873bde927e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23b02cb5314463f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc09de141eca9844;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb86c5ad82c667895;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h160098bcc146b540;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d6f0c1d8fa35662;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33aa9186ddb41494;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7de043b0642cf43f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39ed1a8e05615bef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8db4f2f192481b79;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4ae0dd8d19f82d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h733d107b26fd6152;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3374c81bf573ca27;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b49eb05343c94ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcec041e427f2e957;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ab57d5fabff3c09;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81669e5e23d92e30;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24cc2427c66c5df7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b473ad9c1544e9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4462c734c89c1e89;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8381b4a6d629449;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f746f9d773c8b6a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h82c74ba316908f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dc095cd96d1803a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee881782891a3ac7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3b2bc75be49dbbf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85b3e1df06270926;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h509a24e0b83b5db5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51c76b5563e44367;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6def39411e9dfed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5858f2d4e6e8a0db;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a5905ae7f3d509c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8df67ce2b3b9e359;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d49af12ca51d34b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a1765cd9030e760;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46cf2ed173d619cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8240718b13f329e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h786cdb159372b0a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h714e01eaf5e7f88b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbef24d8a9ca379f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8627294ec7e8610c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha176a2d45acda3d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae37aa65762441a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf303e7a4f5ebd7f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h507c5bf166daadb4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc281dbad61e3b9d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdfa8fba91cb179c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab89b2ed5e48468;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6325e4d0da22f8c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25cac75ad96e2b73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he71748a9e4b7dfad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45cfc865298cd591;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2981edbcb9d62ba2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2d4d27b39cb89a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70d71699816ec9a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d28ac717c837b61;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfdbaf84e52b910ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h232199f55d77ab2e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51a5ce6c1cbce152;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e14c4c0cfdfd111;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6780cba58461fb5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha47404d32df7087b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h849948b46cf55ecd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h635f0cf0c151f97c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78386d2e536e8621;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22318bdcb2eb53fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80e8beb947575d29;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3fe540691030c10e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74b57c174fa6a11b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdebcbda61d937a2b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98323f9cfbfdc594;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4828139ff1b6fc0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde09cd0546fe4416;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31147369e10f9fba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7f29997a1d1ad88;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h722f8336c4a802aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedbdbf1e71a458c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h847978b1ae2c80a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habc7dd485fdbffd7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he53cbdbf8cd6ac0a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h540ea575f9a99206;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e0666850f043a89;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf672be387632a29b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5e7fd30aa60208;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96ab31fc8ce7ba88;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had873fd0b9725f85;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h226a2a088230c3b1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea6dbe7207b070b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfde58ca5f9cb1e27;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3bdc221c72611405;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb3fde94e4d10ec0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ebe32ca15821fce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29218f536ee5d742;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h60c2fc6d35a25b73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36930406d9b832d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee1c232bb0c40b4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc216575baacfc38f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he20831b3241f0cd6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5948d1c9bef92135;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae3d2e4bbe6d2dfd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hceabd87e866d3f4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3df13507ad133681;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd67a8d2febc2c970;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77bfe399cdd647f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b0820621bdd84a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ae53fa14c312c85;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5dcee38c1f27988;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h582114be20e1d294;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h75584a059b202a39;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbdf48b61714272c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf41d8b6392b6152;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9107b1456fe4985;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h575954d4549951cc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf68c2e3214812a1e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55c181908f64db5b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52a9281725382f69;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h440dbbfd9868545c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h304e765cb1fd7089;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15d21a840e9d2c0d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb27f20a53e4a89e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31bf8efddaa1cce8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f18f1afab5e91fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8da7485dbfa848fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8281f7de9177ba52;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbeafdb02f2f6274e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h551f99abd7be4b48;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ba2b69544e36c51;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87e7f855a6e1314f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22531745b2ebd38a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37a064aecaac0d1a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6140d9b6a8a15b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f6c3a93ab3c4479;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f66256fcbe21dea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdea00a41a63dbdf6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77f8ea198aadd33a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85f15719446aad36;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72309e173c62cf29;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f8259f2d8ddabe4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d1c4c532ccdea2b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92321fa435e4b7e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb34fefe1ab8ea4de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h298d8121241feb31;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hccea0713847b4344;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9ccf216d9658fa8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42a8c9329f78d85e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h702e9807d56d3518;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81e4b681bff74a34;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9280b1c169a1a394;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2260b4155c2a38b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h228b830bddbc5788;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68137485a8f5d5db;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc88d3e85827d83fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha5c879924e0527b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd868dcca5681a19;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f224d7cf4719d3a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e86390342a39968;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76516545a58a9a52;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3825c1ae53dcbb4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30c9f3de89a600f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habfa3ec1fdd2bd1b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef93e1717756baa3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b79e9ccf4c46bbc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9e029c8ba693303;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38218a12adab2c5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c1da8e5776932e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h359e957767062d07;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf177a56338d34230;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7377d6baa3657889;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c0a28eca0eb57fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23b4cd910dee0228;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16052409cfe0240e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h118b26219bd60b19;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c5377a3275450ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e6aed2732c37d30;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c444288991a7567;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h109b885edc330dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ea6c488c5a63775;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c8e7ef3b79a83e7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc90d1ea7e347191;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfe89e846e01f3a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc04fdc40706bd3da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h720a8d97a29e95fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5baf375154a19a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h958199228e09324b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fd9eb86f1da4e59;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ba021487b6f4521;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28f2757d6516b3c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d656868e5cf555f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5aebe922fe6bc72f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a75c52ec7d0d9d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf27c62e28765ff5f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc99498beff3a23a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3f644f11aea923a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec00816431bae0d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0221a6aa2d3bf80;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dcc979b3063c767;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b95fea3bd4a1dc6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdffa8fe93cf95a14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba95d7abc045c91f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d1b5cf06eb40d4b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1ed06f81e92d3a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc8fcd839f19639c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha66154361055236a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc5c3ed218101947;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ac27f8214e486a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c322f7539e509fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h104a3e71690be210;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b5f1f0e09018436;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72a1e3897b5888a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d6c2d07a49f7bce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e6cb48dba23ee87;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h665d2f287bf63020;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h496caa935aa6a63c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd654cd8e7f97349;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4cac999936a36328;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84b6c1fa3ee36aa0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h978c5fe0f481f545;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6de8081b5a90928b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd7cccb9fb679e091;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5399830820c2471;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda9d1d203cbd3d82;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b99eaab7920b800;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h964fd24209eeff2d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9ba38735f414249;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc993d2bde1312035;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94876e103f5ed6db;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff25bb2fb5d89744;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a549d206b2341e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6bb110dd0d914201;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h137e12d1c4486944;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7fb1b274381c0409;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3bd6da7d8c3d0456;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35129edfec275020;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce5cd67320d2cffd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6002668b8d1fc5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd803deed1d9bf9df;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb88e826100c0aa14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e061ecc53187735;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h646df95b139380ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62276877db716b54;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b44a9fd54e63580;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a73bf0520e72044;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72c46c301dbbd6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4efd3357817e949b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f05aacd4e863fe6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8323e98ba278bec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h314362cfe9a54595;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c368afe659518ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdee66f43e2664e4e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4165c70645e1d432;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67e2ed56faf8b1a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67c03615539bc33c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f6819b47cd3c025;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdff25e0aeaa522c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf62efff5b6b86612;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58c7004050e0881d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58d0935c06138d89;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5be149d7aa838b42;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha00d8d294c60b5c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heab4a7a4a38430a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2c3424118d7598;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h671caaec68b4f009;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h661ad8a7454d8453;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddb940c5c6b816c7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77b69280725f27fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc0d7518b0210d6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa3bedccd85c221f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba63d2dc1672eb3a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb60582545e58904a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46a679a1ae6229a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba519697f0f1cb36;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9af02b68a8fa6ba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5328defa25f48831;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44ed63932e4ec84d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79ff1c626b7a2afb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he96c240028a3e24d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ec7917ae2da2810;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed768fec7f9f197;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80fd9c25e28a5fe2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5d16d64afc77a1b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb334827b22522c48;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd327ab7494d0d6fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c9ca7a9f57ccd31;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f4074f190867b02;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae4c195a6ff56e54;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46e248bece92ced5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hebe6772edbb5a041;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ea4546fe64f9d71;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac8c3935ca1742ec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ee457a1810fdb9d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha255853b81b432f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf64c27d79116b34;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf7c603e7f3be919;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf03b006b27766923;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h284d3df5a9aae6f9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80517e486fbf2e88;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7fad4d9dc726304;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c88c9ecdda9589f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h783eabec65894c21;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f2825a385ce39bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd57226ab447382f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8531abb893f028f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96ad271cfc803a69;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49a42b7bed9159c7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85db92dc95cef82b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd545e17109b10921;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce9250ec060e923;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62b14a9e64b5b55b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa6a362452ff3f36;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3771c95d773b15a;
        #1
        $finish();
    end
endmodule
