module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [7:0] src9;
    reg [6:0] src10;
    reg [5:0] src11;
    reg [4:0] src12;
    reg [3:0] src13;
    reg [2:0] src14;
    reg [1:0] src15;
    reg [0:0] src16;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3])<<13) + ((src14[0] + src14[1] + src14[2])<<14) + ((src15[0] + src15[1])<<15) + ((src16[0])<<16);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffffffffffffffffffff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4677a775136fb0f88c1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2423f77a4332b6d42ec2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e417bef046f0ed5bd16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e8a7fc5b19aff2337da8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h112dea6c1086535991c67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h64142d33214eb58fc180;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h91484eb9a01a679308ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h166c146180bae7219c6d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h149001346d6e4f712a39a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39ec3c13889fe4691730;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac770268e98ce5c3ecee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he8c1fae148dc3f3a367e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6922999780d6294dbfd8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a0f8f423af5156c5dd6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfad84767ab5ce0be6dc4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h144b80e8b652bff73fac0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1401696a5a2abb8d5ebb5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h76a196f211f97ca48faa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1faa584d28fab2f96ef86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2feea3fcf0b780e2286;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9879c38b72849ec630ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he632464e5b379dbdeca0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h183cafe3bb20645e0e2b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be232076d46ec5157103;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd783a4c321e798fafee0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e740f3a9ce5c870f53ac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h53ee7f5a28897087f86a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a574368a980efdeb956d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cad6d386cdddc55ab365;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d76ded92cb394c79a1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd0a895deed8079920925;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7e5ea91306f9c6ee4ee7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14bf21ea500dc10cf95b1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hadc226012d97251cadf5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb8e823320857bc046857;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d3c5f904c5541ce8582a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c14cdbf5bf7760da3f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ccb790d3c1ac77f2490e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eba3f99caecc07adcb6d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb7d165932a5a8134ebf0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haae03d496a9ccf8e8603;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a6c4c8cbd140b6c1232f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hce81be34a21e6753dc3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3dbca475eb7cc0d46f69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e239ad913f303b9df6b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h59f98ab77f42f60ba63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16abf9a49e288e9924966;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92ebd174788dac5b4586;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h33881c14f6f1baa64bab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f84faffb1850bd22f18b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b6f580820e7cbbdee2d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1994c66a5985f3c55cb83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31993ba7529a5c1d4a9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f2fc21356dd27e2e7c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h97f1cc999e19ee0f71ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e2ad1284f8ef4a6e8dfa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h164a770527e6ea104b7ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ef1a61a5f91a1f5d4c6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b139fd57879e8d2431b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fcf3538dced689535eb8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h201ca677ecb4afc9bddd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6ae3dba1c18126971cbf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h73a248a5c6d3e175c18e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h333cbc74aa0121237f81;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21ac21d7749a0eb0ea44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h179ba638fcaaeba137e40;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16f1fee6de29ec959a40f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d98a770ad32a5275960;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h413b9d803aa5a692a441;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h81807b97eab1b3902e20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ce21445f9d8aa299f430;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb18ca93c0393157a6f76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc1abbc297b58c35e2d0f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcca8381f0bc29eab995c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea6f5cc2e040f0a11154;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10564a5fd3cd238707c91;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15de355cd39c959d77480;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf5e8096b9adeefb610b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6e04d68465b31cfdb319;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h636c9a75a41865c5fdfd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea6517a6bfb8d038f5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he2597ff284ef32c54097;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17808bb4dc9d778830682;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h49fe0c484e24bfdc596c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he6afa134cdac7d300ebb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfbcb2a396981bd7495b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d3328e6f0135af64899;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b7d29184c8adaa348de5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h62fa48a7fde821681e05;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c08451106aef75aaf68e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h67388ecad60a94632831;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ecef80ed364ee59cae0f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf95053e0fc52c13ef9cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1537fd67f2d391f4ee7bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h34617ab1de4ef7e62032;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2e12fba6b2bb23af9f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f343fe3d3b43a1b452;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf208b6064b1ebd90243;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14197b9886ca7570069d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b09c9c40aac74e4246d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11112a4a8540c4d16e7c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae184f5714d62a1e9ff9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b85f70ac11b2e4e753a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6d13b60f4fa8c5fbc2c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde9d263e7db3b8be5f65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed885088f24b7065651f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31367a15325442e8b127;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc0df99434ea8cf17bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3180e61cfb02516ee7e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4a5ae5dbe0345b0856fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e0e389072a0b32b7e1a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d5dd3d2bb7fc95a18f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h128c25a0f1dcd37ff2d9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h644fee21710f6f404ebb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11cd5b39d4e2b84c5bb39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea8314608efd46594e21;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f46725363fbc8fd6c287;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114296b7ee6794576730c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h699db160ee111e82eafe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h677d065f8ecb3412567;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h186f02878c4df24d9d2e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf7ede7ef283224f050b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f2b3bdb50406b3b074c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc77d965aee9341586f78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc5b52cd1a70fb0d526e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c305dfb71da2e49d468;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heba4f97c84298cdafc4f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17a31115520c1aa4a6621;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8cb833d5473dba14f6ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h36aa1ab6fc12edd38624;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39dafb7107ad8fab44d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d51f5dc612a94cbfdaf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1219f8ea12e9672a0129d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h385cc536f38a1c27f34c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10cdc96336ae50ab8e216;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89a52dd10b17815a74f1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c13bfe269f264e79c0a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9a9bfd9f14fb62ac16b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c085b53ad9903858f61;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38761b43fe8b58719ed2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ff0961fe3e00310361e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15748e287dddde391429;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h502e439ddccffca884d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e116c5e5c5f8515d2ca5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1587f4171373fb1dae9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h96d498a0685101454a5d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf598daff56190078d5fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b44c3a6721a2e612c85c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha02570a4a14fb7079776;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19d0e95625d46a821e68e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd38451220597e76f82e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f3c4222ec132d54695d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcfd59e9111a83792a3ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1818d414e1cea2733464b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c0131883f5fd8f4f2d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h93d1775b32ab8e40f7f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b4ec363d5e7273e0a1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2087642db3a5584645c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18741488b35c29ed0798b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b6bdb065c34ee5f4e2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h461cd91e889d2ef8fe58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4a47fb3ff8ce9c131fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h72c8170d2b440bdadf8a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1519aa079865c17e33178;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ad5132a275452afcf03;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1450ec3abdec4b580907d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb08b8e6690626e0ad7b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e945fa2e3f6810b71844;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf8b313b918509a318bdf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e636c563aa0ead4417d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13891a1d017bdda001a27;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e7e7a722318e139567e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d9caa70047c5eee6134;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b5995c15413626d380de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1879c674a65fbadf7857b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he4d09c91db7c2899a1d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16dc83e7c4a3bc868135d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca50ff2de96fa419c7b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4173ae56be38b9a30837;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h182e5bcaf3a00efe665b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4ed4d17d2f68c9e5a133;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ac63c00cea1309321a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d4e243fea7ec8c37667;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fe89cd5fb73a417fd239;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a912ea6ff79b7786d79;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d0147a29a50d7f22ec25;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h25bf836ac8d69c3a7e6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aa03ae6d5fba9f88aa55;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h71507532b1cae10d9107;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ec05bf8423fe06972d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15879a0dc8b133a3673f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde9c42100871182024e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9226b13259989a2a2182;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf61d92eaa5a5743a73e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c5fd52b32e18afc091c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h182eba42e9328f00bb67c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h316fea66afd09d01ea88;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb49d5c155d2b8e80be76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc9c5780c4dfd7a239c65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1693dd7d2404a4f4e7ac7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10eacd0993d32710be756;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ee149a68ef03ede3d0bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd395a59e941fb363186c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h157a9c833a21ffbb30fd6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f5d04d2862378077b5c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h78b9b1717dbe5c028c7c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h135e4701462e8de545d6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f4bdbd83d7f30bd15c1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb9da308a847a0fd0aea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a06530eef03f1c4946a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5471d25896cd8d715e1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1416465589498d0436bca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca0306221436b894bd09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c1cc489d6951109439e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14770d70e2399062f4541;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18734adcedd31c41e12bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d7d6a930453d69185247;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6ed91b4538c4b623f732;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e57db3ff1d430460b94;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b7f1d60ba5dfb8a85f57;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf96f2e1987f1b1dc4d9c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb73e360b889fc8b1964b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc16608136679d4d5fec3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h78e70faf628b3b3eab7b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba54e82a9fc7e9b35ee9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd00748e2b88f59cbbf5b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h85a9e0c5410a5b789038;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h91400c00107417ae512c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb6236ebabebba2b5017b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb5d3dd3e36d0b279208f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha66fb5c4bee3e7c852c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d2c5afbbaf7fe4a952e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1261699b66b1e8c0a453d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d9925287f6b0c26af76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2eb098fbd734c4cc9864;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h707855d1b3cdc666f52c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18a712667f04783dffd34;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h619157a234f9e57876d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e478aacd3d941cc7dad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8b45cba6b0568b1d80f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2369b538b6b5b37ab107;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2328980b1eac4f78f5f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192275ab481c3637edd52;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h489bfa582de99272b1b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c4eed5da13f22e482d4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc10cd25d01b7004ce4fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17aadebe1d2b82cad03f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17659934e0847a27f55f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4241ca51b696bef6f867;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb8f369bc3ab0abb5058;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h157ebd631d764394273fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6710890b220f50eabf1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h47cecbf6230fe71dc8a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h161826b26840a38de8c30;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed6e5bf738726390976d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1095abb2a46407d134d6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b2d134326c58482ded4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h386784d01d7a3b99245e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd9f797735d718e88983e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h168dc938f13380bf8e5e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9a083c87b161b5f76f08;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h753b2bfd39e3b8c3fca0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8fff39117792bebaa51;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd9a1221a45698dbb3fd6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha3d356e11c7110874c2d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7dfec65bb896a26f467a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba888eb80f66159bc37b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h33bc4b8f04a6c6935232;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h915de305785f4d15a951;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b9563b4fd67bff4ac6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18db59d37c9eaa044c134;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dced1b8f95f63b396138;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha40eacdd973a0f4ec4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19be393495f7d9057f09b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h154ee38de3846164568c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5c92170f01394e5e96d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18ad36ec3b595ccfc7a8f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4566315ddb97631071e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8a76c2de5475d14b3e5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c49723bfd6c0a859014b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fbf2ae5052e011561fdd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7bce298c92a20c4ff595;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb649f3b7721d6417a82;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c21af605570425c23751;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f457c75a4d4a78f13afa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb09edfa298a2a459a0e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha97e215e949f7808da01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ac14becf106ac1a0315;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca50c1feb3232bfb571c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdde83a49c4dac60434f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7abfb16adc7b984d380;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13fd752b59bf61b174dcf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bcc62fcae0ccf2d7866e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17547238e49d6790d798;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdb512904005c173cede3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h131161167083ba4ee982b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b55cf1b74072eb43bf1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b4f99d78473f9640652;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f66bc8093e2ec49fba2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d1025705ae3afb9d6e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6dba33b0db24e8bf2808;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ae551d9aef8c111fa2d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1866bcccce0e30a7736db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h137610c86aa0ccd05816c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ff2358cebf54a3fe9361;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19aee880583a2310a95e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb2beed7947602d1b41ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h97ba6b49171cd39e543a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f928774312747d8d66a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14660b7e04fca2c8facdf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h100922166d5d026283637;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7f179ccb3c588558c82f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb080501009931b79cbd9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9b92eaa3a5b68f65d871;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ec305549ab0238f916c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17fd80a8ce2bd44536383;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f5322f2f9bff9b80ce79;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c94316a1057edacc6ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16dcb2516263709760a49;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a5c99ef2b9db94b132c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18641eae56b52fe95540a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h132923dc213412f5fe5ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe30c91ef517f5ebe45f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h279da15eb9e0f1af46d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h102e5171f8132bd401aa2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h139ef80be81dfb149e23b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4bc9debd89240791b851;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2cc6dc5099034846309;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h142422560fee249c6dd72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7deb6757781dd0b04b67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ffeb3dfa7cdc55df986;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1df29ab7e3139241563d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1124b6308b8b07c1af3df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54bdf2743c6d09b560f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h125c43c9187326b13fc79;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h41629898ea271a279624;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha009f3b7e51eb87c17a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e28bdb53ae514f67fb7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h50bdb1ec1279036bd41b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h84955abd7de3a5cad444;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf8e9c25001f430e21d2f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2283b61b8741af7c22a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h376289fb9282d7d23b4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac0c47fdf988e47f4350;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10f93bb0759a2406b2819;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68c2dd253e450a49b7c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed6f66741dd0d0797ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb793ce1094ca5ad7b6e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h64fb34b47a1ee37e3098;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha6c32f3300fe7a8f9985;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19c62e76d5889537681cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h111a0bdf5130f75327df0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10a898b430cea2b8af4d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haf6ce400a7644cd59642;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5876894e397e9430b72e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he48b9d9763b123ba5044;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2da9cbb4975bc43599d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89acc00891a683cad719;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b9aa259cd88f21d86476;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h97a84395242960d91bdf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14ea5dc9673ccc37a1f6b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9c3e73b4db17c39032ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h197b30f5cacbba5505105;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1412b17384cf799bfc1ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68e3360f3dd20e312042;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bdbca1f75d3a21a1532c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h183e81e09caae1e12e172;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af6691a921ccfc1a4aea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hafd14fee0d472ce7dad4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1440986075e6c4d4b2d1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h93237930e99a034a7141;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb881f5d94035205c21c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f9f5461e35aa47b7a686;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he253deaf0e1e85613088;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f93b45972b82423c9058;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h157ff7f9c492a99fa5efd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b78f0d477ee00dc9927;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1790c84fd830409856b28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde95fdfd189f04432ea2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha7400b8997feccea6ba2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c0ecce56d1dc4adce5b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12d8c8060bd9dac26a492;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4cec3dcc0a336f2559ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6bc59c71e83a189ee80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1502eb99625e2e326348d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13a49f220067df27ae794;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192968fbd33f7fa6ba9ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b2d17640020e0da1b3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h421e91308f7ff1680025;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123ea4d5ed5fcdc030e68;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e2ea2b6057530e9438c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1282ead281f05f842a024;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15fe986e338aa8195036e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ce7724328579b601dc26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b64ad25b461211ecae06;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19bf2d8a66eeef6cc1425;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6410e9fe706b69567938;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf277f451d595a27d90a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h984a3a86666c2d66352;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf6a5bf63adaac617ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1753f0d4e79358e9adf5d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd5c41cd407bc1462e9c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hacb07cf85f79673c1e42;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e0e2bee44cdf84b4ff2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d831e31b6bc81856cf6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1840b96bb09b4bb2cd0c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h69b516627927df5742fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1111e00da492464be9ecf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4722bae10882350da060;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heb586be9ecbd1ce7cab6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d20e97c400e3755e057;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12537a3645ba98844b4a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h45a66db266900a9c7116;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83618cb54b87c1cf0e00;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6eeded8a8f44be548b46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac04ee109af9b530c29e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf4c9fcdbe5cb1480095;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5440e26260d5bc322300;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b85df1d675e7f92e5a4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed37dd77b00e9008be4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h804cd0cea5a9fc2b4476;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h793fd7c86d55edbe1144;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he40a8c215ac19dcef0c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h47cba57d20fe03553239;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfbedefe4c4840c6efe96;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h163a37aa3a93df6440795;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10111dadfe54046846d98;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h244b058a4e550a5922aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a365e918475e24320865;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3abade4954b27df0fdbb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha7a8fa794cb9a62acc45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b469f3a48991be635c46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he40a8e62d2d71ad87efe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbeda82c6948dbc40ee71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha359706e487ae49712ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3fad0cffbdb49fadbfc8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd7d81479bd1611326905;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14fbaa8ceb2301527e545;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hffc4254aa49ac7f7f2f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6dfa63e1516fe35e35d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h132ccc71e83de03d5bff3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haf994abd8c70874795d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e4198fed9d9b80e1f65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5eefd6cae3f1133d7af4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5e20a61cee1a6f19adba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h183d9d364596d82b36b99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf08b80efa6f5e75b613;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h61f534feefd850f3a2b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h87ed5f9392507ffceafc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d7547b96874450eab4c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h167ba725066b4fb12ae5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h193d8d36ebda22979f58e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h905e638a8b0e4aee9c45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h198f164cbae9d37ceadb5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1622a3eb296d2d3d36384;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15034ab9005505f0a3e17;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h156ce2bad56b7b3d0171e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e169aee962457fe65564;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c4b1cafbefad30e55bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9a70807a820de90746f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d3469121b4911cb56b60;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf1e623a1a834c88fec9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2cb6549f59387148b546;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d90dfa8d6ee80d5ae04;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14ccaee66b222759cd189;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13640c521e5796aa0c22c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hee9dc97d33d91175b10f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h37a39272285c19c80547;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h824dc029f9a5bd3483f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h244db46f4421d7f25fa1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdde0f116eb864c4d78e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heaf0799f84f39dadbce5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1581167bec450fe117037;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h445b8a2868c8d7406e9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4a3a4e583e10a7e646d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h685a364ae6b73aca3d01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h86270d6d88df2aa0a6c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a8b2463a741ee462af47;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1443147166f7d7299b5a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbc528fa735a0f199c753;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h58ba8910e88fed9dcec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0ce3585adf22dadd865;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2066bedb5a32dac4f4c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17e13b25706e80251d994;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2812cb80faf9c446453d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c0a2a79e11ea8b6eb2b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c314a9760c41abafc1cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140e5b077ea3e18f007c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb89ae63098f023a98c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h376dfa2f4db5e487f250;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3f663eaaa45c81f3c97;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13db79804475a7900e01c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1146a8f38c221c6a9ea4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5bda350306c939973e8e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a9e2a6cbdff69bdd5ca1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cd8fbe1538453291a8e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h162331041a530a745cb51;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b164d684ee41bbbc8aef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h518364ca7891ac3d498d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h723d598cb8aa1dd1db2a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3fe56849c0646a6fe4ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd9703c947d186091edf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcc7b07c06e68cc427904;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1853b59bf3f02c7a94ffe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1826652e202fe70bb7846;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf314692d9ff7a3298c78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h132951d447052c95c4fec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f508198c556bcd0c31dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11b6630391faa00babc59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d862ee2923adc314e123;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18f789c79a014142a4651;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17042f5c92bff049bdc76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1758a9fb6874c15ea533;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4ada9ba5069415a2660b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1591c212d188d8ce982cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h775e2245f43b7d76712e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16f08e90764c57a45c859;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db6689664fbaf7af9298;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12880d8fb5c3cd573d4c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c1da907f70680b27cc80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5175ad950c2891f2e463;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c1f46c9b2dfddbef709;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1643456f92242003bdc15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h36802c948cbdc69f7a8f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h181f5ae4c62c9c61e5a2f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed2d7687abcf7cec190b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c032cfef69e67722e782;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7dd3469b723890977489;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he97096af680938c2b0cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd734f608eeb2414df3a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b65c5248c40ffbfbd34a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hefaf636cf02e563f71e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b2a5677a726831008847;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h414a3e7c613ed6e8cd5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd35a13fc63d2eb8bdbfa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1256ca6b38ce2f293f192;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d149ed5a53894f8f2bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192c03a8ea42184120836;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7dbd19b3e9eff25b0a9a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ebacc1e48eadded16f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b24afca6f0cb2814460;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h665288163f3c347f70f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2c49cca5e8b9a8479527;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c29bd94cd841365b3793;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9e1cec3cfdf459cf4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ad22f871df5c24c4d032;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h180cc765c8552dfcebceb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f621cf1d5b34924ec250;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1345b4790f6a033d734af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h195e4d3ebb595e74f5bac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc98fcfcc75804fdd3200;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1edd37938dc172b6b35d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbff63c156d20fa8657d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19d38a302cde62bef8b85;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f507abcc01ff1b08b1b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17cd69fd6382490e7d8f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf4995a2707b2b9ddc5e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfc4137e87aa16fb9365c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d2347d7fd325dde0aab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13149c8646a6d6546f0dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148b1947a11e2bb6b9d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he3e953767f316232cacf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h108c77de6d3fa89455feb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1118b8e2859f7ab377a3a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f8a4748dadbbfbe8f31;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e8ba9d5c20147e6170c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf34dd18d2bc94adaf6f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d3064d7ae6921a049f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb75ec285ff4e958e6dd9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd209266ac2611f5fe1ac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19286065902b0ab49d0f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4b7f2ae2f135006997d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc61bee93d2056be0a875;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21f595930a4cabae7de1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc4300c49a43ca13f966;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb2f6ddd6caef593330cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f960f3d5f4d7609cd28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44c6100098b85390e876;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ef57c0e3dd3720b5ddd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf9a7f77af0200cf2e1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he3feeae3e9c16805bfbc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb033ecb09b3c46b6601a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7fd6c5e17a3540309c48;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bfc12191bf46750190d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4fd9672df9ddab4045b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19ca9b86b95ee0b4639b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc98ca7ac11f9f7c33fa2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6aa59cb518336be696a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c6941d7f66fccac1550;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h99575064187dfc23f4fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h269aa296f3a7f8406971;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha219cfba972cc9f33e46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e534de9c3fb5c6f49e44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ad670238e668952bca8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a84890634bcd6013979;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h163421cb7d802db2f11f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c79f1f0c4b1fc54911a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1181cf6dc653b9b1bee0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c246ce52ed451971f1e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha7cb4c797c6a3a725b33;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12481d31050c4a30d0327;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4ec58ee01c976739d84;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19c73c777d1bb2d460c2e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7146deb05c49e3268bee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd416db0c629dfc19c824;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6092c14f85440b850ce9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1989c795309d704300ca1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b11b19bd0600e344f9a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1993ba857a492aec23fdc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h79f6298931a49302fc29;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d356810c5f5198dfe4e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h47bf8dc6b7ae6e2a7aa3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f3182e763cf51ef4045;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf90b0831821ac612a2ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9f9b2206fdc171f0a862;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h191a56cddd9c94d663bb9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd7af7c8c61a03853df16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16fc65b358633d1534a82;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c1e1776e16f1dfa985f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5261be1c46c0ed092494;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14312c1dff207a3bbe899;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1370223ce2f7de6f08730;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a4b1d666101f80783966;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h190689a5c2b2ba6707a07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3233dbdec89fb05be7e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c56db32cbad4114131e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a22f1637487bcbae282;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haada3d7b907805f34340;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e6ce91a8c76805dda80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb0c5e862bec5bdb74bdf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5dbfb496810dd7049337;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c7c868688355c990949;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d639117e951ab078c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb447bfeb436ed7e97e00;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1504a01bcca3675835c7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h32904d95f36c13e809bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc42e86e3b6763de4726d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9b1204b3da964a46d56a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8c05a6c37683349050c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6266f9039d2c68079f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h88aa37c20e4584c8f862;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha962438b7bd03e6c0b73;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a03ddb0a2376baebdb7e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148ea409c4f9e71531428;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12eff43c860564805ca0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15fd63379e9e8e52604fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf9ff5734a8c9cec39eea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16920ddd98369afd447c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h50e84a09e24c6fb2afb6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf0627e44961cbf70495b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb216012b7a4a3e3bb109;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22152c227bdfd27dcec3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b0e07e8b8e9aaa6df56;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4640ef86432ab618c895;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ba4bec559d512da5fb63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d951bfe0c20ce8924187;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h165568291c7a10700bb43;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b0a6743fe6623d15b273;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd0231e1bc79b9def1910;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ebe679c650ab7f3e260d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13c57f90ed31c22410741;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b09e1cd2ffc82943c20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h164b5b78feb0d0137f9fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13e29ed6a5eaff06ab5af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he8c3d6465dfea70946e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h126883208ba012109dd8c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14dc843509d13425180a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15eee4d21e8429420498;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha95dd8595271c5ef70fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14064079d9515f5257d77;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10fa3016b32ab8333f07d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4d27a376541ad4ad517;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1455d57e34c0348af52a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbcb7264845df5a936816;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d00187d1a98e4600b1dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h174c11804053f0e1d1c72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6d675000364ba89dccf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15440bed828f6cdca1f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd44e6afeeced7a7aeb1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9bceb795e5283548d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h414a134d65a0e8f3e2cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15dadeaf43e0cc3b2d74c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b27f7712e7d0bf370eba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ebfb4c7efe33fe3f2f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h190590ee602ba9f6730cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10cc1e22af24c38e8b13;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9da6075d978b56af8eb8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f552aa82d2bdfd8300d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h759c309f7ce9a4f394e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12d4f378626902350b47f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1562383c80c2198a86b4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5aa8a663fbfceb1f3fa3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c52f25dc55c2e31176ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha943fb65743d2b60c5e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1398c93b75c13d7ad6419;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heefdf1bebedc6580b7d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5d2d1a7684a6721d5412;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3c0668683a3b780e3322;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ca547a55e66365cf4e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ce560095fdc9f7decd1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h142fbd0ff93f13994d379;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196c2e94d9e498b776566;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8df001cad2d1cdecad4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1240d7a66a2db29a1dab8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1856aef974f71fbd24b74;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b9882ba4c1fd52064f30;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b25d8784a006be5a1a9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c0fa57e37316ff215c87;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c33651ade8194765941;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h144ba4d39630abeb3210e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfbb13977c1b53efa4eb3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d687cb9856a9f4231443;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf2febbafa067d9be07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf19a7b9c0954b68d8f18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h328570e5f53ae5b82a63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1242e22cf7ace6a600ad7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18ce3d6d461dfa9f05356;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11544d5aa5b5d4a37934d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha0acbc016e5d5d364e3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he621559ccc508bf42104;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6f227fcd2ffa74689fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83ac01ca5a59f56702c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c88a4525d457d1bb964e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h162101a2706220246f1ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a96c6149176ab891ac28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1feb7faff54c7ac77fc15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h406c6758734754bb0fdb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1822749ead21da190160d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d6a68d337ef29003cee8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h799edcb703740d3fd90b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h67a58f72ee04377f8991;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9325970655ec9a03a50;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h193a3210351b6739efbfa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcecda56de6131dc36717;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ccfc752d157aafebdf89;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c1588bea70b38303d98;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h41037d35e57eefbf222;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf3059bdb3652b3085247;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h65eecc89ad96f9c0a290;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ab393416d5808b2bdd8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h202589022420c6a3cbe9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dbd07f93adf7f66f1863;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h27499a767c9c9659aa45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbaa1cdbf4fccf272c509;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124ef31f70f1d6713197e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e0483923f6122abf0c70;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h32642cca30c999ef0d4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d182a1e2d6acf41545d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd16ad3df41b1a5bc4bbf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h97bfd434f4789f5ee60;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11b9c68748b8b36b5750c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7988da329ba1d069f149;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ff58367cc07126c21852;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he270437249f3bdbf9187;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e25d2f089f0872faa5d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7051e583b7f55846b03;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h48388f8abc483dd5d1f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ae038cb4a2b0f6e1935;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h332c953ba46b07d7b6de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6a272aec42f9089dd65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde5e2cc45284636b65c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3750048decef7330a8ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3f66359602d0c398a52f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha3d0c38b4ee443ec1b5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h118a997404c03a6110091;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h47835524402129d5da15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ad56bf210a2a005b5ec7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16a05d61e9572c212b923;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha07494f0df30256adbcc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba530dac91a483c21dbb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h160c57ee12fe4c9821ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1176497d273c989d28b6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h191f63011e6b6175cdc28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16cb7b7caf53f71b88cef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d806493e12bafa4b87f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1beaa0ee2e648af9db798;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d9cea243473cad4d22c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a27f05af76ddeb396655;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19aae30ebc1f65109e1f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb45e0b811695f6a9e80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf48cbcd0de429fb7eae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hab2187a3545f97ff4b64;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h45f6666c962dfcb886ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h137406d9a86a0b150fc55;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e10957cee3a329563e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e272591c924793da770;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd9b1b65160e13782a6a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10ecfe8ac7cda70dd20e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6bbe703fb71e10216315;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b428330812dbb9268803;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c77c4dc9c63a1aff0c08;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h56af5e24c4ec53eb3802;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb965791e6dde8d2f262;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h37bd7ceddb6c2fa658f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1058540121e2bf7577f52;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c05fc940f73336c0bc29;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10946eed7c0b1344e70d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h37b015fd8f773a828185;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1536a51934b74b7b35326;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b0e9c15f6b0739f8ae28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10eda13f6ce52766b5a70;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19773f48cbe51289839b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h165dc65f73f794ceb2b8f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d6f8d5746af3dc1d998e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13e0d3d44ab0a048212b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdda8e575195fed7c1d79;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f5f02c26ba94064137e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196243578710f5d2a50d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc92bb0b07a917e3b1ee7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h163502a482bc0a763f491;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d269fe2c3a360c096347;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8ea4ae9a2e03e6bd8128;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h113aba8d3a3369fa435c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7e3ee58c367b4560162;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f583bb828c7bf11c9bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc2f61e51f830a6866042;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h128c21461b84a64521b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e16d41c5adef385b5eee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1986eba4ca0d69a6caa5f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e6952a3622aaf182541;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d51319c1c5a75a2fade2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d3295c1fb35516b89be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1722c6a0f1059b5119753;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe4a9737240126b0ef49;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h775ed964e88d8ac1e175;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a8e3fce4f6f60d81428;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14f0216fb0d36f1426039;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dccb6419c2d5516b9011;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h102c3f4a73d96e75bdd96;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c7a5c3c5782e7fc5a8c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18dbfae76c1335dcb2f68;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68966f3682432c17a73c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8c0f166f2c56719eb125;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5fb1b952abb8989b212e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h340c0f2087348ee0217e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf75e750f037f07eee06f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e595c669436ed8a1d22;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e92f25fefe1cbe39a5a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2a4928fa733eea724797;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ef7e60a02eeeab47c95e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha6f45f7e102326777196;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1daf5c14ad7946b50f359;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5966e2de4ff53435023e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h121f237394d99c0011d96;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b7ef32696b4b3304b51;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb933552c4b3dd6c3652f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f17fb7b80c8e9257935;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10723e5ba9b86ce030e47;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9bf4f1559d477c286756;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16efa9a7d1cf30c17fa5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0ad241b37aec8dc0a6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1680f4f676336080b9791;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c7541d892c8aa80d959d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb07e7cd7d3405c5463c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5391cad832c15e72a0f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1094f66f2d602d11a05a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h168f0449e31e4483bc510;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h186db6355d3885d8d8222;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eef3d29958e012b09a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd095e9cad6ae3ceb1ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h160b952dcf3f935b89259;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196f72d74f9006309142c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb7195dcb905848579b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac1cfd5ca8941b1e1b61;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc153f0268fcd1f0b9b4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31977ab0c3b663b71798;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a4362c77051c56a05edd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d6afb99934300cc7dc6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h87539b4163cc1e83bc26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7efd6cfca96c503bb742;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4e7a9d5d67d180bb22f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143cf2cd6cee65ea0b77;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1234d74dc7e35958afe1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1521975fd0cd880c391e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h847bbd6612f60a38dcab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h117834d9fd9d9692b2648;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbca2c3ab686fb7e4bd28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8589ffc6bc820443b529;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h106ff196daad577dd27d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c14677a7ac603746ff4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd7e83c36812edc796117;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha9248b0266a9de7b624e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h75e039c04522b1cc69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16002e661d3e57f370d0e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h138756f7f1cc54583f333;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h125a5b068a96f53cb44de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13406efe018d0eaf39d51;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12bbe4a63b357faeeff5b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h112011c3b874897430d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h263bea27bc7b5216b035;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1289b9b8509b6f63042fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h307a104a2524ec7342b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha988edfb972d159c8ca7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8f0cfb1720abc3460de8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e22cb0eefaf8e2cf732a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c60d385ff258244c906a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h65145abc65c3069db4e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd873f090b8bc636c00c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h182bbd19277dca2e3a775;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4868a980f3e5e246cf38;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12fb900ae95a731652e55;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8dadbae28153d74771cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h141de5de20a8a8e637bbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143ae82deca96b135ef4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbad5b722bcd6a04dffff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h383fe36e83b1862416dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f7ea5c65d7329bacf45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11b3d09c6b62e09d4a259;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb28473d87cbacb063ae8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he50d59c8f6c0f777dd7a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192aa3602e3d58ceb0162;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b1476ba5b04d94a60849;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15179e20cd2af649e017d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd0813d2e89bc084db5df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2faaf71f094b850e87ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h130e9db7b3833a668c6fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4810ac3c5fd275a5ba64;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1739deea1bc11268e6e36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf90e9bb1d994ed8ae9ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104572667bbc62999f26f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcff148a05e81ca906934;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f9426d57cf7371e94c9f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d612c692ee1821af7a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h595c3d604439d3d74516;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf03acf4d38b852185c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6672b27767a5ac51a2ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19a284bbb480f4e3490b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h93ddfa8b3a8d77aa13bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14685c7987f115521ac5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d487dcc05ae8bb33f0ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15256024ea44fce03554a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dbcf7cf321b7cc1cd2fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c841b27471f5edad7a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb444f52b9058ec5a97d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e4a0c2900e9ba04f467e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5026510e0ed7dc97edd1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1602b977e5dbab941c75c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fca45c068e83665c49d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1956f675c64c17f90b567;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf3788a03d487e60a27a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he2709b1a4f0a1de21b04;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc8f6d8a6c70c19be9124;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1746f8712b06ed83e3bac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1683a2dac8a40ad091869;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h90e92cfdc39b167da8ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffc0436f230235ea5dc3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h113b6a56e5ee47b9224dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h87f782b1f0acd03100a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b7802b33d964d7e1e27f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42f47d61d344d1af59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he596e8aee07b68c3123b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39f71529e36cb843ee68;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b12d8c1e94edf40cb1c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf495c53622bee080ebc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1349a1ab3ed90b206e1de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h53ccec18c87894232786;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec2f2f50dae8b8d45bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0153054d22036d76c2e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7fbcef052dd0d85d7fb2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h55583bbfc2de183e0515;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h118f9ad8c06e5e6b5129d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf839057b2f7d916077ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8dbf61231abed97ccc5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbbd849629d4e9db9cec9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1da17c3a1b41aacbaa25a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f618f58fd981419800f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2c50de2365bf31557607;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he6cc60b715835f7e2f2a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb8ba84dc04a612b8e86b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hadf0c823171ad79f7c2a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fa656ba6558aa95c8a20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h813e2fce54c2f90c3fce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b5c1b330d88473f2424;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h147d6a3dabba23ae70ef6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7b27eee377511ed6cb0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha1154eb54b36824010ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8ac783f093898eda373c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a85bf98bd64c09ae699;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he2c6e7a27044a9eee877;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b4e6c5953780998b0c53;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18729baa7c492afdd5e02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1108d4c6d564811c7f052;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd86d113adf7edab1faf0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a2e716f319ee668e2419;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h151c3d28b73180bfd13;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12fb25d7ce03289831cf9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hefa6ba83adb0cc435b71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16453294f4ba286b199e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3aff90726d3192a522d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b72c26777ad32d1e150a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fc36ff069353cdd46010;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he10c99b59f92de508845;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16612644a802cbf5e7f80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192888d65f817485d02a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8057e2d372997df55e86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123e495cc3fd0beb89a3c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e1112922683a228c06eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h847feed45edbda77493e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12039cf603b5fcdb4fd5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6121aea1f44721bfe67e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12cd4d97e134ac476e8b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af42d99558434ace974d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11917aab3c41fadb275ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f6f08139726f274313ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h132bfcf1ab534ccde2cc7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b14be30bd93ae9d1f0d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c5c25e3d074a7578f209;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea871b5da83c970c4d10;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h792b19305a05955f97bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h172a72be2ab1795ba7750;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10046c9f889622c26e0ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haaa75ca5cb6211b7bb18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h397d69bf317edc457344;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h187ab2deaa7ed2bcb68f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cff161f49ad40645db78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d91c48ef5cfefe84e300;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9613a29d9383c1d0b45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h142eff55d27a77c6495ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha671005c854add80841f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h59836fe109deec0ccb3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1714fada7b50f5d6bd36e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e51669946efc4427ce29;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he55f3f0746669f99c8e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd7e1741991b932f18980;
        #1
        $finish();
    end
endmodule
