module gpc1_1(input src, output dst);
    assign dst = src;
endmodule

