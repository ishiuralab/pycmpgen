module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [20:0] src22;
    reg [19:0] src23;
    reg [18:0] src24;
    reg [17:0] src25;
    reg [16:0] src26;
    reg [15:0] src27;
    reg [14:0] src28;
    reg [13:0] src29;
    reg [12:0] src30;
    reg [11:0] src31;
    reg [10:0] src32;
    reg [9:0] src33;
    reg [8:0] src34;
    reg [7:0] src35;
    reg [6:0] src36;
    reg [5:0] src37;
    reg [4:0] src38;
    reg [3:0] src39;
    reg [2:0] src40;
    reg [1:0] src41;
    reg [0:0] src42;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [43:0] srcsum;
    wire [43:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3])<<39) + ((src40[0] + src40[1] + src40[2])<<40) + ((src41[0] + src41[1])<<41) + ((src42[0])<<42);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f55938a775f8d884b2831a10da2650e798d4f66518cfc629d975ada95cadbd09b401ad78d4029f1246dc4b5abf7e91491e8a8c28e2a09f30692866c1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha579e1d58e6bb1470f79ab440b7ae44fbe0859cc9c48ee63450062a6649268c880f6ac09bb9ba50a49ea8ab09363597d94b30106f17fc6793b9a09a66;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb27f429c296afd7d7ba6a6089730df3aa7aa973f3b7547c73458da7cafe0bbb41c2668b431f2312c2967cd9e5f3e4bf303d7387536e763c6e5f5679db;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf5f455295f0ed028ca55b40b3b38ce785d343df068b03080c5c65940c8ea3e71c5026b1d653df189953e9a49bc6dc561a26e6b29acdbf234c2d20e50;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9642ac958728a890b0bc534e5d484107b6b3688da01492d6aba54b346d5d8c97362172ef15012f2998dc37ee6b35a1e83773883eb30bcb62e90031a1f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf94ad45d56c27072717a1424b144545da11624dc54cf53a23aa7c8f42f1d5f5e3467d241ff78c9f82ccf4bfcafa5161e3622c1957f5aeb3a2703ad36d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19715afc17453345b8515b00ebfa7d38b7f16c15a60c4b187327353d60abfc73ddc6af6bf1c03743176654d91afbd2439e25211ca9c152ee45138dc37;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9359ca5b9e5e49e485b5759d14772b07170a7cda86c91388e7fe11536ee44ff6cf9a3452e854c33a0f4bd8ac6b6a3283db2249f592ac4ab8822aede24;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcadf6a7e1bd8e52e64f2c52badb70e1cbd3e10b4e43c55031bbed7a75b5f8b5e08af242988662d147593034a89b52c12341779e8903848f79ce0c074;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8e17d3f878d74f5bae0dec38f37ab72faf8014947d30ee90900cdda7dc38e4ec0e0cbfe57f3116bec81976b14560527247eb8adc2fc37082df60d7f6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b563cf07a6f46a4e720cb807eb068fa3cd325bd00e100b0510906262938358218310d48f1440514d3400157886d2c0759db2a117d3fbb95001952f78;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfaa2e06d7e0b0608e33c8987f88340bc74a929c7a135ab7a9b142d6620184ee756c597e8fc86d770916ec41bc5a4494b95558c6af1a44a2cb23620907;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h277e93fb4409ab0f603c0341ae7e8dc8696aca038c377a6581a9657e563972cd3152c78d40da80629d2f0cdb4e07a082f51f14900dce8daeca25306ff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95b48044b58ee180daca33ed85798ff1a52b77ff3d0cff25cae952d789d29af270b52c2e560fb121b34408cdbe861b9f2127ab1fba365942523c41683;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ecf409912e39993c27bde950f3ccb5f3d32c3bdd180f7f00ceda6f432f13c52b4edacad0ac2172bcad90ae5b68b501786b82f4a0d0299d698a4cdbcd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5eb964df1d5dfc315c157cb927180f4838d8e781ce33b70a3a00166e8d83bc845657acd9dae2c191312a86a6e8d3cf4193b200b8d134aec2740f59cbc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc729a21d1010aae3c49a572367d57c5d4a34027863990ee9b3a636a09922d21d8dcfa592db9d73191839c110480afe2d3e6e7e1e8a6de972b4221af96;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49b5c239bb2d8d4f308ec76ace795b318c2b8eb52cc909074ad666d58882fd43624f0dd8948a9d88ac15040062ff9b1f30ee77112b36ae97b1455db7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbfa1b45be861606de5cfbdb873d888407455e7d3d5ec3094dbccbd0c73a7d3877720d99690894f2a07bd5f03ca4bd1e1680d45482ae4661be7db2ea44;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11e454ab9c01144393a9739e8c32b4cf5ab80964c61b7b6e47da58d195dfb02296789b55830485fe6e77e1a8292deff10b4ba6eeffb6085b32223e65;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd03ad8a0f0bd5dc915cf2dad7f22e86930d257d133842d9b7d17a1801d1349e8875d355294aa590cd9ea8fd2da228af7eaf1c18950c696a869751cd73;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6cb8c289cd2926002335b39b4eea0ef3aeac32c20bb3f76f8a264f44b8527d7e5c6182c92799a1536d4c2fe65362cfb22a6e1fd69b3d6d993be509c36;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h377fa46cac95f36f0b820d08a03090642edef149f233bcfbccfdb1dd6bbae7abb1c04cd21f5cb391ffdae05373a7485b5766d170750697eeae2301467;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha384e1329ca9c43ce6f6bfa8080c0790351546ef77a8234d6bfb74c4540cd19c5e279315719f36cb67309b77d15c4ef4fca339ac4856a15bcb07a7f1f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60e3a152be05d7a51896bdb9bb4eb6e38b4019b623aeab5e5ddec37d47702f48775c90ab09026767db920095f864e40ee6a5d7d2cf968de80d76d0c2f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7eed8c785a463245549666604ab01876fdde872a08b08944ea4c0368e5ed67a67c268d09a792a9490a5e11f069699d2121941bc521c9765d907181ea1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73a31c7957216bf3b5b7fcb5a1e6525eeac74551cacd82031ccd45fab449d7831382aab71f137eec5db7e208a8ecfc339d279b6afa6ace54602ba1887;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3507432c046d5bf246fa6ba4e19f530a5cf4dc2989cf202397b8190e1e4bb6d34f0331fe70fa5dc9fc2a0b975f44a23df0bbb15e6a0d94bf829620301;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h271aa2d72b79450e3339dbebb29aa2c13adc215433efdb66e2567908ed85f39031678995d575eecf7080f52fdb983095ae609c884c01acbf683532506;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c5688b12fe84166c36a7a5ef472f2517c0a84297ca0fa00756f48812f48225df4f9596b66dca6369c78d48c2c6eb184c13316aee17a2420e1529a228;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2975572c53ef7747af4b64e2312ea15fb6b161ce400b2ff46c7983acd7f34775f33c86bd13d97ba9cb2586351fe16065e6d84b4a60a17db0580e303ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h111359c6dcc9d43e231598c81116bc1cc8128becbfc2eb26fcb82d08ee5dd46f104e9796bd4290301fa6942e6a45e51156ad5ab1d31be3938c8674668;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c321d88e29c8ef2d1684a3d077d9f7770c5cb2bf22e02dbe4b4887eff9a05d8aa104759ac82465ed3d7e0b33faed2a2827399e31844c37b20207fee9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4d46392c20dfd090cb29e12502685b93ae1ad88bad9d5b5da390baaece42fe4aba39851f5c500b8ec4ae9355a3eef4e8a910abe909c7ec96ce6ad255;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc701a78c61354815befc24fa09ea6b7f3407a5a39aac26403ca6309760bd3c9b5eb8e219c9a10fe788e39713a74963be07fbfaf07c6ac2695ed311ca0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fb000c3372a210c900e240b69c6cbcfe9bf4cf70b27641208fd450d9dcc44995c9e13bc4c24cddfe34461a0a137bfb45d003e46a2f8eefbe4931a5a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he431fc83f8a693e836840f9ad766e3e058275ecfa5e8b21784f018a7752cd99e919dae640b59c84087622de5f935a77c3bb6f08580fc23f5310e20a92;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haccfd8286901a06f25bfa5bb0fb7bdfe9c8cb665214bd4cb9185921d15daafa17e118a2e99645e56ac54491d3ac13efa224a8a07d24e851a090f3d46f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ff8d8b7cd0beb6472ee1baf47e430b44990442e615cf0247ff8e949cc2d0d4d2510cd3ab25abf76766dec6f6cf6442bb828281cc9bb9e4bfd89276ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd00f0d98bf6e549d04eff1385454a433499c6d2295fc80fa20a2aa326178f00b66fb9a746063390409fce917976f0acf346c82f7d5c060ee657f2e67;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f71cd6c306793c20484781e358652da9e9aba7dc9cf87ac4abce6c3055523b4b545ded6ba67d2e63a915bc2576fd4b8b8e9f718b5e446e213fbcad6e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e9cee40bc283f3523ea2a908f262b9aa03c956a80be40620d508a8033745200f9363ffd493843b8f6613738275333920b6ff9991e140c3c027045e0e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he15636bbad5894117a02efe4b8a701606fbd66f3de059a66aaa9c3e481445971d3f7550da5d624cf48f551a67b9c46461fb8cdf0f985fe43053a8d3f8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb134ae15577f8049ce1f10aea6e0d23b1afed92500f9b6b1c3ce320994be2600fb8ff5c41ff51f0af3a59d03de19fb25fe597ef381ea48d6dba1ff89;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54d57c9cce70392fb96a7971af3ddd51066e4a7fbb05ade319a962090b97d0c1786076b8260bcd0a0c6505860a05a5cd18cea1da1f0842de6d6d1ec0b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85750c4dcb767f80ff338b4c16c6d46931c7449d2e809ae748a4b5fdb3750c199a261587b45803e2b3ffdfe19ea3128f2d116333c9b1139238aba1b38;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb2db2aaf4200e33979d867fcae67817d939f4953e01d8bf321ac3dcd57da7cafa0e42cfba80eeafa38af8b4d60b2dcb57e5b21bca7df91fd39cb4451;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b83ce109bd33d687bb3e4337fba8f8b713f04238746f1218547fe172506403d2cf28f08ad3484782fd65989dbb345a00e58076512f40dafa6216cf53;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10fe161bb46950cdfe3b18c00b2eac5fb0b35802972f22ec9f9dd88816a874a47167377ea0be1abe01ac8630f49968e8e429930842b0fde009bb4f7d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38445a4fcf46025c01a40bff64b23ebef3b8331b23dd9f78a366a9f6ba40ad44f2a75267f5f9b3e35d162559e969e58ff2630a6db58c7e946ebe0974b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ffb31e6f452c60007567c65aa903b965b82b6bf3984d1adc1cef44e6c60a6fbf1c87cdcec1bbcc01269eacab28af712626262bce43982e87b5979002;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f17bc5162f56897acd357e396286155d98831b40b8bbf94cab82028eb3a7f21bdc45d38c347d25c69f6d828eb6682e6f4caa646676102ac484d68981;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc54f77f9dcdafb07d5bf70a38dc25f9dd7d68e640482f3fbce68da9fccdd90bb706b90f87fc2720cdc0f76c012dd482a2462725d61e1ed0665402608d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf312a85855072e77a04ac63e3bbb1383372c844dd6b6e64c62abdff2b08696cf97e63afa93ec3520bf630e1cf0f150eaa083291921d69efdac8d02898;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha92da928d9554f420aa3e0f8880df68afce4f50f56b79376e8521d7faca94eb010599eb1c7e9e4d3cae29865c17c3927e9839f0d3b14125a3808a07d9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c8c97621f83544df20695590b7e636b2260e09ef3c175923f06d31ff5c409310e0f97e9a0ba89f34289be1a518c2b38c73a87c17d4000eade9568962;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22478d9ae775284586ad834d877f7f5371fe4b08e9872bc6d12e6fa3a3bf937b462c714536cdb5a6f4ef92bd5d42a46e90fb832a8dcc761b78630fb1e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0831165f9a539d6772d3f6245eba53f40bcd8db5db13380bd9daf1bb63c5e6909c4c94fafb0d35337f89314c02a49bc073ca03e351521bdbd0382904;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41532f4d3af7579becd249550bc9809dc2a3070faf811e77c4b29c9267d95973cada683a72307e85afacf76c25197dfc38aea5d0be0c441108869cfd9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5210c46b8736f24020a70eb8efe1a162f5392dea4a8a4fb3214f1567b0e01030a7ebedf4172fa57650c8aeeddae21ec714d5930998e7b5432f7718888;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12ace47b67aaa3c19cf56e756c20fb11659c4528e95f3a87fd0afa7fb7efba5028bb1be9cc061771b98a0062fab707de61479587686098926eaff145d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he1934a2a6dd0c5a1cc9a16f0bf0b3c4a162864577962983bf3c0ff0e401d3c7faaec025f62ffa527671adb3d897b9b0c8b0167b090a91ba2cc96a73bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8d583e5690b7e7ad57ad9f2ed1e38b8621eb9f937e08216724a468062fa2258dc9a5fb779718dadc24be3bca1cf3879be32d63aa17535fc2f5de2dae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h810a01f5bd92cd7ec69cb6a423f92b779a4d389a561fbfd81432d0a21581b1b6d562347b29cb9a6ed290bcf1174f47d3ab558bd4f997a7a83afe61eee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd78bb3cd5329cf0dd68015cffa6844075548f3012686bc3170e44cb04b8373e4300e6ad7698c895a50b448e20c47d4ddfeabb3c7cdb71e0b2c06b6517;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5518d12099303737ccf848fdfb42cd660b5e1844bfa5ddb3709945f936f8449039c2876607a0cdf12520835e90666226235b7b06c99d011b3bfd13376;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75a07d9e79905b53ba36648fc1fb609987428386088b6c54235c3bd380c86b043e1b6a7a69d23dd38a956e3ba24f1784ce0fca1066930eaa3bf3ae43d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1eee1054f0edcec9b6fb87b3dfb0744cf320c1d2d3a9083d95b01a5c0585ab32f4007bbbb1420521aab1b3bc4a170db30602ea2c66c559eefd9882934;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ccea3d37aa73d9b4b2f196b4fb3465de2f29ad08949a1a14598dde8d67c8024524d3af1969e7fff6c1fe7bfee51afa6896bab669ab8702d5466a853;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d68644ead769162524daba4bf1147f87bfe60415f523ca46d27264b47f6fcd7b8fc9cdaf925780bba9cf1bb94f9847e76c766c1993981317fa468912;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d28901fef51959e538d449bc9a9d0d7431cca131187cdd63616ad5488828d399203606c63e896563227cea68ea7588a664710dbb99518a8426ec686e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f352fffe236b29aad768d751597b3a8b9c53fbd6b637528c735db96e10b8278676c9390f862bc06122acc4fae720a608d52725f8205c8d8648e82b1b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd6b1a27ac02cff8212018fc960aa9c0a4b57e1e4f394c53094c9b68790e531c05ce23f0bd17653e171d13a7ff9c5785abd6980fddf5fdd224166a5d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8edd28137d08c903b60d9b649dec8026fc1fc201f85023f616791c28586f1687cb584b838fbf55fa62e4db61c98dd7b8aa3cb9f1a6f1a59d37e5e564;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdffb65d0aa275b89d5c4419dc17ec85b57b832b9010b1e95af07a52c36eb07439aa7b9b863059e2d109671f5a43eb628d70ac716785b5859aec224df8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd921dc0f1f3b5fe088fdcba101d8fff178284ba5c785781195e45e1352a33875e0ded6fef49b5637e3e81a6b9ea559e9826822188034dffaaea0964b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee6214e3c4b240f64edc440a39ae0754c728040e8188e08bcefd66023ba0bfc291d1b521dd4ee9c2f89d2ab8ce4cba81f3ff0708707a33f1909904286;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbc992a9e686d97ba2c5d041a674e7ca94af16f684e96f60c1b7842ad2eea0b23a4c90865771162632dacb3716898fd4159e7cf269e8915a0f6780322;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he44048a341047c9234e8b7957b3f2084ee9c707fc48d568a2e17a5df3868cc51e7ad93ea51b270d419918c0c54886aee67b3e9024cfd2de7a3ea9b5fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8a50b2cefe775d2a1fd78cacfed1f8ff49d2846c2a3116c44b9fe7d638b2cefa36be9485a3a61a509d7ed55692558b5c1cbc9a6311f4748cb2fe34e9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ad1ac6a7cc2d48fb07fdb8007f3870785e090f212b99fd0322e935065fe386e553a148ed1d961e6f0ad04807a9d45cb7ef91b0970541df04f7764317;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f6f5eadfd5107fc7691c355b8c01b4903afa4a4c9a66ad0a58c98ee74bdc26d5d781734528b1b54a8f827c3db74eb09bed86ec7ff66f284e6da318e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14c0e10373e7aad8847ce109b48a82bd5a7b47f8c52390540e1da5ff600dd9ccd8a22d599d7fee68fa30a1335948b4a1773893e7d6481c49bde379a28;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd42e32f3f80b5f57cc2b9a8ae58a66dcb4be779c2cd60adb82214ae3dc337ed4a79496cdccd6026168327aee681688c25fcdade7c7496b43d1fa0b8b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc697c4669920ee37ecc352e05bde4f279d37fe301800a184994c816f6a37ff25ce4f66ca80abc0de19bb13c957b5be308fb8546e8ad487fd58b25e58d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he1722f255457e79ff982c6f0878767edc93abb0eed698420cb95b051c272ec77572e2b06130c0f0a3e58eca0cf7021f5f9d4a086e1d6552368db915d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc334c0ee174c2eaf075bcb941d32fbb96303e28974bb99e339f0e21f9cf25bef1f90ef9299928d6f5f7b0d07750f86aaf9a532e0f2d38db4cf341310b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa2ed1ba1eac63185d87f33212c4fdadc97cf610d74693d8f62ce900d4f401484be6a410321e88211b8a1500702e9f089f8a0898c67312d326da791e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c4eeb75832bd9799d3105eb7f64ccd4e4d26e621be9ff7d4763d69ae714e9bd2e2d8752b9661f92a94eb83a47907e7073ae840dc502d7df2839088d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc96e91e9a7b36d490e01be8bb2cb6b7e0a107ba84af833b1f479a20891d53cf9a33ef3c5350995da6f2985c0613f020311d06b3001fd487c38d949cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h448c91f3d2d458cfd7fda821c3f4af50bccfe0c59c3ab4ddec8d54a595dbae35060c9a5c97d481d598f0a8bae0cd7c28a90e3e9cfc41548aa0b8acae0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heeed17d2dd54edbb7e125b81788103c9c8d1cadaeaab54a35b791ba902d52a60c3031713dc3809e8dea2dd266b82531d67df137a4e345f24a537400e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f8714a8a0a9a7f6f6aefc7b1493910c6fa106e4ef57a28f08f591e44923f027ba45b7a3a716de5c304db98aefbd1225ec24b7c70517c1099fed2deff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31be8985ac615bca6811d6ea2465c93a479d6abb89b7a973583c98aff643996bad130db590e00b8f07e74359e676aa41bccc9a91d60d571bbbc4eaf89;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f051041f11c303bec3f9a7b64272b52c7ff8a000270e7a445acefe01dec4a9ef8af3745fcde069a9e01879f561619e980a43a9ed4d52ba70cce57e3e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h198ee117295f970933963b425fce9022361a5dc0cf71ad4c86d1407451d11aa11f21308334d1a77b73a728744057c6bad1e37bda0202d9117d93cc7a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97ab03d6d7db51480cdfd67e3385dbbc1b0f044cf6dbdffbb2fbcb6041cda0115a8cd2b87ede6e1a78de62c9aa8326472c50ef947d6f522f73c492ca8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91f0b59b6bf8e2b40d8d4f70d6f149ca0dab53be8975a7884c302e5f69dd1c024ffee663a4e9bcdd0fe748920c434c1ac100b57d0ead2a467242af29a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fec6dc3429ba70d160d6abe54c62102ea68865d43af33edb163e4ad11aba15867fe2e421da0e52e353254d406a39b0c0b1f337d673d15785ae82840c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbac32ac744f7b4ab8de486a8d4c9c01a67ebc015321d7b71abbad0a0d18e034395abe99b86a525299710ca0123ab96a6291be94e28273c5e5b93bb770;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb62d32652695d3d1e47ee7c464adc1fa6ca9484ce9b644e412f9482dbf06aedc914d66e99a4dcfd5938d5e6defba99863662c2f118eb9288f5d47c74e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bb0bf1e049539bd22dab074322268610fc396358a017b44b76a01e3ddf63324c3eb031dc1e11b3d480df543ba99d4f41262626ebd14b24932d098b85;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ed8d537f935a9fc386a71b21f7d1362b838e3dff1027542ef6e39ee2dfbc901b0f3b0a5680f7a1c45868c9a01b12ccae7e11aceffda6a45a701b6c1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a01fefdc69c862316317711c84e9541cc0d0366e26e80f92db736a0f6f9aef2c3f1d138b3d14a041d5081cd3b7433c32781c63f917c23040e663deb1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ff0335a002c46a84e46723331567645ca7514d359a814e3f5bc8c02b571c0f35c2279de843fdd3e6081173d94d63ad752c0bb2e54f321a227f8fa972;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48535236b586d1890f8d02a288caa1906545969b46b540598c61bea512e8ddd6a2c0382a668ff782919514264ada8a737ebc1e01f1ad01ff23bfc51f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he98afce9a9b376712ea15e61566fa4175b37d5ff90bab9d12e061ca40b039c973b79bfaf357298c9956066ba33ed76157bec6a0295e11a0ca533c6876;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22a0d71f4c68d6b01c1f667e12875d316112e4f638da2524c7d22ac97f51e369efa03a6dc1e2a78d2e4cc10ffa807a892a3c92f4f3801a51890fce559;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b52dd86596614a751d6109812db15fffa67a14362c986e901ed94f33b9781f356b545d1ac8a29341235bc0c96d4c058377d99dddead171214c7e20fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h880a6923da5d9bb8b97ac712d7a8e3b765546305d983fe60d23d518110be30c01d56d5fe6b5876e0c708916ef4ae8a52e3c7914074f8945dfb6f93e51;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1c19fe6ae898b2c39fee867a51c0d90fe37e1c6559aab6c41a6754ebd2ba1960abf1c6aad9db42c04b8f634be7fe3cdebdc1a3935c18cae029808071;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdfcc3dacb4f1f2db85350c0dd986d02ba00b56a280493c9b710b24ac221e07adbccced525f9bd36ede0eb148b081aa88376b3f019d7f0cd23974ef8fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h750555ea3374fcd2e33fa8bb4bfc73575736099718cb6a39c2437f741a41ec798c425fc1638f194f131d2b58edbeafd544a44412c529842ae9817fbf8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7642c4b75d8d62925592f2b86e306e7e180b082b99404aad4405403f5d2900260acdb43d2ad50f13da9db3408b82f6e559fdffe567430e464dc7f72a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49f6e31e70ccf25c06f0438ff79fb24df317c0479575abfc8574e7911a165d2e129a7dfa3952615165286e76b63d699719c3777f4081e038653e89284;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9e3648969b3a67357e3cabd0eb615f4a0c49073dab87039872d20fe5500ada3998e6d26b353b2fed164af498f29d79657d912df27a3b331589a6c50f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f9e23ddf1bdd47df7b182be8cbc12394b90aa213632789efb5f492fdf777e6c9cdf72a006ee4161c73e58a726a8dfe65aed34da5349bb43b6d8335b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdf90f7566595a999cbc62343ca761806e18609aa6063c634c9df305d910df174220c1c237ed37e4ec58fd6459bcad143cae6f466888dde81102020e2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc42c69d87cb150c1682be487e42ea421694e00740a47cf23ad4bcb3ed2be6a0a0d431f2c94c777c2092227abc6ec3a268ae111ada85c24452479b231;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fb3a1b9267fe60b9d3d00ef30fb056da4e5992d1363d35a09e2eee1e5a6d2d43600dd9b152521f554f26f0fa28f16b10f3df9331bf298b80710b1b85;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc58c3ee87f4c4e52d05e367bae2981d33d5ba2a14ec3b03f76d5fc6a905a30cd649191219210cf73cc9491e7ccab10f0ac53b54511299cc54df0ebf28;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd605ec915dedce43ad6890e1b4dd0040b6631c05e629a209bc0613445c34ab462394ae9784aa6793b4b9c57baf5409824338b911c59501db0cbda8305;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h571a21c8a0c368e2ffe4df8ea7c8d25342e198c7d7d055ecc5e2eee3d8d826be9f44ba93d62fc0a76d7502aa11ed9597e0256e2a61cec19678085adf2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d9555d5844db72649970b0717405236a5e8d5ef0374cdf5265b394d5a1033b5dcc3ea85e7477a2fa3f9d7abcd163500c6463a178a8d981ff061f45e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h169ba790b6c35deeb5e2392ccf69dd792f4bce450299295620923a208beaf16ceee6409269c928225b415f39fd3dff21680e341a97f45a22d5b8390d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefc24f17b96c99d566e1487b0003eaa3903322ae7c2400d3f3beafee96b0a6c7648b2bca223effa7ff731a673ca9fdfbec60f152b9991f5e9d40d658;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha94a3343386bfb242ab494ec782080104c411e3102b9621e6716b62c101d5e8443ce5d2bfa7736d863bae67f9d3337071749aeeddca6804873fafc0ec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3034179a2a2831e38e998be8b1a0e671588c8bdc17854fe8f9f08020ad1dd3567375d37073ff6f8661e0a88382e7483a7b0a75004e210e2ca056058e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67cbd8017c5525c7613de4c043b107d6e3da99491d6cd5b0e0473f48d843449a9c7b5eb8163faab9059b510b7e96fdcff2c82357fb07493393d643b76;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h904446e424647af43a90495e4586190d8b646fb7632d70c7e7d62c582abbe43e8ec58429d2b745d2fcf0578a36c406d977db1efa8a9e9db9f85424a1c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbde550da712ca3464f63ca5aab28ce0f01b30681ff5f86bb59e17eb11231fad1b1243c5f46a4cb2cfd0d2e9a36db8137c5ccc15bc7d378d307b81bbb5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb729a7542ffcde39c14cd56c92e85990d775d7a5a59a85525e18892915cf76bc9e4e9c960e19fd720c0bca6d42847b5cfd662940f3243adf2d138f40;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86ccb716c88e2d616caf4589438276401d5203088621c0f6221d91e8b7b8ef81c46718dca171c3fd5bfa72a7c56c5715ca16467c7a16a03971ea7011c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1db56b54dc7b87181307ecd99248b0f5df79d1b1dc34feb074b53ad9e2b8e8e8637a493690edd22e8641b6446bdb34ac78b967ecae705f96f52bf1ac7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h981b980e5feea4e4e9ee818dfe0aeef6d4405debda4b83df536acde058eead5cd74451a6b298c7fa255c884a007047142df981e27e6b6bc36457a6ffe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9dc3f6eac1ab241e256d545ebf0b89e8a94aa47a13f53ac90aae02e75cb090545e20477f9d1cd9de455fdc6a85e636fabaa3bdbe70402ce8257eb13a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb368fc1072d02d9b5a86e06541dfd2c7e698df7912b3b23abd5b812d4bd10833b7a7420179ea474f07fdff4f9c077f2951b1f3fdb71a4f3aebbd1572;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1eac7537b6d5b8644c859a2253bc1ff840de18d4ef53802d8ca402c96d3b715083850043e6eb1eb1729b1a8deab2e991c964cd5baf0bc8de5090c6a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44755febe9e46329431a4805db65197f375996c934a965de1d04c0550090fe5a1dc18fa9998f746ca2a5ef65589423f65a57759617231a81c791acb36;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc968bf732efb58905cbdb7fd946061bd563f0454b1deb1921bfc2669a8b00a8fb7cf48afd3ae4c59841828a6a63185448b94907d0521903eb951b69fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ef932c2dd8d5ed8762a73eb222aeb3347233ee96e9f23c95f7072dc05f3edde15a821d534054a266e8b8abc975eb91b547193287651f0a021f454506;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h425932529fbeda8dbdcfc22fccc00c44c6c28c223c18353515693df2ed0afd1046ce0a9ecb4476b82390902e2b1d41376a79bd001d791eba5d2c96ef3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b9722a21814e79663c1f6f37b7a7a1ed07876891fb119ec15ec619e149f3d777fde7c9d10fc9b6cc919c611b83df03805b5f65b6222a6c31c88cc673;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h426f8d2ed6d36bedfccdf5475d671aea2991c0a0c32b5fffb0cf3d42e8472b29f1bad67e021923584a3b68aec47a2887f366ff04b5b691a87bc36d07b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34b253313cde2e878ae9c552f5acf3af83032471a7ff43f907f8601891270db4e2dd91e1e72659d2150fb5a29a43cc23207efdf85c53566ec48fcb9a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h632a1f634a5463c6670e26a18bd1434d3f4553fce90622b76c2144cf41dd7294ce7f1163db9366bc3eaa3d1f9f46072809ce0e342b0e3bbfb7e4a1b59;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75b6dd72d18446651b6fd7c04687715bceb6b4121589ac2fcbd680d51ab6979455528ebfd9d43a7ca1b5164cc42b3e739173c7f701334e8174e026751;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc784e29a2bed614563980d81bd0c61a410e614a2c945f21d682bfd3b1b1905bd4e4fa902592dce84474b11eb6f679958acf9d4a2e4015e87acfac9791;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe0c28236cc87f08f090046d2119db9cbb1e1789a2e784b0ab40dd4fb45030579ef7fe314d474c154fc157cc380264af27b58bc229d799eb2d55e7fa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2af91ecd099446ee14a1b5c5c2fb6a435d58782a7d8997212ed54932a7485d2cb6a595732fe9caabbb398b3890b777397f9e86d5cf90bfc45166cff1e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7581ec5ddc6281ddae0d34854b08b0037aa2ddb984c29c9b5595ff5846984297cd6d74c0f8a3439f39f7fed96bb7a6d9639e06698fdddcb4ff3425a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfca8f614caeec3196bd0fbf3db12805185bd65262b7a3af042c6f5dc1eb0bc3645e0e41d754d068deb4de554b95eab84a9772f35ebf49fd1a207ca73e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd78307c8ff4653fabe867890cd07c7b820eae3eb5997393f21a6c7d6d10523aa1c3dfe5f432dcebebc5d35cf15d6aae067d87902becb2c4e2a48edb7e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h552921a48c7b5ac51a8e0c8da09f5142fcc651893c8136128a8d42320dcf93f841fb818e31cc3f6ce549c6b7d3edc5179e9b0ea18aeed5a002f3c4967;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a1d4c1b8a519c001229f8f20cb04aa6ad00e496ad22deea8b924f283dc60a22a4db43ce6d18498dab79e72ebb684df374fcda85d4b65d4f8d7184918;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f8e7850115f59c4c5f8756dac04f70b67c3e529ce3ff1b3a1fecd5a5b731fb48f5e1d397b3645f64b5ebbfa58f1cbbd445c2570945f216134099aba5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b7ed869d07102a243811b748bff80f54cc263011893a2e56574bf6be76bfef73f2f2b011a0a80b3340147ed74f1b078660587a3c4c3a821df3011744;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c8033eae6eaa202174c9ce3c2176baa9a2e03cc76a5e182729690d5c78469058c80b5cf4988d40be86044dc32df3af6e9841ece047b09a4717dc45b1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8ad44a4fe6211809018cc81f349faa811769b0ba3cf7ce2ffe03e7b32558dd44dd2ca08c205e1ac4dde34dda1f3a740b7f72280eb7b72a121a1d03da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h614f51ec88e227f0958cb2c80518761be80e1665e6531693ca1d249e99d4240852e2857033cd5a4745967734b5024dd1d62fdc87f9a8124746ffe324c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fbd4614cf4492d6fa8ebf66eef669b5dd7ba24227af39a1945e5c95e4f49e03a2bc6f084d68fbd1d74a7a03a06163542dd8895ceba1735c5bf9e9d3c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41275945b30c04713100bb4ddcae22967e1f3c768ea7d7703c53655466117d5e4551dfb2d4551934b3bd5c7a7319cc0feddda29f69bdb0912fb3784ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdc2355505c67b1d436968396fc3c8141c86f6a6f2959d850144a67d4311a2e43f27f77d7e5f50ea3783bbdd65d057aac1c81cb412737a29c648493ec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h127b5df693e108bc0b9b4c2ffe067ff6e617abfe00c7d219a4db528c8d1358c92d5db88932c013b2f6e99b085493840911764970750c2fa24679077e4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc421adc0dd61aee9b969ca0bef4476dd88fdb8bb32f63b66ca5cb09971c8b53f58872d24ebfa958f813fce2e653d55d03e5920243ba5a495e367dd17a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he285412b65a7cd6011529779161afd3cfa49978a9d422a777d9a13e028d0fdce757b8d32d4e340723fd9ba7da80cd0ce43801d94519ec31274e77f375;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10ac3b3fe6549602bcee24a597d60b969a4554c44a13f3bdf2709c5f6394551112498227fbe4a36bd6846211e9e5b4083077d7ace2e1ea2acc7a5bb35;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a9fe126d1ccee1de2afe336d6e185524b04d4632f4a4ee0fd7a3213b6e59530806e0c77d5ae68257ab077f3238e6fea32fa0fbb8763b36a3b4f0c309;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd62c8d0a95e4276dd1a06a59a39bbdade5b74e2026f83b42b554d9111ee807d2c2be72c3f668435a132369ab4624c18c3e192caa6b811f906cc948062;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a5131d70616c958df8598655f921e820e3317938fd9ae025efcff8a3992191fb9bbc3104e6340028ec23e17c490076cce6989eafdcfd74a1f4316370;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f485d988b69fa11a2e2f3a50a61862e9d34ce166f7cd5d72714c98b2f2734fcd0b1d8f9b47ecd416cada5d041cfb9576f139c7050ca8d994826255f8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda952a27a2e8eb19f242b547b9b6a3296d422e42dbc90798619376526ffe65f16e224ba16bf08ee0b419c84f4d538d2485cff87961ae977a9e66f8557;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd9220c5c52888d6ad8b0b7770b8570b5b21cdeb8240494e87991cedd3673123c9bad09a0f8abc232696e7130241f99e38af93012c3f3b5b4f59a49ff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd8eb9a905cd78c8c2a883d25d88166badbabfefdcd0e50cc6d6eca2c0701ad3331c02c5aa5686ef5d0062bd1725f043943ee772411685333f0b4f409;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5c93745aa9867169daa3112f74c7e43df9a61c9fa5c23849541f145faa54abe6fd429d2d067079a5b8624f14615b58f9d739c43f024734b277c32341;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9745bf4405a518ce4f64f9ea42ae9a3e62de3aa2132d5ea2358e76b0ef8bfb1a6a4da698996e91971842d59f67a9ee9597fd29514ca9c8def4a290ce9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hecc29a6bad23fa5b5f72c4707372c3244b5cae5917145f422c0e9bd1da1492cea772166658c5caabfe12fe9f96380503cd099121ebee4faf22b3238e2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55092280e34770c8282ac8d400233077737d882365292f9c1db8c5312d057004193bb700bb54e46b7ce2632331f9798693472f12c18f33af51f7dea41;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf228f6037c2c87f3cfd2ab431f222f56bde6de4e6137b646964fc21b1c21d691cea0d2d5917e78567935fc35015264d0aeb6d35f374f1cb43c605f2f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha052a1935e30d509dab57d1260180594ff14b87a411b77c17c9b2706cadcb57c4944ec2a79e5b787da2bf6b55879e410f8851961d0d8171ba2df2312d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h630c265bf9dd5e2a1f2e72500fd049483f7e2efb9572e85cf39343b2b2d2f3c1f552f4601a2fdf46bc656837bf1c7757190c25b7b238471832550431c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8902ed72b38c1e70c2ed1b97ba9540d0c3a355653bd8e5927974271fa70686743c29238698f928e80aa1e6d59ae674e99c2c87fd1f0fb74fd497f1f83;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c099acf4a32d75c26b067db6c8e19d8d1d7d2bef289579a02dc8e6f14fa5c384a74d25cff25b234c18a17b600107ca8facdeded8e6287cc5b64b1b8c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7a7155c279ff270dcc09d1efaca4664a3adc27e4a33ef8f7edb8ee120b97afb333d9df66347d591cc0919dfb7f9191c5747660dadc0bd79fd8d4094;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89f17f7fb36161c1677ca6a3363a5123937cffaeae23785b016618abb1e7aabe7aef5bcf6aa6119a209734d202e05c3a902031df0a8fac52d84f66aa4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d10bfafec64a620f6a456a6a33938e646b41320e5254d771ae7849a7ce853e8d51e87c26895eb9f548444a30d8eb04014969db29cc2582621ffbc2da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha74c5764dd27abb8dbb465bd3763741b360913ee75f23c6fa4a5baa89e97be38aa3969f06993f488b63907e85776a77a4b2dc2558b1ff8a1809b381b6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8592271a681f7edd176b3b2f1dd2ebc0be04f0786a7bbdbb57edb18d1ef18838aec4fe1d8604535d3673975d9a16821c9975a6a4776cd081ee6da14c5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd629d84cead6af026ddeb1595b4ec484d1c1d945da34e2f8509a6ef30b868342f9d298f4d6205fbd0307c8d9129bb68e2ac341d8d8b0ecbb3cf5bb63d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa2bfc16462eec2545b10efbc10bb3721b757ea01356bdf304d8f34da9aeb52c9f1df54ed229da4a49a2482cb49a93b6f3de104281e854d7ea70b90a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49ef6009ba166a2f0edfe816b72e5b7e69e035cc420ecca955469c4db1162d55badd4c5760321b0a8a5c9ac46af879145398488bd629d989baf9f3534;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9196bf34aeb11c829f12fb65dabbd4118883eb6c007193b2347b6ccf46dcf4308d684ebe327c69ffaa583e09886b314190ad4d5e80db2b4a04d6f00ec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h833b576ebfbaf5b624e1b25ebb818ab6a12371ce0858e90e15d898d9dfbe793b0c87c4f72c1e1363e56f245f18e48c9cabc1923bf56f8812d3059095e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43ac32f3366ea1f23b3b6ef687e90aba10a6878f345c0b17998b1e4cb6f0c9a74c29e82ba9b1fe8f31329e9e7869476be469033776e5619dcfaabe0bc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h923e53cf968ae8f240a857043923d28258a751d5ef5e50ca508c4c2cf4ffba5cd50e0804a83aff7aff7b0a5f9ed1f5c64ece2e779a6030fdf57f319ec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14d174c1c2da441bd94bb5e1ebedfe398b3dc9a18bda15884cc7fa95d952f57a30b2a24cb7af1580fbc6875dd28ea97cf9f92632e6e4706835ba1dd09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbaab3773f25869b23b73dae105f0bd15df195c0aea85673a08986a8a57946f5baa0588dc3daedf44917a4d1d0037da093a255a6cbe6f8bc238dae6ea4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7886fcb6f2e100bc1c7c7d6838fefd1650f6c0e96b7871d3ae2ba387c296019158810974472423ca35f5bacb451f8440fcc361af54ba2f5d111ada755;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47a03dd5a32211f42fb9c8bce297cfa7863f8a58e339fe84e2101c722030ce3c2c361c43455db07fe62dd0953973dffbc068425663dcf954c1dfb009;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h938ade23deb1f427efb55e863e66a82f51764a536bf0cdd914103824fa1d13b80d40991c78b551b83b28bb783191118f47bb67c746210f933d2e2f900;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42f0b1885bed42bf3a74c920819468c3cb2db9762374283753a189095bfe5d87d40227095dac2e8e8d0205050f0f558a87d2e6ef4da9ed1b5bb9394eb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51b5fc5001508d23fd3b9f33200286fbcd9a8f68ff4c82ae19aca55efb6f5992e58ba3dae48e1cd486837ba308ea4f1803c44636eb2b4910eb6f9b923;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd8dbe002b1ceceeb1ae2db1214b20a27ba1e0152ddf0d7a1c9d193f4f4f77f07671bf154db75349a8195b2d666470f0fa3041acfcfa90ef1ffae05ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h186f388093f4c93d0b92a2d0ef98ca9ad5465e77eb262f0ec031c1c5f8cf47379814643bc72be4fc65b852d5d82e674fc6dd8e3598e91a47e18e7f426;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4aeac647534a8b27a21b02b38d13aecab511695525e9b0810871a4ae164658e5912d8e45f4314b11c54782dd6487f10a093d57afbceb6d81c743168e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h789b397dc433d920ab98579ab6e3c6f915d96569d4b853433f2006a31671be8b235f5a7f3042da67915a24bace4eb40e39e39782a6e6d92af1062857;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h747d41e15441c29641391348607292a4330228bf7d78a52012b6956f82c623edbe2b3b2e35c143f5fe59bdf8ed7827468fd392e84a3827059cd6863f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc44b79a10e5c1c62274f3037d3813ae1051557b458babadaf7bc15572dccd105f60feaa7101c070592fd1e235fb7d08c424db8a383261b743bc157a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb5f1399295b844dcb24db113f75adbb8d9a45df47405141af4ea581269336474937bee9892fc08fdb653bb268633f003833e894d9a204ebcb50736bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7671e8dd3ec00d3dd89f4cf4f19191a5e114088a69650700b02944c74586c2b257aa16fba2a7fc62e4c98bf7dd4c959b089ae7cd8b04edaf3aceb2cf9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae0a8b24966448272b5aefb8280afcde9e540b5b9d8b1b01cc0db6e273fcc4060e093764f0116f348e79a8befed31c76aeb865b99b3d8ed87450e8253;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h203432cb8e01f581baa94ea7f160ed39ed626542d1aee774134023981c8eadfe92a9528cc5df840bc8b8ee430b7e8de612a314be569457aca86dec80b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5150438bbaad94e78aa08c191dabe9d61190f18a102298ac6e1d03d843c4bbf5ebfc9c9fc6c01fcb0388ed9d87a55f0f6e3573230062e6c73b14c35d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he958687e0596a0c03c6423391818a93146497ce6f45c55ce7d93dcf07cdd993445e078df2dc5b890400d0ca840ef8f6456d00fdc1eb74f314953e82ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd929e840d97d6e38f7a9d3f1616dccd5af411ecb2a15172975d313e421d28e48376735f3ecc156a0aea5c13b39ea3e39d5d0ff2dd234e63587b6383a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a2effed12395f7aef9347692cb3c6007f0f63a84b43d58845b33996301cbdb4eb0169382a46d8b8ba2d32fd0278ed583e8eb8d48db13aac4969127a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61b9feef7eac7dc402a685ef1d08ad1f30253530147d649bd6a3deadec88d60febe52ce0d005ad800897de240624ab427d73f2f80416c2d28180d1561;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69da38cc5c62ee6e94db7134d4cae8240372fc765800844ba1b2d5c2207ff2312d64badc502e941a4206895a67f5be7ca8a834482aa4bc313a799a50c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7f03a8f5ea95db91cbb3b3473ed40fd143e26c70fdafbed34379835e2b01743cb097673652b71737ca88dfc99fb465e7b5f3e628bbc6b175c037a204;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30c13f85e5ffebdd41a1fe5e22e3c93454495af8857f7c768cdecaddf3a7d811853ec1c27978387bac63d39d57ff1293ca22d6e661079a506f55de891;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48685e4333c57c1e1853bd4f5853322c451f5fa311c29e6476177e2543152e2bb90d6dee125d1429d709903eca841998d3a0a65eba6b9db707b98bda2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcbcf7dd5292ad1403e269f7832630916ebb09094dad295b280cab9d5d4da09f50a24a196ce535bca74f72fa9fbfe06e5c7108196eaa1066deccfa5a1b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf617d4929e79057179069d8d1894f353e12aacd4707049052c7193f8b9e3aa3a909a10e651a9e354f08164655593d3133cbca36232d42ddfe0fc6c9e9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e1e91e06bdca4d0a4b42f1e06ca1fb332f5af48aefcf2c508fa5e5c0d782e46fec7e2dc658e0923e46ee1f0da4fd625d87cb37596ff330ef8e55e6ad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8b9eff695a0889a1057ecf5c692fc546bfc31be21f4d78a7f2ebed10b4630030107a3415246e0396225b102b8064d2ca802cb15309c215ea7f45dcc4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7bf7f65f0297fd1f744d0ad2a1025a54d55f77f2099f80b8f8a8613d709d57721bd2ed1f35126727fc0c1594afb40726d59d937123855925be5ff43b0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heca037a0b374b28849a4854f830006739fedc21cefc90aadbbdc675b0dc5effa011706072eb1cab3644640d36e385e234eaf6561c67af17c2d801d993;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac9329c6323334a931acb26a88e48c3bbb666b18dcfd797a33bdb2ebf9eb4100a334e4a72023306fecfbd411e020359b28f921a59f7fa934f0e26e56e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e17b13af8f888c3563a444aefdeaf8c55757104978f3ab5d65b022125a703e10d6e1eec8d78d79055bf661525ac04429123c20239bf6383f9f1f51fa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18aca11bf24092070e0fdd9829fc4cd5efc8b576f8e3bc3fbec100e52da0c3f8a000887745468f0c19431e3590ff283bbb41d7a3ab45472c50734deb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60ebaa1aee37159a8ac0de82acc920dd2b2e00fdfc0178b30a15c70c5e8fe463383ac772cc77c979c0204972eb3108bdb0ddb932103ff2a88d60e80fc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2814d95db2cd91c9a02903864dac974f06f40e8e54584b1edbd52867a5dbd2014d4d01a803752b345fce06ef9211dde852c298af4fc4243d50fa21eea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf91467d58b32a719658ec2a13c6f76b00327425096e7f16666d6865d60304c97fa663d39ee6e6ac2e127b129d6b60af06cca7d56da847397e30a7c50;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b2c1b719aa1b2ed01c4f0d62c677b80967d842b971cc689948348e799646deb7e82ac9bab608b089710ab287b1dc6e991f14a6efd0a5ce96e6b63c02;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e201e02930f87e8ac3802687dca953f7cad55ae24d18c5688600de7de663a3b7f2baa9a084a3b0e8d1f3a89bc68d59e0d4d238b672322e91c78a3941;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0ec2b25c1061f68d60a568c51b601a641d9c2574173c9efd785cec839450a4b52ce1b345113c4ec8dfade37463ee09115d9e77cf001a8fd565ff18fe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1190d73fbeb5362e52e7955d91ff66ae48e5fe3aa71964fb4c1b044ca5adbb2010588a0a2e60f20a555147612153382d68e39928245c917ca9dde4609;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h755906ab6bca76419cf64bab61fc8714ca74dae103f661b2d6dfcc5536c622f8bbddbb1b9064790de5dea1bc689db65190bb65441a8fe34d88d06f505;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98f7499269ea0c225fd4a67990464f406d02ff9f244b575bf47b13f69bae8031935bea7817afb379a42dce751596652c66c770ec73b91951b566cedb0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe4b2f55182c6e71548135753c18047c97f84b592a56d4956ff6695978d52a2753c598228d33a3e1d63e414926900a8b37bc8ea77fdc77ce57e1ddd2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6b13faefa85163180142515395ec53e1c231266b8bf21533fa6f9c0d2968dd9fd234818479d42c2108868c130ec3abd30e8d817b2bdf8705413b73bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4ccd0296918f428692e5a2e875c8485b726dea9fd4f5adeb39efd50eb4ef09fa032a2d9a77c9bb7a5798066a683bcbce6fcf738f1aa86c72fc247e3f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e0b17643e5add396279285524497c158291cc21edef2a9761efe22806420ae8d96721282f63a23de71149f07211d5fe0919822f0b6688b145a64070e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4273cc3844306f2257acde09cd3d190e55e12e2d48a0c48f955f8ff48500732657f8f915ca9462f86364fed7cd933e6e50a52cbccbb8cbddc8131b51c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda8ae5cf12af4e6646492fc86733a7a340046936f49b1ff472c7a0f9d33110cd60af979c2a9dcacb0de8bdbee18b7ab765c289673591c64cad7098580;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he02ea74e52c43aa6f1657e829dfd8f0f6a5a98df6be653bec94c56f1eb677b8f3963c6092ee1dfbf9a3889200d5f558319cb46bb46f444e7fc41a3e8b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha069f6320a023add341ebb93875c41bcefd833e67ba70aab6e892bcef6db9e726545e1f772c42b57a026dc0281d40b9bee20e7e91cb4e0bcd2c6db8d0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h635a53ee17d9b2a2f25c5643cd995f073ac9691ab91fc3fb47ce66802be123688ad5621a08e58fd8e384620ff08535b458a9c2968b9baba7ee8570977;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d3f5cc893eccf715a84af1bb37a9989ec96e979b47312d2904d464b0b2eccd0f02b8df3d494d51654be00573c61870bc75dc3c61fa70e160f47bd0e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b374ef1610d28492ee334d4c93591f457ffa8310496a4c6de051b70f8cf6876d4c2fca376fc28474eb23afae2235dc19d02228cf98fcc820433e7604;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b0dda1e32357d0785b427737b4031fba967919802e608c2cd9a53f6a4cd476908ece1e945e686b28075097fb250f00e81509bc2bb8296c45930e4aa8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hffb9b7994755c91ac90c4c2fdf7ba203033822b1d10fa3246ba86dd68610c5e36789d0e0318e46e0953152b89c8f99860ca22dbb062b2d2a0959d738c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h274e9af7cbf65391cd30029df435b5f2af9f1e849db8b5c443b22ec41ea9582d6224f2ab16a21fe43a5cd115241392930cb3919ae33025f9386dee863;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82639862ce12f7184c164a3d9769f860d8c742b401779aab28173b4d062033a8ee824aa6afc8510e3d6fd504d0ccbf900ad4d7946e6f4528afc54babd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6684bfdee21a0f6096086fbfc71ec4c3c088872cf0aaad3e5feee322f1e26aee8810e1bf21bd171f474d9e2c83c4c4338b3d04e9539e7622e3577ed4e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9c2bdfb93d481690cc002290a3164b9e61a7dfc26d5f1a094a940718255216b10a09ae0e23d6237df4b85d7e3df0c41d4abcabff2026f99ad539baca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74e3a10a248e375f059ed12ab79ed68511e341bcaa2748c2178bae1785803a61e249cdc5e8cd1679f0e9b7ff3461d5be2ed0b8ad21e8d514a9a549cf4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7e751fc68b0decffd5d7b53e53b7acd80effa4008500434d8cb02f76701fe7810ab04ac15908726dc4e94e54bb23e6885d9032769f9cae0a1c81c748;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d3c0419912857902cc21873a3ff23a5a268b734877d84f244dc12c42473cc4ab111953fc5e05c21f7cd780e841217c5059c1eb5dedbb06c88dcae6a2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf377b31663cece0743ce39e21f969085a0a78bc45ccf193679f645ede74660d87d88625bd95cc23415717243792de9ccab057fbd36ab08c2e77dac9bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d5e408030ded7a614c09777bd70dbddc11a5da5961d07b53932b959d40f4b513cf3c59d115b3cba3e345593e4ff2e756b32de1ff0e6d554d3f234e26;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72014261fb3a4306f9e0f22dd93354729bfe74f23a6bc9687a03f2b6f183a264faf8b86b9b7c9e806d608adf11c363f2ace264d3e6314df55897d1c32;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78abf14f4ad8eadd2100ee776f39b09a7b2d7fc15922966dd4a9a36b3ff9e8860ef0f2de70e8d73de1acf172cd552761c93578b652575af8843ebca07;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc868bc08b8d833e6f2f3368bee882e08525b4cc3cce505e6ebd6c9a861afab126a23467652fd7521bc11e463e5650a87f5daacbcad3f43ab4c517f722;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2b62286f710e9e2f9c5b7db76086cf24ef2c9921c7e7444815a218a9a438e9dec841a0ea3ef2eae6ed71613f598e68fc92c9f8e6027b102f5e6d71a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5fc2829fe07f98a63fb5ea441bdc97c372de527c8114c998b90d74a002d60c71456af827b8c64ea84d4bba9635d82256b350e893a39c9fa1bcb201657;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f20a8d79a35e9466b90aca7c62288438772f65e31c8fc395dbe591ff1b2f39ff984999675e72d1cff4978c03ad1000a4ea9e630e4adbd783bd7a193e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5e58d6339d1b49f54a05e78b0034357bc0e44ec12fbb55faa17c794ccac400fb5783da270580d16448ae034857d66dcbc92a8bad93a03fd9a2849ee1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32a73b367cf538d694289182b44a13cb0c1e88cf080bff532e53ea26330a53bc2285adfb92565a21810bd77abe06961111bc5e1a7555ea943179c32f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd666d06e09a51c96dc373c0d9a5653b35dfb9d63695ada255a4017915c2b33fe95a3004d7b211505308976499c1098e6ad39f12ed0d23fb852d21e4b7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b5b6012b7e565fbed92c8fa3a42ca52c7fb8e38dd17462160c314c3e602cba92b3262c1f3952309e414cc839d2a645ac4e4b5ac250c93691fd7920f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68f74744b4596b90c95f2e351e84444902f2196503f030b8251f3b8fd5b0190bf6c6d04f3bf6a67eac96c01f0315f5cc0a1695d48bee093836059708;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb280f142a70363d2917c5c91f110ee0b5202b85883d42caa7b49f995d83b4e02fa46a241f62d1be8b10c1fba1df941366e2695ca47dc97b448ccd5f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c3211ceff436ba1ce967a452c786d4811a0542dab425dcc2f91c2a618b4cba51780cfed011d1dccf4ab7ef80896c0fd4d99a54a45f18ece75c8c2df1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1633f78dc898db3fb80e8a8df4e606ada548d2789ae423ef46274f05789ac3fa7aca4205dc51cbf5b1a9ebfe1cfe6d6112dfd774d5f59e4d7197672d0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h729d95d253b9a66515dd3eafb7e23c8d8668b077d0c7071435e89bf3d1ec7a1ab6a7567b01ff6339428accd21442ea5aa3d1c4a6af0a36fab94fa547;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he43dc813e2a2e901ca484ce8e2de40648251b78b343926eebe1f71358f8ed9c6eb16d27c4edf0fe85990ea34ba9e569e7b99220a71fbf3c0b238c461;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a1890fb93c5c311255079b51d39524b0af8b510c9c26d0e8770176e5bd452be35f141fc02149dc6cc37f69adba56a4a4f32a3c8f573ed922aa5808a5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c2e80b1901977f40ad321acad90a12659389c754b3f325056a150c374a38e12f13525b1a15ff09953d4521f4327607b9b168520de232557463849355;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9be57551bde3d66d810a304bea1d06ca643509e228150cf02db30e1547a80250c587a1800fa51851ed804ffc4c0ecfa57e3a1ec51c268555f3c974bf9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd092eed31ae2e8941c73281bd73d0411ab3b2191abe133dd13ad3f616caafbcac55e44ad79518203760cc1c69f207aa44007221096ab3a4c3d7fbe8a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he1f0e37a507fac17139e83886560c1d4be39763bee64099c7e717143de1dcf28b6ba502139235dbef149019817c59361fb64477d89d3c062fa8cc3c00;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9a1452aaa782783bbb902ac79dd5aee81ba2e176a60945d68c3cfd8de0071de1ce84beb18ca2bda9d012444010429c06ddf871bb3c64980c3eb6ee80;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd62110d31cccbf4b8b62f4f8cef09d1a5bc2ff3fcc4765392c6a383ceb2f81b36187e26771909a63c8f087ecc4ff1bc1ab1c29438a8870bed2d13001d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb62e6c3b07e058a9bd08abf8a255cc9ab1835a9a584086e6a6b31635f523ab110054557b22016dc5278f4690a65136a9a16050e0f54f3c48741f9835d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3ac86cf4821e9dd74f03de83b4dcb769961df297bebe902904bc41dd20ed34e2c5ed530e69af4fa7d4ef189de1a621aea9ee0657dc9364916d694c1b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdb5f154fa002446a15c7440cc750f28e8f9a5391217dd255e456c6922cd7b3a4b5bcabae9a7cc6b843821eab910da62d5101bb9f9f666d99bf8c27ec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d37f97cf116e9e6a510ed0834cb6731a55d2937ef0a4ccf01a554808a10a9fcb2be93915899996c68c3226257c562f7f4c19c870ae22a7ebf8d6a111;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h450bfeaeb3e0d697c8f2fcebbd4dfbf635e18a0df6282c6f5d7ab698ae637b2dd17e63a410a2c89c7fb67434d5f8f4777b97e11e89cd53bf4a68e0ef1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95e45cae45166e1125257220fe169853489342e6b4edabfcf7dd81d1866f3b4f03bb513b57ef992fde16e25e952a06284783c9b706b2dcc99f8751452;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ff3932ece29fdb3549662238e6ec37514c1ddd9649b4018c25b3f443fcdad5bad4791e894c04410fca71588fc3dba6d0e83893953039f31aebd6b85e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc87c4d4543cde67f419864b66dd6a4d24f4962b4c68343bdc55ede892eb2814ff9ac586fe94b46da8c62582a17599ddf174829ecd32540334aaabaa60;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd95ea2acd9cebeeb791e927f57719dee489b3ef0723164afbcb8e221662e988bccf667b8e6eb47d1b42d76f9ff9e09106a6a1326a698537e128186c8f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e98f320979e3d0fb19e3f1bcee433b69178b372b4428154e821b1ed4156f6c4ef4dea3b91a82ee114303c08d7458c6b254621b69d4c6faa5de6c9d3c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2fb709785beecc69e3aaa7676c71c66b72c1b68ce985ac98d9c05c21673534df11b168d844eb422b6ffec321b628d3a01bfcd0e60d0ec160f8dd043a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h749b8fa4401d1e1e37107ebae7e582be6d5807ef32ae893d4199048f3d515988e9f4ac837f71ce8f0c7d157ba2ae34d1356e3455fcee966f5156d06b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11288d330e990e94327818dbc8bc4c94480b385f72012f8145325becbd7051e7d2923455659cec33c511895341eb0ce6c7ea0ad75a42043cf1a258197;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40b6e83b7f705aa6ae1a539eedc4c408f8f844ac3e93a929eab686c5734b1d80e8a86045ce3380208cb2e53eed6bab5c042e2de44a5f90f0a44e338c8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5ff3f4266f748a4cf74b6607b199132d9f6224245eb243d460005153ae5fb6fa1713dac2cd6503fa60803e7f9480be3a96841c8b53ebd49cccf8b61c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f8ad784a5c7b658f63ef5e86cb4fb57330ea359b5c923cb2bdb257f0759eed3f2312ca8adef799e5d3ccaadc135bf8d3ab181f73d725ce9ecea332cb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5bfe6e9b707b5dc2e1dcd3815747685d135155f456c1a4684b24c1a8b5cd667abb3996699e6892026ee37c5d0131d8ade25488746860c7571310822f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc97812c32fc3ff16ee7fa0670d874739719900c75bc79c6d9537c9fa98c7e642ba65efe7a9b7d5a4ecf1412d50f8d8cff16ffc40981bfdee101bc3c75;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5b0c9abe415628ebea042a83e13d718556c5a79308869935d2aaee26c21a3d5b21c5bbdea69a7c78ec6e07eb7b223ccc0a2cb2be4ad96effa3f97bc1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9594e862a760d42cb74a3279ac170f7cf050df152d2aeb1a35f99e807828cc4a7ce9464532963155f4fc103ce37bbbd63e1255d993de4a7aa4eaee098;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a8fd58f188f16f402228ad832ede018e8b2684058152c74cb7a682eddfc4b6f2f214e7232dcf7ec0fa55888219d05d3c8eb6358ee0a6d63563e0af97;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h906671c57747ecfcbd5e910e97a635565ed68cec473f27d8349adcf6241816e8a9acd5ada3928fdc7fb9b394a2462122d5701034d6c8bb9270fbd4606;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h243387edd14a230828e712b4a316bd811b6015c55ebd40eb59dd0327d8ec7ebf2ead7476a00d3f0501ba8a77aa725c59f6434833b7dac6b2bec48aed1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d5a903342cc31ca31892bd99aefb4712b71ae1f8077763a0912c2ee673d9b6ed46eb4efd2c17b40192f99ad9fdce0e885e8b1ff8e5c71a058ceeccdd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42ab372e8209993a0eab148587bf0c0f89b5f1caad58553c6ed053a373239caf1e0447e911f37c5f0ccb375c1059ce66eb1201345c96e80c46077daaf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8aa23932d94ef3b3877d68b6f3b5960880e0924187fb88bca7f20a6ba7e676b9068ad2dd7b7e8f8cdbed7ffe2a7ffac3992fb1a01250a3b2e4c4d801;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79b0f1a348cb4cc1da8792a8709de27915fdedf81ec71699e01d266e5c601d977857f7e948f958e481ae645f46757a295ee31ee572c7306c868367cb3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e11acc5569166bd1f254c16ab2642a5fa2411048fb8a9a9597e601482eead837c7292dbf52f6996aec7a54d3591adf09c2fa75abe32f0549e109e9a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe7749ead4b7a99740c16e2d0e99fc5dad86de5676bb2da3bd49829936d068ef0ee69d7f2e92e9fb7105d5d58356303abf4690122884cb7d9bd73dd23;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9323e658b97a7e0637231abd0e0a7201c0a96cc94b0df2ddb944b8b7b8c97fe21305d84605dd5813a6968393ba6de3e17fab2bb0c684c864b24a6a2a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38593bc4411d325d537dff9ece3d6b91ee892fc8b06a44399ed0a79e94137f7ffb943e8c5eb6b55dbeaee8bd0b945e556ec7febd1d635af4b86d5c8af;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac3782cb00f60b682f7c8f354957804f7eafb71760aacb1143a04fea727a59e466cb320611507b7581c5fce5498a66ee2b09e61c8c540a91cb23553f9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97bb06d1949250fa3be1a5e1fefd0c2778075f91f900e0daf9c82061b8a5f89e3de69ee583ab24b63c30f338d5e56f98acedfdec891ba8de068783f00;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5c93a68086830f3a49ce83cfc7a5112d1f32b2511dfc90a8b7a325219cfeba419bab6c80a5614aa777e731f3dfbc833fd1069bdcad6466b8b540fb26;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8cb1a04363417a18f6db824001cd53add209b1bb358d3ebfba8bad669b5479f5ce5504ffde88ae987950c668e3ecc1d8320d2c95a1fc62ddac66664f4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h257ee28d9f785a2b6d7201588aad1736b8518d6cfb4b112eaa4ed06679322ebd05c9d70f33a6231c69c5a981eb899466d997c7dc4259f6be4628b13d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e28548150d4a7f27189ec9de56a1928412a4ce38b3a606a7344822aadc95a0ee497d874f2efbd3bc749cfa29c3b9dd2aa20f7151c7600c773cfbfa66;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9ecf05fc688d546b6ac3a33e29b1af4afb51257356d6640f7ae1937c23097a6263dff3b1b136f8d047b1a87a62820f718d0cc8d647493aafd21aed47;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5635d5b683cac6ecd6b16f5100203f3e6a22b479b214a2c508d3bdc288da364ef7804d13f406d0ec974c5bdfb40d650dec6d2176b7d32086a93b82044;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h490cc13f5416ed89bfc47224dea01c5e77ac680996700ff866d4c79cf0c4c36da2b3182080fe0cab9dfcd32af117dca23b41962987c806563baa6a242;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f3df1737a9ec7dd6581c25eb54dbf1da3f1eeeac698c7d77f98cf7d2e425e318455bdbcd7afef8ea938dc6a60ce0159cde25fdd1532c78efc3d78018;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd2dfd06af44f728747d076a47d99e78d45dee38a222fc744507f44b9264f5dc1c5c59b9294fa35a874d890cfffb5409404362fc90d39ee9d3adfe224;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b9bd75dd3bd63f7d5a72bcb3c4adeb8796abc1ee8f6f7e32856da449d4ed2d55ef673412f6403588fabe16298e59a34d7336e04a7707802bb744917c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f6a7ff0c58a65b7c12259be29566f9d8c21f295482c7b24c956e7807e373630bba4a05b1f2492822051760e773e095df4db196ecf8c1f0a94e534942;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68aa248b236dde926c6f39d3d4746cd8819e8731e578da7f8c1ca94124c0d78981cadba0f28519fb17e8e1bae533676c10a5f195f9b3f434aa1e09871;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2420f6cb462336bb3398aefb1c411f24d746c9f5049eea5af658260aad0a8a5ae878b04aef47a3a0c24912e93aabd2735c3a56971846bdfd470030c7c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b9f80beb0e414a91637765d714fa81ad330078324dfac766368cd704d79421e49d1d63166a155aa9b9ee9a0f9dfe1b2c43d7524df464bc191070687b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe764c10dc7d72463fc243bf1a4027023b8b1ba46696e0082e182160533dd01eea857cc6340874ec5df0e5b5c47f5786457eb9376724dd76036047b14;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4565f327f09014194c09b4457f50f47b05c3313216de72de42920b52d288e665eaf0b180c9d0a71ce3a1a2a7ae07dbbea3483422a70ed6afa5c3162fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h506fb8d8d26408230862d28e09dff71c83099e7fb127d62262f1153a09f67060d2fa010e9e36e576e4936c99886915bc2db23ccbcf32d2b4824758f26;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bff88329f2ba69822e482de67173cd15581cf25957c784448d6bd3779c03a6a3266f85349cdfe170348e8c2576e5de7fdb53d7ebfbe49e5e6f03d20;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h424bb8d74f06fef56abc6b96bd2ca4c04e3938494584ad4fd178a2be9a2455dc8434dfe19526c5f1b545fcc870f26af2f67eef0d9ac8ec04d5f41d56b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bb6f695554f59a2716f91d24071ae459cb91ca12675009d04a4e63e105b9c0c4287bd329081f2e79e7e8d5abf0efc88ae6f80da180031d65b9ab97d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7c305b81e94f6fa7ff48c185358c80a0d522bef2e4e6b0fc4b607b481c3e584356ab2b780610a6c1bb12d51109e035b588337c90bec3f080c0718e99;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ac5b822ecebac2b643b88d7daf4b7efea05b5b9db55d71ae8ee803d62a3e348d4f2b45104a3a081ae30849446bae4e8bd807929ca44cb435789c2f13;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c61b1fb05b5e4001c1936a802126723712a20c21a6ce17b11a2d5975c92e27e544102a0ad95aebef3c9c77305555eddd164591947dc09d48016eddb3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45b131bade92f717147b615394e3c23e5a5d693b2376bd2c8f2e1075027cab08ce7aa07950c3f5d582f2b73477afa21ce6805129b4edc64d62a982bd5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a7b5f32c61757f6ee6bd9f55394d539f9c60417735463adb2b6d2eb10fd8e8854892bb4266f182823462d7e18ed84e8fa382179f4a09dbb95f2380a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0eebc8dc20fe86286855cf79e8e9a6d024444db48ba87d5792370c632f8953a12942cd56474e3540a00eeea6cb2beacd9648b02f6dce1f441f50616a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cd20cf9445f27f20bd47c0c454b82fa5674c3b3d843b0a92c3fb3e27fceadbe9887f5fed7ae42371fad2fb5ab9b4bbbf40439471fc76331fd1d0780;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf29d3f3671cb95ad656195c6b3231a5497f3ce16aa9df2cd1a7bb9da3fa1017bf9c10e874fbba15e4e0e997eba7072c95ce7713dd5bc8d09bfab75157;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91ee071415d1c4592a1bfa497d289b83f7febc88402d433aa394651718e0b20a1f6bcfaf4b2658c1b77c4ccc83d642332fe40763caa4c732cb1209992;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'head0abd6fae5dd227ffec5367c308d5127768023ebc6c7756918126d7a312defb026c68e797c3a9377ef34ff70ec34bee06b4bef4eeed8c41099005b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6eba4f2c0bf875570d5df75b090016a49f3835401a2af284ab7469cd9ceaa0aa5d1d1c31ecc7c215db0773be207b1c4df6f635e099177122ca419c730;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he40e04544f648264b59779c2c3f841c7aa30ad1f217f14090932b2dbeaba1218d34709c1688feae59b91c054ebce9d9a534f093319ee7de93732fecb5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he674a569a348f48062ebd2f91686b3b96bac51ff9958098d8519738cfb9b47d469939ef004518072eaa1ffddc5ebc348e6f415a6facb8c2fa961cb1fe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h673e7df62ac62645e38c5857e19ca86175d1ca8b29c20b9f3ff8ddcfc617a3054a161fdae7d233746e7e6fc48883debf8d8b9851636b2e41ff18bafa1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ef9fe8e55847ba91c4cc9fe17852cbc0df1a5c4c474e22e9012a6230e00c87e53c87e7234c3992efab6e19591bf5c2a7d592152aaacaa32199be4812;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50f631b54a8e7f7818760365bdd7a1891f39261020a9aac483f06b6be8588ac1bba5a967ca799438992fd81d565193004dc3561b26be5609393c8e5ff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ff190c43f20d0ca6e0d40cd7208ab31dbf12b828d109ee7b997c658aa4553dab61a9151ac984ac4b2d79eaa3b3a5e2c983f865f943c082d91695c8b0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e498b68188a42d74f6abc2414e2f5c3922024c353767255b3cf5526c08a023e7c654e4f134199364a2893b86a69a8c9ab21017688287a6b7b403b493;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae3ce3d64f76302cc7178de17be0b8d9f494739eec303f61fe7f18211a1273f8dcea4183e2bb3e76ed277fbb1a4840ac8a9c42d6e2b1248a34750c8dd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h746cb2106f89cc4fed726dec7d71116d684e2fbe2279e8c7916462d657d8b93b01c1ca81b81a04b65540ead17632e67fedd35d69f91c4bc3754c25706;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d7a3d868e18544a4bf6258650936a7b49b89c62b19d1031fcd08709f42c78b8ff1779be94b4433b3caf9059a5b150369be813cd3abf402247931c95f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9c2d0988189ea23ae30abe01d4d69649f1bbf3715b29bad782f6c6343315808bef26b8ef7ca3582b7b4cdab4fe508f2201c05e00aae776499b549d51;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd89e1376ef4f88e7840b8634e647933ec9430f3013c5750e090bf8dca4efdc7c954b6736c5d96cf73ddcfcf92e333598b95023a753cbf74466baa05;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hacee1db67ff5fb2f872f55617cd1b6e597155c93b43a5c37b56a66fc6b95f1b30aba804970d1657fc423573358abb96a3b4d1a608d25ce721faab3fb5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h678b232e9dc4588944cff165f42e969db7f4701c028d00db3fdd7da1a92109a85edb0297c3ac593cc02d71283d63a89a700dfee9a9b7efaa282b889eb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5cc84eff8c8cdba54d708c5c9a791d304819107539d825496b6d336e7c69a1c9681c23daf8d7f293d65b7040659deae6d60dc4d7eba7dbbb133f1b31;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28015aeebc6341a5bf070a31c886ebe7a50bffe86ad5363d1d00ab87b9976297860a5de400bf5b154d9868f0ea3d04070f24b88cbaebe2cac3106f89f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h552303157056b5d35ba5cc393fe2c320a9898695ad3f9c1cd1c6bab4b6f2ee5969a17be45de1b43576053ae05be247af8c77bb9ce9c6db4808ea894fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9742bc7b89ad575aad591b8e1d940fb19cbda7465ecbf8bb53a3c5fe3c929c33f2d793f317bd6efebd9197b06a924f012ea65801c9f9241131e5ef8e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0297f8abbfb84053b46a97cd215096c3338f61575ae4d102e3e10b7e2f4364d18a8cf9dfec6cdb9f99162a5d3733cfe775ad47c30ad25ab2fdd49491;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9268c04b7aad69d1faf3cf74c1c4036393ceccb950d5c76e1a737a588d22d46f5a4fcd45fd929e57f9984bdad16ca98e2dab03204e0912c123ac33631;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf56d079c9576028b2fa9aae9189b73e9874c1873947b9f1be019c3b2b4775b22a6312946afc6da34f3e85a3904692aefc34693c5220377d12c1d42daf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9c894247efa24cfd90955a0c075b61d7e63c3444d60fdf0b64f0ab869f671b08bef6a77593bd1c2778df9986dc83c9b809b326943fbb5e55d4b4a79b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h145a9a448a545610f3c511e3dde9097ec72d85e9ef2091f3a518b8934810395dcdd1ba330618c717676224538029a81bcd2571ba5ee1cd945ea0d7610;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab95532a541af28b3c6a0da008170139234aa02b18beaa7d72ecd4dbe57621d1c6c21da65cf03dbbe31e18cd7dbdccb842e4af63f385fb8af356f2767;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55566bfd658feb946c8619cf8ff0ba4c59e96e27d13cafe9fa19ac83668fe1d0b580a41acc805948996179bc756fb82166222eae2afa083ee585417d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83b776eaeefe185127a596d5e5c1f392aedf72cd1cb3d95f8a3387c287dc79e2555c3b004bb8e97d82e003de19001db04891b0256070b2dd01bd57477;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb82be1f35e76e23085328c01e977763955f9c39c08c1f4412d5bd62c7370515ed8217bb0713a2aa704b2be3e25c19be67c617d38b3af5ec046b597b2d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b9b64e04d99bf3ee284b6b875fa80d8578f58cd40f9ee4f115ac36e71a8086809f95f2e15021e1bc3748aef249a128148db733ca0d1d21ba3cc06439;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1231aeb462ea0997bc32dfb6602c8833d7c47e7e53ea659f2f86ccf8461bc576907e45d1d230b7682c054902cfb118db117619e7f1ba3dfded048adf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h492514c9282e0e65c74e6e5b315b66ce92f530b0b85c779326bef3ffee1e8bbc4ed35a9e88112f05b421df93180b709b2737c9dbf35918c1708301db8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h201266255c9b459bfcb84469ae8be3850caea97b1f3a511680d06be8eb62acc426418ad145eb479b0cae9e0c517aa24cd50d20e0301816039a4fa803b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82524596a652b69b0d463d7cc2a371fd98ce40d0b1d4c0507f3f334c5da477b701cd4b8f3cdc81435413fa9290243e2556b3720605015986217782a1e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hadd4207fc3af7720a3f85ba9d908918ba48026cedd8a2fd606ed2a5d239cd89614f1460afe7af743bb07aecef909cc32145f24a99d5198f732d1bb901;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1880268df4dda6030bf5db2df412b7b5a8eca68dd75d9ae0c2e20a63cc9d095a3a6dff0b81e7c3d460d2207a90f61604425975876349b7448f62e6c98;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c0fd182ab0b8f2cb2258f9630e7ff5f24b2a25219d76001be26884d9fc86773189b0b76dbf3f6e01eda772e0cb893f0ee2585d3f6442876f27144a7a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87c7e9864cf4eb80a4aae967bea5d5f85fea42ef83afdd9fc76aac7c6b5988958e1b0b89fd47e2005d804a0dec12c010353be9efce9d278354731417e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had7c4d7f39c5fc4aef6067a6de9df5156bdd2fe136982ebd998e427660c16d9adc0c21c15136a53d6b1c08ce31b490ac5c24a459df0e5f1e4d620aa2e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ffb0e11feac5b774bcd1ad6250f4e159a3cd83b057787a16f905aa0895680f66531e3769923cdb4fe8b60b3651686a1ad7689e8bebadd7b9045aea71;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he072ae1be4be5d9d170d68803f0e4e03f3a6da6e685a9ec5b9f4525f6f02b325a39ebadffd3dc86cf47286a84e77ea4f98146d9d2da7b0ac330cbd08a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha58793b51fc59251345ec5d071704bfa99e0a4411da723b341e2d9f3512a4cddb7481a0f10cda0d03209bc7e100a2ea9b4f29230c07e472ac6bee0962;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6310160f04bb9cdc2b5dc5bc3181e6ac37f31a9e234d7ea5755b4d544b23275930af9c7532cead6e746908841445a26cbe4a41838f08d7990f4aa153;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f6b4d0d292af52cbcd9c4c48fbf0f9441659c9cf35941bd2a03216c04d6307c199b1f70f2010cea8a43b57b9621f54eb1a26cd3b3cfb27d5e909f440;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf901245271122e2a6e89474d39e2d2c7c49ac671b6539af79aa234b8cd22cee3d5ad2fbf2daac706c4ac67f86082a268a8827ba5c1c9fe1e92b6a01c9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdb63d0e4857fe8d361fca3f87627de47d50fa5e2cacb7b142ea7bdf0aee054b1a3f3564b425da7aa79260f012564810250a7d45f61b03c472a119284;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf006b4c2b1c921edd889c9c9385c2a91df0c666baabfc7672e0bd1ed0906910067c5c26b65c5c782ad063a2866c0e23b13ea956cd004a2e66d53490dd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78fe4daa3609b61c2117d0f5954d096feca6fade4bf67ba69e609d8cd235104d0d2f3c0e28b6d0997164d8b9ccc5a23ccd2376b2cdb470a74ced3a89a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c0ebdc893c70c3375170d05373823216f02e65a2a91b4d416f957d099ce802d402bf4b3c66fcf69b9c360e2464fe5e8c2c102c0b501875e1df4e70c5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3eb60fa1e17648fceca8c8d08a038a65a1e5fca5e17831a408164c5a394f5aaa699d19c02eaab2517ede68bb718e643f1c18d01836d46637dc359f525;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcab23d5a56a520a130db874306daf584827a1573861391a5eeff5775f95ab6a298ad0b60025ba978d9978ab31d6db53d15c8fbaf8d87d9a007263128c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9666add16826ccf1a0b1139b8fb960f665d31a5da38e8ab113abe7dcfaa2ce194f576c3ed788ee79e3c2e22ff273c2b90fcede2d6f4be10bec207babd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0753928712b8cc2e8ee11a874c15df9da756436e5f95551a874127bf365efc69c89eac9c41cc66c37fc025c41a96f6699c47a42fd57a5fa0b2274ccc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc329f427697d4f37807a8ee8f539ff4ebc40e5e081715c0daadc943cfbf88d473a33e23d72dfc602fd7c8a074fca03c8ab4b58e37d2eb2fdd98b12ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h586d354b1612dd783feabe7648d520c28333ab9febcd0fb2a03ac07e1c75e9cff307ca1e6812891fd8885abce174374d55180d1e8002475a7f29371db;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4125dbe57ecaa099a46b8e29485e3f4c7bc0539591335dc089af2416e240844f7b5a0c7288a59eff6fec014c3f44abbd35a4465fe46a5dfa900212b9e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c4b6eaeaad7f8576bce309131bee600ab5239b00ccde3416a119e3e774cfd58fdb47744b41e52eed0036ee40f2e50ee64e478f955b292e49bb21c76b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4134ee097004fbc5c15b0df010511e92cbb742ff21386c64c97eb9aaa32311e7f9cccb3e264036601d8005ecbc77f6cf984b6e1584b99ad6e120e9878;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8c4dcef18c875a4681bcbe19a7be7a4ddf27adaf6aae8467b9c9bef3aab5f38744cb8d76cfa6f3e766fc8c2bb145963592eb6b5612e67b9c9a1f22fa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4705d70145dfa9a9572c1a8377ce2cf794cc1fb6f99af717a489870fa275f855c36957065d071b54856daa363f248e80122c5cc5e8602bf24d63b3469;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h255e9fa7d1350b1ca55ad0ff034c713c5f2eb6902c60bce4db1d93227f3e2bae28a0a075ebb1b73b1956f1b78cec17c7332a6caf1918e890a449317b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45dba7771355ec9cc1c50bf79ab454d1b18fde8faf5e4a728c284aa3ed6d42c07878a5f6cd24e81a8f0cb634bdc41c5e514a75d0d4fbfdbfb11dd7f59;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d831647f07675a069a5d5213a1edecfc1c30552eb91ec7ae014f07c5848334a851ab16897227d8018f25d7708ff8462d15a205a8f1da28bdccbfe6ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h550e4bb3d864b861f82b07c92b21a59fe937a86d55b14b367520478fa93c454477413ff84f0b53ffa6efbf9b634af38a32e0173ad94828b1bd6121ef3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he816176f73775b6305447e54e8482afbe578e7c06e046686941d8f562b591d62231f9b74f537aa3dc630446ba27c98315e8940669d8614df25ae32c4f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f86002e84772bc64711a6c458e5cbea81926fe971423fe4f6382a2d39b8d1b723d0a9a27c107155e011877479c637ad58c0bc614bd9fff5380c8ffce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9f22851e1814d23ce064d640419614c42791a3dbf7a2828522207311a2cd44c81d9318008e473e6105671cb11397ecda29efc8711efe9b0178bd4dfe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7b98abf8babdf60ff3cc5c828dfc27d5380c856b1fc844963b6d703e3cefc09ae79836fe7a3cfff433a19322f7a0b566c783eaa13cf99a572be390bd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26f42cd226e56e68f556c350c4e5d0db63509d5cb9f82e8e5707030cd4cc07f879d09588d3e05233c2f3c2a637ff6da459fb45830fc2eb80b94c574d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2aa4f6d94d1c56c01676394abd965dca80278bdb77681ca0872fedda48ff32b3085a3e87afff2be7e9eb2f77bd9cc5262427f6a28b3f5ac82a67bba0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a4a358da476a770688d5b51940ee5b543ea8c69fb9b85c8a0aa110b4f09f5e7f50cda2b16bf033601214863108fd43425625b9e62b4fa4cffdf842f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ce4725a5b4bc28fd1906666b17cc202b1c1a4cc1d855da07c930d817f7c614c35cd24bfd896ee4f8b6522f1b3f70ead62e6b268d1d766cc9c8acb915;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he91d13eb55f464e2d3bc322b7e56f02aa400585e250d709431d87b78191e8a1258ec8eca070cdf92c6ccbacab1eb1f29666caa1835b73ed5cded93e39;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb1a2992560f2388cd0ade7276b406b67def087eede11d7811f67d1c62a1739748ce02e2473fe3ffbf9b823a10c6c84695279f220481d180dbfade8c5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b46411bf92d24e8e2b2cfa89c714c12470e539f5c5c8c4d23004c8e0fad63b9969b5efc03660c1acbbdf21acf6d9d410389f75485b1b3f0ef9e66be7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf304db97e2d47f7c455be079477bced75407bd0f03fac9a796481e1fe5bce0425ec13ff56d3fc1052499f6e9eede9d9533212561eb973d84d148a46ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd0147b6246a2f1088bfc0debae50325807731f3d0b0fe220c31b3410d0a952effc52545f6ec1d40494301cbca464c4cc7b7e0fb3feb87b06eb82650e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd4ffbb3989d421ad1acbe0f342db8b9102e211e65ff93d8e8e2b68cc791f6cf0edca84f71ed353deb4175d7ea5240845459123b871832a35e3e6d000;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6390b48d11a0ab7dda25f2cc6a36f1b8a27b9ef22160226e634f3011851010a86785488558a5cc1ff69d1af9c2cebe4c0370028a844db6b4b885f8fcc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3474cef6dfbb65fcff714eca5ec21ebe2e486c711c564a43764030d10991effca1fdb8b3e3ca270c30d1ebb4d72273ab9ac6a6f4ee0b2ea8764c7df1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b7d52352dbb6ac8ee0c0146eb5ef89e0b4175476b8fbd6b09a583b5cdbbefb2847cc7b0d112349296f361d3ddcf107c4be84e048cdc7d2a4052c36de;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h151fe265cbff5bc7a5644866ead02b06f7f16868b8c50b84c56b07f2674c7e35d5a281c44b170567e6859136b81ba8d3628c460f07ddca0ad4fc4d5a2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h156ff7911cef99d51ce00b59e260aff29791eab67738a6b886e775c6ee9e9658623b636175d14dda337b3d5f34302da7745c87d9ead5b9005256856c2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha65d515dd6531b9b03b40b7b5c3a0ed8b4e746b3af6757ac741b962f2f7a6e15749936cdc184c3734268118447678d6da45ead1b574705e3ec0919b0b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h382b063938f9f6fff2f658f66698cecf577e4b768657bd2ae6c382925dd2819a720ec18a8d430084113b28740c11a72601a8dc2a14c36b29d270556fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc386980d81d4b66859a306675d111b8e7aa52d6223cb977e9b4c2b6f5b77525bae40081b7da242977fc0e75843803f7d9ad081f7cc0a9e258d714d3e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca861b2cdd052620257ecdd00a053fa59e5c5f4eb4bc34fedbcf27f01af0f302e3bd5adb5c2d8ef41992b4dfcb00942c687653d0756d753d47b7c3d52;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5826337ba71349433be48b2a49c641a4cc7e446ab76531e80911a8b5f28048f726969122ec9faa37e9c8c3c7ead4c54130ebbeffd7d2044151402718d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h639f212a6893e99a544c1de9680e2dadba0f60f7db1bb812212dd9763e31a26f9ab2d1eea1eabaf5d4d92d68ba84b05494e15612cba37a7b9ad3184e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f0aee890f4768ddb7c991d8ac9d4f65d53425a3b7f4544461799a2ed4ddf8f8398ea5a7c91d0fffd226b5e712d02dd76fc787636b3b8cd223cc1b5a4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7a46e42adb2b68674a64b46d47c4e5d9538ce6bdc927aa0978246beeebc0e57337440c9f919c2b43ae824dbef2f9393d9bb78b455a3da55d094a46b1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf25c326bf46e0d1cbb818c32b6c088bbffb76d1df7967cddaadf31ec49f5aa5467b9c41bef1e7b595f4b6d36f562459096645f7ff5850825d38d13899;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd679c7cf9b95f63e6234e3bf19a11f194e277b1203231f932432d03f557e81109ab7e70e532e76f122a1af0881faf6076cda2f893d2ba2b3396a7846;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3eec5916e9294f9a4ba4691ed19cc950e1fa021e9650e66374044264436b4438f6c87b15daef1da8b6fd2fd63344c9b4d07dee7d150f09a3e70bb83f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99fda35d4c3ceeffcfb7d3ac62f5b1e795516367fff5a6502e058d2cca332a2455b9f76b803e69d0ee5b847b5d37e219d4de3bb77e67cfd762e40d5d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7677ec9d735fc4f715a89b971937cf9be05bab1ae14fbd40fa5470fd393cb7d22d8381b893312a00374330be2f497ceb2d513cff5e8af4d0d0f33b389;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7520cff73bf9421cfb29643e345ce38c2deb22e1ea82019f748e6b0ffd3062faeb854f32df280e3753f865000ec30ba8d0917312c7d0e450f15c1a990;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6cc833c10df07f711f58bf09f7b4b29f0dc69c37d85ba8dcf7a51e63107363864785e229df748806dffcc956a59b2c017678316472e1c95a3ced8c72;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd2469ffe9a616e2e493c939c80bff27697eca9798eed2861c76d3d7e6354f56e705ff7a03d586d3a4229f43b80b2301d3bd80ad85f9d27722dfc3eeb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b5a81d2df4bce36c371cd3430c85e3f534e62293841e4131188fd1753620ccf46031fe116263a6d8104fbe0dd6ce03e6290ee1f632c9581b2929dec5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h840178dfac1659b6049b4e193eea3b1ef1e7e11fdc1ac1556a16224c30b30f362e8b103d70f997bf53139161e7a06b24f0bece174c84f22c3fc8d0e79;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcaf729114a9f8610975d10c4ed1d37eafc04ec8d4e7b55ab4611092fc3fdc57f748160798030962a87e4137e46dc605b38b6ff5df6660a81a00142819;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb669f3c4c6c586ae4886fa13cef792ffb938d1bfa7955420b173a963cbfe28c7cc3330720f3bc260cf8ce2d8271f7060d70bbf57ad5da2cb63fc24b09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf85bf501c0544be99828f0173b1b3a2e6e11d48c4e206bd0965278bc1dee557becf774183c2dcc17bbd46e8f12dca8570bff6cf950e30c927774dfa1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba48cce823b51250aacfb758d3b32bc4a60e951adcfccadc0286faed5247ddb3207ceb27319614aee038a4889fbd16a3e301b758623b5e09539e487b1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf40d26dfb4b3f77f7c5b5e8e0dfb57660010f47491b66cffc40fe0a7db1a439684a6ed2c78c1982c9934e48dea8e252dea45a3b10376db5e10d20533e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92c9b31159e60fa496b679b32caddf3cf79edeaae359215e85aff207602df5433ad05d3adf54b7ede1d131e9326948794efa9ea1340fd79b918fe1667;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefb1e173f034d2cb968fcdd0c70a6b1882f04e8fd9365ab35f4cf6cd4388673ccb3982c26fda2ba6de1c5b3331d8fa83e171cdcc8c6b80a142a68d350;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd26f37f0e0b953c7fd10d74d7fc23b6bffba5581c04aebfb30ecc92838770724016c31f511b9b31f213c65f82353472911fcaba0cb2565f90ccc6a4e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d1c72035eb06634500b7359006d8ef5ba7a7353070681443f861ccf062e56d0421103407bd15e9b2af201f8c0b9820e3a47486b0f55ceb0b2dba94b6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c980d750c7fed38be67d6d2a73e558727e83ced0870e779633b2c766c1042fae2570d167134d0229ed230f37fa9e660ed70f7720388222251246f20d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0a8c983723f23e6b8ed799cfa4d95d0e20e9ba6675ddb184d8b79e8bca253db7aa587d71792e8823e5371aac01bc66965b7d3013cd2221c0ed73d6ad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ae9105b177676635ea954f37f3217a2fdfa30855ad357386b76e3d6698f68a5e216e4a5a4e7e93b55e15b154f57942f92b4a04aeecd9052c90877be2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haae65f97431c1daee22beacb44238905f3aaf4a70b757173f75b8b05428dd43c837225e20e4029915481f92dfb4fbc2d7d6478f568587ab51e3abb28b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33310484f071cdf5ad846f541a351d58a0a946e81f3d217e6d515b15a24c7696a8d2fdd0141783a052b7df08f74cf05580a35a2014e5d091386c651b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2da199d1c1534524d43dcfabcea5d31e698c128d10d10faaf94f5b7074b66869e23339cbab540b340f8bc66ac7531b44baf659509106d2afa1ca275d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbc14206f944562f64c1bd58ee78b039fa9365ec5c20eaf35b7d2d3e4e860bf0b16672e4c04c8db8abed772ab6393820d68a2e25a61eded377d9eb495;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9996a5d4bce20f2ee8f7ccc83abc7ec5c16f4d43294175032c3d0effb56fa8058d681a53976ec0f75d5a09890b9d54496074c037a36a9bb9d07fdd042;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda7d1d2b3f04f4724208b21791cc39eb12a8cafe058316033a6152b4b5607165c1b58f97dc6316786875a6fc3b9f03088f78b59fef0eda4b284601376;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e9e1e55379dea815da154a3e5bd1924adb8dfc226018ca6bc7a41ebff25a4ca387f678d58ddab6357bccc141dabe919eaaba8c741082eace60a13736;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he17d1bcde69899a04604d9089d64465a3fdc41edf220592ff05d0dd942a82817bcd7ab543043588ec90da65f99564173cbbd5846717234d8c22e0ef0e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e7f66ef8f2a54c9808dce4601ef565c4f957e9a680a896a7d7cc90d6a4a904a29b8e9ecd26f533b27233a1fe8e01e19d8c1edcc0d3bbe4a611c4bdc7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc8b786c4e82708519d4c11690c288610270567fe2bb813cca9785126b51ddbc1915f08b7efb474d97f1b87d7488a964c6308d2e3cc79807df9d591a3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha92db7f885c4f23616fd88983eac679dda8f93fa8eada229a45cc3f80a82c6e8948b94c11286d0bcd6a78562249f60b23f2d812a1b3d45c71ea1da235;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18e434be24d3f375add564111ceab46bbcde562f17bed79dd321714fb8bac64bbe89cd5ed02c3dd47227f2bf02e79e661f21977edfd3ad62dec7ea54c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c172bed7a0cb12d11126d63d4d2c3ac57f17f4e022856c119e751800d3e7a8931643bdaebb70f84f7232177ba8078ad143bc89e7269ac60118377849;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha36c10c3fbff7623fa93b0d789029b26f7e6610a0bef1b0d98f9857f0ce721ce090437e497180236d42a68fd7ec6dc6a77734724dc13998bbcd3918ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcec37e97d7c7df6885cf3c1b140722361f62fb92f085cbc92e188f230cd90551444bfbc7328fc98aeb47206e2c8b34ea8a05d138406667cd4326846f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40e86e0dadbca79e5178fcf48231f1dbc76ae37744d6ac1635977e4a28d35d1e82accd1db69e61c9f94cce0072e186c849c5e507a9ecdc9cd6fe38d47;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14c91721b1908616af54b119d270f64808e77ee23eed835180d32c2515f52b6f82c56285dc7fefb9a43e1c763011b1618ef1a0f7d8868553dc18c88cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2af2fd829692243b2f273bb2d3810e48cf16703e4669c102f373d027c4108fa37302e376b9fd81d5de651967ef7d0802c2fadfc362ff8fd1deb1deaa5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb236294d6f717acef60879b5846ed2ff3ce0fc1174b762ee1848492f6a7cbd2d5db9082a3f4ff096638077404dce9b4d9c78cd1f4d57ac1bb71f8666;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51e1bb24b881d1ac1cbdd61debc442dc7f5b4e146c906f5ad6aeab3ed96165f16cbb3b1afd69b4e5e808f1015f209c69018fec5b843ea3fdd8dbfe911;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff480a7ff536020d981731ae621d4ac5b64ba6dc08fec167cd324ab5eab0c1a2221250d334fec67b6094c7f8e1af9cee830738ec8689a580ed83910bc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24ff28b2269e241b80ff001df290a8537bad9ab8f18d8c6173a772edd4ce98cb78ca6763dac663dd4b444e801eb1c5048b7ba046ecdbec632ff2e92c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heacfbd335350dd4855f6878e151a48dbb033351a1eee6fab21be9d26e6169b61477c19cf3ba455a77d0317847f18429ab6bd6dd8ccb620f41a68b8a60;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18b9119d0de8ebbd6422980c799faa18f16a16c1580b4973c86e8ee4673dca7375b23538a826fb566dbdf2ca0ef466d5c7a5442a152a70f3b3924d17c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67a01e186a3faebf9a3dfa37e6bed774755bc421910d017736710b969159ce2275dc242e541886fb9bae3b4d572657573a6a932da1aa4e9fa1cb0f2e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71d804491cc3c4117ab5eddd088c03252350d5983a7870a7df6b461b2a24595d7242ed629ff9d3706e74e35f353e5ee4659faf3639afb793921ce5ebd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf7b0851b12dca9ffb65ed05e0546459de4eaffa7184bccdc42a91b147d2913762d5f44c5c24f4d07163532edc47074ba87f8559e02daf2e329e3331;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2c25adc249958e4ae9be63d9d5d3a510a80f6fb8af0c3e3b830094f06d67fc6104961a1452d1c1a76e460ad376c0741bc0b68b2e703823236cfaf6a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7abba8684beb89a6fa9500ca6a82f33b5f25a769dd482c14d8a083a72300ed8e1759c86f6823917f9c305523795a11e05dd79880551a9c0a5f7502413;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd741cbd4fdc8f5f57a6d048c3ca613455185866e952b98e676e379dbce43bce782ff6d04ca01ee0b0bfd4fe05195e41885bb34e6992360b32009c7a4f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h423e61667c48bbee58f8d09b84879d8ec1da45a1e4dfd7c161d63559562fbe216c15f445d6b8d2b6cb550d8d59c9c5449ba6d5917188f9eebbdcbd81a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5835dcc388398bec686c525bb5082f163c8fa80e7315160abc3bacfacd0b7a11c9dda1f2f19f97adebf2fe02b7fa72d61b1cbf6b0ffd05efd7d722061;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h398056cbf09a516b2114c0219f4c9f29c5d520d7b5e3cd0d5614b593d003cc082eaa8f8957a5d3383164b16c41ca5cb0892b752bbe9ddaf9913cede50;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf89dd9cac61298bff89c4465433724c3d1e276081883479240d45caaa0979242abf489b8802d91ddf13140bbe81ab5046a3a994e3d3d2f4aaaee35fe9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h976b042c5853b15f5fbd7a595c7a7e65319a41c3f2ec34872b8effea2df9f72598d4ffd3b60554ce4be7c2a19973b925badb4f78d870e6b637a7b0bdf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97909c36de53329fb0a92309954da891fc366e08a473c531020e532213756a73dbc95f3fb7deaa5331d9b7ec94bf67326496c2f6911fe79f36f1c1332;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8eb233d437fc7589b0f0df60ebfbee3f66bf349354dc1685fbc2d83f91e360b7f5a6dabbdc6c1a82596674172f12ea45638369960324a4bacaf759e7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77ffc9db8d2213906030d711f9d2e4b81e9eb9bdff4bc3a6c24c875542510b13c25b8e4b648b77ce9e2d256bbcd39a7fb005a3481124e7b9585944610;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0377cf5049b2d7ab84e12737b2b09c9dd33c8d3798467dd663dc973abfd895539de9940f9ce723e09bbac34db78c3058ea368289dc93df365e5fec70;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7323a99bfeae5b08c1e27c77dfa1e3c983ba8cc772c3c36a4077bf7d0f8c05060a6d4999ea9d956644ea499054b9f5a793e7e189d001e2366fbf0888c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9175060aa21554fb4f730e03884cde13ec31bc1090dcb053051d436d7280a61028d733eecccacbf0e1235fdc5bd23ad437bb172fa22714fe8237e4008;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14555bd13fab8b90451e77b2fae3d6243f688d1e470b318647fcffb98cd1c76d1e40bcebc23a32452b6de12499dc79075049e4c5f2bfba4e70f89777d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d5ea22fb420aa96b38b9c563358a15d0823999150385f4a36b6439bb8d270bd8c8488c92141dde702ef98cc0c22ea37e95ad46923e3c13296b43e4be;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64250c06794adca941384215478be48cdb16f2134e794aae25b68880ffb2d4081f6fb1240a082b4f28f82c87428a668fb6a9ea17ef2f164844b64aeb2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had605a1613c361d4ddb570e8300a157163ada8d69452c91356dddb41835d7d874fda44423b188646f96c5e62a94484a17f157096063bcb0a90b54c333;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e6fe120c49a69602dd4b25f047c77138275cf67b6b8914a2b99ef0eacef45442f85517b44d6ebe90d0785c07c0f142f5ac889e19837bd1193e008dc3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd67baf75307972fa49de553e1350d56c228c2bb1537a2050066305c7ef94e76ecbfe209a92474cae82667c73b39753a72f276baeb295f0cac7622493d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb2b122d950155f15773fef7a6b373a1677ab48ac1d524803b184aa6f9a3a350f97761f6c5fb6f89dafa68eb820b8bd5b5c3323ef313b9c3fa2bcdefe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b68d97ebd76f1fd824c1a390a32e9579b44fa180ce08988f382aaf71dcc7ad1c705b6463b7ec7d445dada9918c16d1eb95442b4c660a1c6a0c414508;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86f3afb3cc1455bcf6e183b1f359987959d42e33a1788049317dca80a5efa33355ae577309eeb596ac564a06b5a45a5f396fded3f933c478e1dc3de9a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1704384344b1ed04e98ff17e98d63936d0e4556035e0f529db896b515e897495d816c568c2067bdfd521645c78314e8f72fc29e64e5a234934ed01db5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36b4ba20ca0cdec107b8fd7ad17223ce96f98f68fe579c8f703f4fa0dc0ecbc8a256f158d0bd7935463474d0ec86ec2653c8276f680059b89823e4926;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6db9d99408fc666f04dd05d72d42fa24eb1cbc677d2de6664c1128f0084a5a732da9fe1b5ad77f4fdca5f5dce478e2efbbeaa1ddb058c6d21db3ee8b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h177fcec4f10e4f538b1ed58e051151cccafc02420de2ce92c6fb5d0756a5fee24bf95bdf1931b8328c5188b6fd6cc75fe7cddd03df6036e78c7cd3ace;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a471b104f1c45b2742c5ff6e0ddaac5099f5b65444e027d9199e51685e35ad3c58cda7c13bbee50d8ed04d06c0db5cc2c15d9d035737de551069e668;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15fd5ca1be557f2a8b1db0ad70e7f28e17915281441bf5e9f6b83666490fbaa25fcaeaf7fad38ceeb64f7b6172ddbc025b7ed56805392746a46b2c7cb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac196c375fb6108ccdc8b1626973c42f501c2f538acec9ab705c80d4194e5b0876dfb7c22c893aa25e86e62dcd4aa559d0ecaeab5f694fc9ca93136af;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fc03019918dc760b3e2045c5cb2db1cbe636c2970ba265096d8a2c685c53bfdffa69452c2dd0bdf8deef802d1a83a160f9473512f70fb365c91697d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12b30e05fc720ec8582b9fb1dd4e768e558273e6f0189872b33058e084b7a9aeb411bb972f76c31d92083d65105af060868b61d4b92458591d6154a3e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he1d1d56f4a7b43fa4a437f415a4c461dc5f44552cc133a9f9b9c6ba16ce8cd854b47c59e826a23fe950b92995b197d3931720a4632da56d09539d7688;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb443bf17657f7361c105447337b7160a42a42f054d3853712434ac036e33d75f6ac852f12b8fa8dad4d536901c9f4ed03071c8c9591183d94687dbd9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa8fc5bd4b584b3e72e64b64465c5c06fe6dd0cf5343f883791b3303bb5e0bf32120dd3455c8b1a812400e9e8be47fcd5e81881c5c8fb9d72f76332bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f944b3e067279d70b4922c93834212361584bbd119efa59c31ff24beb8a37327268afb270173efe932ef8bb3131246733557bed79986b3b3b8db33d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e1840f8590ff1886b931b7b1e7a6ecc824667434acc1e26c180122a865e0641ba3ff1d3d98186e533e283bf1091110e6d97419811df5e56bb8ecde62;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10ededc84e8ed8c94a8917c90d1722273c44999fe44def547a5d6cfd65cee553227054be37f17b2aa242c3870c49305e987f2e749d4e1e61dd1b16383;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d5e177fcd56cf9f6cefdbfddb1d7300975d6c9dfeedd06d9ecdcc35889956df92171ce54561b41730238709772ec3ad1eb6593e8de2391e16a969c06;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4625640375b128ef8a868fc6915a5bd187598cb5b5911fc6801afc9aeaf6eba95b9622f9725bf2512ae25f55e7c08193737ac469e09f7946d432d119;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70ba77a1b4c359d3f36b722d9a0fc0d10321b55aa35f372bb7f2bc8635006576020858987dcf72db58eb96fdc6f3db1039067d2c509c4f1e79be91b05;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc97bb06e238d1c7da2b1770dfa722b6ec03e2d066cefcbbde7ab11032e7c63b168f6e9e5252dfeb6c52cd8a3b94ac598bdcfa57319fb1f6cde8d809b9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75a3e0aaf4029c9df7895ebb752b39231af6a46fa648ff604e447cdf54e591733013c610d3d2aeccdfffa034162ab4157738e5a5a059cb915137b8160;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96e93e1c22cd998982c8cd8fbfea0be8d460401717a83fbd7b7ce8e07c1895375b17f8d63b509879892a2402adb07724348caa116ca85dcd88e6bb39f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5abf9dc0e529beb498f8d024d9218e4bd6e4a77fb0b8226fe04072c2528f39aed4da868416377e618b61e15039d092ee383e8bd6169e752f33e5cf407;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heebd9039f1fa3eabf524f660a48eb9063afb5e1a1f9dfc2db230b41fee263f87e5b4edfb2c3d660f6b435bf80a3095b10bd7b7079b167f13e38314dbb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bd83a9af1120a0d9e9c53ba210aa07d1db5c83516689eb972c49e08c1b68ef1f648760031d31d8955f5b82896c087a2fa623ea241dc254d7390aa25f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he73707cac20f8b9344707697c648043007995567ceb0e765be3ccb56089535116a91ae4021a533f1d41eb93c88af76d3304815add4370a942a4d474b3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50d2e3fe32e81edcbba172729e0338aa696fa3cedd45e81b5baaf3b9f2d3b3e9477b65b36672e4e75a8c14cfbe91d6fd999ce643dd92f70d6b5074b41;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c6e03315eb1c484407b017b072e7ae9b9bf505215ae6b0c6c6d54fd38d087949a08b140e63e2b20427a6b2e502eeba4a96e04ed2f4af6b29ee618d63;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8efc59cd9ef645f7d2ad13e307fef19d061cc240ffd4b411926902aeaa59c9a85431a1d55f990fb5fae3f3459f72d3d977e308eaf5034a18d4448fd04;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h148a8cd8c3bd6f5133459fb59b216833bfcce31bb77a32ec63944e2e4fbb1a0a3d33d5f5d2f99de89258a925edaba57879a118aff8769bc3a4a1d2951;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ed78450f1918e52f9cf34404a836791f9e90b50764c427996fbf2a424c8ab48d8c5a6be49b27c556c6fb0a95e374a4d5497dd28929985745ea6b665b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6236b2b1363dd3955983e22977f263d714e0a108fa8236a3ee6b4b1b706e89e020205261d196e9c13fce5969983bbaa8b52c3119534bc0414f1663a4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3e982b2d3e2deea1c938e503268d4b23b60c1439d82ffe1319e6fbcc816d54c1bd5f2538e3570f648f269dea50db7f9673aec928ea5541b343307334;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h110c3e145a9ae6ca449e6ff34c7e055d657e36c8d2386df8cb8560d50bf94e4b8705f2c41ff01453e698b776cefe93caeab4ae71a5724478321af53e9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ccab7110ba30919555c6338f12945df906ecab131e1f4340ac32246625f1d5866ce15349115e5999e6b91447b5f25ba538b9b3c1037950fd5914f3ee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53906cb1b88ab3e9593ee6664ce85fcb209a619d052c658d4d3e7aa868959d760a589e441d7737ba11eadc786465a064f9bce47b6a8649254c56bbb2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdfa317b5c20620c08d0b4c91f57e8b4547ae1a00403e91830f830b619fbd721e97020b26641cdc40a3a4f29e95b557bcecfc02c7b5abe08c620ec87bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbca4701f73832e7ef497223f8643ed5098139627896f3d9c351dff4235c2a0597af4b670d3627a973c5e1d59f752e95da4f9c53fb9ba466f44cecb17;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ace3754a5027f8872c7762c1fcdd4aa801bbff23f18dcf09d71b3a946a8617e10fd73295290547fc9ddcce13c2611db0379e5507b599586ff9039df7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h709fe84bbba070bea371600017286011941ac6aede404e796d9f81dc51e7202a9737bfc07bc8fd40d5e1f199cd4bdb502cdf3efa5363a61ab095c1275;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h218be999003e2e54d5c29a113d664a75083acf7f6629726da7beb26f9b50acab9b066d44a4437f45f83ff9c4761384df3cf6944ffcfefa1ff5520cdab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb3d455d03804e0267244a2d24ac51c4be2f1f417892908f58b6b119420515649fb6af4f5a7e680b2f8b2affd5cb57e175742c7746752c67b42084a6b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb198eb0d6723637a2df468f4e7bd04b0ddda6dcbbe7a1469a7fc3c90dbec1224f55ae19f509b204bbed5bceb35ac498de57bc83af88d700bccc52e109;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80cec7b9153df6f4e6b2b11083b9b421657edb19587e9d8dbd3b2789cd8897209664ddf17e05a71d3472d6d1dfcc9d496abcca73ef23ac39cd39750eb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h547fd8abf10d6fdb93f6dc666391532f3d7bb85e4215608dc120b905fb18ee2f986fdaa52b2ce9d61447a3b59873215bed914560801ded1a8949bd4b1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76250a94be6b8438002a30c515af87510ad542474bcd52a8b1485f1d649969d43b76796fad68496caddc0cc7e8bfffd59cff107c77577e9efecc12866;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc67de405f59242d09672f3251118230d90f10126749573c2412261787323cab48867a66e9e405484052ad4c4efdf1281142d9dbb32270e5f8fe519493;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdb466a01d9e34123386e62a2f43de314153d31f277cc6e039d6e7e9b2a491207d538e8a6f86f874f9a9aa085877ac6b8eb3a99349d8b68bf7be44b65;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d7bb1e64c4971f49b514de762d48570668c70d939ba25ef7f41eda19d6578b2439de67a2bac8fafca86c649bd709407862ae890e0884f0a6d331ca2b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h899b998115d0be2020f66ad5f715045637f77d69d6a90b8751992c5ffe6c13279e841686ae765eaa7007bf88265f38982834bd8281fffb7c9ff90fb9c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b74f4ced24eef7ec8dc538aacd5a1cc95aa973e5e71cb114363ee6f1327366fc583bd644b7e8daf732ed0670fd7b34a230cdefab691397f67a428aa0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb4aed3c0ae4322e2af6aff5e4bc82ce2294abf2b34254427049472599975a649785c3f564a09f7f06745ab5d2434cf8cc03edd914a83631dc2e7aa8c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d85d0c9372822e507d4395e025647c555ea25c19ec3577f96636a4bb5a8b49b733d7689098be23953812df7e5793065e13614dc3131cbbc6ff8c5816;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h462c410499ade7f2c9c1649d5f1ca1408eb523a245a99e91ebab0e86c389c31cd0dc94b1ba86471f67ba3015df3c37772aae2ba6412b586097c9d7745;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb186dc061b0b3a07aa87dd23d21dfd7116ff2876d46beafaf3c2f19fb800280c0e295d218ecf52ffac5d226789fc32ced4b89d4c0bd48af0625edef95;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd0f129079089a35a1ae55378bffa3bccb2204fa9247ef80a2fcfddf8da62df1352e75f4d3ad69802456b13f147fdc762a61b6cb1f109af72d80d7a98;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c90ce7a2e39fda3b646360bb465e27092d636d9ddd351ece355f2d72e2756fe31f95410ced56d303cb9a7d5fd581ec05bb42a38e0d66748c5cbf47ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3592c3c2c61e540dff53abc4ae056fa1348b3bd476f050b25ee88ce6f53b1662f9772436686780f2d36f346c032c973ac688745ffd6c011165a3c8408;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h824b74fe0ee31bfb0cb943eb6a96fe9610a17c495838fa1d6d1d156c48b181157a63c45c9434e991365d20ecbd7d6c2a95b57bec9e7704e50823b70d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf97f98ad8c830ceeff69618d7872482bb3ebf539309b9439374eac6a30522dd39c957ca726f1017f98cf95f9147f5bbe62d459372d767c83b69140777;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heab2aeb1df6fd8ef6fb4116af61b3ca0bc218252af9b7f8e2a2d2d26e077f180ad095fc4e66169ca0dd978b16d2407140576c5d2d89380cba6bd9278b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he1896bcafa494c7d603f281c05f1776d74ef7d1a10a28f4f46037b308c3487ec3e0675cde9d3fd0086263f9928b3467ee301c3b7b1cabf5fed84070d9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c7048941531383a9eea7e3a9e371a6ca7d912f166e3a2dbe149e12f7726708561163e152c6bcd0fb6f48828a7870864790301953bb3ebc015081d066;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98de9aefab52f993ce38d23253470f11285c744971f839793084a365adbdb5dd57aa4e709c051e883a0ee1d22eafb5130e153e64a979dfb0316d9f261;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8368329a9e21dded99b545185e498a3ab74f624f73cb7a751cd3296cc8579738933399a8cbc833be0d5f0b3859c6a6b33ca8f2e8d6fd1469dd3fb9591;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3fae8d67385070716bba8e76f11b940fdc3d10cff571dbd1d47b5f61683323588ac1c065db44df6976df783ad4abb59e6465f1dca7c914335d91a182;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99054d3f4b4ff5673c7f3ab23e54611d71e3acfdb047f262f54f6768f32dfc768b6b9d4efc8287f6f1708bf13fc98a30b5445409f92d76916261f4b6f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he53110ed2f0cd6bbe7380053c9bb8b513d87d139211dc282089e4d588ca086d3a7d81ea1f76afebcc58ed7c1e5fc127d1ecb65a29cb56f633f5bbd2f6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33424ce52edd7c0fdaa926df2975df8d50384b90ce118f8883d184fbde5732f840bb75af78d37fe38be127240e850189ae45e6c7960441dacbcf34d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h407ef7f2c1ec9409ee993d00ee481c1db75570f3b5e856a43076fae8ea0600c8383df98fbe84a0148a300dded2efa134c51774a4761f7b417857139e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1da97a2fa693346c41406cdc2a3b662e51b814a329697cb8e4ae9543d30b60399371e5a0bf66c587372c3d31dcb8decd9ff183d385b830e5113a239f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h769b26b08d49ef018af4467fc2584c0944d43be169dc871073c00a39099c266f04fe946eaa186a05044994d91fdbc858eb904e93de29cfe85ec629a3b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h404f1f8e86c1a957e48d5e6e365847db8c4a8aa39fef2702cadb1c47194d57584610782595b1859daa5c385fb94cd8d7147f7a1481e55be9c4d7cc6e9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha021aaef804b8a070d515e24451564bf6f4e3582806c14420b61dfb98f46b4199a25a7e710a27dc7512e3f20f81ea56af0bf8fb8c8425a6ac2d39f60a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4f0328059abeee176b4d5e89c541c5c924235e0d4094d92237ed6840f72ad1c6f0fd6b6b1ccf2f0a2217b854015af81dbad836094cb099a35423535f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bd6aa1dd6ced6e51e33882209d9d77f92443ba4ef6c4123869b9f1f032dd6b5a608baf23688ffa2255883fd3a038b1ea37f0881662a5e92e8cd3f4da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h23e1f078bfc96f64bf8e3014fb4891748a5e354fdc00b9994e4f9c595bb2107645c6e07628023b855c80c2653abbfe7f0969aaac734e36a5f446acf25;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf6d3d33d497f7176da774d9da341d6def46c32f7ca04e6566020345fa3d5842131de77eebb9fd1bf3f71f74046649a13f6271b14a1807972698d0ce6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47966e9c04df4ef021bfbd004d7d600f121e636bde483ccc499acb4d742f1a2036af015c8172ec2ba2f900fc1eaec299ded1a253d016412852bfd707c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h169062921d85b9e0ffac5387662a52157ee3d4bd0f875ea6d7d975c462e63a2a1b9a717c65edd00f9ef614f1a007aff53550a4d7dc13643f25b1927b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42511c51f0e38f8745f9ab71aa44132fa626b8b3d450a72726e8342178318ffa2c431812d9b1764fea03b677ee4cfba6c252146e4ba9283511b270c8c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40458680bdd6b55748fda4315e48d202e618df1d59857c7dea4cde38dd92f1a3ee8421bf1cdf0f736a69d5db3781ebaa94074a5d2c95c509b53139fe0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6cf2d2ecaf1d57a2abf9cc9b6995ca51f396efb684d491df443dcfe7944b02e3fcdcbca523773a9054f7ada4076e6992226af0c08a49c011795b014a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haea3622b163969501c514b4dc76d7eab286abce7ba12c8695fe30192d2c46c5896a315420ce7983ec2b12343463bb5c57713a5199fb15fe6106b27652;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f820a79c7215388b740807e7ac8a419be6adfdbba2ef2217159e89988d5e3d1e7d9f7b7ef56a239d7699717d4f8c7c2eafe6229ffa72fb4307dd653;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d2a13d748e8842514d646e5733f5ea742bf6946327b02edd4fc892b0b40cc955e0d1bf17b215226db1778f4d9acfa3d69be8d7887956585988850705;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd8d586e1fc5c80b7bfbb68e9ac092521d22c928089083d9f1136f458a71f2ddf53b6105b785bb00e4997a5b502e5d65b027d404f34350003b8c03e3a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdac2ec738fb47a02c6a40ae7cf55d04d36ea65a258a42d8fe8cab6b5e78aaa29db57555f42bccb7df0e999e31f5e2c0d353d35daa19f4c0b086e059f4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98056971769608e6214395c39719a5c6c87bf9a1f2f4549a24140672d58e8cf63456135c190d0d40c659c03809b0884ef89deaded6f97dc01b47cc716;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h207fa56a8738a25ad2f30b255e04a865087a18a6fa2f822a523853d90aedbf2b80f4672b7253e987ab5eb192c3acf19b7c0de77b0293dc8dfbe728307;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20bab9b3c3ca4cc8c616880f18bf51bc946a9dc7caa0db50a852607cba5238d8a62d5208ceac2ccc439b336167d90b34b16b00b7ed75fae4eb44e7a11;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb71707f56307a7ba7bfb5472a47cec0e53149d446b9171793a31efb7898449998859dda0a60e6d735224f7be8744e5ea3e82d722105165ef5673693f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h569e7a1d42e1780e618d616b400fb2f5aa208b2a9027f98f7b3e577068ab009764904507500c81c48fba8a2aae702359f5d2d1487396b1f90c9ae39a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7420e3d2928325c88089023c2cfdd4f4e855b9520eaba748c759f9f6c2838836fd0804a66aa30c2033c2988265b61f9bf2071c9c700a013e25cd9d83;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8daed6c84fc9980c683d17775d65ba667a63c06d209b91953ec7a9045d28aa826dd5c43faaf8140d31b5b66cdf847e23341eb24facbaa3aa9c604c1bc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62c8c6d5cb3d02bfba0f3e52eab6c06584a96f694282e2bc43984e4c996022858a622ebdcf1b11bbb088cc1e74d9da77ab28c4f91e875b0bce25f3e34;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedf9cde47e5a4d2d6906a8e1734794d51ba71a739a823f113c90a733189bace1cbcab70d13f75b43b633926445b7ee2fe4b4ec1760ed9d07543f74473;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e99424db924507bab61fd2ecc2c8036f25ddb2d757de79f8c7aa9360ef6727706e94f16a781d44f3ed7e2d70b4afbe0877cd25bce5e0187449f4ea4e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4cb9839c9a7e7f704adc1b9cd40bdecbd10639d0649cdb0b028c5203e68c10b4c09d06218f04ae0d2b61354ffefc77f6420f5a3cdefd2e9aec478cc1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca8d4a203a25e7936aff6d38e058e5386333046a97ce9e04beee917a206f7b2b6106dade9e6067136901fe873f9ff1f928697793f2d411cf4b6db1153;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42880b27595123847a7c72b6b0d77589984141de13a96f6bdd4f9c2f7ef05b58a5fead819a62eb8a18dca099aad680c6b9ad9bac715adc60586b6af27;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64084f736818dafeb8d41eb28d510b85b0f3efe4e9eebbb44b7d2b591fe665507d7d39e3fb2a61ba51584e38de4ac556a39f677f1c248cd4ec3b4f6bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1bd6db338508f627e8ad6692ed9acd8c13283af597685c6775f11fcd6afa7833d933de42fe3dfa0e2bafa178948a5efeda0edb35beefe67aa992f4211;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb98c3c91af680967ad04a42f141f846dd41df613543d5fd03a9ed342464e564b4164772c92df5a204debd98000a5f4da01d66976b8ccc0387600c190d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc8daf53374e38a41522ccb7b837a2ef98122830278b159842198c9e057531dbc7fc4a8e8a820315c7bc3452c3d8a6bca3c3e9eb5cfb560f287d57947;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4b18f5e052bd6aaed253dfe9567f7d670890fb97d42417e67a2724880062c14326b1807e2cff163922ca81d8aa010abfcb7c30c78c57a218844fee64;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8776e19ca41cd8a8bb7e00e5850c5aadad76611f63247f3bbc069b7427accba91c6a1aeb70d908eac9190824fb03e2bcf5415b1b256d59e6688cdbfba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd14b1d104f163a9a43a9a4148d10f102300ea2813958cbca917fb9f0f861656e0bf338fd06b25f028e5dace252aaecadefa6aa72bb28a37ec2d75648d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89897880d40f862617197e7711fd39b148f9d3ccfe9561f65a0ac5f9cc641a6d80a2f3dad788ec0f1523244c9df06f554102176d4640e8eed470e620f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf1cb9c0ee1c590b793bdbfe31fe33d8ee451b5d953d681b1737fd9062729f3f23abdf211dbfeefd26c47073b4da3cb01c579788c77f9f56c293b7cea1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19e79d4a30684509e1243c1c068e018acfd83bff9ce4f48b8084840703dee2a5607bfa201eda191e66762ce313a0afe7c0df77b883a5b63dabefbfe8c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80598fe93cee2d5bcfdf2965899599894a16b08c52d99af35f03dcfb49ab6f99bca80f40150871e3f82f851f7c35ada200a3081b25c684b708c3b2473;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h831216c932abea3b923e2d6e011343fd01d295e0940e2f1fec98485870abdaa27d802e72d354092ba0183734d55c98e1452dfed4d64b9c34b6485a851;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1f9b07db4794debb087348943b2f6333d1e5d6c322778e33e49f856a495a12c6eb68cf682c774e8ff4bc481381f08703ca1b0388b1c274105985adba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8396320997f2005e985fa4e44136681ca2ca6d2dbf1df180536bb4c379e3f9adbc55c625728d5fe9a46f6f1d1a75d2491d5d5dad2a8c1e0bc59807c3b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h303d36aba41a9e642e7072513e3049e1864693ebbba1f8fe342faabe813471099a1a1f5ba13806bca6350ebc4a780c4ccd4d4249acb556e061e8c15a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ab610559bcdb379710c84f8dcde39de9073faf00cdab9f453494f2e4018d9b6b6c8824cc05fb0ec04ca0ca90e2355ed6ec67a9b7cbd91b8a718ec3f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96837c2ad0539e7d6eace465ae0df2bc79d479b27fc2d69c0fab6e3e6efe68a0eb6ad3b7954180b117a458fb9756dc165bf5c576a49236911ea2b8e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3ec4d4c4e2e6047afe5e57e23d6089b2ae2d8bbb6252fc31f08b2c66aaadaa49b7e626786ac46f7e76a7ea321e5a9359764fe08af669e458395b5b96;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d42b7faaaa577806839ae17aeaac1390ac65dadc69af034d8697a089b62156b54a396337e70b9f893210a6a2442a1801402fe32e34f470bd3656351b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc95aaeac3031f5be822fe11d37fcfff98663a2a2245c7398ecb5fd97e74aa97978bbda0fdc05b3cc974e6b65eab233e511dd14bcee544e4cbadcca8f0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h584139b1c22af34e44c835a251c2455bd0fc34d21b4b3661ff078bf4da62ed1f22ae65fbf860484cb9d160a15e1d580cdacb96066f2d83a50072f3c9c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95ac8ec7f7a9c653bb3903477616928c9b6631cf71a61b72ceffb669ac719e667a7d83484de517f80d4907f3bc0e3a39f02a74b80d1b2b337fb8c5c28;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hddc7f3ee6d240f335a4f0eb522583536c870ab3613eb11730bf998d1d6d5bbc03d8cda78d7a48b30dfe2e16e2494e35f8a99017999ef03a2916b50af8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64a905b299c6c83dec81e5caf053d94a7620948d2baf82c1a2874894a6f69e6f389151e0014de5399d34071e3acfe0b4ec0f650b076aebaa5956fe35d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9e376b5e9476a6952207b703861650cc4b31cdfb9b2ba0f779c1f3d41cc694ea9b1653600c46f331aba6cf286366e90b01a94849b8d7e20f1f3473a7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7898ca26b61c21a4a40e01c78c7f7240f790b46e2fc254a7c50ba426d8924901fba460abbc6c23b87afc20608b0df8298f52a3f43ba67e5124433d65;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90843630ac271538b8d4eaf87228352a846a1f47638393302761b0e2711db0706dfc011243269dad25ef02b4b9b4281ca6ebe5d22d579aa43a396f161;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb55efa207cd077f52b176d092b568bdf148df11d48b9f76c4a3eb932d9504dc1b90f600b1ef6f4f5ff158b75338f63ecdc8abb3a081f61ec0ea1778ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h251e0b6162b9e019b2f3d253bd8e236eb451f9bd33651f5b6222a4829e319cf992b368d07aaa9d1ea770e559b960b5b7ccb3376eecb365890103d9986;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4ca212d93485c16831d917999e641e890d2b035d90bfd0f7751cc3d55bcf989574847c69de144046c1b7068ccd316e7a620616942887979442c703c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8204af471e1de113f32b6843e5d7e842acc047b463ebd254341b7d8ce02a3f7a78490a6b0c22b8bd789b200b4f5c1028b58610fd57874fbd099b1bebe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e6d639d540f1f49eacfd384088ba452f762d063cf36dc5ae9313cbf39b939baef13c1aef07facd5c391665a9990e0397ed217032c8c3df0b4e2e5684;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf212109f3036239d032aa668641755cefb2921a1dfdfca20673a6effb8c1845eacb0d5a78fd39d4a002a4f2b49bcf43ff52c1be06369e4eb49c1660cf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7de9aa822a4b28a1d34037e96975751adb94d561e79d978184e67be1374e8847f71445e554cd108e77bde8af8cd71e58f53f6563ef90e2f51f2c3c827;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h208024fa7a840699104cc4e6e8d4a9aa478c321deb98b6f9837cf91586adc8b3057a868f4e21716135c1d41ca007261f778d25c4316a0c7645b95a85f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d34607046212ab06098942918e2a6137a685a71535531bf774ab9d567891caf6c00d51440964c72305d7533ceb6336729a3a0c512211cbd1e550ef7d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59c5404945519a4886b3bf569497dcd87acab41cfd441f8faa1533dc9bd732689f4b8ef1f6a5e24d50466db32b289908b7fb87f293ddeb8de260594f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27b4435f84590be64940a725b70434794d238fcdd4c253e66522b6b90495f25a081767494b81fb00b3b8fd4d9c0e09d4f32722afa80e8cc4d609c3f80;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7aa288ef466e926af29738210753b5c38f141d2f0f5123e2948d0c6837790e1063a800413b9a2d9d5f495d7304e56d6bb26d2277825d7ac207041c6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7dae0b48359c16159cd7d3ac491f228ac7006ee3714a5c70657dc993c312fcbd7049f728f277c9fe8681a74929ca279b5e8301935e70b1bbcdeae786;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50ed532242129937e0c5aad5d5a8ebab814630187ea326544c7e66e7b74dac6e0e96d699e588f0d386d3db4fbd8a54d00d460d15b35b814132a901765;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9132a1775de6ab5ad8b31f2abc2e7f42520ce0bbe2140d12044ae7df7d939824c7b6e7ae636b662348cc7b17e63ab6624fdb1c1be1ea238e7d6db3447;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e4be9b52f95ad904982d982a14513441d011dccc42ed2c34ad78ac86d095af558662e699f0e1db1087c3f0330510d30a8bf3ff4906e208cb4ee5fb02;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36bd3d630aeb000186acf6e96f4dd10effbbdeb9492a36bb94454d907e4bb9bf4243f84b75152eb73b80bd1b35f944bcf89dbbb79d095494c4408793;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0b7aae437d4d9797c6b8a6446bb5b09128752dfd0e9328224fc11e65662d98698e3d8aa29f2bc650c3249923f8260ec77253fcf5aec482d5c8c66129;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9db999a6d16b31a6d8501ecfae06a5fee0d6c58a56683be37d7be9f87454f9207a600b09c1bbcec0c3711e1e2f7995de8afcae94634c0d29e0dfca681;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h727a01ed6e67a0208542dc5e3d168e6d834544cb3b83a33f733eb41216f1ca411552980af8ef14508877f9f716ea99dea2548baeae9ba3be9f70df38a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f41aecb6a887ec648fce23851760ea5667ffdd0ab554add58f753f9bedaf73bf87fbe32c14f0d2ffe026208d9c022c3ab5ba57b3eae6f2d80671e2d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0cb1d4114caa0ea52a320373c6dcb01a81c23b2f9470024e98759e79b353d2eb7805bc47d89e5da439d137a15202f904283e9ec55a368bb91208ce90;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b06951c618be3a0e5a1ae70f7eadfb10b7b28e461844a1b04b41d758c8053f095471f0495744b0f8d3c79e72cb488fa2d997e218f67e8c27afd77c38;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h335d27a92846c759cefd86798b631e16f01562ef856406bd33666ee67a34d324209f3a8110adb3c49e00ce459148e9ff6921876335982674da407c02f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66625349e6f2c5c22c98b313f9a8f4b84f9219c012ec84ed84c73bd25d7cec59b5d37bc85f89ecdff03bc1c022d5669ff11f7359516e0709ff6398f61;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa913c698020b086aca67ee9df024c910a3ec3fbf0516d48b2da73b1fa0090d8f21b0dc69e1d52f7c34394918a59143291f65fe67772d4bf153fea7ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8423c42161fbde4a3237291ebd1137ff3fe75643416e37ed433273854f6b9731cdf58c4c165c618971ec03e5b731b04f6ad806bf7a862bf933cc86bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64b9c2c1be067fb5429338700db5f3e8d88ff1c44943522e90af8168ab8efc8243c69f7efb8130ec530e743a828061e31f245fd66b7d69d6a923fcb4e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7ca6a6857487975ed21087dbbda371af6b9e365b4de6d8d8c453ccf347678884f822268cfc35da3fe3d53db25b17ab0497e6d15b03b3c7eeeb75442d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b9b1854238fe223e1ccd9d6e2e2c5053fef337ab4d16a227dbc352f9ed25881b0fbb6c972f8464fe1aaed7d43f581e1f8f414d718c9ecc05abe59abf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha157bac17bf1b771b2f7d47448f73a850f85567222fd87fb59d2d1c0f2eaf576553c124eb2408d6966815fe4a16efde9d1320f98e97048dfbcd044ec3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc11c0f78ae2387d5a91078a3fd92607d0e03cc64886b298a283dea69e7aa951e8bac0e9ba663ec0ac3691bbd59c61878e33718886f19961d0beaf5434;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7fc3ce1518b4833cb7e6dcba8d7cf32d5adc596d8cbced6399508e545baf7212d6c836689abd35bfd07db7d68ea44b555a7ef75e621a591b0779800bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6cf43b71047e83148d21e3632796ad90e9771ef1d81bb8098a629b8da3a888f4c4cd771c8dba5f20d2fd655409693ef9e1e77b5042d8a3b73a0fa0462;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb584b7bf9281d1cca148a23176df71a192321025d02387b8dc0a8c08436086dd7490154cf6bdec1dcbab6ac308723833403c335f752f42ccde6d0aa1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h404063b701f9c54bcbcd696208ac9167e97f7c73eade16ab2da4b1123d3c9738a0165b0952857ecf57d57efaa4f6c580dc3edd3245aa896cc3220bb1c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h872317814428a97ee32fbf93accdcd05342da1b43546b298b1406ba47cf4f4baed0fd64fe11d4c6429a01f8c2519196cd8b124657b64d6b20e1cb5376;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4784fa94a0f0b77faf518d4f0e1e56751c79c729b3a1431de1dbd664848b677525dc4fceeb8b6a0213bf7d1ef0169b521e2270c450b63c8f562f18be1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c5c621cdfe51504c6851ca4178c4b83076d5fd07ad41541e645c3b41ebdfd1174002b7dd1fd68361c3b82aa743a20e6f9dce7752c63052d25dbf36dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h291428ec62c39f441abc22d7035c76d7e80455c6b59db4f042faee64a2527be7ad8ac194e81f98601f4cd4804cccf2c29005fe6dd5d3f2ca5bfe8c31;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b7bd1b9cf1a694c7b3f49d42ee0a49d10c623feb5188b5e3b2991df29673c5f94605ec0f685b3bb26dbe5ca77c63171b89507b07b5558a2c54aea66d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc8af26f5f62955f7d4a7ac3bc27b955a3e2dcf254c944449186c340b34a0d74480d35912ca6763d963cc598c51fbe974a61164080198ef8f4eb92fef;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb098f10f24f59ab3c20f746e5ccc8eea849e7805a02739f2a380d51ac0604e4225117cd786fe66d025171e46e130635556139eb75f256a948aebfae27;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfcbaccffd01558d61cb01db6596399cc6003086a96a74cb939ec3859403d2113f0d923d02883988840a1cb1a858721014a062bd0a5c09ae8c92651dc1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h372ae1f9e969040794be623282e2ac22e5c88565ce038da23212dfc160cb76aba720921d26d77599f911ceb8bf0c22c76f7174a0a7ca8715072916dd0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6cce78ea446043c351c45604cff4df6be088f7aa86682ed407ee26777b4baf202db445e2838d8ed65d05971174e1926ac132519006906485ada93e8c0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc559a6f26a68cc0c639ee2270d1ea2fd7e5483bd99388dd28762075f105119ec7258846376413526242252e477c939945cf1a4e3227eb7f26ea84e56;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2dda1d456e034e0910845e50618ff5fc7861d4ebb157948e4fd32072f5061b2d931102854cc13cc58dafa3f8afba45769c623ba31c1d35fdcad99d83b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0232b248429623cab443e23d3a53a93a1c846cd578afd1dace2faae321aedd7a6326c2f80cfd03da7845d0249a97fd1ad02a7a2b9342b74b260d94dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb2e9efc3161b702bc90a0bf946cca828aac1148f4bdadcd62e462a691b0a24716640c327e633d107ccc6f5fb9d1423bbf8c2c2def7d4e7b12cd0dcc2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h920d8f1ce95459bfd11a5d7c0de6f7658f3d2d20e39d2be6cf132751388823d9b5554b0ae0235a67b7fe90950cbebe36cb369e0ed70e9ae7836b2a75;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56cafd86d0f94392c6e7d851d22a90d46ab84a378401b5e12b419cb214e03aa8872ffc3ee71dbed71a2a336e2471b8279dc281d7ccee533688f33854a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3dee7a59b4cc6de676cbaee54565a9754c339baf03d01471ebec6ebb46c31f878aa46b796450f09bf9913ea22c0aec696d7c1edeb71cfa9ab60c2dc85;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4cc377bff53de200e7730bce764c1e71b77983532036fd1225f643f5a645627d9c134718feed2b19f8bce4db237b5d083ae79f9cba1103c4f5d4c987;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72773d2285fa7f2e75cd6ce86b56aa3983d3fb5ed22a218a3c3ef5786fe4c60c0c0658e01f228b21d06de89fdde82f654bdb6bb03f520c6d5e408d978;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d3117bb24abe3e965f9d48fbdcc694906da14052bbd2525ee9805f34cc85e17fe31305730df2e5ac0c5c2064457cc8ea4375412e0a2ca3a6dca59b6f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd223e1a02b0a73f8ad9372dee7d4e70c260f89ddc1d2bc749a83679a753dbdf7e8f9bfc6e4795a1d2f7ffdede1448498998e6cb8bdb07fa2a3f1325b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb036260a4ef6f15966ebc00662625be375c5b011e315411a0cdbf7c2f4220178a3a3093e3fd5f03431aee38d89b45d3ff7279e2fbbb94302474a7a964;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3657b55a12f287795809d4ef14633c54fa3d6ddaef48a59c4b2ef5e54c8b742edc12e442047772259cf9a6510658b956071ecec5c6190563dbc85f570;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b22dd3e7ddbdb6166688126b73a29bc5bcd8dc47a6f39c27e52e18076e9895b1f8caafd94678972a724d5366881c42927e7f31a36217b0e3aa63665f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94e8f1d13143eafdf4db7647effddc301f1874e08ea832595e91a76e4fac27c2e41fa21e3bccf2f7fb43cd4d82e3ca37828c74ea19b8c226311ddc443;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h785c80772c46e0115583c87f93db7188f4e11b4a14a9896d1ecf126079a12c4f9284859a46e2e3a38ea6335b16e7e0c56b6c0d985ac42b957610d32f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0bebea4aea5c0d3d79cb3fc536a52cf190f1a46b316653902e59f21387349ad9f2d8c753a6923c14aeb022c53853cfbeb42f80ed41b9f5e0e722d8c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea6e21b8ffa71dc9ca9f325e4f2d40ce29254d4bf9f76e0efd2e909d484298ddcba7bfc2c00944051822ee713e6acb6fdcdc6361a0d5397629ce1b646;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb13aa1dc022d75fc1579b07e1980a542569f80aaf95db1d3de49e1a0bd137fe14da6b0fdaf6a275c3c66ab4c317a8be7d172ec319cb4d5942f5bfcba6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac786d1bf9cf55e12f99bd15c07573360bb6b9feaca1694f53aa7c4758f63d30bea7c027af84d9842f1eb81b8f2262c36d2d651f10b4a62e3e86dc95e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e06a8ac5130f60b73fb0aadc53ec1a7409322c62227a8fe8b2b7eb839bde7db85e8ddd0b76f324c577720751bb18280004c5df51e5a789858d7c11eb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e1c3bf0ec53a9976f7e9c0008e418972bf879ef956043510d7f3d7979ca0dbe586a28f2df42de94536aed539b54d3a0c0a19a150d903b2ae6f539de0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85bc72b7483b9355f1fb97ddbc4cc489a97e08b53ddbe050c24d568f2852928f523ea1ff0acbb186b23e9f13ae1e8aa62e9b3c3d2c167bfcd3e548394;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h139d5ca51301f09406e0eb61db49b2a06443b189468617985ecc3a8b3dd59f6b922b63e6dafe2c15be60b9c960e27e8ebfb83fa35f4b7a8c8c626000a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84d2e4d35949e80ad316c3b839b485357b47f344e70f96656d83977da33ee32d45a9f4250c9042ba7cb1d3e70617fe896502758325ba06761bbbb5465;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97d0e36d44c43a6c81146aeec12bfb7dc609b5dbdaa97ee5e95d72b684c4c2b11696109caedf0e1f24be6e36231c32a16dd11aa4e592e98e0b778605c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h298f6189c3f6faa33028a95f93d0ee3a2ea96bb97331029f7820de234af29d54a7003a0050f999ca83072dd53c188e9ddb4539d0a46bb15007ca4e6b1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78251671761c69bae62e8f9aff211066b5d6c75bb0a887b32f02a9e3c9ea2bbc6386437f86bce1a9291a52421487282cb780872b72b4c4b5f1e606d5e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43796a10f35d23143ec120ec31a49fd1934ee8de6c69d6624c167c6aad850d717d8a566c265871dc01ae0243380f1491fada4ccb9ed39e6f9e939a469;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9ba186dcfc89274108029d0a91101dacbb90d74cdc33acf6ea3d39873d30193059b3f8bc33908dab44b667e7f2c2fa9160becac766093a2cf5482e08;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd15db5aced5cfab19f8cd24feb1b5f1c1a3dc18e378b384fdcbb9253c347bb2260f72e82cfae89b3e8d76e0db5a29fdc719142723ea9a706a26ff7e88;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha126a375372cf36e5810e755060b3d392a2140cc828aedd4bb8bec55f620764b0dd77019500323ecc3fed204b7d59b8e3dda547f195edd7ee9f7f1992;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf276389e1433fcc7a34f5d8cbd3c4f45284d7b807da0683f811e7479fe609ce728f95f93823f542413bcf95d86ddfd740cfa34fbff8e5827f840116a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h989ba48c0e29076511cac86de47f5d14efc93c4067a7027c3657ca68507733d392135252924a8e36eba0ef1406924df5d3d9fa342713c8ca0d9c57e6d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9a5b4cfba8719839edba531cace23a5070982768d3b10c41afd91fef9712f52e5743a39b734b0fbb7cb5720a5399e6d7310464437c8bdb315519ad1e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h973a25f3e0cd529d8e84307cabc0ebc9d319f57624d7583ac92e60e9db037bd1d744a7d33d158602ba81317378a29e19860a4c1b1d6d59613d6012e5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd305d6013cced7440b779c423e9d918f3769dc51f07a5d2775e3f22730ecbe5e9a7bb6966501ae0434a484a254190d36128f82c87e84344dd049bcc1d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77292475cdcac6fdadb109326a3a7bae186062da5fd948d82a972a72294f2c50f6ebeb08a37def6ad6bd6ddbf631b4e1548f30d8009e027b5bf1ca37f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b1be032eb1ac093b3760fff1f7664c7949a92e4826aba9686c2d5550504bcb06f34f6cf23878c4ea0e8d7dd21e547891b79b5022626c593d4eb0b866;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9364da8a0d3165c1567171cf290fc41bc6cbbb7ad50218c419b7803b142154d68327ff7969de290f00e1aa14bb8aa4c107fe83b4aa521a50493c7a4bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5992d32b66886ab344e93960c8b8652310e71a576f0c1f094556ae6260b9972ab00e30f39746fa0365daff54ba0ff88618efc4e0f68774bb63207fe1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24f2048adbbf26fa21db77bc92dcb2016a056c8c99776ae8bc1550f6265e2ebd81f234de3c2bcdb425b335db4bd81ee5dfc1b3e40d678082709b7d891;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc93bfa32222ee62123a08a5a658c932fdb1bbf5001e64f469209f78953a1419b88aafe7fd27208c0eed1b77c1ca328229a1e05c6924c529bede48bb11;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9551e67fddc5064da3dfdeb7b0dbf358e03bd641c4f53b8bdccc02f2eac02973fd6e30beb0ca7f22b3dab584ed866d13f77fc4782cb12f06c10e3fac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86daedd5200b99d6cb55a0657a636f7283b4908015d974be83ee666867b0db9672cb87ca6e5c1cb1f5b4bfb7898d9244247ad27f738c81a631e9de213;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38d6a6cea0d6b54f96dff5c801baf7ac4f2dfe98bd56a5a63587fefbcd5c324ae11f8d7494b7c9e50d63721456a36df77a524b560cfa324190d8798a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h595ba2e4be15abeff37ea509487ca96874eeb158aaec4ec798952e474d3cafb12ac3f373f569b97f66aef8d909e696c50b7bfd0ae40d63b40a1203ca8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5c4db86a9b200eeecfb5f6415807bcfcf34de2298b903764392c8951172abf734322443320f78e569af857d427fafef34651181269bfc93ba22937ad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96500a68d04ade48b40cab3d54b65d1d76bfeae13c6175fd62bfb392191e9a8072ee8ed423bcac3b22df96cedcc17993da0a0b71316d3125a8fdc26b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4cd1278da439728a81664a9bfb696dc653313fb5da004fab7c47a104c2097c21b1b8fca0ecc582ae73f9ad8d23815c471f2b01307a929a843a2ecce9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2e7c5a947944f4dec6085b5c5bd9e8b27f2005b4dc3dc09ed4e134e26c592ecf71464c94f3ef2780828269e68a1fb72fbcf3ea03be5b158ed738053c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8bf6e651f071bf042bfbe4a6f80dcce17c56509949833f367634f483d621497ed54b9ea43f65c72ae370a8dd6df92803040960095bfda169da666e56c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2fc1fb7041dbf4ad4e9a57a575676035e71ddbbb355ae9f7f0483c29266b79bd6adc6928df4dff8d268d25951cf7ef9354d49a047c291799730e082c2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbafa4ce6558d6a70762fe000aa0f947a09398ae4d567fc9f38f93f8b28fda866a5ce89b1d1955ae1942eda5e5d17301278733f627a2e76196b145ff4a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37c768139b780d0d088fd96f7896dc67e946a8c358a8e0b4161732f4f5e8ea9d3c7da04c982586c50d745f27abd0f0d39b26eed52149f0643d21e1b7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h322ab9b97b8adc106da6ee0d24b7ba98e80690c7c79fd63bc9a628ef8576c8fc9438c9a76b27e34c4c91f88c0dbc0650ddc8aa2766d487542c5a4ea36;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7558831132215c0066bc578dae7a102d37299296f0d0150ae6f7cc61a5da00b8d8caa93bc91c4003c1ebd5c66650900b6a2eb01cbf9f20a03bd51019;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fb8f73eae09047582a9c8d097e1da97cb372d304b9ba21ed0c6058145ae312ef35c6d369fd69da3ae8f230605788654144b2f0422b5081af330bb363;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h561010c50697456c463da2775aed7c4f4c01a2c75a4b1ba3a53df98c09ca905b4e813c429610c9ee9073e08dc69665b4314a4f5b97546ea5272662768;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c3da3f9de2c7dd6520faa0a36c7cefa72f48a4db714ee24108441e6ab689490bd1cfb54d209e8eab077709b43340d7e1f7b861d025d534b806376e0e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb54c61a40880b7a85e35450b8a7f9af9cf89df5730c8f3e430ef95916b5b1a12856e3a4ff4fe61144641c7fe5e7ef8f35e18248c2ae3b4e0acaccc91c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d387ca3a5ae100b19aa00f418837e9b813449b283e345663958e2ab5b43a575b43cf1504b83ada2bbbf999781bd6082075358325a7cf0fdd21bd7dd7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he74348f602e8ba50a300c8868c4ed27c9ff042173c5e0d709ca58736d1844868e192df744af24b7e6ae1087bdc2d79e6c24f02529ec7ef477e861e7e9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4908b597f22e3193d52896ddeed6625c66d0d767d38aab2cd35e1845dcef5f054f87c4ce77785075c66bee9385d1337c0f0704ab1254d79266e058ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb29b0b11fb08e7b29aed705dfcdb2c42f45ccc867127604bb91fbe3e210b2c12f0a302b8325f7acd006afbb57a70d74a0ef4a4fc333398233571f6807;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9f459f1085b49359c9bdcaea0099a1693c5073c64d9890aaedf02cc3e4112738d95220e265bf9d601faf854d2501ce885a7c8caa4e603ea16f0dfd19;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h262a1db4fd3db9370833d83f27bdf3368c2e99a045d8dfc75608409789892fe9fc9174e320d8c24908dd293d8494b4aa8039ac55c6ca79aa20cac5b4c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h759447efde87df6822942486dc8e7cfa49f4acd489e622153177cabda6b3778450e0b88eb0f21ef0898a0753aff0ef24067f6cd98ac02147bc369d4f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fbec9c08ac82a9405316d5a30c962cd0dfc8df7a79f407d16dcd8106a4effec809af8dfdf309072f218b85b7be9fe59eb68eb4ba69a441be8957b8be;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38be28306e99c6cb89f6001f2725af2e2e1ecf103b510c20c1767ed58de39db5fe7dc3e67dee37193b71940bbd98f0adc1ed6d4376b826379acef1836;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h109c41219c1f034aa43db3406d4501f792ad61232b5b13598f44109b2edeb4f4a48f52aa96ca0c52969bafd271cb343fc924a460e1b42546fa0764303;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd2fc4888c8c861b11b5bd3855c2590f89f8ee371b0e95e71c23ef07cd5b2ba3647bcad1e6225bae10cd66039ab2ac89b3d405270ff65210570c64e8e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5097d825ecdf66d036df2704e09ea974f872874494ab3dd93a66c6e3b61baebc1c3ed20e0bfaa245375b5bb161e961f2f9e4ae74b979ba31e5006559;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b096e16ff63e0afeea0833d4d294c5eaf3d9630ab435470f37eace1c20922fadc4dc8ca47482d2f4a0f0acf4096ce93bd449386f406046dc658ea547;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha97eeb8caf931039981c01f02717c765c4efe185451c79f9cb5181da85ebdf543223d7d5820a1888e4e58f39049ff374d5139406130d4895617b3f7c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12a69e3e1fcad10755f19795abbdfe20a6bf949bc8a72b46f967f01b53eab1028bbe1395fd3ea5ff9d3a60bd44078fef6bf175a3f0ac30070fd8921b3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdef3f613b79e9ecad11671bc6ddad50cd33011e547d16687e887bd3f2a4c6234963ad17074028511eadd402a3f0efb034e5fb803dca513159c80879c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76ed34be7e9f8675365adc2d06861acb2e42eedb96c0f630061ab06761500799cd81b57e08c4d44690be721cfd31c4500ac49d1ad1c643e4696b9cd4c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12209b9ef7ea0a9877b78c967e2cca399df793514b5c68c8ab798b7feaeed50211dabaf4ed5dbfeed0f5af6996b65aa40c74ed184ce044cd3f69ed2a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3ee2fe0c6f876b22b183456ae8e6efa6e9457cd102359121652cba8ce8695b66244655379ffee67d091d6065039797e68d1f8ebfe191205131e219e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda2e0f863a69c8cfdaeaed88c7926f698efb6d7f918d31600befbbce16191a87fa09b0f7f8cb9de62291d56735a4a3a027c17f5a1f620355a31153dbf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21abcb1e6fbfe90d8f73db87d07628b743ddbf5156f3b1af21a363c4d49be2c2b590453b0a72deac3ea7a8b4db4fbdacc6f71b105b176ae6759e7cc94;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbaa6472d58fe693bb407caa9f4cceae28c4a46fe62c0824dd348ee5f89d23a9a0a8af5024774d5ca5296537f6ddebce0af049ea802457b2bdc8168c61;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd38906d7c1b22ba17db9c359ed6a25b9b05f3963f496da67067bccf85ce51fcf369cf10dbac28f56e0869a066d2d01b4b6627aa7387937f65a22e1b9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e3f238f18a20fa0abe577a697ecc2be2bb2906082bca390c4d03d529d1071dd9faff14508108294b84b702e9ab734790a6ac6493998a8397cc82f3cc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54cca9a414300ad35de2a3c8e50818836d8b1217e2ec18564539ea463932356550da8812474c937d55bdf6b81c0f64497621a972af97c7af8ce36ecdb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9dff570b4bf79081fefa58c2bc7f03935916e7031270686a497b12bcfdcc6666a4a83d68a5b4bc9478a56097e6d5f37b2e9544f7aeeb3ab12ea717f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8533d15fa0c28a9d7a0a6e764a19fc211f77126f6e22061bb799f64643f68db9366d718c93b7d41f9062fa7ea174607b4838aac2dcbab487924be2b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2cb4b635e62d183064685099593df6254db8f41343f277845b2a2dca4df3db8b159158c64a6939335c125c4a135fc65b63e7a5b6e8a163b899ff1a477;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hccd6cc2cf5efe23912125ee30e04db2bd188ae0ebb3396759af4fb22b663e8bac215202526347fc93c94ea5a4bf6f46c88137ff27f430abb245679ebc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16d922b9e0014fdeb19949be279145aa95d6cfaf35ba652b38742b77fbefe25e18fdae62b81e3efd3fb7a2b72426f5e360c27554885a3aa4bcc8ad437;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7bd77eb77ca801bfe919cf7e0173b80bf1b11feec551fa45087ab81315bdc1eaf463126453d48951d37869bb309bfae9c26ff5561422708ec9eca98d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8762ad6ee19ac47277ba6318ec685e819922b483f0ef2b5d1dc9c3fca4046fe044d2abbcad7e9506ee7b6aa529066398b51f106753cb12811216fe474;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he08e4586a0b6b9e4f0cfb93a98409e8e6b82ae37a904d4a8033841f2bbd17118c3e84052360784f383cee00f28ccc7de084d12d26e48365b685b5e462;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef2fd6974bc5c249bc81d96bba6d12f6a960c96c9a219818c5200c598d204a21fa7ef64ca58546e1957672a7d4c153997936b9425fab1dc0b0fc345b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1eb7889a562678c790a7b8a052c89f6e19385aaa489e154540785c63cf6695a08ecfec4656921c79994097524b5abbcface5389a9cf37f4881ef7463;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c5f6d3af48c381defa97ccc0f50c74a4acac21bb33993339bbb48302a7b7fe79351e0e9559f52832c6e3bc90c7dd554b2031ac92cf15611b654a512d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h633eb1cc71533fc9a60adb2f9ee687158a93786f1a11eb77385561ce236a4932cb09856e6323f38123debc71f2d49541e8a4e7c578f8d03db8fbb7ad8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hffb73686b9407e9c87b695f2b3d02eef063b67855d10e7695dd6540f2a7a49be2678f0392f3f68c8aec040cd290a81ff908ba5a02ab684e470b52aa7e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdfa4476a2a498ec7739d8be368ab5ef5a00dc5b43dad138773392392307362e1d174531c79abf0603f44160c2df61ada43c6f198d4f5fafc7d8c6184d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7a2d88c7a1306654c6c68605a668213aa22aa42a5ea9914e845ecd04d47eb199021e0e3242c28d3809b95c9a96c3d88353faeb2ac005c80891ac4058;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7871b7e6acc25bd65089536c7c4b3483d710a65d87451bbcbc4a0de42726996da5c16c2e39ef70b8510d5cee072128ddbf9056571a284bd3b0e45ff99;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha513064a0f5f90ecaf323a67a042c1eddaebbc424b4ed0f9f0efe98289eedf02366e8d01213984a7036e4aa6b46dffbbe7040b2879b07b7afedf69d3b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc04e9052a68b237cdf1eadc6a601b56eecabacace1f626977697655d2ac40c61261af1e34c1874eff68246c02474bb9022412ec575e072cfdcc171713;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2aae0ab2efac7e3b52bab2b8544abb5c3665fc32a30184f77ef4c07d68ad4efcd19eaeba2c98f6d9e226846c317db87e80112db9eb9373c19c1bb9fc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8a3e4700e9d2fb43add0732def90e2d8bfc8180fb398ec7a215069165b7e53c33d047efcb0e9270e1022ac3e52fb41f7566758c3f738ca4315d6db34;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf69adecd6f22cc3e1259e98357485380355e6ba6c3dcc4813f1f4646aa11bb263ea99c0c59a0f040941ac28a4409781b8664fd374b234124814d29bd1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a16c94dc79142150955d5039a7a4b3a201c5a12114ec3d870b5571df84b6c77f2ad39d32d2e80da6879384e7cd80e47553e2d42c8343d6425b291863;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9aad3453aafe7a7fb82672b0034fd0c7f4a80e3aff7fd52912aa5c9a126112326f07aaa945c4bb5504fe334c29d701d3fa9af3888ab9661d315901484;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6646213a224f859df885b94111d8a4d490eea890cf0fee4f2bda18d10517f43074136e73656aaf51749bb82744782c456be06b564e6a894011812467;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10d53bc1d4a5c0ac715c6d8e065fca8ccace9ff312dabffe43a50911debd44e6f616e2b793d1e76ba7c4281ff1d0d9da67ba40b6fe9788db446d9ce8f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed90470845d2d79328ab394b138093a4a9908fcf50223d36e6a28a4e0243219d4db744ae3f155933241f463b166760190d536ae0f389458435affc737;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heaf8344b1fc99ec7c579c18477cf947d268a0de3f58f2bb92ffa42ae030f0f176a01667b059b9e6b44d92720a5df878bf722424f3d7d5d887fce8e720;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb15d34de539f6437a7c701d6c49e0ef4642ea0460b67533da8a63089fd35bfbbe534e4eab98bd40c96a2c28cbb3804563203cff22b238954e29e75269;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45e7f48d0379957917395211b0d01d93438ece49f038a8d62bd37d70b344ce82d6396db4062fefbe87f47d9e736e7584445c3ee53af75cb7309841c60;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d0c222dd413def367601e36116cd3e65498d2e87f3fb869cbe97580c1cce846e274d980414b1c5fae06cc73a96ef4a951de6c56a457ebd9dbd795f95;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57fd293e838e98fb4481798656e8838f50ed12f4295d8dc92edfe810e0c62afb5cc2503ced146cd70430424e6ba208b5a9005f7b1080b4981f8f2203d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcec1481c39b197d7fcf8dbbf07f203dd6f8c8ee08b73c31da7e194ec5eba081de08063a563a855c857db5f5ab05bc9ebf13e7c0944bd081cfa4defb63;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61d96259cba71c22b85590fd9c4a0b1c7d7d05a0e39183f5e68231d2d862aa1169b1b049a0337c58d321b454bac97fe29003a649eac85c456f4029521;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61bf7c245c95fdedec714e0efb7e4addf785aee5c046d99d928833907c60002990874d4d05f3c9c9a7a555b0189066417c04b147d95ae493e24039c3a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haae62d60657e0458d07330c438a827dd885bab3028596e6ae8ccd85a3016c9de8f54410d5c49707200220d090def5fbd704efa93b00c06ed0c0d02a0f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57b9f8bb39c0b3c988a1f87740940ed352180674351599ba29efc4b6b090ac1aacc2f59a6f830241d7c4dee4f259e534eb22a204f3a3ac0d403687b7f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf43f3e9450164d40d8d0ac1c98c95965bc025e2bbd69adc22d88684164b7d95ff4b5df441c737c60e7d64263287da260909d859769f8c0c908651c89;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f9fc08790dffdf7623d49c6c7904c67b0c5b05acd5b4d15f9793b16b90f3420bd6f4711a88de663895ca126b54ca0d46822e188a1e03b05b98b169fe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c6d450f4c5845ce69235955d2bfff9835595d4510a69c15d824835335b3064d61306a341c464f7d20482ec5266a7b62adc6bb5d99991851889047639;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ae8a4fc1f51c1023088998c9b244b40c6d4681fde2fd1be38ca5a1c3911e0f91f945d82e26bff75f00b65286ac334a9c8560bddad64feabd4a28d9c9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19cff0bbe6fd5c8c1702dc69f588486ee3449b3cda8b8de77e028841998d76d778dc601706a0ab52a4d8294b3c47ce91f8efeef8cf4e5209427623504;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf72c7a9e80693e57b26a9166fbbe1866fc6bc7a6741c9882a1d3003dff9695b1d82b73448361038d9baeb392a8a61d02b5cc96751150f76ed2d0d4b50;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c8d46f1b97602adec946bb9768b74750d8465dbee3448e8878ea8fbd836d4f29e9875e1821931dd745ec1885872fe461767b78e605715c609d100e6d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96b347ccb751a879aa2c742aa6332d99a921b3f9ca6057dfcfe1b355cde732572175f5fd624475f64ad8ba208c9563184d97bd47c0eaadca728c8a521;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7ba022d596c7c296e4864439a4933956afa55ac684b6a606535624a9f46a7c3e2c8dd883221d4572c2446635a443bd43652bec7cb5130a3dace19db1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf018fa4b62bddddc915119f2e6a931bab14ced9bb7a34f6af73cc77f1c0bfc1c47e6c14f17062b513248d5e032a3a2c9eaf9e0af659bf8c2d360dcb35;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a23c7ffd1d47c67ecb52a7a73c133fc6d624ad72ddd07dc1126033264080c93d894b7bf610ee894e2708bd1d45c592988e67a1da231f93c9c420a00c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff130096bb9bbeafdefa5697b8de2f353cc0880397ac2ac64daddc99ea1919a8f8465b0e6265dedb10aff330e0725c441b0bcdbb2ff16952dc1805e2e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcfb1fe12dcaa2708303bd3908b4490f7dae3d9c9af6b413142e46eaaefb6a3479de01406c7695d054c2327344affbf82f35b6c263a8abcae297375c0f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50351e376b130ddab70d1ec0ef7f91182630f79ba76fb00e60f589a20660249de866cc4f79b408904fe21dbfe22b8885977a4e86e48b8e6e39baf7b84;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53e3fc2f7aff387dbaf31e9dd01d7c90dd08c9d5edee48e22a0413cfdc8e879ae33fafbce1d687ed47b87cc0625aa76ca910683ef00826b359d33a184;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdea48cd206150379896326be67632b1674e32511d3ad38b9e9e35fed1450a002b868b93da1c58a41d4eab2d500799648fdd2f52843e4c27afffa6f010;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc342e6903c2b90a813c425c1401d5481370706d0b684559094bd2332f94836ff4a807cc3ef54ffdf380c06ecbe72ed7faa6beb5fde02e9e3134f39709;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdeac96346eed99e17bdf1a843754f09dcac13a4483062a12143db8d7b4e06942881d5f9d4d45c442e593b4d4d5cc09a25d4f7e498caed28785b091446;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57a43424e7fc9cb59dd0c355096fa779ceac35aa4047fa7e9936a85ddf876544a88fbcdd91e4c36f41639c1e74fe41c36d727f75b70f2ddc119f9d38a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7725073aa767de9878ef55dddb5d0fa03345dc0850eccebc3c96794661adbbf41a1ed6ec0ceb398046f4420cd3ab15b4bc626b61f46dd6e14b941dc33;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcaef3477d117f793805f745ad092fdd7713952ad487270dda96a6e8278cf0379773ae71e614085df0fcb7a52f4b87bb650169944b98e68dd04f758135;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7652f0f197b5c67c4d3410f13e7a3ca99fe2a93dcd77512071886f8f54d48a7d24b0bc30a99b84bebbbe6a13a0713140a1eada4316de5fa5ed46e2bb1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2733c3823565f38ace00c795bd9b38a9bf16a42029e6b044226cc8fcdbef04ae352a4100e697a57d75b6c0e8fd2b1ac2a03b7a4103361d4cf5d6d9ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea97a96d0a5682a3f03d257f828c29d0f5dd22a60b8553fda602e0dd7de2cb6734e60745ee69bccb107046549403b5855d483d77582f40c4051d338b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8abca9351566c9ec0b458835d05f6a224eeb93366540ef3e8d227014ed15283413bf9cee12524b887ee2a0e7d973c707a8d41250bb0b876e2ae79127;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hafef41a0ee9e23e4a37ffc37530aceb4a4bef85ed948e7d37de22215b4aa30de864e9ba7ef989eb7cae6cc08fb7614db0539508c5d0ce75b447ff49b0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46eecd9176e71d430c0443f620142e47c01d3f62a1e2a73b115ae113884a0edf2ac0c9b9b9e7310b0ca108eabd221c97c9381275a95bcff74bbbba3b3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a7e0092f9a041dbda260ccf37d4e3bbd606b9cccb9caba994991168c8cbdeea64bbc537f9f2bf166813ba44d669cd08acd8d507556cc93e0c14d6442;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b918e8e9e42a74d87b3ea50864ee7f6da4ff3b3fbd2061d2ac28a6e6443859b157a6fb9199b0145d86c2755f4bc400ff06029728941d557f2a83a2d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66ca5e3f4c3f2ef7d2ce79d8a119418c98ca900efe0515f6dacb045494e9155abbb1531c5695e8c17ce7785df68ad19035abab7ee09a87b75a5e3108f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb346670001b7b298e7a11cfa2f6c4800317fad44211cf3fb171f12f1907fd5831414e9057ab7b9d1e172afdbb33d98c0e7def196746d64aab8ab1c9c5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4868e6b8e3249d5cb4940d5f3e105dd3c5c71b1ab5bd926fce11a4ad8d9f799e51a1c4f7e62f7da20d68d4a7434f01e057c1ac6cd46e92596290dad7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3cd2d3e13921edf5e682c318730ff98e2ebe0d2236fbc7359dd3dee0865be1495210f593c79a6a81956738684f7cf74061af29df674948f8d2860349f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf23402de822e2845c49fd255f4f8341b753f8bccd627f2bedd4ef87e5ca8390cfbad749b90f63e36535136f878ea72ab9224f33af30c108c613b7cd0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0984adf58cc342070a8d052e5585899956a63ed4aa338ebb9fad1bf652b9bc8271556c9f978c6add03ffb9bb992270da06ed96de377a07e8e42985f8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd35b1d7412d998a013260f1f48afb0094f2ce8dc1e2c70ddd25ac165d2855c0650246f4ab1a1815a7ddeb03d27f7add2c01bfcf7f3116a1e4006bf9ca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5dca3be47971b0310e4051af140c9f5e8ff95a2bac6bf8550223b3f18cc6d5186dbef92b34ee35a7d3689b1d673df56ea4078ab0182196dfba0c18270;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdeaf50aed13973f79c3ea0d919d15d3ba21869de4a4b34517b06deeb9b6684e26e011e20060670e90e5af7ced14491d7c48537be764680ed9b83ca144;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb828756d3af2576e0fe13180c7207d005236cf8a96f142c0a910871bd59cd5e4340590dfb096b9ba9b4720d4845ae15644ad2036c159c849d66ccd3e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf0cfe5d9593cfa278e4704feb2b85bb625675a6d61320adca7b67008171d195922444af02e0a345876bedbdbb137df8bb3d81ab2ad1dab3e0a383aba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he51e4b998ea66e2bc040cf1e84c0b2cafab9af018fac614825514e1b5e01d2b68fc818613238271608b736fe0899049c7d6fbc8c35fe50a212d6d1875;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf4b7d8112b5e414281acaa1f062ae0654080f5712cfdcbd1a4d228e671d4f5e949abd130b66d12b448c13596e754a9432ba343df2b5a0ac02dc3f28e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18d67e5979e467cb56f20bff21605b0e1ba1a33c9ba3eeebcc4ec0e870c5bee2c137b092ca0e696ed6f8992d91663ee2d17b58329827f25b9f1fb1ea9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefd5331bfc96f1927aeb098127b88324c7657acdc26c8ba72562084211c9ca8e96a8698bd34c96e594d3fb580f9eef46bf33146ed4a2b75ad7ce2345a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4dd6c4c5622007e0bb1c36a350f7cb67dcb6e3f4219767864ed289491072af1027a4bb86f4dec81756b2f6b99027739ad4dfe155bbec2ac0d17aebe74;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38599454dff99b4bbf3126ed5ca50cc67cab28e699313bd2ae4bf5e913255e77e4d7275bd6cc02a8581a44b097312d6bb292a6313924a4804333be022;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f4db4fb7448f519a9ab07482090b73eca9e9095479634bf0e3d722d65c3cf6efb2e63b0d454c22c3e62967f4d05a32491dd0b3bfd054df158622cac8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h825dd74fb2c7059e079202268d5dc2e611054ef323d21a54197ad2859c375fb51a85fa8df96f08f2e3dd6558feeeed2ee71e3d43f8422d744b28b044;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h789dfa3404bc277d73477cae754cee895dd70890aad6b958317263efb98906f2333503fed5d47f551326a3a6ea3c95781ec11f18d246625ff0da589bc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6f92b05342180be45a965faa815dd7822692bb655dc76ef6464cedddcd221e9c7921bf6301559f1425328eeae7437633bba9f861fe035cf3634a08cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f206d64fef8a0e51b0676920f28a77858b8ae089f14b08e35fd7af264dae5bf0b887cd7a55c6cdc79dd9307fd531fb3a321bbf1ece7f6a75987489d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f51a3a3143416d554997f81665dbb337e6062cc55f1fe56f1d5124d3a3c9f4c80d60d7ac5d55e2af882690745ab79d703e083e92e40246b1ffbb3f5b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd437f41c6b6c6f7432843073076b28820c11156dfc0d4da4b8e259cf80ad9ad35741bf7b8b1228b76a2d74705dbdec48cc6e91bdc7e74d2bff74b0292;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4649eb8aa5bf5f929c20ba64edc2ed17caf88b86f6bab70d13afa786f937eea8eb2dbf7024acb32de6a10fcc8bf1eefa8b82a76c49330df92f816ca08;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e614d7c033a6051264fe251ee39e3cb2897be4021c2f7fa70c0693f2117ff1e2a6348e62b7f931fc02be4bbadf35d2a1332fa409ed61289359c2bcb8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd87a7f00e7a5b57583cf4371e449c0a6294cb128b99475a2fa34f61ff6a3b0123829792686d363d866608a28fcf1384bb3e7b6247a125bae3ebd2e1b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbde201b9dac615d8f19ed13c6ff4fe42b6b007bc88b3d5294fe20b636e93c2abbfb57880e8ae157e7af80fc0a460fb3c81ffadb910721f63e93548a2b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4eacc1b7d2611fee8dedb18cb9b34a1c98a2c0cd35dfb73d1548871329beafa1faacdd8d83318e5ad9b80071f812fb66e705c576d4f4e5562fd13ffd8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfafe16b3ce14a1ac8616d1424cb1d3969ca7e90c1d359c6b5c9524df0f364b0c20c84fb04c285e903593ecc7e433616e647f821447d388d0adc450d5b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa42bcd60fc41a3ad694a720a2e0728065a1fd5ce2c74e8f5a1064e0eff5f7b30b9173fff1f93cee19f4b392e762aff357946c0fe0cd23f59e16c9ccd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h663ea7d3c4cdfd4c9f1a3db7310992282fcc4e7042d2bdcbd1e311c1758efd3189e88974c9f77c47c3fb6fbbca4247f4697176c947b3aeec49ed31b81;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdd93f08af049bb721b1cc51679f464f9773797fc6d858d5ded4bdf510749ea3c47cc5f50a9059bf30c927b827920cabaa08fdc6157e46b1fbdd8e997;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc25193e032337c65e7eddb8011d500a5af077b9f2fa6c772b216b8c3fce6d4b42a7dee318f468101751e36a9a2fd38902ff862d005751ad268bf504a3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a7f9b3f1545ee9a8b2432cad2e743110b5c073259b1babca837c50246e569dfdadf407456c887f682135f1df2ca163e9ad721fe9f27c37a12608614f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hacbfbd6635fbc23bcffd5d2f750e89c5875490c26971f059a21dbb24274425897bff2271aa9731f583f9013baf68d4e749d0f528b0e5eb709815ad820;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb9c13a499ea6aaee31475f311d40742a927a4d7acd6149d4d562f7b9464c64d4d48f08230e0dd996536b44cb38e1af67f4704ebcec36eebd70516f7d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd67ee5ba2cc96389696fc04a863e9926be1b5a0f3daeb01c6b5ba7d652dc3c83e5195ca2720af21f92f8ddee6d5eb525e59f699a72782fd64381b181;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b7f664d80653c5641f35bcadb347937a020452e24c72825d2b022018d9fdda181280f1243f65fa7f579e0ef1c47dcad602d006d17a820cc1467e08d9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2439e4641cfde4699660395247cc69bd732d40b8ce557c3108b4c0a5ee074481c192f154731a330e526beddec87533b9b3956a6094343ecfad4daadc1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f84db34cecf2dd797559cf83daf81705ab794198f03c1d1d8e255f160dac0f7c09b5fb746af307fb724f275806866288ec110abb0ac18cfb4c82b114;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf47ad88f78f83f095fd861725eed24b6416fe5847dfc1e2d6326999130cbf12635c77a3afdaaba0606b5449b7673cc31cf5e1197118c5d1149ef6b2f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h594869541e57d7b93285c37fd9fdc9899aebdca1a45e1db09fb3cf120320383f8adf0f93bc8acc0e92d893035194d3f7a15cc75b95b46c13011e561d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed719a23acb7b2a516309332ce58bbc5d61f27604aa579b36b5bd6aba82687383ca75c42e4af47909e133253fe0b549f402a0262fd250c08579a63cc8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7831c4e2e5885deaf83bf135863026aef5b72856a7f7c3e9ef6a1858b0e8f3541695043dc10b59e468e738b3bdcd4727422330ccc680fc62afb1be31;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd771cfb4bf0af911a3e35c4854b90699ac32f709d46d49ab0e628de3396fb14b74af7d5135d481284a1f97d28b15390cf3b683fa30e8546cd1e68f621;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22006a0433a3668bb419a096db143d59cd5c001e2c660d6a03d859a86d9e2a2f208d4b2271a5b5c5c312c9d1e45f6ac527bde62a3238a99e988828cc5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he1e0ef450bb77b0956478f08a7b77e281ca860912f4e510f0b3a39a7e0d4595bc3984fd3e770ea096c66a848227ec9ccaf632c9a45b4ea714492aaf78;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc77020052cf7605e221ff3fecd8c69fdfba8c9ba222a15fb1de58149cce5e3ce1ccdb76fa8824e3dff3420ab352909d4204b6c2348ff4342eb8baf283;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2549ba7440d70fa635793ca0332ce60dbf797c0cfed021804544746d0bef0dbca168fea0b3a30157369cbc964369def6d550af1cf24e9834f9cd6d36;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbfd11f246c234bfecf7837a39a8c83aca088c0a78d571af92def26b853583e49d6b3f38773aba09adc23390d624c6fa4ec512e726f135ae8845d5b150;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h212e63ae291d2c96e85df2d52bcf1f40766eae1dc32f4131b94e527f188a55f003252c8f7defb168e5727c3e30eda215e3d0add8ea7aa36233e530f9d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83ad2d101b91276c2116050a8f8c2fdd3448a0a3d5339e62b85e296a603f0f55c8bfe1d0d62bab904f64945cee3a7abc861dbc0932e212aa0eda45f98;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d1002641b8b82146784fdbef06bad3bfcab5caaf35da23802dafc8a3ddb4b0fa382bebaf48f40cd59fc4038d51c2f0180c24919f798e2e2ce4868e13;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd407b842fa66fc6d88552980a289e480f093cf618a080d6467a82a30bc996f0f3751640378ae59abe541f4151020e235b1dc2c1e557fe2e3a6c6b130;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb49255bc00d9038b9ed6381c5a94995be290797096d6219eb2589080a484fb79eb989e3e77046f331bea767703c658de20ccddce322357dd8923df1e2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cf4d3ae073961ed843154e937f17040d11548ebe90fc1843e2bfd735ad3f6fa370f007707dc6f145fe52acf675f6380633327be6514acddb6413f25c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf43731e17787b8958b0b480948dc0b67bbf407c17b4ed6804fda18e99ba08c8fb26d736192e23202b9b5b3fced1a226232e41db628eb6cfd3b685cc26;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0324e1a5d120e53ee3e18d7d558271fb38d20742c96f4b236c9119d8fbd440fcc0215c1e5741cc1f28a8c40949cc75d690f436d4d5b8256a6e4e3cea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8539ecc56c4954b014492ee9032b2ed6a23f648bd333e94058e39f704de4935eb206153ecda892e5ef50b1eb8f9820c267575e6ab2c9c8042e3794929;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2568161e77fcc22f75ea91fd7dc4cda3b213a689af1fba7b9293b80bfecff2a97c40cb3515195d2302f11c329935e4b2c6a31b8c907e621f49053f52;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7a482336ddbcb8ec897bea1b91bf0b1daf4c6cb4db8672d92fd43dde126be16ab359f7cc3cac4ec52c5937b6d1f0ec8f808cb33b95ce7b9ad15d9a51;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13a316a29c6bb5641afe6080c5fd927399cb46210dd2cba922a3e875e02b1b4b1e06b2ea6eb8869d4def13ae79f3ec86dae8d0ff0c59533421b3e1498;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hecb0cb8c20168a0a5155aa598c09b3c850f67d0a5692016ab5c9acacfbde77454f33933661487883be71510a594a629fc1aa6729f31244dfac971c6ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9cda14ece74a30edf587ac347b0622ed54685f1ef1e948593bb6a0948b109de24de9a6b18b2d8a4a7553f6599431e192bec0192b295c324a65d32f388;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb6a1eb2046404f6ae8646ca8d86821e8db97b0eeded8d087cc5d9b785bb47b22ef32cf04814a3bf39d10bc17b186b0b7dd3b095ff2066512ca9f5ee2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c7d5f3800a8b2bd02015911cdd9c2a2d70f5f5a90c787b2f6acf4d6e58b91086725806c511b8530f004ee3f3073a3f2bc9a3aa99b9d4bc9e94bf8b28;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc24628e8f229a61258fe3c1579ed579e39580479c9b345a94995663536628ec220f4b38b0e09c16c33ca9d6ca638fc3a4627f56998dd9e9b8f79b6384;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe46398c0cb3dfdad53254a1310969cddbc359cbfcb3c9cd3516d81ba9556307f56dd6d03f8fcbedbc28f1b4be16a625a9b8d71abb844f9ab35522e18;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefbcead4241cfd78ca419e931ce14bceba9a48916447ed8b0c21c787d617fbdeca1f448de98636abdda80130b0e5c37f0b1b4747860be0223192d5aa2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ff0f0353816e6b71bc485a8154a9e3db05a26e46a20d239528c793cf9f55d7aff1754f5fa288cd4c959ea915925751fd3d170f2d850d62e87f3b35ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3882a65f2edfa858f5e469c905d19ea92e6170f24b0e35d153f207159245b998a844eb6f3bcefe9c49c27bdf00cde3245af5a82a559d4a738c88c996;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ce517fb0b5b619cc3725548f0ef5693344bac663e84c20a3bbe9075d2510086c3fb6559baed642e73a4479d146f3231e2ef4c19e465f37abffdf87e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d916358037ff2fb12ddb60d46ae77209d168bced5f9d1c9e76102404eb8b8614ccea9c5ed529674fdff1b5f38ecf9b5ea89923c5f269f0cdbc59fcca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fdb9d1d8f4f19a3f53a426beb822df2c83f671beaf7323e744bd7de2d149a6a3af837b4a349aa50e6dd4d93bd197c531557b48dbbf34513cd547ffcb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a398519c7a6a08b400b0a8d84bd248d42678780747089408982e164b264333b7be6ca680e03465ab51cdbf016ac37e6d9d761b19f474d64cdeca15aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c67c2c222a1d3b0b196ac3ed95f9fb03fcfb92ad68cf8d77bb0dbbba728b820e0cc6d454471652ff548ac3fb06af5145f646c1b4a983f08ab0ff1d89;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0adc3b0e1ca866987983a9671df7f82e2b71b816903f094badb07800661a369998075f1ac74c0874e76154b8f2d647ae34f255511ae0a34b7f828b3b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac5d8db34b3e36685dff62b640a0d71026ac3a7e2de5e9aa4b70119bf6457636d6a38f500e17d052548433a5eafde905adfa0b02356058080e82a19c7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee5e2b4fe4331ff369359c0dc33b284592bbbe605c159dd950b857bde0d262501c18164faf14de4422468b25d710c9f7f5955034933edc6609ca35cf4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53d3f98ce38497af560c074fe859a254c0713272357ad992779705ef89d6c7fcfb90d740a7181f89eb848beb23d0193492b3ce3166a8cb83992df474a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f67bed2a21e1b4eee3fa4f923a3ffe5c96b297b6adacd29ae77393cc7c1f7fa2f02036820d128cd613962755b13c66052809b5cfe70618aea5ff43dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ab41579a692d21aedaa58682e1a8d54a39d8ad080be655807c3f605daf1db4665699f62ee5f558c5d8be4b1f5d1cb70bdab9672d6408e0c17ebd2df;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1eb54ce584dd3542e8e1932762f6a5bc9f6199bc395f7eda884c1eddb26b9933747cb69445e791163953efe0a0bcb7d70b5e5b10a33486b429766ebed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b37ddf5c40faac5897f267138ff3d44a15203a49ded0ec7cad78db003c721910c6fbb741cd7b604a2129d660eedf1c3325dd6a838a054ffc85139d63;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h688ba19ca8dd49f6cbe063339080b49a4a40b121b19cf5fd6b200ac0b930f9d2aff14b0f97a417d91c6562a9ef09820c5178870a59aaef13d4f703c2f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf196d578183cbd91af167a35e69c5e8fb6c3c4651b62e731025e5c755d40f9373091eea4b8c84d3a4a8c8dd993092c1dead17321c293f2969d088c2c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7294b11614bddb70a295d8892e4364cd3551de80249d4efea6db8ce2ee741366b22453dfc530f40607f93e8470425b5f4a82f31faae1084a0d5deab4b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27eb0dae481c978058bd2531fe076229485ca34b35d11ccb810c1983bbbfa4290dbe87baf2b4685abf2bd93a2a553dcdcc1703db92993efb73f1e9cf0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a6c85e63c4349376bcd215ba2251c36d1047f2b6d65147c5b10272b53858bae9545eba38f67b4cb780dfa61d3a9e4f0ad376a798a2692e046dd13985;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he728a383132018c5749ab8e6da06512ac8f14f9d0556d2bd95a736d6501dab74388240561890b61f3ddab6d82dd84ab2994d5c5a4fff099ec72683da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd70f51fa80d9e5599d3e1b24e00aef62d569d990571997fac01300451dfef6d2c6a58469f27158247510b38c8df09f6f2a444b8310a692c9caf95537c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22e73c4f06aded51c3a64eec2ff4bb19ed0d23fba91909b89c0782b2c9a472f10a8737186a0f1877ca06c0cefaf5fc6051822460db63604477dda5bed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf1554c817536b2600ed43a13b3656d3c6acb853c27fbc8d187f33a1b4fe8ac4e130a198a8e5d0a5c017ca13bcafd237d38506379485c647016e386a10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd28241d4452339db6e50e1f6bec0a114b7c348f8d64b7d69f6e5f35a313791cfe5b54a10bdbc81a30b6a38fd8ede2472eed09de7c382bbf27f5fdff5c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84e7350ed0e0715b6eb895bc0551954768b83b51341b09c8ef964d633687de6cc141262316a606fe6d91a3bc459f62971576b2b17895e7da90ea45a2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4bf376b7acc3db30b39e9dbdd43a695a44eea1a42403f9252c656b2b74b65533260e24d4d6f61cd11bf88afd50dca952a472bddb6fefa5c0b824d7e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb3330ac99fc78f8892c39f17234107b6fc2d822ff9e4544716e18ef381c780364f6e77f8849ba91fc0ca8aac56e7f092491ed11912aef748b20e46cf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h444ac3e2f4ee82d85d2fecbd89150cdb9a85192506b39c6b16fc9e422b6f7f7a60606a613728f74585ca86056a2ffe580635d1d182fd7fe3f183f7181;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he19ddc8e13bd6b4d300146f339dcc6cce175550dfdd1f7a1cbf3de66abf453ba46cb6d0b18568dffc0c2f1ab44b1f2ae66375be4cf8e32e1a65c42959;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4cb3dabf123d5da6b01cf6b672f48698055567c20cc6d9a39aae175c5d8e52fbfa045dd85ed93faaaeb038a0fc5a1da685a563039898e58cda35bb03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h266053309f54c537cfe79cd446a2d0bb57679ed9f6cfcca8ccfb773bdc62e67c95ee25b56c37d669d33c6e7064930d3705bac42ee1b41ba09256cbf83;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22f9bf89a8505aba77a6a07108370b968cc4354005f31b8b07626271c2d47cc40e9c92571da357bdc05d97a0777e8954ecbc9d116cc4be6b9e27e16b9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ef3e16aa132b1fca94759c55f0c3c0aa547407a84e342ee02f05d0655832bd2e8bec82aeec85437bfb319557ebc198834c3905348902508cb89a81a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a6ed832cc308d4e7d3231e84036dc1a22c4c3477c7fc7a019ef1d11a458678b13221c66a791c8c6e0dcad9c41a0acf8bd3a9ce77b6b4610f7df62a79;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb812f639fc644e3060a6e74f9db238e91ad6c86d5b2d3c5629a40cf3a8bf62e29075570b5f7fe1ee268d42cff12a22953cebd7d2b8e469f8868d986;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2f1b9b4b2fcdfeee2782a00f9c8593786ca65970b660f463b9f5adae7e501edcf3c3c6c528e0a7f78fc7ad3b4889bb493ed0fe8bf62985a54fc2608b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h338b1c1c3ab3583479870c22cad79553fb9a18fe7eef83d86f239a9887df2abb871ab4aefcd8a32a4a234798aea808b5a662492bad9b24de97af7b0f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95403fdac1d792826e680cbf3dc55e26318d8e72253219c3c87b7710cbb8bbffb8610924c2554b193df40e90efe37352bdedcd1eff5231efd092c3a9e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b831fbd5ca2b673e280de1cdf8a0b1c1dedefda239139eae5eb2ca03255449a82ac6adb2f1ad592c6006d697301b94e639b3bc1d299e7f5d8751e9d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41660312ca650d742e7d1b7d4515677dda485c70ce10cdd1760e15fb499638caee4f140a3aa61501559bbd035ca551a1a4d2a71d942f58eda72481a86;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19c499a11b4698e338802f9b698f40a5bd00b751daba956600acc339f03fd78ad32f4d072805b7ee6fc8236d14d6397ebe16e720b20fc12a3bb078765;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h212179f9b722d2277071529896789b389d0e8985490f327bb6e11cd29c6e02f6d014a9e76ca3ae3182b031b44ae5a429547e869616284312184c3702b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h687457a65796181248b33f6e8cabac6823004204228983956dd36a8d41e911f243bd4146dfdcd976e0c0136b0e234011e9176286ec85070ba812dd46b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd076746e438db56e39273da4033ae5eadd272255c915bd87e2ec494f8f4ccb55c6e105d868d1c8e707cbe1351c4ebbe08a9be21a860ba49a0183c0524;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d27ebb3e41c9ce4ab0a96fb389fb94dd4e5c2485e9607ec12606826da2608f4cf873ccc02d628bda2f0aaa28e342e2b7c8be49093653038fae0db72a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2eceb0bb988c1be0b09600f2855da76712bf042616a84b5de666d4a696019fcd978413de21ca5f8f1ce53308a9a7d8108e953a927954ed194dd971966;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde7788e7972b9063162bd517d491eb1315deaf1ecbbe4c3ec9305bfda8ec86e75a254c8a925961e48e34ef718362a61416ce2aea8499dc871b3717310;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h965f288404f707e12ff23f55392176feab38082d407501ee18ec62058a6bb28b2c1c91034834f255b7387c8f9e187180b836033a1d7b1de800d30feb8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb97f346a1c0ce95759dfd46e2585ac15063d4fee814767d46b603000c7118dbdc8242ac1f830d207a7faf1d476005e87544e12393e30cf9f5941b96ca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8147b337107e1c45a3b72c1e9382dfe5c41497be1cb23642ef4e1363c6813becf8c9cac46ec2c97a4679033c88b2a107604d6238080c269e6e02daea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h847f4b83b9f936cacc85a3c533d9404efb47aebad91767c1e4c60839a459c44fbb726f5b97f01092208a3a8da55004ce6d1a9ef830e6dacaa5ca208e5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f32cbf8637a3755683acf860420b5d8e2d150fce2d389562169dfcc28d8d00c0f0ba9eebcc826da44148cfcee95f5cdd12bc132e902b97fb91c8540b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9b0f1824b89b25d4e72e879bcf6a800a7fa746e913b16424e777f1c2cb626d60e18b8eeff6d23ae094145f037565481ef59eddbbb96980af4953bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c7c0023b900c4b7adbd4b6d3bcc05ce6a8d27a8da812f5731fe16453b8e704a344e6c6023318a49238b2dbd518ef3eb4455f3a6ac34675ad6efd16b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h239e21fbcd01e6d2032cefbc8f982c66e5ed9bb308fc178c266b7c52025c020ea264fef333e35f7f46d2aadb327fe16da4ba9643ff05fc8e94aa0e96b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0a114b189524a37d4cfa9eb1c9fd0bba35f86383e67ebc22b71b6ad063a9294695aa634d417143dcc0c6dc24804672dd6d303fd77355733a94f37faa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52c6ffaf874a1a62fcebe79e2a0977d5440d82c0e02b225aadb23b06e6360403d909854d516f642fe2d1c1ebaae7d826804b2200fbe0642d3b8d7d046;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d68ec2004eee9adf2d64fe85ae1d3c3814f8477db5d41c1aa39f583c90cf6f2a0f46a7427c21cff2d01693f78a303904f0995dd14bbba5f075765c49;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc27e32535a7eb221c68a7e2ea1766dc7dd270f98028c8f515337ad2599a59ea4a9fdad1be767bcee9c3f0de7f21e1f32acb62df9f8529dd61cb255947;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f89c5113af11e64990f325de49083359bd6437dfe6f25b5c6dec75c2c861ade491e0c71f5e6d0509e4108dd2e16e6a8e45af984937f1b165aafc9420;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40bf28dadbdc61348701e259aedab8b530c550dc3241917f29bbae2b9f3d6cea9d9d24ac4d2137f16a71421c43f9dd33adc0f6f451fa6948f59bd2430;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd403fd938c3f0ca02806985542b581eadd309cb77268e514a08edfd56cbe7fdb651261e9f1e97e57bab667a67a51e1670974c0f729678fe4e6cacc3e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha99530517c975dc6e5bc77cb850f45cc0692783d146cc7b91e0c6b0f5eae62c9ccec11075840ca8c3eda5e83b990a8b2716ce5e40a2d97bf27d2fdda7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda0671202f5463e932f124dc99053e5b41a5ff2e89c53a9bc7464387a153f01613c6b5cf6ac3ae5c8a9d0ed04842a8472dd454e6fd82c6289d4610f94;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf4c8a32a4843cecffe219626491b755c024228d982bcec3bef76ac1170d13b0da8dd662502d929ecfa29d61cbdf7aff22334456e65bd1b0d585c7474;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf933e87ac2057076321aae9c74c71c5028d4b82f319e882cdff82ffc7b58af2d0c4a0f3a142157cccb229e65f169429ec69e084ec5887d84f9c719c15;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19a7900b62ece0cbee5fc9c9f5b594c48d53b0ec8fb9564f95630a7b626a6ada3e5c070b14e553f1db6b02e103285b57a833325060c33f9a61303be95;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habb2384caa963400d293fdfbf8b16550aab71a17bee5e9eab60c4649660ea4a591dfe1f8fcdd5b29738a6176fefc02b40434e0e8212417fc29a18a4e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51adda4400857410b4c903a442604976ef3f29ee3de1d6a39422e71666946c7294ecc28c18453942bb4f235b677ce3eeac4a5a5a051361cad5bb2d9d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f33ec839fa5a5237a7c48db97dbe38f06fdc733897220baebcabab845242f4d6c646b941eaf4504061aa2a4828b7c8840432261f1117b5dcf1e03d83;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7caea71b2e0667ad6a8835dfeeee06d832ac13164f005f2d2a2018d719c5ad093fcc346067bda2472718bc39927dbd256d20ad6292aa7b7c62b435c80;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1fdbdffb61dbe1094e32bdb94dd24e94c41f26e067d7e026796d98180b02aaa803fcfb5ae409bbd6955a45d1f62cefd117e3763b9421e6d4af3279346;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4923af80e94dd8b738e0c141b0b0a47b917e3a45db49400f4abd3d37784e58ecae7fa5054f709bc2847ad872022da54c3d7f7f070f4d236f005123f01;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haac64e8f33d500edfec460b79431d3947f313eaf735b54c0b9c9a479189ec5378fd403bf17a5244053cd13e5a8a7fbd0e14272364f03196e0d8cd9804;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9536f4b084175d3293f2df01dadd07bf43ef34114c23b2486e2c011490c07290e2a44cdd3c1a14d743334dcad11b292dc9c3ce00dd4d146eefa96013;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h213614db10be55d5931e83e5ec37f20aa288941bc634718d8c186a67e569e88fac02dfc950f68debf1b047760dff2d284171f302b2a0bbd7169f80e7a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1dc44d6a159af1611f4bac7bcf0bacd7c33746c91fd135c5600ad4aaffaa30d541ab0589201011c85e37025f6570f3b686d4ea97207c8167e06e7a88c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9e091c3f74024cab9878afd952fd840ea87ca5e8b27d4207a667e1da3476dfc43bfe2b74ad9bbd95ed89f97c7f4d3a8c6726f5ff212bd0abf1dc466b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h953449cbcea645af6165fcf3a7b3cd9ef35571f458863caafad309dd29d790b80e6ee316d496353564a1f1529cc220e0234e207e15d349fd8c29a024e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50818631d9c34af1eb728d5861d6a8c14a828d359b824050f93539c68af427808213492aafcd5c32bbb6571d636a8c405c1310bc6bdd3c2134379767;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a9c913daf001c2df3b7d17a098104ec5f5ba6cbca19c228be445ebf0bd710980874b04504b762835b0fa040df4bbe8f53e2acdf7cc67b8297d84af0c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf943a055def4b600c0cf630e99a14adc5f5211b11867ab8af404f1b99329992293fc1d9dc32c2a863ded4879816a8fe61de30687a84ec6ef70667dc88;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19aa5725de1e30251c81388c8fdc86102ce8f0e384ad2558210fdf86eb3a3d162d1f21cb90acbd11841ddf6c3a90de75c647c89957bd530ceb46e0f89;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee6b8f9b2382b4df6bbfc3751d7edf35b033d8607fbd221bbdf09c90824adcd6c5435314092a60409d3c4a530acbd4dea610774a7e956ac442d95612d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7909f0671bb21a5f10127d3c6c8a5d0c7238fff47c0f2bcc21dc315d1eafb5ca465ab63b6675aedd5310f82b77763fc83c5841f1f90cebe812aaed12c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5a5b2def81c938c889b2c5448597ea774dd4cb981a751644e0cead6d5764a03f04457a6a2a8a6f1047200d54105680b8a0cfa4c731b82af6287a917d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc9db57a0358ff9d27381134250072e58dc8f3ae814246a7d0250f3e0e5b8bc62cbe3b695fd3af28617db4c2a150a13ea7166c612164a56c5d6307414;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8a6092171160ad427c6b71bca7ae25809a7dc42a4cb5fba37a15aa95631f1c4b32eb6270a4382bb3d6332f0d970621599a7d6793e92286ee5dd618ab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h430525fdc6d3819f28cb45e79eb6979cd6a9d1c68ea56e66c1ec37c693dd4358720c28b2d4c5ba8794e299227b04ab51dbf2a1c127b582c98c6e24333;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c0410a09c097bb2d8eaed7ff699686bc654c642ca87266fc28a0a865ab1619d490ea20de45051d5b0cf34a3f171c74cbb37a8e884cb3d3b77aadebfe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h186c84ac3f6302e60ffa604ac8e06b67eb5625dc040a48d84111945bbea68cf54b3eeeea8ce3bfadfb327e59d9f4c591928e00f221f50a23fb60ac823;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h629e9354ba377be6d3b8b7cfd7728a264d638ddee132b83f2f8c026c5a35461d48fe5f5d1ef15c391e13f7ddab8800cd4811d31f7b62eaaf3931a0bda;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h738d15382b1efe355ddce4ffc490ad84f8a3d4a31c5780d3ab6426f530e593e01c8c0e423110d118fc75ebf3543e87862a3513fad117bd282ef432825;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h965bb76f79d27974115cf417d299a9346980b626a16b85d792bd6611539b11bb8320430026c4ab32f426616d35b71fcec03ba9adf66f07e6ed96682d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4470b9d521415d559c4dc46273c46b8da9bec61135d5e3751b87853b255e6629e0373314ffea59624f7e8cb1eabf418a85c7c34491a7016e8075830a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79ab5be78b2b3e6f473fb125460ff14e5a61ee84f7d7770e3ba6192cbb35efc5211dc7b8f303320cde410901f5d6788807df62f3396b407b9c9c71a9a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73ee868f540dbc05720783126a7e00bcfdc220b5361bc118490ef167e2dc58de109ef4f516effd7586a6fa30aac6744fd29b2625192237a59d7480999;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92561779605e39acb0858fd57f123cdf1fd876ddae5af3c5e69b3c2735669f1ac2ff6482172d1e658beff084dcca4b47acbd99ff83af14fce36a6ec13;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42fc9bdfd8f76a169cde14ef99bed3f94dcd480bea200442d0b8bc868208ddf7cefe0acf90daed8f76617f9727ba46aa89a5d20433a1871454b1020d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49b58fd5516c3a76f083f1dcc209c4d1032b5b365dfbb388e08c8d4130fe2258ed8bbd1aff3eb9e25080748decbe9f82227c00255b2180bbc40562a58;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h477df50f8a1c1e789d546d9353959a390c5abebc9a751f2a4b361a020319da96ed98064ce06be0d6c185b84f69234a921b386782d553605e53b10de5e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4666efb816fcb01d6501be6c7bc747d9eeb89455ea01068877cee32e8552cf553f390fc2d458f4e03f887dd5b1c5f044966890b2d42a8089cc9e8c3f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdde0ac4b7b5b14b4c67d8d57b36b04a140a5a660a117e16d9c0ac588cbadd01403e08afda09c3a471ba1720a834a6bd9a41f407ad1ac35158e773050;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52d03891a3ddf11d73f8d9b4042232c578f2d8c6fe75542e6987ade63b145d73cc92258445299b234d2f78ea5b3c66b901c4f3236ab587956e9919dd6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfaf2b7df02820052946035e30e1405c40b4bd0e08207351e080d046350377ae00b05b35000b39ede75ef0cb2f9b3bf6a4dbe913bc08a775ac187b6f30;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94518c887f2621779ed9724e7951a96185b34a3fc688e44887dd1022d501a79d4a2c3d594b1584b925a21fde2f8afb50b9b4257d9345b68a68162901;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58e597e8dc2211bb21abecfbdd6c393d8594bd6322cfd8072a66820d985a63c20ffd940d0ce4660ac24a3e60316a353586578b4686d7128223694d482;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2589fbbb601a4a23a5a2a79b1122599735f61a80d42b13532ed37905c8ba33d3c224d95c085ec4c781e004bf845b6843e0a51a60d22fcb26d59b4eabc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfadf14ef20781db96733ee4a2c6f027e528828552be33852081e860485279e8d30d4e507602f10fbad934a817f891c6313447b9d1a22c3115c7b37f91;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f14b49c36d514890bd8fbd2ee75dd7aae534f828e2e1cfe06b7dda6fc0019b0680c7a6654e9b33271f25d6a6438a73fdcf7c1c11d7749ee676e1a9c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5043463b4c2cc9304ac2debf8e04854cd9ae025456b05f016d9fb948171318b2907a506a85bb95221644abda33469dbce0272f0be333e3be1473c0cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc400b174f61b5c2dab4ca9e6ebb3d5bd1e7a4b8724965948a929a0f505561cf036a0ffb240eeea8575cd2721d679c36d5c8480d21fe398d600982f3f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a0b7aa41604994279ec3c0df144cb110565bf0d378ed064165989920d5dae45d700372fe047e6fe93e2f97decac1e4f464f45f102e5c3fccb1b3ce54;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf76d065b70b7a1de888c6a9e7d43eb6d657cee369405d626b273a0bb42e20b5691b178895f9bff8cb03b8c5ba6eb3706a442ae0c150b6b31130f2bc4f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22f77407b79cb8bbc6a9ac74b4af2a63404ef6209c4ab45a65aa88bb15a1aab78a2931501e941a91ea1db455b86a2bee90b91792f5daccb231bc75dd2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70719acd28cdce406784d166d7db9ea21ae7b6a02ae225f2b71baa430990451ec66640eea45e12b27a40f6b945064850e78bd28443f54b6b503dece8b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6809ab0fc635aaca60ae98c7f03f39a76e234104f32452f8fe7e8af74158688dfb9bd50980b6db59caca304a6c5763fae60b4f40499ade851336abb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8960e5c6fcf1582f01b15071521173af734bb81c9cf4f9d2f14385512e6b1a9491647ecd585fcefaf904b408b126c2b2c2fa77c99cbccf7df0397f3ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae7c43827158ae0f56ee4fbbbcbb47dd71459b369050e9f96a20552d7d59eea77379bf1940f6cd91253d1dd9684d44eb7b104985c2ac1dec75b3d10ca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcda97d57a94ef93e5e6b8059970eb680589641fc24c152f53214218b176c2e22702cdbd665d4cab607ebb884eb64eef313cce85a6000824f72b558bb9;
        #1
        $finish();
    end
endmodule
