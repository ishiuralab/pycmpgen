module testbench();
    reg [23:0] src0;
    reg [23:0] src1;
    reg [23:0] src2;
    reg [23:0] src3;
    reg [23:0] src4;
    reg [23:0] src5;
    reg [23:0] src6;
    reg [23:0] src7;
    reg [23:0] src8;
    reg [23:0] src9;
    reg [23:0] src10;
    reg [23:0] src11;
    reg [23:0] src12;
    reg [23:0] src13;
    reg [23:0] src14;
    reg [23:0] src15;
    reg [23:0] src16;
    reg [23:0] src17;
    reg [23:0] src18;
    reg [23:0] src19;
    reg [23:0] src20;
    reg [23:0] src21;
    reg [23:0] src22;
    reg [23:0] src23;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [28:0] srcsum;
    wire [28:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8653a8dfdbd65ab8f03f3b2c639d28ebec9eb8a3819842bffa297e5dfee9a61ca40c63c475db7343f1a7c4d8dae0e57217d6cf75b9db07528a07be5adcfa11ed76800f85e6bfd53e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9aa1d7a9daa71960f31a0076f05cc7b0d0375d97e500477a9228c943926a30de49d8fd809728f5c31f40d9bfdf77dd796f1cb5ebd5666320542b57cf23e9e60d6907be933ecf988;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa1110e7e1f12ae142978aacec963f140602aa904941606da48f9ab93d06777a30fe745bf9d066dc894f654e8f3209d0f2f25eb7e1c66613639ece46162767647117be351a596ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4425e5f818bfcdfbd8ab250affe43ee964f768fe7f39b7007d40891d7ec17f8e8e25ef56de4b01bb44166dca9971b7ce8b8353704879fb0a0cab4d9cf7b3625659348d1c7c623ea3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cfa31387da37207ba43d657b3c9342c4742b1529198752f3c6f8452cea3359986cf58e786e6f6ca1c234b6a4eb6827e840b5f7de929926ddfd8eb20a167aef8d7f64e66dda491dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85cf5fae8d3ab764998b4556363e2339e0d396dcf30117cff17864b4f6584879079677beee0b1b4d7d4753e60ba3692e5303c4517d0fe4ad31ea792a660764732ea686a0c71987b5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9684d15fa9b1138c9e32d2c977b9f4b399473b0849c9197f2de8085801787cb8a4f605e5f5bad220542e3b5a4415367e6925c24941608ad3b232b797160a10e1213c226e70896a7d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2239b152ed52a651fa11a7e6ec29a1699264862a38b99c757390da220ba73945b5a06ab49cae5c14e43a6ed0f12b9ec74f48c256d2998d47ce3143801a8d26e0fc374befeddba375;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf8d64aabb5b38d4e7b7a6d40cb380e1292b5f30267352e8e2c5dda9b70574d29a25bafc6b6daaf5cc37cd5f3140b28ee84f4cf885d3f92c5d5bb9107f5e83039bb8ef947a92531b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e1b3a320623e19abc41fbe5bcf647cb23f5b3d575b2e700b64f7ffb6a04490f2971c650c0bbde1e90e52bac1bd8c5c6ffd84e025b5ed321fb31bb9f6223555d8cd8992731fda784;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8dcbc59bcfa930d8b11a1ea83ba42965f45efb05140e3f7c717e9c675d784c1b636595e8a9597b6bda827380fb8b3288598c26ab46f94f2e0cd45d5f1d7a37ffb55decea5b355230;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d7b12dbae5e4b4843b26947ee0188ffaf480fa4de50702596d1da540580103f7825605bef62dd3372d18bf02740b4684f0f8905a0cf2d4ed3940499bf7ac8b681cba2bbe1082bce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4b82aab8656697cfa064284027672592add9352206aee09d71ab20acbdeb9f381b831d545ae530342e82e7cdfff7c0b4646cce3b932f31e54c5a2f27ade2d9106f5bca6cacc41d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfe51246b1a321f255853b4db6bb353e5633f27dbe9acb112e0678200a2ad0393cf44f4746172e5062ce26d8837cfad4397dbca891c7b5ca7dcae05950ced46188442263c21aa8a3e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h128195bbfe8b5ce12f0f1bd01fc25111734143a156eceb264fa8740199b86c3bdc3883b7592988310d765057b74f993db395127bad2bd5856111092479ac930f184b4c286b98bb86;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5be944c65ff117043d5c730109115012719fa945eee083b21500ec0bace1150dc060f62bbf7813c81ca8521bd88cb2066436ae3bc243b4e07292d6d24290ade25493247107d8e86f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h195ddd9692ffec084c3dbcd93ad7060df7e6d6eb5adbafa896b0edf856a2e491c3251dae970847d0590f065386de986c32ca58da55c7f5cc29204fc7279b57f874d3dcd4079960ec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb8bddfb5195832056f9dc84e5c972ce954b9dc6bd08427b6f1ccf7a9e2c7b13f3b81ba23a71e4802f5c742cef454f16677b3bf727db962b8d0b12515b08cca74e2147775e5ae248;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a87f31f46b56414bafc8c93b0a7f761a764af0cc29b39274f7d710edb5ce305455e19b160e7113f2bf8657d6ee2f9ec8173158f136bbf4cd5801658822c382897701fec744d27b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h300777ec1dbebd4d66bb04848bb026b8adda505af6fafc2522544b42fe89cd9984d0a034d32d0bd300195a4a58774d024da7fb80eea5cdeeed3e4eaf9aae87d9c33f0ed6e0fe66ca;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3be5f98b5ca52ae469b430fd8334af02e00d4410fdaaeeaa089a5f8f4b4b302acdb3094c92c1550dd0ef17f46fe5c901008326d3336f17e15f8ac76a2d75bcf382fafe8ddd277516;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hade48d2949ec394a92a98f41960695afe8178e6b154720992435709767616152d7fd36a2eda718bd9ee161c8d40a08e5ee569956948b2140d92c48d51a7660a2d16a809d9990a6bb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc94acef9494d4828d172d942adc45bb65e7555f48e887f3c57f5814d592e4d846ac27ffc261539694dd4afe8c9a9de4c1d16412bae6432ffec0dd3bf9d931366eebf777fcfa351ef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefea2f2b77ba0d24e594f28a0736a00105df4a50f9065236b89fa4b5166379f99098386c24fa31978605d467706dc26d13545d70baa0ba99f10d6e849d2126bc37e27a6293b533a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h225b4d3701893cfb299d2ba96417a1f1a7db6bb80fe5715305ce0bcbb7ffd9958c0c16816bd2fcbbd8dfe94cf924058f1eb797e5d4d4d9e632fe0df996304d48d4157a0bcdbb8465;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73273638fbc0e077ac4bbf1d40c48bd84abc5b5bf5f27d9bebe53d42903681258fb9cef00708b3e046875608331dd7b98489fbc36f22975afedef95fc86bb45551b737a883008b7c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a3e964d9fbcb2a3909e64ad1bc181c1ba68842ed3643eb28e1ff25c8f5dd0e5bef8398c760bbc855cf22ea3f532b658ff4e2a43d287a10e018429e0f503fdf9b1de88fc3f9c8d07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1c4878f2035b08f5a0831638c7005f4db04a0d1162c6a68fd97d34ed8c890ab481ae5c906c01486388c836395cea4d310939ae8ddecd4f6c73dda216d75d4dd1aab0d70d0567e27;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he107db3048d78e83c3952a4c5cba8e301865f528564e4889da7f4d4ffd9e4d287205bf201e64913665dc95e028dc72b0fbdea79ce2fadba77d07fc7cef2f426d8232bfdf95004fab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5aa5ae0fb2450306ff55b9bf68243b04f69f59fa1f0a662d9fadb7e907a6ed9985f6f4ee950ce7329cac91e82bd4a668dd18508dd40850d4a8a0e47f4a4217747fb093133ecf391b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7d26f596519a40ae25620ef11bf60291271756fc6fbeb442e797207bdc46127f3e44f5b8f70066a77e8095682c2d9831e49263f0313734cf475b674a17e86c04abc4c6dc961a45e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbdf134582d77d1ecb0350e67b500024a802ab20e99fb38af34e4515d0b5986e8b5bdf8af23a976e27ad2043be33f747858cdd22a7bb04574c61b61fd3fa124b8cbe342712e3fe7ef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6093855767127e6d07a3bf8fa77baed9dae1cec95ebf3a4a82effa0c7f9a08c90c5adb7f2c86647f9c41a641d0e7e10e27f9709e4db87328f604b26f28b27580bc1dfe97a977fffd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1120348ba5447470b97214aabfcfcaf42729914bbc04293ef558e822fddd102a5560f5c7dd890ef872dfbe8c2805709c8b7701d2734c92598bfec16a1580ebeded3f480418f23513;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5a473cac5078a5c7eba2ee80891c7ad8d860e33dae77c2d05706981a12f85aa54735fa559bacde6ba36082c99236ec707fa5528252752a73d6fd0e31d77553dafd2cc800c711a26;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd816a663fcd07418cfda987b4ef3e6abefc9a08d6625514ede4d9c5e0e1bcfefae01b42a462cf1e0add67e06a6e89b20505685b542b4ec5b762b954886e7896b7bff90f4656774d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9a7239529559b078e27249bc79f5ba99b9d8e0662cf6b5a394e401515a26992c1e036a1863b736b8ea414643963825be00b954c03d99758c07aba688a64dca2f4f97de5dc96b7dc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h256b4dd224a1271e3884601076b363ff34ce9699095017fd39015b77698236e4cf99e900aaa0591dc4d3c247d4276ae5b3dced8f609dd564f8ce771e4d003d7aa602631eb7d27b43;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h525661c0af12ae0afafab1a02f4b9dd066365acbc3e1bf0c01eb1b296a817ac08ec832517317c59a6b5fc16b90ca937e4dbf89083632c9d90855724c9c520455fe87739f90bc1078;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3dd137c7e6251e0994e28bea185806ded8006415b61453581a915b0957b91dbe669217b9815cdc2177f0845387a446401b678ec3c0563814b64630ccbc59aeaf25a47379dbd1562d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f63ecbbf1acc38cc6e03abcb434bbc0c5b0a2feb456f1207a4a2ba28a5c0b091ce7b110d043df40b167f39b892c291ec26afce832d35b845ca9c2ae0cc6ca7e85daf54c824606e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7fca40e7c337c4d1b54403d93d922acf321e4f86246408af164b5abe0712e0f7c5282c852ac3aaa68fb1df17ef929d054f74df8d9d24b7a0cf70ec8c72b57fdf1ff0360124c6362;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f6090e5fad76cb64c18cce2fcdb42af4e56b9fdf56cdaa67af0ae227dd8a8cceb36988ea7e564d772782b155e7d1b87b2c00a3ca628c1e021dc55bb39166ea76b856972b0b8c6a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he99215780f2cb63c928d99b34bc5e4993441a4cb06430d939bc19d2a6177e27408220786155285620cd9267c0cc7ef71d52b2d0e79bfc6ef892ca02a86bc3d959da1dc0d42bb3e39;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h431725e8ab83594ed1989ef93ee2b136bc54371b339ca0e735359445682dd622b6248acc641a381d5e7d0b7a6a3b16124cbe1b363315872558eff8d9dd4bd21efd724e67e1589d29;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdffca493c981b5d2851b8d7bd4d2a87b2df04fde23a9c426199262bfc13d729264e4981d675e34157adc82c09bdcd6301ab058baf3fe299cf243afcd645dd0d9654f8429cc1efab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haad78ba2ac010be1d51d12a2635274a87cf7cbdd791ba48d3cc33ae19790c5fdc97b2d9600d710db17146ab2591f9062a3d0eed47c24580f5e3a4607b9eb2ac5eb4263fb020131f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b637f533722e9740509597aaf12b2678316d3c05b1994194cab5b8c6e6a31cbe5aa1e09b976b735bba6f86438463b75ba6349a7fb3a19506517471ddcefffde5bb17c0421413bc2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13fefd9d89bdbb7d558e10991ef4ac62c0b26342c6b60e94ea8dddf33a67a3e4ff70471c3e64af82fc4ab477ad3bb8a4e1f762f297b376dc6e3903181f4ae8797a8d23b8038a424b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e44bfff20657531df4f2ab1dbf2579c2f9d9c0f7ae3c4f903a2127e09723dc5f40480679d3ceaf177a719964bb9414eaab9aa72cfd6eb52e56e420b2f3bc0a87ad30f5722f84159;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd61d5b9a8f602485c2b62eb35b4556cd80030951173eb396500eb94f1fd959d5e77015167a6d1c3f63b718dc27e5ca86b1d1769f1c0a1ff8235589f7946a06e36c11029d5d34a198;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2f7dac34116b364d69b4938054d5f6a1bb9722fe357791539c6f2a1140f8a6cdeb72f1b416f1965aa17684b536733b987efb91acef01206d3bb51fddc011d7b64433fb1d3c412aa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7fd4744b24d1d7fccc604788c774012f05711d98d3bc3e6e058b736f7008145cd96077b6676d7c696c7add2ae876cf71a04fe6ca716e0d783ec2a1130436f9e81bec98c0541170be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha83ff329009b41fba44b60080ea539bda6e242c1dda031b366055d9e5e1436e4f929356e529ca4e50ac36a90342eaf64b0d17c0376cb123b76f39d08521ffc3728d65d436022c269;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcff4023d27fb8e96e4e0fee19afde8205c3d0ca18a34d2acc042f34883c9f1c352b024073b0fe51bc9c4d84870ffc6f1f3cfb1cf1ef22441685fcadbff1ecb9c31ede8c4b9321513;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4a3cf404a21db2f60abc01d7023e9d0be4bb11e9e7cb2ab0f3137132fa656b64728fddfd33d8746919a0a21b035ed5610c1d291d48e4951c7ca7d326c5e9da3a4b733ed4abf64ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habbe7e9b29eee0944d4d53ccd05e0a1eaad8a8bf13af0026f9cf2e3902c4c27d3706aae9535da991799a411bda4fcebde1add9568a2b322d06e9d6923af58b649642c46e090f42f1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55a2a0e216ee2deb1ad8e75a278707845d67c3761825c07527bad6fd887fa0ca98b378b9eeb22335add9289b3445a40755f01a5fba381211bbd0b70d6b6eff2dfbc6e54b8f4eb5a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4ac730cc316f9e43cec7c3cab56cab963520263bd1ecff17f4279739ffebb00fc62c3ab30fb50a3e7c40c6ccce39c33769310fdcc12cb5c2711ac8dc2526a59e451a572c6642bf4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he04bfff18164644f958a534ca05574817ad40adca9860ba48b3dc889f5d13286db9db48775e4b77fa1d69c862e8cea1a7ebf94d4516e1880a2f4a60410024a8edbc0f6d65811dc5b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha06cec6434ced0cb933392c0048071cf0226007c402669dcd2953dd53437d25bb116160660c208ff6ee56d32ebfd64cac69a7fb927535eb9ef816d726f4fa1f6fc281ea0e37bc3e2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83e42371782f8e38a051ec4efb7cb2fda21992d32439d5b59e34ff254e0603bc9d94c6bc493b4f631ccdbc44e019a1a786c24cbfdce071d7394bf857aa788d0bfaae0aa1ec0b233;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffedf9d798f8d89f720c4c2207d32f0fde264c72e5630c92ba37c3549540cb82e6e600b32bf31cee7f8786b2c10f7940dc848a65156d16974034e2126edcd24880cf8cda53ee9d83;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae349360c738d8f81886793eb3e1a4aa2dff4546942cdbf1077032852952358c02830d6dbea2f279efeab31a2ea7afd5f96b73cfd73c45d7481484ea34e84fc436fb557859a5aa40;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde04580ef6d80bb75f99e578ab5bfbaaa6a9bbd697fdac84a45ad66f900b82884de100021e6385c049907b63cb5d91f211ec934c45f5551db3bd7913e610841131cc2a06b8c044a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfac2f3814c2472d2e4b02b5b6fdc421aed2951d7423c1bd072969594de03983c671d5a38a22240417df5f81e133160d0a9ba7bf03d8121d6ae94324affc30a66fdcb215db0747c83;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h169a0e5b4a43576975c1fa80c7b29e66470a411918c97e37df06c10b3c6553d925845527a2b27964e8193b3733d6b0810b3151f01df1f92156a12d734d01d917d2583650bb728351;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11cb7205bfe8e1e461649975591187e25cb172e507a5c7b0292f83cf8407a5ea75d6123062cd5d559709b8cc44cc3b000742cd2cf0c7f50792d32234295fe852c40e499ad1078251;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b1e80d07d1ed0ee4beafe152741033dfa06949f7deb3a25790c0234bfdb2651c28756d575a3b713423499c4d0a37a8e207685974a2e8cd1b9ea93be04d77b2f0f1701819086d2f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he32fc794ce8f9e3aec7a2b7af9a5235cf37a5bd9c3d5d3d3ed8135a6b052f81c53d92bfb6e1264df452c0534fa881f657beb607e5014e8988811a817daa8adea543a2f4060c7fb2c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48a5729f1f1519004d12296ca094ffad22a4fe7213d4fcbf074e05d6f776112485b0951f1319c3f721a7f7bc716b3694e5f82e122f7bbce6bfb7e0371962db62bdf67b27b22bfabc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6a65291ed83cfb0f7383dd0145237163b9db4c8d523032bf5960244e47251e08c7b27c90207df9f2857586bc5f6e2f2941cd2316cf5cf2c582240f3d4fde2f4160f7124b2fd8389;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21abd4ed4a780bbb523e032e91cfc88c76cc2de24e364257e57293065f853adcbd623292b39bc23da781774ad2e72a921c3e60f6b16e955605ecd97b10b901f179d8ee0a45eb38b2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cbe0a09c665b41437d4b672b26a310f6c245b8f1cf357cf60ac69d8865e692f923fbb9835a3af1042894a231b34069f04a7c21e9651abed1ca3f48ab6ec846b2e3c7bc0abbce6ef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9180edfb3e80ae647b5631f44c1a45485770add6884ab5923d3e0b1a1b5850375b5053b3d62680fa2f60a400d3aa3573ed2187553fd240b5dae35c1db80576bee359dc5a0aab9ee1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h225b62ff92dd001f74a7bfaae5a6ad68c9ceb24cd13bcd84382fa7eb1744fbadce6d76b5bc0d08ca108516474288c40598bde7cb5fa0a9d0c170887b0ac977d1facf2548a91068d3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h679cfeb6813a45b3855111b109640c8a3b7fed2cd29e854545da1037fd1af712521d969cab04f9340144aaf0a8bc41ee696217f2a41cc761b506c3f3294029fd600c57c2bb16479a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc46b9607345e74e9b9e2fc1664bb0da04a44df41bd2ef202437b609d1b95d76d5da92591df1d9210aec7ba6ce5a5068c12ecd2e18aed5746fb4bb9644a29307c49ea4291afc64127;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5cf9cdc51cc17060b08b1d3b4aa90ea7cc99d29345a9eb5211487c390d0430b764191032227a4f383ee37e75aeea317183ed259523db39e7ad89d898cd9415a14ae0902a972fad6c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2fec57bc3d5bd444d034a93cbab8ef72c876fa6edc95d4c9db37b79c2b12fb53972c6b4028e20623e50e728b45f49e6f6986cc24358deb98e25da98fb8cec57213dc27498b3fce6c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b223dfdeea8f7c4202b0874bfda3d3c4d427a41c416fe1f367cba0fbe31a064e92ad8df4e11bc869634e71b4c112a7cdb136b589283c27d6cefec1308a6accd4afb90ea01de1c1d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b9823fb2867c332fcaa9f55c920d0e1b1eab2d6990b29e32712e2698344f13952f482fcdd45f6b75da8a9738bc436f52bc163de653afb0520ec4f64a6f80832e04af835d18e47ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h806e7af9fe34da848299c7f63cffc52eb3581d7ce057211414e77f9cab4e8dbcd014a7f2ad25e4f01cf2ca853582897d108f0b4d95ecf3cde04c3dbc37e76e5a54b847f847b91223;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde34727c6a803308eacc29dfccd8cc3450b73ab07160e9d19736dee2ccedeb4f507b4bed8d960c1cc34e26a4bbb0aa3a4b0dbe3c362676239480d072d5265f5f05dd6082e910663;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c57d9481087f77481dcb793d8e9919a46b9874cf29eac0b0469b7244bdfac7822ffa436bbda916a8d92dc353853bb4d6e816fc7b14ab5d8c5e805f7c0d647fe4967d87737a5a337;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h767ab25ecb6bd001f06e64bbacbb6a90e828e4b0e4734fb9d40755b5d937aa0a2a44772030ed498dcf88a7c37b9628be2adbe674b95d6d58b0a898f4e50d31d78b9ec526d43394ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdb81384bae0fa0513c226b5a1a2b251d2e7ab8c7d389ac3a7da23d84964353c95f90041c622d1718f1c95f181a14246bb8b7804a5a23f00855ba2eb8e519985d18b23f5131c0aa8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac0b87b76e16a724911a376cb46e15f91eb2572181b5b902d57a8441f51064980882d5e1eeb50c5d3a135ee82f5c0ae6516d595fbe8896548b5e1e2d6f9c002e200947e4881c7d3f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e492e158320ca5dc4e4e59d44ba581527411a2ff7dfc6adc04d215c6ae9594cc15187b88ddc3592dbc3963fb102f9ff2d4b674cd706b804a6b9d0f19e0c034e52b26444626ca949;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdeebf277a56fc95582ae92bad0c61e8133da0797e95c023dc9c9bd7cc1f1a22bad5a282a2f2e03fc66b59a0979c128896cde5ad7929232c7c4c39659562fe75ec7f5baedabee4385;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38da045ce77862cb190fd0bbba763a453f5ff304455c9a8a48df7fad28fe0181edcbfef3d500ace745ce71000a9b373364b2b81089e334c4661d691de5d575136922fbe6b3c7685;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79c695d769309bc242b6f3ad7bff5dc5ac5ec23790c7228ec5a010898a887d5fa1f9da6b601d57b027303e7c3c431c3dc0d27bf8c0a9ba431ff67e27c71e4e04522a24bb3f664f68;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd873f66b186f2da928b6d8c1cf7b4f8cef3fcebe3737bd04c75eb1a692b34d55e2def9791d2784f99b89520b6dd4b2685f1018b588e36a5b423892b00ad619c21bac8d4f08dde09b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca99e7d1e20d3692ee9e293abac28db39cd73469734ce4f703c25874de02414a7a0850d0c1cb5cae99d7431d6a27bcd53070b158051f09247c34275d6961abf5deba1ec5e49809ec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h544f9e4545992d9ea39d3d1e4e684b025838cd043808786efba66daeb65dc00c819cd154e39fc995f25d6743515a20f0dd463bbf2f6fd8ad771e2cd8da0885e898b1ca7e07ca22d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2fc31bbb0ea70877daa18df4e6de1f803cca5e8c124d94c6b5dfccca4f9937a44e56b857e2da51ee3dcd64061983c26034729ba30fd588af1846774c4ca0b65a59144e2625b51be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ee3d650f68c9025b3f0fd979767e26df5ad646c596b15b5f25cd97a15fc139ba3959b1ff173fa47f7df32fdb79f35ea2dcbfda193b443c61eb46f548df6d0fe5c77841fb37e2ab0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83e32e7fae52a41d4ed1b9e223f0b47072c846d82262a907b2848974dfd4811ef6412a460230f5b45f0c203c47bf2dbf41c15283982325a0245a8ef73a52bc085b012fdbcd295e74;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57d264468a101bc853f38e94ce2cbb957691eb4f032997dda79083f58e0d0aba4fb02018c321e588d08635f27438878d4c59658ae818d6ce73e6ec1a39176384c8e9151b53fc8bd5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa3bb577085cf89fe08a0830a6c0ab3747a8c0f886830ad58ae70f387df21822b701a9d357b61f61ac56cc6ade2574362d76a3754667f7efbebf440ddd55327d1b77ca4e92b2482e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9c2e5db86dd2862049afa32a9d50e2858302e3fa89a1876184bf737d2ef3f61cf0cf338194ac9a7c6ee0034fe4f613d15896aae09a5943282d479de0871492f3d69dd591f44863b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83012b0685b4c4fe7867a04bf27212fa8359455a45735cc3bd07fb5f342f4ee807cc12831677f9c471edaafefef52f40dc435f268dc969eb551185cb58c2f04351c3468077cc3728;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf078528b8b4dc6554dbc48a5180fb492a7cd00c72d41c11329c3dba363853b3d26f04c7b2dc2b5210bdc1e29ff3f6712962c451e026215da4d345f77321daddd46090215a977cab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ad7b6d03a69ec8830784534248e5dbb688e0755f4e12618c400112784db19a82452c190eea977c7818ac0f198680f836f613475a11917ab9ff651ac26bb0a07252981b6e5e0234b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfea5838866f6a4f9c3ca4dceca677aacf3bca1276f9a13e9e7b9a5283e26ea7bc39bc8031ef54dfafe5e4ae1d21ad167590762975732c48a0a7302eab4d9e47521333d63f19f6fdc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe17eb2cdc67a75aecec7f3b44f90f354a0ab6ee8ee5f479d3cc63c7a158303e233199402423e5bc0e11d7e61be5671c1368131dcc8b39ee5edfd534cf1a0fd6629d26040772d0d4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdeb7a49c809d2a5052ac9a67c4d4a446f520ff7e70daf0f68cd8cf0c40b1fbf0e35b9e538cbe038fe382f2e0e8d4a888b8c2903aee89e42991f0b2cfc1d2266ff090802decf8050f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc78453ef9f097fead83dfa4bdadee5c5567fd1f3e993105140791b4bba3680700a46f74c9f99e21cd90184d2804df2f2c56168f5543cfd6f2934f2a541a2cb7fd81d0f4ee8243ce9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc42142f81a8d4a70816bede587fb94089b943e3a51948b658833300525709ce6d709577aca268b9576dfb62ac77b4471ebe94bf0288f762cc2f689a5cfd500f1f30cca18b94f82f1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h258f28dbd275e5871ae97c7ba25565d1ce088505390b0722a46fa8459c8c092e800974104a518ccfce2b2e27e99c517796bee42f5ca984635568f2ea386015417b3e3e3a4b41357c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5bd2fb8d25d4712ebebab02891c3d1a7e560c8f862576bbb92826dc6a37c456ca3a66963cbd15f4a5e7d90ddeedff9d24271b6fa6d017a0a9c932ec91debb1fa52f4a139430786d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e8b427810752430f0b685280533ca4df2728f72e4c868757aa2e691f1bc953e455db76a6293d2cce11e2fca360ce447773ee2dcc344b2b8cb0063fdde0ded2fe80c55e936826960;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a92d75fae4ab963921e2b8a2bae1f9a01198d6faeee1aac2d85dc734e83dc7c39bde3bdfce4fbb9e4a9184a213a1ecb4759c547164ef25620d1fc2b5358e2a16b46d2a23dbe5541;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b5129d7d99d77bcc78c152a88c275a68212026b11ee564b9c4c56464921ddef8ba5b0172dd1536f10c609fbeb161be73a45e60271539057fb40291ee75feb7742d396555ec74e8b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc962ef925c7e8bd1517d7dcfdb4c0d9ca381bb7c7fe60c169426b0bff3ad7b93c9d6322dbb0192bd0b809181c9707e29b186b8c64062e0e6339c90ff3f6f392ed8cc961efe419be3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf958cabad99f85f7d1ab74daa4c2d77fcabb736de18b065b06da7888eefaf98ca12fdf139636ff41c80f291da608daa1f3c515a1772ee438bc2219a8b8dd4adc23ae7d210bbd72e0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc21b329f2493b99be600f39fd31083918a91ff0b2afb3d5d9cd9ca724fb3c7ca4a3eb68d3902b5439fce45d640e527b19e8deb51fb25bd384a055730e85b85056ef54449e569b452;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f7b57223043fb9b1c8523fff2f7e8b4b6b9fdb5d4c120f61fdae6210cada31439c9db4060fc6aaedc838d406082f301a1551795ea74c0a6eaf9de28f26e9e84914ca8a80ecbce33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f6dae74b916c5a84e62dacc3d9b61bccfd323d9d495af0ff90576f2875210c70718b178d791a675ad1b9b435d408195feb680afc173c78d4cca096d8da56901a5537eaa42caa8a7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62a812c2be60e639de564202a996ad310863186a87ad5a1710479f6e78f450b3f518a36b4962a1f1018e18ee5ffe57db0b7f3bb1a9c3d8fbb0c5108b2d35324eb12a88bd326f1c69;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h726db3c51324436608e67d400d582d375571ad09cb5a919f8b15757f22346b516107387553d193461656c872729578ad6bb5d4e86ad657413be50886a2101731d26b29b81eb8d9eb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e5ff33710daeb490c1c28a0b9d888709dc0db52b767043db3c6f7030c8ba486992b03457393c39b6a08491dd4f6124f48b43f6ada7300b3cfb8380406fbacb5b3a3ff0611f519c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1b97c943a83555fd021683bf7ea5c7bbd62000c3c958a0c542a75ae75d56549c6b2a94081fb1058a221c8ebd57670f79455dfbe18c3736f5685b1eead4dd17c1da6f2dc0b37f374;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d8c12068f0fcd3e712642cf1e706fa0e3884030dc0137c9b08961effe126aea0b16ea5312c87dee12c7c24b7a2776b995084cceded9c1d6fcde0aee8b31a6dbb4d47b9402e498fe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61453e4565d944cbef86deda3dec3393882c0147c29e900769c00ec004bb848164c21505ffb417a3fc2a5cd76e0f1ce451e82ccfdbe2798c8c34c1bf82429df06d5388512a5dc73a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heed5889940bfce2d53f4d4887813263e8021f5fe35404e9911f331ea0fc68d25002b603a0b860edf98b76101859566138a467532ef1dfb267799622435203a67787f6c62366a4255;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81681cc0a3dfec0d729c0d5663d9ddbf72811d3fba6cd81febd126a97e468287b935e3fe80a874992fd58400db2efd8daecdc688b635e742eaf0ee468a89d9fb7dd25508d9ca6c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h998b0f04b8799b1badb57dae68ee264605385151ac42375bb96b491c7a975734dbe4f4342f2ace714361d59c0f28d50959039ed1c3cd04e2461fa545ed757241bee6abee32786112;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h809c91b7d89cf36ec913e812454bd6542837ec0edbeb305ac3375eecf5b04f4250df447ff2b5628e1836565982c9335a5c075c11d2559b137c0b8a20e50bd3861d4d4545fcbda8e3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e4f6db5c55e8976f44734f09fde4c5894da53210fa59ed2d1ecfdfa50968b2ae44c16a68f7b19f509460bc7ab9d9a7d375a22d9622f3f44a06dd2ee14e3c35899ac6aab17c9dc33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ff5f57dbb06f09a13d27086feffa8952fb9eaa57139eda799ff5e7aa4d610f1890ef3ea8403fcadbf6ccd869eadfa99450ddfa76a6931920bf068bf60347699562864effd488670;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b633f89f8e9bfa7c854e7941ed1e80c37fb938bab2796bdb8af8323d5a20c80f8a1aa7215dcc19120a40bfca96949dfe679cb582d20b30fbf43e611b0a8a3dfb78320167c8af8db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfccafe86077ceaf22c6b68d35a8f87e29f4d90d025b33af0fe8479cef01da985aa3c2aff1ddd41479beadf7b2f16b8026c3e5a66ab7c5c8e5433a2d8b6414376a40b193f99d3f9da;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd1dfc573377ab934dd9d6676af2603d035308e64d4c3cc0592b082b8354e325ebfb9ccea3ee6db7099a8651eaba43ccc1306c3077e22e06cfaaef9dbcad05fea3eefb70b93fb2c7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0d8d9071ab6324c040777a7521fb6e0293ced1c8ecceb41e27fdf674b953f91322bf95a9960bb1aa7c1873391a4061cc9ff7ce979a6ae640cb121c3bddc5acf1c33de2eea7659fd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbffe78a2a13753a10c55daf5d6fced52aaa2611be28eca8038184103187dbde964742680a4ab5003855142a30a006761b12f6d093b5b01c95f8f14092340e6ed9774e3a5608b47dc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had14a14e16c94b24202f5adffa0f11b673465ebd4eece6d900f2cb7a33ddf96ad92d9188af34eff77e437574ea1fe5a3d8acff7087eaec796cf7af93f5d8b118b32f39a6353b8418;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81f96ba8b91a3a130fdf858820c4ad232485a6170e6a59e793aa9ead037ee04c7e40a1d277dfdbda3f94b26f716519e333b5040fcda00edde074f15222c96bb0469c94e8cb357416;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72e0ff4d55dbf555b88a259e554e28165e971116a9f54298ab8c344a0457e5ebbfb688ba61e0ea9041d7106e189d7971a07aac833badb930baa8bd40470019013aad836d20c1392c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cb29455566d0440644e29b86515bf7207c7e404239ed909b03b1e58e8d29eae3cf2b930177d7203de0cd3ff4c7e5cab46cd554fbee1ec0e63bc7ac87912b9ad9e02625d69d7607d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h217be29a82b70eeade599eda909ce409e81765c1fa842b98718acef0cb7bdb9b5f0d1f9d3fe9954ed5f7f55fbafbce66acbae2e9f548f38812544c84bd13dabb341fcec1855bd54e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddc5b7c849e04e20a37d508544ebc483b17cfa7e25a9a592bc59245cf0dfb58565f3091bdb88a09defa7a31a7b94c89c0d71ef096496a8a63b6504e3cb03670d153131855f925b2c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h573d554381bca49ca26e73d542f2745585869b7c49314edd5366678abd003e8f24dbfcc4c04f2e6f999b8c4e06ab9aa85ad091ae3db66fe64ab8c448477d4891fc4c5fea62c17fda;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h981f5b8e282e83c750e3072c3d58ca5092d555f3f15dbf2651425d19427b5c5a53cf45a8ab759e96f2c4d2e188cad9785d2e3ffcdc3e2e6348658562f7f2ab69cb9c53fd2b9dbb1e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc34df8347f7b4e71a7ddca9fe8121d3ca424bea04ad85d1cb54379946dd75a3d790b7ff8221337b2c7f8852a1a854c39853bf16207a283789f86bb244fde93df50c06dbb1510fc43;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h332ebb30856a29ff2b1e305a85fdee3be2210fc4daf26be2d857ad009c846fd41e74b64fa43a2eed9b039c23cf908b54be827062b87fd85d2436fab83f1feb7d2985dcd2f5936526;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e68c7aacb32be10eaa62e0feface369bbfbd3e64edb20e85cff5ef5e2a39ce68e6e116c5da5fd074d5877e64c344356fd44c665d019d25bd27f4023f017c86c47fbd47b23878e0b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf57dacd7728a419ba6a7dac5e89e6c15004dfe43c8b334b37a7f5a61d0e5c3730a9984f52970abb443196cdcae2db400816bd0786ed091aea5445533d7df43c82f707e08d9ea0e92;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35b215062005914294463075738daaee0742b7946a8ec95964d7f4f386350fbd776ec0fef5ec061c8b657b1d663741b1abab4cdb756c886d83328ac4cbcd7a7e6c469d218b9525;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5290c7bc931d66a0d8db8cc364786972364d2915e0fe46e624e942d460ed0bd74e9f885de607d48a01513401786f43a0f90d177f3dcc40045baacf3cb138bb846f58a7e3b010741;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97d2ce4895ebd361d7da81e9509a067e2793a266544fd839d0b5c2adcd6451886eb94b27dd758bb9453f1d59fd26b996ca57fc59f92838c593bcc7cd1d502c85eabef71fcf7d4417;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb75bf722cf1ca6af670629e4a309656bfaa23398cee4713ed0d568f1ff997e4dfa073c8d10165443a4a946648c88d5035d89151ccedc2895a598cd8bab990be327f7071ba36a0650;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha511b30768964ee57c3ff089f6ef570fb51615aab29b651b98c2edf5bcecf0c71de33532c278905483b1ca7b0b3891895ac1db4115fcf8c24efd3ffc07a9698ef23118dee5f25797;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbfc1cb6ab049cca3ddcc9903be187689ffac713c072834750a21c0510ff94b5c17e1d7ba1844039bcb481d4f751717c7cf15310e2c13d75dd5a07b98339a78a964485f582dcc27d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h329deb3d5b47c514cb44d521dc95a764762b7f05d83c9d8a6893dcec57e086e07552a6dddbd5e8018b6f574c86b5e83c917b52eabee64e35022f455c21b620a0eb1f5e53a25b327c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1b0d81484e230ac12895fa4b5a5f968ea2d88812de47ec2b016d0094392bca7e0f4f1cc394bd466df479d0edbfeae74a4d20630796d0c290be6d78bd51ea78f09989d3fc61acb86;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93390e145a706a873abfc1ccf0f47e7b2d3560fe5ca1c404185f3026e32e9fe78aef997675703cdd80b8e655dba87b6268c964a6f60321fd0eef94722fbd29e136502b9669c80dea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8fb2a22f60896c78269e86b36e0e00b91d163794942eb05670c48b42378130050b4ff4717e7c73b342ba83297e1a775af5de7173e687b80f425bcfdfc4a308e960778b9d1d585d95;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1daa37a44e6272007688fdddac8652fa79695705dcb0c0dcb798f9554930d80578f87bd213a1c79c76448547fe139bab3dbbd6c95e54a74419e0cc58979383014eb584aafab364ef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8de87900660246a640cfb835afe82a53b412e3484aba563aaaf8560848cba837cba8d414610255d84b22f043a69be75e88632b31e3935cf054c3984632079687dd11a837059eaad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c984065f963dea3992615c2f24318ef6bcdab8cf4575f2a737cd86e812c47074087e05f2f1b8353f084814a4b5e8d537e9340fac8a12c0b2956b49661750fccd4e0d3e5595377c3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb74d0d85208793beaeace52def56e7d3f52f149395c284a4bfcdcd4c21ced97bc222096150398e96663554824fda4d06a66395d5c64bab4472f96db53a6a4ab1d60f83d1a79da858;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56c4675e362e0a6adf664fa506fe4763c8501ba6dcf6b16960ad116dad9b88f6a18887b54f6d4036b94b6f04bfaba0d8f208ad1d608b3074dc844a39818a745cc03243d2e24217c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd4cfd79759b9f169a46d1d7aa00f42460214bb75c597557238b5628d9655503aebde8b57488fef7b9dbdb6433e64e20c600399cfb522b543728fca099594aba51dae4e820cbc53c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a60d2712049ff1a15055fa769e709cbc2c2b462e44619964de20f51854b1b01da2f9cae466e52a16ec844b8cc2d9a51f557bbf168e00cc515f835d16f0ea485b02f7fb30e604103;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb192f5925682baedf3de16e4da31564a4d00583d89ab8cd2d3c16b7ba56582178bae3709a609637da7bc936ea577698c00074fcba33bed653bc519ff66e76fee01c6fffe059867db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9dfe7ecc4e4a7727ee3f261f50e1f6a40502ccaf6825f9823412c2f8f3cab9d029c702fcb06262165cab254b4275d4dcdcea13cdf2e17addf746a58998744fa17f24184dcd7734f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e9a2ab8cdb4c4c816aacab133955dd1acd407eb8fcef1b892d8c43c540d73bfbb4e82ff0bbc9bb0985e0219f3c75ce1f46409bfece24354345a7b2259e64b5ff9fe17ddbbbef906;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6cdec9a0f5eadfb3076c3b15f2075828653e1038f2d952d8040b80631a9d36d525260bcf415ff6e3e36a5d8e6332ddba09f4fb9ab745d80de619b02bb7366c2415e15311a9d679ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5321a0ff4716f9b90e2f2f6895355aee4fa436422e2b6311bd3708ed3b896e7dcf3b5be360e744412555fc46f7510ffba933eba62c09ef602df44fff97b2914247ac0b5256271cff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b1282572df7902e019915e2a932672f513f0a27d69c6b999348b4f27fcb860a1dc90e1aa1528d0bc9afed6293a4abf5bedfe0fffa8d61881c18aac4741d095872c436cc7d0ceee1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0edc5944b43433057c2c25ebbec27228923f79a435f1a522a7c4583cd6970f4d062586d28ca1b209c5d59e4abe03c733c139e4d79fa1d94ae7a65a4400581106ba1aef8eac2847a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7598735386b76071bea7b6f6a9305413f8771d71e2655ceefdb9f2acdd3e6c0d5780d076a8459f7e774561ce0ce16feb5c769968e23dc11fa912220138c873c95aca89beae31e75;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78f09ef939b257ff065d6c347c4723358d1e57cfc62696533baeb746e85d2f22c1b20c363b13e6e58649f05ff71e4a68fd5529f2fbd1f80522d1f56b59bb9ead0f4a65396aec30cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4674cb306d95d05865856cfc389b77ae5851a50c20f9bbf7817531cb38cdd085a898d1d24d6c9ef72e5130a22e4870b657f24a5f6c741b28879c8cf7437f1741f19343a07845d583;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2aeebe229dc5681070de70ec50655bfb500b9d3b327b7c8f5105ce7692442f756452299eaeb305e9b958d965b9f3d4a558973c87c8f3f35804c98444b8f29700d2a8003c43574681;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc65e17c510461b1b242249fc9108711ba25c409ec55cd06b6647059b406ffdd81f8ab6a913fa75338acad9958003411e4a9721aef32ca53828ca62b0b510fb64616db7a9dad72a43;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a21bb0e3e7e73324d930340bb769e685f7f922e9ed9cb90f5246ec90288e041ccf2d5ede684c90bfcff957ceada26e3d956c5614086952be0ca1dad55d1a0c5bd049136caa32169;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9498daf6cea328b6f14475ffcb55e711ab1fc0dc993003caf2024ff9b4019fb23e1a77229e319cb60a0e41bff3ba33ae3fd2f65b56df74af44c4cecaf83d7cdb5dc599a15ab1cfbe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha520a4d896ce825991db6d252d5991cb44f9b823e622e801fc050e7106d8b80bf13d299009afca4841175d13d49a6b3eae9b8b760014c0d0ec48cc4f42cb6f9344571cc49cda9c0f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3735cf9557b8045cd7e25de2b551aa4f2a64ac8c7c8ab1aa845b7516dcc8e356c08445ce2c2ddfb4e2bf3af25d9409f773aed1ace7b8deb7b71b9870b7306e09ca00a34ca235b424;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59db479b87c09f32304b6b9f02cafc5416f08ce58a9538e000c73318e8a966de07e0622400e7f8a9b3ef37c7e9a5970412ba8f534229be79e8ef93cf9b3e8e74a4814bb1ca88973e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2db080f87fefae67538080cb656657504b9d7a1457a38016bb57799c52935198e24abedaf6db3d1e52f676148d889c736ef0c7a0b01e1e521d3f8f33f40cf1722e96db5e05ded4a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he63224b87e231131cc31150e8de6c62d355ce0b8e809c8deff94ed585d85214b0c84f663028f0d3580e1548bc83740de8a0a15561a3bcb15c7fdec88094b2e0682ece1603cfe321a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f72fb4564331924b71e2e7046883d59f0145f8d64e6cc93075f9b160059d87f8eac27c5b51a010b7e4fc96d15d5451756dc35914f718542a04570521e0082df788455c8f7a9494b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb7efa8dbde6ba61b042c92d00c9e82787e5c81ce398dda86a64fa810254eb0d120f753bdc37f124b30ee68ece82f973586aeb7f767375d13f876e9cf45e97121f7222554c15e179;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d99ac90040a368d28e575d4d300bc43e72ab68babf99371d5d4c4e16172d3cd1e706a248a7484632cd197c5a96d2d21b2ee6b342b5d39279c83446f0ef1c730d4a54759b21d5332;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf23839b598f70db8f3e82b967aa9ed671470691ab8ed704d256ad57245b9d803ac41e0d9c32de6d8ca1be405c604f6044a47e85bc4f816cbfd68eca14da0f3a8489c75c0f2623da6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f22a3c7a1d7171abce9fb900118f8b94619c83efc28995639ad938b71d496115dd4f9442b686455549ae4a4c7c8fade33295d64a22e3110165c9b2c3550a902e85c9dcd45f4c119;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha452fd2ce093c96909767838cde5abe728cb52716855270af629cd014b4490c08b4f5fd9eb804ba0f2ae53b31334b829db1e9a27923c8a1b806b4e382bf20947466d506253e1ac56;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h962b29141d4148b30ba88d854170feacb8abc80e23b5d3510c5756a073bf096cacd5a2db81f5dc8f36f436654bbdf0996dba277c1fba881a2323f5f362323b23555cddfe2a0f994;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heaa1ba8d9ac92bf21e95e77faa450bd256348233681b5c599d5c8fde221d52d226ff85fa26a4106f6c39b1d3d9c0b32d92ae663ca87c325df073dee66b79909a9dd3b30bddb48d3e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a0a4935295ac18f280475844021a967344f7ab513c0d5b687b9818987c26acaf5093b228319192bdfe62135cb20039158840e4048643483005a4b0ca81e8bebccf48427d7f7786b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h506eef34c2c737c5e442007038b1db4ede01174af3c60c2056a5ff4d3faf595e0be9591794899a67b18eb13320adf903e0e5c01a92be1d7ebd11edb3c3ed1af550ba34b5a42a364d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5100862396944b28777e49d357b2c84b08643dc692096f69842e2374de9f15515e45944600389a453d081b7631800a24de5feb10cafe1c7c755ee71c67708d37b14594d5d8075250;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h572e4928b2f37e522e7ea4fd64953f0b7f6f3516cbf892286ffbdc2a6c3835f8e127fdcd669a9b67f98b6ab3bc7aeb6ce3d27eb88d81f4db0526ba829f33efd74a34d16f9fb45409;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f50de3061da5d45e259f87a8fb3c3ed30f2983b49dc20b1d852887247b3e7001f6effbf6ecffea53d5b5d59cc8796312e269df16a899db62c47da331147e75cc094e7186f7085e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd76660b03d8a2dce59f75c51b21586a1b1f2f8c64c6453ba094407c63b43f1cf1dfdface5ac36ec75912bb77191f248147b1480b243bc63061d25494e2e52c16565a9af9beb8602b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2b9253bab97b9ee170db06543b9c6cc19ae29b6284f65460a1dbe8ade80477835e8c49a095880cf08adefe233ba0b47994628d49e8b0edec426af35100684009673c7f406ce424f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e54601f3a7e49343d0788ab6e84081bc5af8259ee9756a39c00d37a90429c642f3afb27ac95ead7d1f1f6657de1ae502d04dd331ac8a614378791efa3086f29321c784485777bb7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbfbe306a42e60143b09537258170d0128a35a8f8f0b320b0ce9125189c5a5b9a0d9a10b40bbb8ba9b4f06538652dddb19f8233ab05a7fe4e6f82519e76dd9cd9408ea25a8f58803;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb9b1923b6d51898bc0fc0c44bf88d302bebde95770b3b6c4d3c659d748012e4ac12071b4628ea8b9e86412eb2fb2018ddfbd11484e58431ab2953af0ac7cb82284d973421b44eb7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3745604479d3aedaabe0a9741b1b087a9e2b7e8ce6afe940ecbf53b6f80293dc81b9c99fe5885943fe2c7c1e695bc13fff54a4a7eee0adba414cf0117bbe102e55b554d4439b8e4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8a7283fac9caac871fc13905b9303ace9c835a2a4f7e0b21a03b3f3422383f43cd1132e8b9e68d1b4de00c1f09c0864d48fd01966a809dad1a9f2de0c12e52561c663f5968a2fc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62b4697d46279a15401269d49e851e1f30c907f621320733fde060053e980e320aa250059b40f8465f52cee619a96fdc822303db8595669fe61fa2dfb7dac5f6d3e4f2ed5777ca9d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7db4edecb6b1b634c15ccf8139a12aa40934209f42f8dc46ea6c7cba6afa10356a34b4d9503b32c570d65ba2a218f489f8cd07e3f47c9c3ed16e2f83c473ecbca83a9c467d43e23;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3dacce5cb36816649642ec411cb512f360bbbf5ed985f3e48ee137638b2877c98d0dfe795b7b84f010b4acad96fa5b322796e36c0c70c6e968ef322fb472fbff428c9d352bdf8a29;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb62967296f89e177f572d0385fc6ffa374c8257e7b8e98c92f4c27098b47f19db92f544427a707a844be158a826594c4f66fd8005c98aeafaa0c73e5f52e9c898adef286f206c3d0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd888d9e222e10488a156103d7f213ccbb0f0783304ceb42be3fcbf47370def8f38ab3fa97234ff9e0e475c83c4735acaaa0a81f1234d460fcff573fe8f66fce8eadfe86b0232c6b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67d50af39c69fa031ecb91f66e0cadcb9984a565b0c1f4014504d1a486c1b2b464b0c7060c86a3425ede0e52e1a947b65235cb76f639d7f59f2a540e9930aa05d139e9472fe9c061;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2030a58edea472c08d8970fb92c69ab2790f63868c7291bfd3e97f73054455642fcbb2559170a989fc0c667cc57fce6ac657cdc871cdab36c48b8bf690e82ce08c64fa617787f468;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b0d75a80d3fb49bbc95cc9ab9a1be279aeef05ef455156d9126378c0f54c644d54f38490b22658334ee2f83a79c15a51591f941a6e96f73b7312756dae7d235b51c8725ca2a69f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10f2981a285ebb02064aa790d95d93da7a74222f14d45b24fe1c79ca52d46b1f663f5a1f4b4a8249e4f752b3f5696db3dea70174e24553444dc618010fea26dffa19230997664a0c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2195e1db8815f7bf4ca657f48c57279daad08838c888a4fe192b68044a8aa30e6ee69ce9500b2552e24996063783cc7d607efda3eaaec0dd2d3af4dd12f4950cd02ad699e8ca8069;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2db11f10cd4d5d97f64ab0ea71d3c5a9499d90ef87e9ebf5b5f534634aaa048b12258c82ec639c7c217e8bd8a6c11df3c6b74a72a6c6d6e34cbdc4d8e836402fd3028eb06938c0c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4434d3f2f097ed5afdf02e54868edf2471f649cd591405b6571cc2c7790744333add19950111bb8547f627743bb53df3ca241bde7bf8902580487441357cd56b5bd77dd374a5673d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97fe8f02773481628f9fd566bcb8f7156af12769856d1eb871fb03fa86e92b2adedb72d2a89bfcf93e03210fe45784d3404a44a344cef50ea1251689b6ae648c3d9607abfcc303c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f0aac67be6d576b07b4e4d65c3b3d056e17ff4d2d2c89a5ce1803abc1bdc63699e7ccca933045169236d2abff711568e56c09865b3e692289998cfff089728fc2146219ff2c5b97;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ad66149af58a2e8334459b7c664b0dc44d33c9098cb84f2d35bbe162ab3ac57c17a7e732b20aa9f3061130584a4839331deca2cc63889b34b6675ba11ba81ef68eca9d8ee4a5ef8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf60c6b33dc5457cd7d3c8c7c7a45da14a441b6aefc303128a1e8475f9081b829caf66407443dd898ecedac02761f8292f3dd888f8f35b1ca17f9e563685bde1fdc78474a6c70fc46;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf0eaab57f0ab496f7e41a58afe1851c8537c4525143d79fd67da3937ca12dfd27802391cc762f06ffaaec2bc610ee2bb3d238f55bb085ed2907dd48675d7a93386d53422fab45d9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd638969bda13aa6a635795cacdcfba1558d112e2610424159eaec2b2ce54199e4ae2b1feb7310ed88606e3a3d0fb2e4c6704500e224cea781e2b29521e06ceb155526577e0d45869;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1178e519a54619bc40c0833a96521a941135e5e3990b7ffc0d6b0afe2dcdbf4ccd148b66c4e1eb593d78410fbb469407e973a8c18086320c5b4f11d3195a02bb2a1a8272010469e3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2a3444ae8efe7bfc3602b80364c7ac678588219565667b47590b0cfe07df9fb875087ad60ab431686b3f8c9fbbf7c399c1937604afa695d03fced701d95aae8ed69d8afc59e4b79;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35be9b780a75e9e5a2964db54b5711491eeba93b6ea69ac6dfa65667f297c4c6283a8de81130310d57346fdcc40c6e2849312c1c388b9748c66d5f62ce62a72aff7b8cbae9a817fc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf67548a1c55e33e17720f9d43b52dfa16bd4e80d6f9fc6fdba73623003213fc4aecf960dfe736ed8d9ac57842777bf9eeb50932933c6fef5f9062b194e4045c20f722048ce42f35c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10bb8205486475878967cee66c9ee153e8422fe94718a27a1854b83501ac5fc3aeea0bca1eebe225d80c98b69cc4d5033b8a40ec143b06e08c1ad611464c5ef76952d3bc02b620d5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h630e757c36f1db20861701cfa19581535878d5f32bdb0196dd12580dfca0dacf2ba6d5400b02b7c90e85dd8961ad31c1373012a80737e32ad4ab2ef52a477480ebe42db5755b958a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h569313e085c8544415d179dfd4737bb1f047ce8cc8059fb2b35cccb30b3ee7e1871f8517df295bf62624c36c578c0c07341909e9fafef15c821d7f73e0f7b6ebea7b06c67890cf2c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61688181a4636b36ff83238bc7e3fece3fa92a9c5cfa66027c97f52fa39d5dc2b11d25fcca1c78a58677008e37aaf46753ef8a868a2f1f3f5b248107ce3059fe98a03329335ac28b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b2c7c3ae02f6ac924e4beb0fb2c365598032deac061ec21a339cf32809b2647ef22bcf494bed66f7a156e399a719b092b0e5e4d510c5ccc1936b3e3766b2c1a1ad8ca509cdb976e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9b0310ad57d4a51cc1002ebdf03ef886f0135516000f14134a4e26cd9a108fca776e5bc36beca0dbdd59aadb092cf6be9caa3079740d6b1c3b93d4aa31e237755d2c518df00eeb2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h725af2ddbd3db2ff213f6a6cf77e280159d456cce1f1b3f96a85d67a02e47f8df467b4c92aacaf6fd5e66c1ee1ca8def34c4b57c618136d13b21d3f028f0b40e0b2637255c447e87;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hebc1455d50ee88f0a37b3d62c1ee5ef924baf7b4c481a593625173ab47b742ec69451253992a1a880eee4fd034e2e941d2757c7809e6f6355cd7107c9430902c41244acce47ccc9a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8add6ddc9dd4437a1278e6f78b0979e24570e13a4d119ce74e7fa98cf7bfbdcb93ceffcea5d73ac360bb88b080f1a16834707a3a09db5b04dc2611e54c087aab78ca012296156aa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbac5df0d9281f68ff4835bd0c260f3954de7d505b31883671e22276ebeea580699aac196c1c0b70652d37f581216240450e2270e424a292a6ddba589ac59484863f06ad6f2a094;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h284cd8154b40ead04432da48cf4232d35bbe1cb6570f3f3e857d380e2600d08e17494c5064f20e06f5d6714c33af57770705e553911cc970510a40ffde0990ec704b04d7afaec60d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8612b046e99f079c7c0360f5092ba7de0ec0f7ed280ebd4d1932fbcf34895cca64f9d1e13a7d592c63c07eb1d1098da9cac5524605516d93717a5b7ece9a7f27889e3c7b30cf8523;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45554a5325530f837a0ede19e4c0a272996f259aac30991c32300380c66c25a6bf00deac8bca0ab5d0b3ec8fadffb3e16851056ead4e2c51dcb2422384c15cb080bf0e94a3dc81ca;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfffcfaac24f38a5e4ee3608813a56c3eb1cbcd755bf95ae13b5c94bb3d16a8c1e691daa1c84fde939d957c4c6459449d99f847d8787fd9eeb020f0d4811d19d7a6f78309e15321c9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e99a48a23cdfbd80d28574b927da15f32df0ecf3759d282588f3141e2531e1cc4d9ba6d47003d9aa80f6ae61ac2379895e4abe5da07b19694228fff4442d99aa6db9d02b4791eea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f4168f5bb400f3a0ab3321d854453e02969349545dde009330b5ab814ba70e2c8cb0f7b89ea92b639268cd93d630b30eedf77c467c4d2a1a1ff104fafe2d6d173b55db96659c727;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h166a63769c957870d933eea72ac32e8e81bdacd2ac3502f42798535f4ed9846a75c8f65eb9249af0cef3286f125a94bead3e17bba3dedc777981c8154bf5f9537f4054bf8b22805b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2654a6d6a6eef8912a2b24d9d34c3b2f37f33ad8d9a533fd0d65ecb73e601ad1f1e8ee2a51517e961d6c880758ceead358102685b46d2078757495cf5c89c1a80178ab6eb17e572b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3acb95721021259e409bfa6883b98e1dc88fafce9da058cec44a58b35a819bd91fc2ee437da634e55a2e1a1dfc57796b8fb50f919e2751cde2e04be699fb6446ca9ddd1a9b7b61b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a509082a286fbfb9129e0d06e05b40af27bba5e6a0168e743302f7f1be2714de649b12b94420f4c85e4ca02cf64df706f5711235130719fae7ca0d805c8a2c8401b33a162dfa92d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79ff771d3ddd38fd8daaa487c8276ba31b46456158e0da0f5732fa4185a24e7765c85c5c0ea6184bb0780771e2174ffa7c2ce5ca1a542fa229a63c5ec43e60fe2f43da58e049f519;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a89dda330e706d01d09a6cc2de9b448b90dbc43ccaacd1748a1da0924b05be718473f447ec288817520d8e846fd02e5e6953f58a103892874010a7f57cb3a00b53f3ba38debb064;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf7bc586dedfe5f0423e7bc729a09301a6efee7012c7c5515a4c52c6613df93c0785b73b62d0c91a07844fb1ce9c0623bd3ae2705de8bcb06f37c18831e159e0d54e95296457f454;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e990597181c5f3725d85f4fc37b7abcfb9e6885f5f5313d21b6d82345f865e5919046be19010e3c588e2cd63122b19fc9ee3c95760178e3acf6b2354fd751c8a98f0e829f1a637e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83272775580708931ea1d54e5aec4f78ed1f096182e8ab1703d0901123d55614b6ea4d41c035377810446e83e48cecdff884c1282b842d63699c39300fb6d8828967e5f5ea4436e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha53e80274fde10c3d592e94db8ae2e222e4ccb00d8f1007c66aa121ecb3ee294c60d86f522ec807c957f6af3536eda9be9537a8e8856bba0f556fc7a44f5926a6b8ca400778456da;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29d27ddfa882bc0104315df377760c91e7efdd9bf5dc02c7fddd12ab00438fdce1eb660927771184c89904656b94c9c4e4465f66c30e58569baed0c9d7decb0e366f5fea59a2dcbb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55e15e6164cf93e7718fe70a027db35e11ddbe03c0dcf2f82f23fe6d22cb34c1c5a563617c92ee2870858fc24f8990d42ce41be56c1eeeab78f94e94e183d83208488eb720636060;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc4722c25a94c25de030d5c688e99f87d5b1ee54dcb9fd525bfd91bcf66232db696047783835030c0a1c3784c023649a3375ebf1d5a490fc808d6a3948d34f992569f105d5327ffb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d52a95c57c292d1ef89baf1d87bbadcb73cc63adcdfa86def5497be850740ad2031c8a11842e6991a8606e0d881b702cfb6b7397bba6e17bd7888f2b4c70d01f06e08fe91a23ae3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd6be86feae68da0763cc90cde7096d468ce9df90932a59c59d78cfff8705ffe00f565d74e722fb6b26728d2e7d4679d6849e76ed521edcbea01867ed2bcb4302e4491ba87d1685e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38c440656451d16f956e4bf37fda4cbce7c36889948a71770e063b794ebbad6a2698e3a62212e6f86271424900caae3736862bee0ef48b6171fe7d199ad6153c217454e47811fc9a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1cccaf6a8f6bf3a3f376d0de24461ee20804c28f26d0daf639e8b7c83f935695b65b113bc97fc54956b5788c06bb854d63258a79bb01834e35fc2e5f6b80ea8521cd95a652de636;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha332ba72a1024d40d72b3ff9557d31af51265bdc5aa938ce0c7a6a8b67f331086b8d127bc8105da7b75b7be96a34556a4c74efeef4208a8ca2359fb640ffc91c7ef35a117992cd03;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5845e1306d04a1f302d0310592d20d9041157723bcd6fe8303ae64beaae53efa03f348cdcf38219b5ce13ef154f3106908819099a6e00679a14daf9b81205760befd253bb5e7f9b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9173459a097f01a06efb0cf7174b7da9e4014ceed096673dc1c079a8dd0c1c34e990bb9d567ec00b356c2bef4e67af192b1a009ecb2606fe279cf48eb3784d688b36b8cf5d044f1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2037ac0f6e1c480d00a26c7d4a8f7b30b40a9e8556e05afdbbbae58c7e7f0ee4b082ab18921121f4290d900bdee58bf9e024d375ea4b9d178c3b0aa2373abff8763d0ed26d4b4dc4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3bc81c0bd7a465e10de86028614a0038529896582a3b31434121d043d35617e31334ce5139518e897a4d3be8fb99600d798ccaa158d572c8c04e83db07bf75e6fba19dd0f33c4d4a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h972f4e961337cec75b48f999652513511487ea4e2ee4c41c01ae2724506a0b52d643ed14e0d87adc1811dbfb702aab32972c97a58fb54b65dfed0a983d19841a1357bb4a2d4bda60;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h918db052bc387a0030307c0f033d28c1e6f23467742e984c1bf93d39a7b9959cc100ed8e22d6b63b7421f2f6e17bb59a37420ca8660bf002f23919659c04044e5cd9a7d6df1c9a24;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae2baccddcfd258a089e10972968d980f8e6432f306d9abf998decd2a51bbecde6b6e8ecf0221edee9198ca41321e930ae273ecde5d4eb8faf491d66899287d3ad75a4055424c0cb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7785211eee082118230718a852a5b258e09a973a676c2e4eaa1ed92645ddb82786282f64df098337e3e04b6189fec9756ec46983253d22b966deafe9ad5e7bbed323cb5167d03868;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd404089b5f99d24af43f5f132730a6871549423c8fc98adc431c5a0adc51d4b71040dad546bd401ea31e13a6e4f800fa6898addb52a26527a699a8728a6e1942c566e773c3c0b7f4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2be63c970034fca6f37429cf5ad9288bd155aa21cbfb29d74044cf388c4dbdb9ad850f0cf3fc147c18dd4b5e6aecc8bc9e43c119c8a6069f7e8c4ff51682f6ac94463c7172f2c361;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he04ba74e2c6e5f17f4eaa46af8efd2f9fb3db20d9d40f7f350a2b10c6521ebea0ad52e981ad92c93b57e57395241811ec6384cc36cdfbfcc0e56d9f8e51d3310290a22a0c402b757;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc68bf2bb3e0115d33baabd25a7aa3f8b9b82b5c77a5bf715b411a43a1523feb00cb50884b3e9d32047382591eca076dab93eedcfe0b5d18f52c004d1005db69a2c44053050bb9ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9dbc189b00932e1e3d223e85db9b98ab72ca0ff5cfb562e2a2401367df553f67ba2cfb08cfc728ef3eeee6d3d99765a6c6b6defa2bc5ef2f1d2f1e589f5dca75fac69d8d9aee24c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haddaaf05d070bb6494f79df821fb81f03a19d8679640477ac1dbfa8a6eef55b1d45016d8aeb9f6daea4dde57f57bc2017f5f42cec4f28ae394927c5aca5c7d34e5663b1ba5ab9f94;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h853a7274254ae4e334d89481431cce5106fb03321a4ca156cbe103060890a20ccbf36a6690f7147fd0c9d0f0177469db6d6898f8b01edf0ff94ba727e4cb75f4e21ece55b4930731;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1748bccf3d2f7928e0ae5f4a64c3f2073b5c487e2f43333fd1f69b3957810d5a0ea0da1a0adce2f62c6d465212f6fea673ba41bd6c3fe0dd09fdae31a22ec1666a16631d550477ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c6aff392e60b753e09854d1f0fa3a180b512ba5345177ca272d7e53f5ffeb8f1f3a90529eb1b5115ec4b8e6ecc15083619c539e4d603c47c3c9fb9d712a806a80fdb35c7abd2231;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a4a23d16e0ab9a166367b41d08540623b1e0fa8adc71aab367f18c2e437039b836b67b0b292194759ac232107669fd6727d2751299e9e2918229784ecf933887fe8c1abd93c0bb4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee807c20f5a0d3b3647721805f15070801fab1934cf7bf4a2f12c92d5edd770adac84a00610494d4ceef6dbdabc79fb9463126c7ebf6c7213640630813b476bbd67e6a0e835b9408;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he547ddc908391896a1f7805b937439b9a8c6b44ee65dbd75504bb5924ae32417d129f7cf2f859416fc463d47d806d900b3a697d4444d2dac37fb40f69b19b4016f0b4b3b56b086ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cc71ccb8a55b8ea2eacf11c58d141ec8a49cc659266b1b050b4b210a12500d44e01f402d79a20fce9fbb55ec70728dba577723a3f193f35a80d10cf47fc45a1d7b45d2d92b345e6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a61df18bb421f602d5685b289d8bbf53a7e2f7f246ebf89f53e4ad809f354d92b6b9ba3538e7709a118423f2e6046aff1b9140453d1ca9c5f557eabedd0318e157d1c4fa946d013;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bae5a4544e8ac31ad59c832f75cb615cfc67c74c7a0505b051a64cd5fa82708e0cbf48e35c38fc07a51138119e24717e3b226b0a8558d138e0d474589bd8c6de16685e1ec35f71d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb4e7cd36fff708ee7cb748b555825ed66ade2acb0dbb148046191ded78d50055cc954066f2521345a8e98f4f010f3a7c8955dce0adba842bf8699e202bd79f92644f3db31344458;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a06fa48dcd80a169426cbc5fa34e5f55dfe90b5c0f7500d238694ab806192302927ca07354e7b0eed75bf38780118ceb8e8ab245d46c5775c210f04fd8ad92d080edf22a5376240;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57979c14305a6d919e0e060229d88fc97eebe05df3b890e11700d8676f7b5391e60bcfcc7e7fc9dc09788a1206732839876a046c28aae09cd52b4972b041320b1feb20d7ea70897b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42becce0cf850e89c6d533b3dba9fa8384c447db295cbe8da6836fdd419187383c41111103f95b32daf4d07c391fa6e2b959a701d33d0041f6d18aecc12544658d7b62183becc1e2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd41d5e84a2f3ed2e8f3892b8513c98bdfb4dcbe85bd842cf8f508f4589a337ed0cb4c0ff7c83da69f136b3cacef4992dd2f31535b74e557c4a7276f8ecc000d0af0b9a45a7d89c61;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2355d7cf7fa41a030157f7d55224f2c094e227ce4f23f9b067a392ffabd5d072a34e3adcd53261ffda0b6f9c822c5ebf04f8c7564f4f6dfcfd0cef1c5d86ab2310333c2dcffa1b3f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5cc9ccfcb7cf8a2ef52bcf2c7396b5ade661a09021bff476e5746f97c4c450605a79dca08bb82d5700a626b30cb29c0e623a38f7d3b02ac630302d8cac599f31e2fbf95ceb1c88aa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd4d628d9da766be590d57d063283f56076b82a3620fa7611b8d00a240e9eb6e46bfccfa5a483c8ee5df50efb4c5ab611e3d3b05f67db3af96fe0bcce9596bee818d6cbde3199b803;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1572ffa1252e71bbbe2b86465a936a46db69e19ef65dbd6d845d3509ea5b377d5d4434093925b471e0f53e66dc26a395dcbfc3544329a417a1ff8b174a2ee07279e39a80b54bdaf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8641e5b1e83e0a2748324186a7104434f70af1f441aa3e519129ed3d16479dce38bcb07852eb0bd235c1d339fbef6dd20370264f06a2348d8f56d668c55aa92f0643b7f5dee58aa9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h186c36703d0eead5f6a7d2b3ea5234260fd01c9cc2fae32453f418d4f6342a8efb046993bee95cfa03c8bbd3695f7c4769d4a814e018110cad8f0582b45820e8d04088d943f57df5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81e39e1eac6efe7f082732d0a4f7eea48389f716d27226b2c564eaa46d9ce09bdce568c1d67fc2117e73554568df47f6b98dcd6c2bdacc50228ca43cd3328ebe15799fe9d3367d9f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7450411d747dc5ea93177a8c31987ea07dac2977d248418b5921333db1f089c5115f856eb60f9195e76ee6e2bde4ebdc10178cbf89f2c4d046ddeb5f0c8e347da6cfb84c6daece0c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5469add361193770b84d6537dda9329ad6dc70c45affaba290b1bc98f0c4a7113e9565146b9e594569e0f3e3ac8bf4c57dc0d7e4a4eaa4e65cc94f980caca562b1ab34068bafc5b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2fe6125960a601c0a5d7e369ae3be25af6cdfdfd87f1cfc87c198a3c3024692f0b77e926cbbdec97bf574d93975a52c098c9ecb09cf8349a2c822a56734676c1387ba2a4cfd5d02;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ea6bb48d5689e8e04782cb8e80996da1c925cc1532cf8017c44775e865423aae41d0d4cac49850a7ba92b520c722e5169e03fae5d0b3922cf4287e477234a8005fdf7d18a56f9c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82454616f15ba306d48ae344504916c729db4f6aba6ac8b1e8252be49ac7fe1c0996eb015bbc7ff9946a162d5e6c88830e68e63ae3d04c1eb7fbb9a10b24a53ba2a2ae9fabf1d40f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab28cf40f5dbd52f5422c9dde81c04f1cf7b6150de1187d1b1b95c4cafe97476a03a1bea3dbf880afea1d1b6511e00fc6a651e1ced69f44dfb350b2b51264aa0b6c01f232293accc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9570c8cec0658047f73931110c633c264d063413565056ff7a846eb0eaaebd0d8988772bda595848d69f61d6592ff051fbbea7d67fb921fe2f038f5b46527b4db111685dfde1c560;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3c0f50a199ef3a6cd714d479219ca76de1ff2bc899a50ba5e99aa263603260b0b6e80d6af23f328e51fa8de3f0786ff72e315ff4ea70ea06250bdeddb87ce8b7a2c50926a92b716;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h347e79e062ef93c1684c8082fb450e2a4dc9ab112f5ba164b40905478e3901019221bcd9bc6c37d254b25aa56310a9229953172774c9a5df712559f1e23fb5884ba274c0b5fc09f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5869c9ad979db89894215c243f2266fadb58eeaa405f263f1c41898a46b0a984d62e4cbc0358fc76a54335b48932e28293d0a443b92ca9d833d1c42a078c826b46845c1b451a464d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa5566267109dbfbe719b7e9828e421ad5a4ec76335ac80981f8ec66a439d3fd713437bb69f46f777f34497a5ec4e93dd686e735d73e156df13225e170bc33889cbe2a678730a4bc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ad82c49b71d41556b9fd1311e25577c8d82a8b524765500ad1e6645bd14e98226d00afed43fff37d8c9ff7e68ab602dfb6aa0c32639f7c6d09c9eaed0137b4f21c857259f9be955;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a0ca8770de290a6157606186dbbc0da6453b58665f2b2d688af4ff20ab819d6cdd32a3a851c9414f0cebc63d532e4e046b3d11224636e4d333263d818079b5a0f5ae447278a50e7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71665fcd6b5387a174c2fd0c8df231f654bfb9426e4e229610716c54f5b0ea36a26246e14ad1bd01f5d098e4a2043beb475644b1b2648f03d31d44f471505c398eab0b98bd4f54fc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d40878cb8578bb1228e55a76d0cce1d1a69318bd2092c4ea567d15432e519768fcb9efa0aa198e73a39ff206dc5c10dfd8ce02555b21da9227e4e7ebd2ec06a2a73b11acef75c36;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he12697c1467ab6a7318f32ee9f708fdd5b4a5f59304d96414fc076bc210d84f3c1bb69ec236551c37d5f08859c08af5aa34095105039d6e7f104d31b8ca0c22536c08bb31047c50e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2db06a515fa162d974833969b74d81e95425752bea7b9d16f56c6d5b4e7b35f7cc389bfcc238a6ab7fe73effb2e7a8087ae011d42b495f9b5d75097935213ab1109ef9f03280594;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b2cfcd87afe9e812e599fd9af77624ae085a89c2589d7eefc4e9aab40c4380deefe9535aef82668e2350c2848a35695e9218e5ae9f84c543b5a55004be8ff5ba948a5dea4242d9d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd9b03caaa2ac4593aa8a85d47201cd9d896db54deca0082a04f68cb68b0a9d2426474a9beb0ef689914ec0a897246550441dde1f332b09c315b7e3117e8441bad7f552e75c4db34;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0ef50cbb8aaaf34392bb3cfcde9a6f840617efd853743a41b16bbcedc75b662390b95d694753dea383934bb63d28130a3a89c01df2badb0478136d2e9e6a8f0fb5627da82209923;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h198cf18606fa94287ac707ee3a6a63c8efe9390d8825668a1d088c17fa22691d0639ebcb962c390106a5e5a2a130d27c0c039cbfe7f2cff2437b6c0525ea6f3715abaec63613f414;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha085bf41c6bb6d8d5ef949c39509dde3dfd026ebaaad4fd46530214a53b122380bb84ad12f102f07d6fb8d0073ef2b211a0ea2a12b2216571f2f327aed6e4475862f60a8a5c61ae5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd92c49808cbd4467909b492b3f5b349cb6f5e14132ffaeb801221326434b3bcde3f61903b4faa2e16d8789c82d8e9cd5ce7a92952ffb3ad6aee00dbdae769f8d75cae86d79e4afbe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bae93c0d3c859e46334f2921ed532585b3f2f0091964342a7be11f44b2fed3006b3170dad6185f4caa73b5aaab66f326715e8358e5f6cda590cb4d189bc5910ddde5643bc4593ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6def56711b5e56ac10c89d6006794cdbca093099a515290041768431a0b70977d955d6a635ba9510bf9e84fc7a146e06d57d70e4198a0a01bded55727736a953922fd9ddfa0ab9a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb3d8150d065fc11e4ab7b63313791291cd855806d365f08d15e183a15147336bb09f4a980fc628c822386bfa14d12aaf4d4c4b7f9bb5ef51f20113e077a7abad3db86553f97f82e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86ed98d5e68c17a57a30b97f8139381a1c240277fe53ef4f91b477b3aa0681a8b186d93dba04cd3cb52587d3a14a069549d7bc7b27208fe9e0a4f2821a2ee2b759ee4d7dfca6aa48;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0430f84aa10a65577336582c049d841b9148a0f133c08ac6920da041e45afc6005e6418fd5c6538a302ff06ef70a5b6673e4d9d98f0a696f26a6dc42ade8f3f491404aaa85d14db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8bf69ac30266fcbfa301513001bc641813c01395599c175b420d61404dd354da6d6e35232838145ad50c255177e3beed75932c982ee3c8d345f0ff3690899a66224c03ff54d224f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7f66a52d91c2a78c5d8c9a17b777a48dbb9483212c7209ff0a6149946b1fe987bc632abf6534d6b62e204dc4c4df9cc54233bbea9f6d249de39e953a3008d07c23424603f1ff9e5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77f6b7af7baa67cb01e9be448657e2f5497257a6d9e9a6a87c158f2b45593000676efd62f07602e9eb7811e8ec4de2ab2aa3fe47924b5d7cdbd58f30d073d2d626a203332f9eccdc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haaa7b52947370f01b87c1468b37e431a8a2f7e15a8ad49e63718754a50b56e3641ea542584a57cfeb2266b10768988158a62d26a85b815fab7d49d1c19ee9de5ee8b7965ae8845e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd66c44955428d44308083f9946c41e97199e9cadd4f96e1a6ef65703f5df06b8e94193c147641cb80040d4e9b38a6e5569919e5242555428ea20e4a7e97260fbfe058992a2bac1c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda96dd64bf5777b5833089760fcbc77a2dfc1c1d4070dc9ad10a7aa440857fab27aaa0d8875bbd60534171e3d24ff25e7a712fd5f62fa600473e71d62800f4f5dbb646acc161304c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd87ef769d92b76b5f707d3f810c60fc893dccb8a6344f21d796345e3ca109ee785f7e1d763606e0b14fa52b7865463c6ae04906925e9e28bb539a787cc23da6c6f0db8045f4fe23b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9bcc3d2b865965e3d90c9474dad6003d013931eae20143534d467db476029f7171ba5d68bbedab95142a4bb0f0ad9d30635f5ac2d07e8b12d65288f3bedc19c1e194df171fd017ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd45c9e2dbfcd69df7859e41c3f8d829a0dcf312b165636e10326ae11d2db9d8b1f7d4cff8783bdef9cd035cf01949c27d1b82fa87dbdeb2840a9539ec00ec6a48826aa0989512;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bd0cde09ea64336288caf775a48cbead02262e3c976934075e7259baa62db875fa378ca5fc48ec9870c8512f9bcb5e42740fa3eb38aed5e5be1f921297c0fd14074d929c896fe9f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78093edb43e9e93c49ac1e668e11d6095fcef0c75f398471508d1dea0977b316a7b324c102de4b29244432e8336e3e06fe99f05f12796affb1ad16f6d77946a5c3a87c97271468f8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8660e05f3f4d81a0a15caa260d4112fed99a5ed382a1ef744e96aa09c42d7c27584c759c703a3573429d3a7156245b9c6fffc32b49ffdecdaa6cae010d78ac532e94ccff0ca871a7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94b568a445c4d4df6030f3d6e3ff3de4830f5cc6a3df0c373058300e8113d59eee09d213841475a23d52ff5e39e126dee79e60519d4bb44b4187a930cabb261b31700c0e3c8dfe48;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89231220bfdf37e3a9c949bbdda8855a515f0035dd3166b605641878f1cd003d39f75926d975c954625922757d33d153d6162837c90fd8e07f5035819d5656d4d5af05552160f875;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9dc31a23dc069f5d8448735baeb38c588dd11e3ee4ee1b693ee12e99854726c2fdbc3101a6c54a6fa4f8ee6d9765dae8b30b9cf3303bb7ddd6b87e412447769c93060020a305be31;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8aa13ac00e511a3ad8e1a0a875d207791405a113160e9524ad9f7820fd81ec1bb88eed9a69705aef82a08317b54cdcfd165f3c761f15075f7fb37d0474e9936d20924be8bf31fac4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba7629782847c56440555fa2c407980721f8333615a41bb96480252aa0a9df75069a533691ef92ed9384902fe6bb1e7eb741385d7b467a2041191002711390cbe5021ed4948a8b45;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3368f5fa7c6dae769508acaf9aa81eda205c5810dbc50a94de3a2acddc9ae2739978350f3ae491dfce59db7c6ae3200c0598e4262fec241c430c846a53d3c5fb59f85ac42fcddc97;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85c6dee72f658b29d6ff7a750323c3168a5dfd9195854fb8e48a5577e9c8b14786f592f85dc4af44e192836728a20143e01fc0ebe0b2b50e6ff411daa311867ffe91074ac5b52a2a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d2a978fdc911e46d6ee4585745b9dab3504ab04edfa5f1e1afe68d0d8e243936c030111e4cb9c34b054b8abdf98c6655fa62a93445f144bd7dee019ee028efe0ba8b8de3d548cb3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cf36eeff6a78aeec84e57da2c01a770f00bd459bde28b5a6d04a44e49d102dc4e5a4923b90e532b2e767d803bcd406ad9a1e5b1012f7bfea5dad5c14905f023dfcb5f5210bfe91e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he890a7c685247be410f8fad444a36a766f8d0aeb9931148529b8a08c12e7647af6736ae6731936245b1869ad13006dd75c1dc598682ba6a8d500ff0aab7d18a7f476cd9ecb52e022;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5c5bf9ca5db08f2fc1307451465241af7f79656f23f82c4a10bbcfe8d723265ffcd38bab01137f5140e6b0ff969c2efc12e07d82886a53e67217dd8fc6b4ac321dc31ce66b29c2d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd69a25f590ff639942cdd144b80df75534b1f686272e07ba4138412efc854c014527f6230d3e6c87acea3fbbbf4258988cb4d8b54340e8515901dc20988651650e2a42edc866997;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb8dcbfc5dff93c2abbabc339e73070abe50291791801dad5807e680f5e8f8bb249436b5b4dafcd9080792a7306a896f0c8315b1eb26ab240aecc66d0a5f9f5410f6f18264d0d9a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8e52637c70bb6c86ffc21513367ede58a61f8587a803bf0c634a150238e270e837f1259d7f16928ce47db8d841b04cdce2d2db1df9aec9888723695709868b6539bd3d752613ebb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc827bdf5772932d82429cf305dc3be68dc4032b3e8d99e040cc0b4728353279ae09bebe22c7b65ee21f790d9f009d5f4e8bf7cfca84171e377b572c1abac4bab85312989ce19ff9d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h686e13c5ad2f9e14b9144dfa83a0ecf44f484c14764e94af9a5e5e0f1e0a60f04d66097f402aeb3ce1b0f01d0238b6066053a02243695902373cf88d1a263c5448b482d4f899de24;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e833e5a96efcd042541c46d480dd0760de9ccdb5a5f2bd8c8180a8281e87b46838391314546a6ef99032b496a24efa51597097456dc21e57ad287614d129cf6be4f8ecdb1486f2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h523d72333924051fbca1a1c9272a6d1fe5572edeeef3bf3fc5e9bdae493ab5958997e2a0f061d8d942fd41464a7afbf18dfe637fc5b235c8887845f6d8aea8c76abf06a45913fff1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c1059f09eb59ed27368ae55d2b870529cf77114b973e20b6028af94abc61aaa376312945813dacf9eb9a2ea66cf55a5844483894615e244e696974823e7e4043b3a3b13a2cefba3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d67bca05823a439072872fffa7135272698db57dacae7256cde3f0a431766557e8aaf0d512884ac55d353ac5195a75da496692fc9560ffcf0544aa7a166544aa3b81d25ee8a515f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d1d16fb3b949b490653fd3d591b305d8dc8c3831e57b85251c1c5eddb65c8d7e7093f46c818b65b4aba4b68de443cbaa3e80a99a48e106f087fc74d98e28791e5e0dbcf67d75d12;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2891730de10e5bdc56b8f1ab6816927d5f6db7f06b9cb9f370ebf9dfbc5186419de61260e0812fb925f8953982ca79c222af776fdfebd70d5740847c18bf46f245b36a190a74ee9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he29f08924b855a771bf20d096bbd57ac2eb9e406e128aa46275f82866906f82faeff5ebad9ad4bf329f038407e1bc550b81301c7275c4a7683322376192f286c54942c61c7ee2639;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc9cea7c5125359c6a69837b3f68412b06b14d848628f746ab0d9712f8a613a9d7f21576b20d37918c1569aa881d65d1760774645954e4eef127f020df4a005fc3d368701e7ebfbe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8240cff49b6ffd80f6152e7ed98876e84bee13e2f0314ccc7cd79220125fd0bc8e025d2c01171b2e3bf000b570793dae7e4ade3f3358896d02b7033d3388cae63dfb4dfc904ac801;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h614d944cc2161b4d8bda9359fb863780aa67b03d742b9091a9e418292cb7dc636f1d345727d92f810cc1ec5dcbea1fb4a5e01db6b57f0191a8e00db663a26fac1a943a80f63724e7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f360b66cb0b1468a9d8a0347f6d63afbac2ea09fc3e1186b0c8ff897c157a1ea64af1018de9e7b0f6eaae362897b16e21d613afeadcdeae526514714ad71972d6e28cdd0e9ced34;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h606641fdf1c57cd44d651c2d79a686852c92a7547e55e61c076a5ecb92feed757e4956b76bfbe3033a33516fe1acc6f12ddba91595f34155baf1702f8febdea9aa601c45c5d5d125;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1fb212f4b9f5bc2761749e9fc2261dd6030eb46d77c38cd8aab957725ab7bb82532ef2b3a750c15d17f92ac0b78f20736ab6bb20b7a061e9a248b4d39dacb97dc04749b0b2ec36df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1998ea48197cf318028f5b391450dac9b08a50f31cf9b076a31df2e4d99f5d43a97ee12c597a1a13d7c2639709b36564d0db5734710923e4643493c65e575ce22da0d18d2a28d8b3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa06a2be8e2c32281e70fbf7db351414f9b5888adb07ee6b94d8a92a362681cac33c4a4b3b586c4f15111cbfec4c19e99a0185d987540ffd843e7b49452e79915596e53ecdd93eef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4e5448221f010ba45953acea19de3944438e973eeedc5eb6c420f9ed6a91230659ab11db3e611db2033d20e8d7a341ac6be875942dedf7c7738be0907d3dd1e8a058539bb831253;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb55491f46e4ef1f5d0f1fc979d99d913a0173d5a91b2758c8d58ae31bfa66f5338a92864f7706b55ad6d6f8f34c53a65930b40fe604fdfce07905bb6e3fec3b5f31c87d1aabe2162;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6405e20c562d51ae92a9a0069af80a8ada4c156f9f1dc0d21413999ede23630193c0f860c5541ad2c139b13544f63e9a3bca143c40f0318dc6ab164089138824274fb551dbc8cb37;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6625505ad5b3df9f9021d68d9dd785b7cf7c73c302e7d05c981eedf5eaf75f8a63fcc76ad8e7acf9ff0ec8bbb6bd17d71602869ef2bb796196a6b604a28ad231855596b1df273fb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd65a034ae0e5b95a3fec5298f5656832194eb1851c15aaccf3cb1eec43c75b89e0c40c56926ae31d0d8b6903a44d6946566a8255b45f9fdc2be195071c05aba16957f3000e79c67;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b5db3da554e50afa6b7bc390dd9aea93c37ad636b355570fea604b1e65ad919db647f7857727d36e531df3e406baaebec35640f9fb926a9240ea0e63f28c755d973f4ddbebb07c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15a9cbbc5b799d60cfbd5679b8ff4a3552fcd74b547a48ba33bf6591c57a4f5a02afbc7ec33a1e77ac521255d97bfbcb9210c857349bca3149c85ac10d3717c367926f883661a9fb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2127a6fe7825c4d15eb249c4737c2046bf2648b9c94c3effa37ab3eedc1e79b3ca87e1f7178b859ca4434ea441f60fda881a236f1e069a797f39f91028665a79f1ff632090db396f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c6904d336fd2b93fca245340a70f6bfe59fe4652dee2fdc3923138df4887f0d08625874f8355083f8e85578e62acb2db42ca3e1ca66ae9e90e23199654bc727287751d2a082b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7770e11b14cd7d280acfab421dfb741fce1e4137fc22a71bb5967137fe6d73975e9538b50ff1c7d15d610ba309ab0824d6c83d1968ba4e57cdc5edd40da30447b47bfe3327e631;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74088df3a1bcb1bd54d132d74fe6eb55bd1bfd3ebe6c47bf4ea125fde88dcff8c4f40d29bb08b0615f71d3ac97091efbf680e511b5d685bc26fd821a23243bfb2045bb17b514704b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b7fc26923e71d21d168cc80a4e4b0b07099bee42c573870f0de15339f0f8822cb86ce84e99e2887ab6bc4c4cbeaf03b43f00a2bd40feb4c7fa4275aa1dd06b84174d9a2c093991c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha39b9e802e914c0ddaf5bd62f51c5a40127405adeddb17d5655e4c61182e654854eb1092e0f6af0a0c25dfb2b23fe1ac17170469c69fa4a031516d3f0bc166ae3360905b0fdeef0a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47eeaf83a2a6ec8b00959d2de4219d107d744221c3a90a7df5604ef037bd0314783269292eb2c54b8a4c236dbcc0ac0ac623e60f5d9e598ed17dbbecce1734ec2b11a96f877fad1c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8d0b72d5ed2911ecc334a62344cbad90737c85c95978a8013b3316326a01953f4c244e9496f7b5395c2223f6031f0cc173645d2425c5c9a15db853052e6da015af7edf7e814112f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71e066901fb4774180aa6f67446b710fe6a2124c0831dea25f0f0c3283d2f693cfb5b2c917e6e15af1b0fe38265818a967fbafabffa3e66bea51f3224b68ccaccb75e05d110d193f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2fefb4c7689d421383e3c4e2d03b6504be25b025020690fbc9207004be24dc90ed1d5ed6efca3934dd1af3b253c6e6dd5a5f8ae654a3f244a22062e791773584244b4a6166d9962a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha65eec18aef7522a7f44c2dae60dd5adb97e326efe5f2055771ca377415a8595e25f8f8b0cfa253038752c5bf4629243e01f701e7615ddeaf63fec44a0cde91c245793b46cc73ec8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h153b5ac6a2db8a9cf50f7f99bc2fe3e474dec34f5695409a6bb4726d0d0d4f7acecc55e1dc2a92bc2b47699ebab94e5168f73b4e22b6e94085d8da25c517db29358549955c3d2f18;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6610e18bd0611962164fffe03536181d2b4fe54daed8d8a6f1002d9fcb62cbbb8f75c1035501148eaedab526513d0283d7454607df1f0ef01a8152f377cc4f64988a66b03d433643;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h144c3d280e3020734f70770fea1d38a9db7cea4df9e06ae6d052204e58675cd369e429c7c5c011b723a84726fde10598e6a36ff47b9d509c80139b9d0aeda75abb402a0f4c3cf41f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c4db349d669fd6744a4c3edaf21d28622caf0ae3ca8754fac354f82e772d9ac7ef264d35eedc3834edddf2e883063046667882d0b678bc02798e1ea194a19c122df909b440bc737;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha13932098c0234abc2289b8980ea2d8f97d684d5c347637e021c48cfa820410e9cace3fa1063c806268e3b60a9614a18d685fbafaabe369c4558bf27d9fc65eadeb2ce75a8d6f0b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68b1e3f53431fb6d43b1aa1b8844586fc2b8d35236f7af9adda1713055c9ed5ce05c12b925452be7b7fb9321bc79c471eb91aaeb2c68d157b89ea19803b6d2896ff6dad3a2dad553;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbff022877636066af93633f86aa78b5f116a97fa540c58f42af22234e57b91c6fb7adb229c838ae44834fa42dbc08d14b6c2b089daa997c6eea2e212224b58bde3a082f80eb633a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6856eacd0319e3bb5e1df9dbbe0b39c0168da8b7fd2ab5787fbfbdb029b32a96875b48ea657dd4e06a3895d3cce7ce9a8b7ea6e10059d87c5b5bdaf457fcabdfca285254169b531f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb4308193cb31bbe2438664587a1c7263e504e22b29ea78d9e4120a31b9ec34da8fe6a092ad2d9164f8b9488cebee7899b0d96f3df22bd2e7f1f07969a17f870de6af6edc5713b25;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb83ed96424d58bf7b026a7c5ed1b13303a5ccaeb465fce6234bbd1bad14e5b6f70b145503aab02616261b22bf9e571980028d952b63230a4b83c982bafbe4714d774e7d2eb8119ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae3886e216318e65696fbdf1fc32717d24cd34a29dd8710c91b689bf08b46b0760cc2f39fb0b3bc5f7b2ebd5130e99c42bbd9aea101876a725b7845fb086ee62cada3ceb27bb2868;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbdb94576a9bfb57c3d7279b67ea83154ee502a46da76a698b8ba2c483aeb5f62e113e8b407a717f60d6b748349c24dc6e5648baaeb7b3daa392c1c342247d6e80026c7e750eaebda;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d87c477d4545b841b9ac30f92d3b9745699f8cff48eae2d7c29c18937bdfdda2fe847f19f01c0e7ddea86cb8262064ec8d156965f249d420191547fbf0d65119f516c9c89b3d5aa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h261c7a412edb90f3eaa2758d0683bb03568efe2cdf16abfbedcfdb3d4f08dc83bfbb0d7391b0f9bad8b2387a0140cbf54313e5b06d5e4a0e6f4ed78ec863d8078ddb526c8ee72d3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e004f885d581b9610a4eaef86d19f2d23d32fbea222cc8f7a2482c76979558c92b51e0e0d439bd0e6ff0bf6ac9b8d4b4779d11c29f5936625b53b219064b8e2dce2bc090c72512d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c2266b16c8cfe7be8bcd7c94246a04992a7607d585e348de0cca3026d3b8defee978edef568225e0e81005ce917e98cfd44dd43ec5b2161aea2e918ef5a6755daaba4b0f2bd722c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h276c9c8c4f0c016ee5ecceb3b4780b720f87dc2231ff7dbd82c1558d6baed93e55ccba396f93897f3d0d113668c91282f01bef2db238aa2af74f5280a35b681533786f36faa2f79b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62c66e00b98a6b93c1f585cc006031357fae806cacbf783cef9ce2738dee94ad9ed0b8c05facf0e43a79f95296ee505fabc5a8fa71fef9f28b9e344f3e79b82262f45d86ce6a647e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc1934fd6f736a04fbc86cf4fccb5f9337a0178dad820630b6353be5019b57475f26ac7e8ddf42db935aea035ad8058b5ae5475749ea8b09eb1ab6af3d7f1dd9352b2a02de9d76b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b6d3a937e697d9b1728578436ffa32a442c7a02c840ac00728d15f6be770320f2e7b479b79e0dd167ea79401ddab3510a0c6bd20f971485370c57ba6a8a91bceb8ddf638dac1f7a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb00b9bc1849bbb07236800e5b28b89818c6528aff9f942c68ee468a72ce1e55350f014b77adeff2084cebca5b46de1c8803d2c39aac0943547914958cb0ec8e460ea13a52d5873fc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7229db8d461f68b1c3c8817d0f63fdcdc02dd26ab95a05eab36fbdc9a60cb173bac8daaa03a69c6973a5e4b56f91fff6712ea33059573daf0d8da82c2163931b6c8002e0dfbecc22;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9eb6fe10ff673f2244f7fbe34d4db046c21c03267018a70db08265f07b0d26e222e04912940bfc8e9dc12c4f1a966faeb91942cd5792e2cccdf98613792a7865e9f65575a0f6554;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb026f6ad51024b8c66356be67a20f5a0498ae24ecf99b8e07b38cd0e68485a92948b81b196544f35dc1d7944c3aff0794512fe0345591092998ae152007c1b2ee9e00a12b0a3e9a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he066ffed636cb71088d216dd9ea974adfc3d6a67498726afa3e6781f02bff3c452b2df132452ff224f30ec705ca83c0ad27c404a125cfd1afa60e1f0a207a93bf1181b0a93536a1c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41c169876f6240c6eafbe4f2dc415f30990f6173d4e26effb3bac4a4beb1dc05a15e14b0f0c4cb05532645bed0c8019e61e671edfba11319a935a5bfa553ff45811f94439f16464b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a3cefc179f7a8fc003a9d3fa9c8d4c92865df5b1bda0b6cc4e387d1005cb35effc74e10ef6d4f3a535e89aa341ad98f200a9e382b2cb634fa66618205edb096a7c5428403ca72b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf889f50ad1537f06402e8f72eca32dec063fb5c85911e8f911c13cf1ad14746394fe1ca2e43aa99f74fedbba4de18134cb4edb14cfb83a1c332c03e4533ebd92a909452ebc03f31d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3791618ce88c6fe18ef0204d673131dd74a2b5749d7c4f531f7eaad9e3bf422d084dc5151b5de55fbf7c4909324ec15e30b5c3bb957804438d961a28832df6a4481c5b16b8d561ac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb04c0370b130c784270b61e2519a040c02c688384657d558ed471f9e96d8d8c81a6ddc481e1bc653f961564957b02ea044b986083e91fe5d9db525209396360eaa2a1109b9ed5209;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ba8ab6e1cb2947c59b541f86080309a5268df2f97025b23fe1debedbe6164290aebb3497c8d27c20ca07a338374a5976524305d33219ca36adcd6d53b2dd530814bd9af0d3db19e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb244c8476469baf6d5e189b65d25e91280b5c0259782e143c739320a762ca6c768ccd1757b89906667908d2920033dfa8ae23abf512e8d2240b28d6d99ff14d8ca4edba4aceeea9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9bf4f1e3974be8fc15f5689c383ca3bb16a74976ef75cedd933b37eeb3c4207f38ec11512b59d27c8da1aadf3584754cc90be68e42116d2811b8181291be1864bc0d02653ecb8b77;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5cf2d5943f33b11ac7308c4d86246f731ac42da5fdb6ad5540586bc5f5c4a9d7792baac8731bcf463cd76b5d5141d6e89f4fad1813163ad1f4a2f2699289e1d73f699c6de1866337;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70edd7975c14423595380ed8d9c0444e0443351302bc0513f96fb115c011ea08ebea60d59341235180533d9089f6006045a6e44d38702cfde6f7546f6d94f22d29443888a5fa9b07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h699b4768e9201b9bddf28b94fc10537b57ce610371e284948df9518164031f66414e87842be86f42e159250d534d4ecde74d8b926e958cf06cd13e9535876d9ace1f591c90fe0c59;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50379b88b7b9d9e5b116422a74ba4f31f02095bd3f237235735914b39c43a0568a1e9afd64c24cbe4a8bea5d48cff671c2b93066ee74e9460339d2fe6ada460696ab97bbcc60f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdabd06289e96e07c412ed1e95b98d668387bb7025053e02e8f8b3bc180f5b18c5324d55eb511e4398c0e451e2cc065ff53a241f8f85200216cf6c15733ec4b5ba106b2cd84c11ada;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7531ce62401dd66d65949cc418f83b4427b55b0c06cc95960343869627bf30de96998445b819c0cfcc3de31335f0c8b03e4affe2443d8da4bab49b9c08929103678d7d0c835976e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e8c2fd520e129d69dfbff42f33e6c5ad679a4067fe3bfd4d78910e853e0aecf8b915d19dc620c7dd8d1f2eb5b476ef63984267edca92a3eda18c82c972cc30430ea65cb0c1389cb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33420c29462beb26e3263a925bf344a353bcf6604c2958ef2db80e182ae0fcff22e2f60a18745ab725b3bb012779a157501d1cf032375cfca811984b4b39fe720890e4a0b6207c51;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hafceb0c1bc725bc5e0536dcc32c40fb3abcfc81e636eba4aa52cd68ea99b4cf7455c0e095e4c51c3e192e123cb51e3cab04aee63400cb6344a11ced4a0e6ff901c419f556c380067;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd01a6b1457634a8b1460229656d18b76d92b3789ff74cd295a95be996412d58416e7c648522ba44b94286f50057f4b8cf562dee50c9a73bc6d0601ceb9bae46a66cb4d18e772d0a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h483500c45812be25c2c6795894ece260e1809aea52e10166ce5bab1a23c1d1f2527dd22ebb5c58b1114beda516540e1bda8ffc2c042695e1a1c25997649251e9755fe6581dc7141a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h820b2ff2e54d1387fe64defe039a98451a28dc4b767a15a88815c0aaedb7ad6c4e34cd7104cbc17bf665bca32b2ade1e8b067c77bae8956328faa8136119c9caf7e387a049f8dd9d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3235f8ecfce48307fc41bc4794a8b9f804732af4b1c032c02a2822572f0f9e81d1811a304e345976a936062be9e4734782872fccca2a8b51527a0f61bca4e625ad314fc887433def;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haebf30da2424bd2ff363301a335b417bcef456679019cd2efe3da30acccc536f16ed91b4b80cc2aacdcc9bb47861c63c0760f490993a791a60432d0451e729a6be8d92b20377c6de;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0f450ff903cb18ad3addfd8c7b88011d3e8f7e1acbbda4b53d4090525bb5eaa06d94deb2665e2ccee8d4eb21308dd8f116c9685c98527f6c170f0218a51d90df546ffbed6bcc718;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a73dd660ca013ace72485a3d8d950ee4ce3ba2138e243a0f4e1986d4fb92d42d4d3a595c0f7a146376990e003b5400e8045dfad6d6402323f3703ee6bd0bded5ca2f5bbc5b3003e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haca97e713d082d0333b3d3af4c132e832123433d68aa112546ad8aa001e0786d5bcbb506dad96b5062e2a95806b415b6d7163d9f6d74317ff2dd5fbcdcdfc53e94a64946710a7e74;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haaf0dd88096ff76e5dca3f3400c4f59652874cd2f48cf3a72c141061c883ad758ab090a50c9ad58e42761db6f1e6ad9349fe374c58411ee209cc8bf198b643cb34f1aa0e02eb4189;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f34293bde4ddbb90f80c7782d5018718487e7c1e869266670f1dd3055259200f425e3fca76f4a3770ac2c5dbc1d912889c551fc8a505f1e419b17d263e3fa1d40c05ffc94c7a076;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc9cd03338543437e8e625df4de6ee2f05b3cc78dbaeb7c67d5dcfc443ab05ea5db470885125531a0d952d9022b5f1766eea7e87343640d6fe14c2957d9eb7b9181cf31338dda01b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67fbf93973399f6ec037c9d2d51cdbe515298a842fb471e843a4fdc74e6ab796e46e5a4a9732b839ea25471b8e9acaa0a1262d2f8d6927d54211975eab083a9d5b5f0ba186f88192;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f659626128eccb204f264d0227ec729a7e86875593784b1b52c1d2a84432b4c4f306997f7d78b930260f2d54435728e04a8f59ad8c75127137829ae028ba908da6f1e6bbbd1414;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27aefe9094d4b4f7cb0d07cb042f290a076cd5f56f2349beebd90ec66a2f1280ae56d2478faf9430f81b767e5425ec1f72a6e186e1cf54c5f927a21a66580a25c8a2617fe3ac62e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6f1d9e7893ca512315563e98bf27b619f8e02bb3f5935b9aa9ff2a199a84e6c0df5f44159f29a865cda6821f185fc01a81fa5fa8239769f5a701462c50051a7e4abd797547dae88;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he05a1a8d4822cd58ccdad70008831595d3d041bce36328ef17a4bd2c3b5e086b5d236880e420dd81e33d9fad932653617091edb5bcc7e534eb89247ccb8935bb4329b672b87b5a7c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56a3d4a1086d383201fd39a9ba84ac999b76ebf8e207872a767c2ccc34182cf65f51fb951352faf664cbff002557176fe06a36ec72b24a9ed51b3e457c5d3bb68beab489f1ff6b06;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc604da8cc7935202761c312ac76d252e12c5a92a9fbde587af0280f801f470331a78d338ec233d1d830866fcf2c31a7caaeaea775eceb7a5e1adf0837d6cec5182b96a1193222771;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6771bc060b0265caedac2acb63742826c035d19df7307561b2c4e7ebe07b7bf4353a29e87902e65e1c6bbcf74fcc18b2ea7641e27242b01bdb1445f1e11d71255d404f9c07326b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha34b996fad4bed03b0b436aea268df415bc046dba4e6992b7dbb60a77299a4190cff088bc4cf287154e039e5d8c3caba9e5e9fcf586584d003f18c3d65703e634bcb4f71d320902;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1c69d96ac494513bdb7a05a7a572a35e6d68edaf2a2a3f9b657edc551e228772c8a0aad7bcca54871f23b753782cfa9d76b6d64faedb8de30e9fbf030f568f049badbeaeb957527;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc740620f55f8ae22723d0f72f76797a3e8794f2bfc8cc265541b0eeb08af624264b3d97d9320514f778afefd85d8cd2da4d16ad9ec9b760cd4f0a678c56c55c76421eb16bb5c8e77;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a696b2c784cee68a28766618010df8097dc9faa20e39617ed66da3b852dd1b5e5c54f52976f6a4578d9b153b84a709d86c5a042d84fc9e9a1e20b2e2feefdbe04e78a1ce540a08;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a3c6840d39e967ac58951781d9565571b041a5031db8d1745509e0274d1afbb1648dbd44fad08642604404dd05d5f76185edd451c09f4a9ad26c1bc5218f19c115bc6eb2fd1b0dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h971040bdc9ff851689e76e46383f786eeb38d9d61228593f467299b9060cef10a700b3e945ed6fbc3ff7d247f7d8cc00295e458302489c7879243a2fdf8a094f5d06ff032a7512b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd109a93a79af17acedd4da2dcbc2d062a5e2b4891b31c5ecb71bc15dde4c5b42e240c0dc3edd02c36bd06861e3436f3a77f0035d7306e1f7da0fb36c9de392cdcf31341f9cbccb64;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca7fd66e976c1ded2751e66dec47e13b7f8becd416adbda1bda24e3a2d068b520e0d050e6d89325b3b463104025d8c29bb2062b683a3e205b6b4d2c8eb368f41219ca4b30dc3eeab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb77d256e8e50e56ead90ed01433c870ed8c60865b102c44242845e6b9e0391c8ac80ceb4a8abcaae7aedc3467c51c00e34fa18fe42e904f3e50f715fb98b59fa143a3f5ee967ce7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha121bb9bed9bdb16efcdd8452bd721b74dc0cd99029cfe1cc0fc9a4e8b41618dd369a7ad8cb05ad1e3dc289911fb363f6f64e9f27319678a0af045326976598914d20e17b88efc42;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a3535a0f0a5f8ed54f95fdc3a125846c537ad161cbcb2ddc3778f50f01eb017de460fb51cad61c74715321b295b880a88c70ffcd18da8d2d049d8d3070673004dd37c89959bc184;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94422a4369c3914ab10d016a5a27b4be9798e32b97cb7f6daad8e19a667bd36deb36520b4c6803f5dbd213624f0feb25e8a23eaa3b40d25cce6b7b560f1f2aa652ebada89f06fee3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbed67bee13c208ae8431d334af755656590179253c22c38ee145791f5b5888d99618e69879f3617220ad7627414e9545a9797c7f71494326fbe8963161db7b221ed0d7a4a1ab966b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc0222c5081cab516cc5f13b6042742ef5fd7b363f7a7f93b78cbba37ed9b97aee7b374ea3022f0c0215adfe80f2d99fb59302ba196eb7d45df307379060fa2e2d9f86b71fcd2988;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4bbd09f70043ad1c7a675b0b9149b338caa78d4e6817703c61f2a91a9877984dcaa17309b04362614a573ccc40a51ebbbce514d4b16ccf79638a4d6716a80d83f07e2eca004ead51;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb19dab33613ea1894de184f00a0e023a7d46a52200240252b95a1073aa67de291f2b6a23f3eef2b04462bf5daebb3173c260bf2e1e87a404aa4c66c983b5df09c88865fe4483855e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbee8e16c088af899e761bfc39876452d5bbdbfe1a3a68de1c35f24f7a07a7b775a1fd784214fffac615e46e284f25cbeee8046b56987a7cfc4dad84d53dcef97fcb92e995c64a813;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc82c1a2489ec203d1597db5fb03e507f2a626b95d24c30d3c556eb43471f35d73d438beb3e9c389f4d0a35ef4aa0555da55691f16133268f580fd448e105ac2795adafcbcdd844d4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5517ebbb1cdbc5ca5649baa528160277b3426fcd00241518dae1c67fbef82aea7c07fa23cf25075db4dbb00d57d08e0f2e4d7e583913582119d49dd5760a5d9c687a27ca1a7f13b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d67971f5032aa0f347bd445813a0c9516195b92e4ef9d0b7486d945c96cf5825aca4e908b43ea01bfc7087837aabbe8d65a8333c145dddbaf1e7299049c61891c533e76fc1f4ee4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h419f575707483d39da368d9cdb51055f9b40f2be8ef9ba0e25dd5a186dbe0fcb9d17c6141c21ce86f2015eeea8e7fca87aaf7aaee0abd3bfebf59956a333a1328bb8df56b4f3385b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76e7c2b9a71c3038d5be8931288bafb18ef2c443106f25c6e5bb08438f08549353b2faf95e5ae62a5c6ee8a9dc9a6257939734ea55741d891553d3565b6665ce49e6488bf1f0ac37;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69b52b8484525afad60abb9b388e1df4db3a85325f61818b960bf1053efe9e68439f5309672c50f268b3554b90973fe7193ab3cdbdc23e9008a439d329034a0d3747e69978b49757;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22db2fa7152123ff9e2df3254fc63597444f1a691e149ac4d72c189d296623a908e7bc456cb9428148417c72eb2257a6564d6c7822d066cb56e452aaa73fbf52624b81cd99a73037;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d6fead4cf08a3f5b49cab5881f9a889058149170513cdead5caf33dc7428a725b3200d284166f80f151ad5a2507b93ee43970de571cf60f861370369726524f91a73646101a990d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ccce355a27cb72631f20f74f2be26d55c4bff7de434c23022c7d36c28dca0f747a4566054709c1df775edc2d7e0095402c4d7f6744eb82fe2315dc948a41ab0a0c160d47d0ed067;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c4b4c3f9b394836a4a8889124ea9e448c2872f4c1f674a4218001bc92b11e49a1dcbd2dee20f72bdbdacc5d0c314d49426a3489ca667d1bef0b189197d013fd2d8ef65b73f2d9c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c4388f6570ccafa82aeed188fb3d9a026c517a5108cd6660770d0d44ca38eef06d3effdd88224415611428c7037e9225b4fd550ca4f09a90bc3d8435c62b5d402f34ee48de7c990;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e51b39743247688be73c92347dafd960df08f48a5f2f02b3372ea55669510edb5bea471aaa41f231e8078b5df25c64579645f0b363b607d843a5e6245cc25d84620a0914ebff725;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbac0730939165774049ec89dbe9c1df7a4d681f5172e35b1e655650eed2ab39f6e85ccb8c9ddde605d4fc527369e26cf0d7f101c07102208c9715f507e9f1ec61316a132def093f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b787ea3406e68e36d804ef682e5793737893741b8cdb2cfd0c36f389a774db7c6694b10a1620f789236a95814d4a07f28428feeb97519872efa13e4a4c0cdea186e5430e9124f43;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb06f31fcfc994d0e62ac5f230b1d4c1dcc11b99eadfbfeab0b699e86485f42de0a78291d2264997c97d1972d5adc7e7a092416f8cd0a59b705ffe28ec025e9c4c8acb482b8ddff33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8433012896f504c077249d7577771dac71340fea745341c69828d58dbfd22eb2ece95eebc25576a561d568817f2e4586257ded8ed97857941228836517d47fa142cacfb6e9965ff1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47a3ed74949abdc7e45a5b8e73995337ec21673fe1e8409a8271373c257262448bc1b281af28be10d4d25c8d75864fdf329436cf5baac67805cd69fb0dde18f2e919aa363e6691b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h39e61017a00c98eae19232043e1484796c99e507df2af3862a6beff678c5cc31de58f9e961f9e1ace41740bbc1ee727a6c0e5eecbb6e1d3e3022fb91cff8157f8bfe487fd4b4a942;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55ac944fe5628bf6cb6a91291dd36d19fb2b849b442e5559a0fa95e08bc7ee86422f46bc02f241fde1f630d8c214e2e04b7333fdeca2b60e5e7e2871c9490fca51fb1fcc659da5e6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h594f42520f84da3721669a40cf603aa68973de5758be0cf425e88c4aa67f31f4f40cf67f534fd7ef62fd1c37e42fde108e96f88f353f0dccce40a77f5aa863f59dba1e0cd5034ace;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19faf5d49b925e56fe7e89b67b067464e981bd4bce9eb3ce305585fcf449953ba98eb03669015f8c503e44f84edbe2ce142d14bafe67ad71c5e23cdd7234ab8cbaf7351994777dd9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9907625c4b9d5baf17565c5ac254efbaca1eb50c2c9b0db44f1dd67154b95d3afd2a5fa806a26207992d326036b5bce50836ab0aff258f98cb00ca629394c12db713433b7332f8d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hccacc2e2624ca6685418fb7b48cc72f309a0ec153610cbb4cafc01b464f0fccab75b0264df3232bebd75b5ef8f20cb0dae1ed9d3b0f1e9db4898b34758cf341d9102d4a9820bd65a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc19f73d3cf7b582ec8f3ac902b782272d3ed48cf7e6c7f21ece2e9eaa0de12a1a12c2376bf68df4510bf6b9faa8deeac123284b342b6651c58148a5189f76f9a17acc75fa4469c27;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32e1aeb0a078f3fe3f340c5c88e8ac7d2cd7c3acc2c14b5e7a88cf3d13999a58457e2d3a4795d400e1e34bc73168b0eba84db886b575d27fe4303845b5a3fb195e8b10e4b5a850e6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h310be063f378b47965e0e569110fb7ae7e69e8c625706263ec4358b4c8fc2ea9533990a729a1961bce47139cca1aee75bab461387e15e767c28810383a12a5fd730014ba7818a7e8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a47f8f5c8a981fee91719c5232c7d183ee0b83cf943c1c74f509dc2afe66a3d72261c5c7d31c4eeffb3447e8e169724e7cdbd6c6b0b30610ae8cff693145235f0ab5316a3afdb5e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4acb07fb921564034ef3863a98f5187700a2a25be63b35d9a386b495655a53c9e5a71176695e6367c3f604dff2da3d3a5ece2dafdef09dd58958c52bdaf9ad798bdda33f91b1adc0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h449b269bd2b828ed7b9d6f641e98a1a904a2c77c1a40ad0679a95e3ed5dbcc55b2b6b14dc62979090240bb2de8854925075013395fffffc2bba88bd1397d5b33c6b078d25fc2cd4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8b4e7ceece9b04f84ac2a10a792a17e67921bb8e7a5974c9791eb8956be2b8c089656fab800050fbd6e80a46cf005ed36d1bff47800ead6297ceecb88ca1baee3a8e3a5592c530d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h829a63f57272c5cfdb160b526b1e03b54e748cc7e6416da8427b46f40bfea4b2ffdf61fce3284f851f53a048d33b23c8260f777e46751aaad450543177416fda5e1ebd9e660a9905;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5786851153c4da4b1bb0c46e59404cebd61c03e5d317c78e61433e199379f97e80cba318954ee2de2caece452748b3c64f0dcf08339fbd9212995edec7e1276d25c9bfef8cb9b01;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h762aaa95e9b5f58780320c95ce24f6438f9bc65731177a2dc72c0b84bec0bd23c6baeb9f53652a045bedb1d3104f69b4c40501698aa98e46ce4b3d34232b83b834637a992b961d0c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19e3c16fd9a544a91e89017df726e38d2e2f5d64c73939ea18bc38dc06de4f0091748f7d7980a7b1e0d7a4e1db8fce514e0128e183f88db702ef4666066320e7e7a8ac4510f3b39c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90c0ecb299b881beab8a47c0ff9935ae795fbc3734f783fab4cc31b690cb1f2f6c4fb68dcfc249183968a5908b24c759a577585f71ceebaa21d8275a95303e97be8d7819e1ca4075;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79895ab18f7e76c7cda71596ae0ad1a0e45bae00fbf21f03943caa8baf553f11c5584489e9e9bcf27c6423a35200d9bbf7d67a73cd48a9f3d0c4067771c7148c173c8e9f0f62e849;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36f4438384b2abb5ef4ee09a6066f6d9982b2e2d0c538c9743ce379f0fd4bcc426d9d1e76ebfe8999008cff9c3d2be758d4b4c3e8131581e639f266b2c1e1bd70c7bb58c2dbd5002;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a734930793612bcf8a212eaaa7680026920d1ebe2dcd2dd73f666e08ce29ec0afc9c4cee794818f6169e520970f3ae2ee3bc14fec0a77bd603198a69945c844bbef6e532a35a554;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e8976df6e10eca757357431a8eb63c37871f630ff72d11ef68c7a5c61b244dc221bc6d49e49de31fdff77aea9c6d499e106813e1faf5a7f82c03d162ae64dea8d13692617591885;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed55d3d9d27275220691545e6aba1dac886acf74bffb89f20d343f5bb46a1735ee3fe362cd8e864a8a4b650a1dd8af255a8b551543507e8568da824a325fb25ae391dfbca8d533ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96a1a051aba774ed8ef4932ffba8c96f6852aab9e7a585b8c7b9d11be99ff5b544bfe3090300556a5e2c892ad411a5887ab667b7d157b14d3598ed7ae05b47f7e9aa7065c78efd77;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f9124f8471f2194629237f4d4701e598bcaa118c2ea1977fe16e8f41699e99506551905a8ae30cd2074e91d6148df78b2ad9a28d5a1af7ad051ff9185c3510bc78725c98d31207;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h749ef8b19b91239253ef965cd207bf68c1563e50a8f648e4dc41fc5f5154ab7a5536ce5c83db9c56d5db6291a0fb612b819737ce6da4d1d9845df798b06a512ebc842db90c45e3ba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4171111ca5a14c3a0561aa8b23cb7fa3ab250ebb98a4fcacfebb9150aa3225becdcb5c51c538c987a5697700a4faeb06c83bd0082c70be6332f2275bc280a516703da331ac7c64be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25e1a782e68f892fe183107ffee6348c22e784601b1da647dc48b7edc754fbb6e5c315cf215ed86ae04fbb388c1bd95487c19abe4c813bc24610bd6537a00a69a9e7fa3dad5806e6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7677aefc0d901f5b76b072c82a33a1dd668cffb6df12281221d6c11fb664431c5b6bff347d2e2019a26d795a394f45088ca486f879f5793fc84760f832486f3385eb992c4bbadc5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h993ff0ba05ce30394dcbddef11f169a3f89b2a026ed7471809fb26be98f68ef475ee1afa5c137cbe8f4c5696f65af6e2bed610fb51720ba883959f6fb943711a9cfe2fe14bae1c44;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0e24c8519bc55bf9b7ced6efcac66189bbbca6a91776b93699a4128c95aa099ca93862fa37022dbaa3fb46e2a05e519e6bc0c2846afd8905444c6d1139864d8cc02620d173ea22c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2cb108b1ddc774ee51911fa90468151062b09197c8029539679b2f5546bed05cdb1d02c1db304eed5f37d4a119b290ca12c3141fc545a2f813918a6702cb2761d3ae64203c04ac3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf95ac254f99bf39a5eb80b06574c374c122a3863a367f67e07a6908346709f2b7c46b057aaff8e633d31f592205a552c69232fddd19b89320602251cafd844e0cb259848e678ec72;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf3e41925644031d9e41a4cfc7167ccea644e09b3bf9fbd9573ca54764f8c68a941dd1491b3d22cf96b05417e3adc7dc78bc0afa7681b0cd9541f6bcc93093af4bb0676a25496ae3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47a27731522f80517e5d5b623cc9d3c2e32bb1f76aeb5700efb59295c2ad4e2288c639ed83d3d32ac32182199820991fab4175f5f2a9748bc4d63169e0cd801cf17b59b2f8325b6a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h321684f8e7fac203a738f2c5261e6c87a4d5de444165f90b735748125d6d3cd5b066380603601caed14aaa67f62701b5a048b0a6f27941b64c4c10a27baeff0f2ea7e968ddcfb55f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8eb4b1bf14cd4d41da31b0a54b2ffbdc0f1b49b4df9452c0ce480b06e97739feba974af58cdb225ae6c820f459023d06bb7198174a55d3e7c986b0610b28a9bb7cd90b519b1c7ec8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he35c45e0befe68f4c770aaaf8026a5ab1822adb0142550eef413bba875950f311439cc8f8038ca64435f20e202cfa4518ff32a620f61e6366ca281858e8469737cf3ffefcf381fe5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4eb3e8124777eb73d5def571b05a8f636975852d05afc6d70d5bd8e87d0925137ad6f1073dd3c1c8df6b528637b918ca8e7c0c7764956735e1af06bbb3203dfeb03fe118d9bdb59;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e79138cec5a5454af803987ed4a759caa7022acea68ceb02ffda4826e847a89cb714ffec73a060b3053f320d7015d880de8bff8e80e6b55244ecc45b18a2ac4549ca512279d9afd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6bbb6cbb4dc632c3c4c61438445ff3dcbccb14c7a38290c3befc4a9835c194fe3bcd347e64f40e083b685b0289ff36a969dbb70fde9fefe7a7ea1dbb0e3b16f25ff0709222408584;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c025be97b411ef97f79b2c6d3fb6679fc3b7091ce955091a1f70982ad79edb050a39275d385a7ffe899b9af52016c24d4f204216aea361522b489f1ec277fb8dd983834c1f6af5c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b10e04db74f7da43c2d270a8421a2de86bc3c5d8d6cf39ea00718771e766408402c738b3ca425655c6c172d1b915fedfb2c621c2e247e33fd2e5bf6957cae281bd92cc24107ce7c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a1a89d845cca4e715e7821068192363c4ea31a8785e7c18ba24336c3318f038153a51c81161452dd2347b4bcf79e6da2d06cd2df37d665c4a0a4eb3c729ae0a8f978fce2d4deead;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9479a76ac9175076bae7f722f99cd9ab9b1ef6b557af6690604690f2ba30bb73edbbde19bc95b86fe6f3e34368527649eeafa370979f0e796f8dd8ec63c0e1a94f90b806f004dff1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde85509edd52b104ab2b26a4ad395d5b5918e45c18dab50194bb1937dbe2f785c06f374397d0ae7e7d49cd1c909ea65eab6209c395c04e17159db166f0119db5878bc463b6f71e43;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a46d885b5d55da3b9e095302f993f54e871fb5e9276cf6e12d5e35dc21ee551938f00ee3fa31beb63d56c38e8b8d5b087ab4d93041c6972467bffd3f748bc47211330380104ca2c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had495d9149a48875af284df72066dba20d091469477863c128680c1fa230b77ca110974f4cf17f82774fc01c98b23a6214124ea017055bf0022d6df7b51ecfd26188c62084972b0f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc72592677677493c5327e512c211d5efedd08b08df990bbdbfa7227ca4af480d203d1c8f6f1670e38a032522401cddf42c19ada408bff7c0ee70e24b83db2c1a367c3466412ce904;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9360ea1da46796f6284e6e2f07689f0ac0f045d5d19539d1567d51a7af1526cc5886bf738859ce7ab654dfd282f83905caa1da40ced7403d4a87ad579724e3c3196b55c98941c1a0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4fdb56cf5b36b4153ffd66fb933f27b760ddd1013b87b872b954f37b91af36d0d60f6b6d926025302b290d1e60443833a5fccb3b85fb6349e69b7603196d520e4503b87ebec3e463;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1adf92a86ca44e234ec0133ac1c02b065b30a5810624f808266a41b85bb8f23d52efd3f00c1e7d51379bef9c4db97c81926019ed4a5dc7e819c536a01e9f32d1eaf25f5a19ea7ebd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b1e69ca157242b1b184c24bdbb6ef88ccbba7f4d5c58db2ac95f9dfd1a7663df107146a8db29d293a6a39604849145e29252dabb4d51660d40e0215f7eb6cdebf41c2e7e6dea9a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36d072add8852d15310461c8149609948bfc3161e525d3afc8f2b3bc6f20fb1111347845ea8301b953c05d06f12622c93bfb4cc7778ffdf5b188893f2314dcc3fd74ad53894d967f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdef18260897ce76f1569928117422498f0d296f1ca6b050fa486567bc0ff44ba537e0cd7e3dc27d5d03c365b081dfec6145c3696ceed6ba45088fd0088260922deba612872a6347f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6feb71d019d4efe65f9ee8b2108a6cbebcee870ccf0bc283eafa630caa562a921b7de8805cf3e3a71f3b32491af3934e7b2e56c18c8951a701c4a2b01df2c66482f90ce8e1b0f152;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c2f23bad7671d502652db46b39c20ca9319b3e695c1a59abc2ba44f3b6bdf8f66899a1b49a726fb81d8d9acff7117d71b36e51ce0352ca284a791db252629301987974cc72da7b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a972cb48a844c7715cd37910d1022c1ca66be1daa2b8c367a943658d3888a01dfa3cdda44d235d226e0ac80232a3f565b5aa2d08db8967a1199098442dc3f682c07d0bd9b7588fe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f983a1100caa85f2d51674c41fb07e6525e9d079b3bf49219901f7244630b2625e69fa30b59325eda75978a70899b1bc5cdb0976dd75a91dd6469bfe21189fab35822a393c61936;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h518802d0660e7060e27fcff319c7ec670ef05be7ebc28f9f6574dd0af734d40faa65f898ce3c19b0645f43ec2905759b3489b106e49bbdb8e36b24016991ea2ae5a9128a8c69a34d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3bb3083b653e3bf328e439f20f6506d08af217430cc2ee115cfad76ea34fe418c3f97e4958a7a0fb3f6c57d80b7acaa7d62a649feb8cc5a7178723973ab640e4edfa72be83729928;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46ca997a542c086282a55a39a68f5c699bf281913dda1beda5a3d16dbe31960ba31af3315d7e5b4b59f86cdf66bdea89d10a139c4e6f7b34df42d9a3c4a34acec8c9b58ec3943c57;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a53eca4bc5eb88325be53bf78c03961854a18dfbf7a5ebc5d227cdd52af5b859fb4b1bebc95ba50f4d18ebd548f32cf8a48cba9045170568d4735c28fe03f05a2a29b853d8340b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heea8eac91c4dbf43c4a358493063b8836b6ecaee1a6204098df98667e7153b55e48a7ae14d21f7da295d0d039fc9ff515166cbbf1dfbb8f08da9faf170ab605a9fca7117a32c61da;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfad6d42c9c25b37e558a1d20a1e6afdfefbf8e2a724d257931da40a85a77d9f3925a5f5e2e75aa6209f2e17e58d59368d73bbf17bb51bb6f12eeebe9844865e93b1f5eda000dd637;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0ee3297900ec70eaf811739c3d2e60cd7a9d1c1a49f297df1bc35ead6101fcfe1b184b4d2af68c2af0d9c61d4109df5755724fe0d160a3b22a742c24565eeb87472148fae358a0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d4310c34eb7fe1438924cbb7b64288d4d40d2062c35895487a3ca46e60bc52f6d76e2461919e146cbe9eae0494b6dfd9e208f3864ac26bfb36d08d10cce6393b4338c6dfb29d1e1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54f88837aa0525e12d15bd22b051bdb5389a208b0d868e12e29be923296ccd6e267894d3656d939e64cc68c8686176a5f833f663fc78425f0646fd719041a791a74c8b774f90547d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85a70666bd116d81b9af1bfeb7a2341e345fec178062fa220c03fc91d37abb8a84ccb57cdaf5d0e78af7b2cee40b7e07cb294ff565ac5543a9d183049f0f932d47fc94fcb6959f7f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5eb8c3498686ac197395c8f6f23a64adacc3d91c4980b0c4bd4cd79b9db2627e172b7c78fe3e4c05b5b788033fe45a6d847fa72558a7c2a4813c58ce74f1d4ea9091d76914520b5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef10e001592a9f131ce6895433263ce682daa75b148830a08e1a270371cf1cfc21a0bd6acc962bf7e078d441248507230d1d109f83220298f35ef9bb1d5a8b5823b3cad02bf05b89;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4de307050b885f18db0965bdfeac7c6bc3f1aa365a5dad08d6f567380eeb864ddf73fba121bb2fc3f29b20cdee5658582adf2bf5f8b28611ec52849149f2363b2f74bf29e654015;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc1dce3bc6d4e335b0a947673d2effd907df71f034d2e61dd0eb30c9b25ca8b809a6cff09787d19b496e35415f480c5380a1669b69437182de86b38960f332fbf9d39661599ab3c3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0329985dcf978d7bc1bbaa699e74d25ebc3449ebc986b8eab96875339348ff3dd520dce35ef79ff338aaab6094c1501ebf6c525967c1212b049bceeba76e903d0f9010c6e072e5a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f56a72698d50093986940df9bdcae280bb093e5e619bcd2d168e8ab7731779f7981b8763f02f0c832474928feb61e46ad5f4bf736f22845ea56cb620f1ae3afce5446a2918e6a63;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20c34720d2c9a21a8336ad191c6528c46bdecba1f22354580a52194dc2620f4c8a5eed18b54948023af549f397417cdae22e41e7ab6c7d615facb5449ce9895155e5ac1c0dd732cb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h288a2a221fbe861fbebc4fdf589a3e86a54e3b3fc3d9c005dff747b38f6a69bbc4317d7f107d804756e16ce45c0a171f4fcb56af9febac88b49150463290e0457adeb6e337a7665b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d8217ec7f2347a6271a7cc942a3a040b6c571ae78e0d1db9b5589e103da7cdaed2fefa6b72ad0f3a35505d95e2149916eeab64abcfb12bb56d4992d0950712e777d5a382832d923;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d769d1169b4be225757ed94a51085e80c25822fe2504c260f738b362afc8d84e50c30a80b16b4380e11abcefc38c712bec94ac9f3f9739ad32dc8299019ed71d35cdc42831a9e98;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0f90169bffb23321c9d204c65aa4e3efd1a4ba6ed96f35de864633cd7aaded5417a61f0df8e0654c49f591f7990b9e141677435083dfcf83b0cd05aff61c165af04b8f4b0995dc1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h781017987569b727626ab8c9fe6ba02f54edfd175267556925c10ffc5bc491a19519def0300a7ac3d4ae4452bf18ebb0c1c8a4b505eed0fc9bf15725867ef6c5c968d9d37e91f8e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haca01fce08d38d130189c97a34668b7b48b43bdfcabcd5526f6507c59c50e4c9497952fbde174a5736782fd4e88337d3fc7bfb87077f4275413c00a6e671787828f559723090c484;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed195c269212694d775927fdbefde9732456c8f10d3d7de2637816d56c779e7a058cf6ed8de4c6a8cdbf08f0a595ba5e9d39e1faa702dc46ea65e35444832a56c4dc4628f70e2970;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b790718af3b21034a36094a8379242d146997dd647ed640ac2a719082f560ca153a01e4da8c6d8832d54e52e531226e2f2e66386c0b27cb95152c05eacb8510b715c0396a9d2d94;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec91ba8da077370b8e7217f4dae1c6b503bd01ee609c11f5176aef6b57938ac08b7e5e55f80d6f2db2c3146f4865113da6746dd2ee87253ac8e3d693e834b7804d9ce39f5d551940;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd54c6d26eccffdf5de74113d8a91435aaefe9304c254689bb115b23f81e7578e10cce6aa53de8edce1022040c0bc53fce10787d01059a2351f6122a6a1ea4e281bad02eed03b24da;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2d398f719605f1f99786e6dc428801158c383f711a8a5c86998e1b0b90ab624d20f069a044c14f251d1b403ebe82d8cf85f659fc88829b7b7d2a99c731bf0d43c5f461d45f0e6af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36eb752db7a312144aa7dbbbfdc89f9e138c2905bc20dfbf6b7c22894ed58fe16eac46be69beb8c8a38b930d4ea28d9a2ad896484c56a594b747c46fdf2fce0d3a4c7b6a34c728a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c9dfad87bc554d4867775ba0e02e35a28c9daf6d44a89da31856a827ee20a8c63a0c4d36343fe59aea8d55824c2169736015577e4fcfe595760f6c0d5de10bb71064f1d015df300;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9352b3b9722557df02e0c384581b4960965200c399efbb2c0db3a48acad8e01eddfb4ba5c92340404b692875c182225cd632b5f613e9a9efa78adae0e65cb73308d7333c03af813;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b675a6e3f17eaa13165025b7bf178a09d77a14230d6c6c448fadfde4db3b9de84995bcc9f477c43f530d4dcf52dda915b4fe4ed8c405e9677059ea73013c70cd16c12991357ed1e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6516c575f11a148884d912af339c03405ce5426bc08945b9b52b26c0a78fbed87e731b1e20777fbbf7987d2879b1691fa25e3f0fd35d5f52aa2a3c9b8bd2eee438eb10f4eadc9c86;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h294b2706e903e99d6fe2238a9c3255bea53552de003a4c7f5b69a31810f6a19357e20b3e3422c91a10299764ab0e156108b3502e58c9bc7adf8f2a4a4ab9ecc0b03b46ede4367c6b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f2be25a475a184b0a56a28ff59e4c77de5771c3323047a3266035ae3768ddd386e603ffc5b881e661b0e1e30f1e5ddeb3e4eeec7790a0ca112fc2cf5a5a663ed2734a8a82ddec84;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had3c424348540892e780648cbc6321a95e8f7016a6f54fd703dca516391e17f2db99aac10ce4c9db94bfea1a89aaf3c5d5b1a3b7610f068ad901e0ca0dd44c2ae9fed1cee5e99494;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26d9868f4c6a8cc50364204e9b023ad2d610d313f02c343c3b4b9b9a33002f1da0c262cd5e907ba7a090f9821fb445de8d81c1a0edb4d409d4f82bf1bdf12bb54171502e0982504b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5bf176d191908b792e672693d9b6faccfb6f7d55f7108be585787299e61af7c4be04ac4b9487d670f4382b6a8ef7b70bfd38a8cd5de0650457a023a3b81e26b98576015bd3cac15;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h28252d9c9154bc856455b021a046624bbae1ca35a20b58f657fff4df7162a86b530d1d4a829a6db06f4a9d22fde77899a391e393f937017bd285fa9548ddf020887267b01130c97b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13f46195882d7f4ad765ecc4b9bb6936cc6483a31204e71e72ad20a2a3df946be0a73635b93b4fb16021389b7d7e8dabf84c8c543759b6b437c9abab41723380d0cd349de006cb61;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4ed02230c719a7e3813157f4868b522a03e1ae6159f3bba38dc2a3413c50e7d3b62d9e50b5fc6768494d5953177fba2597976bb8487a7b09fc2acf5e6f0df9b7e5912ce4c9cc82c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79fac7bcc4a929cf82e1e30f63ed09579ce4f49a9f62d44135fc692d72f420d4b8acf01a3a9cd8a114bbd1729876e15eee49a3c6de89c3acb14e211b862f8c415a4cab10e4326eb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb950f9c15951181386d89c947579a7ee4390fee7ad14b67f74929f267d82d61ed51b0328f3784b40921feb3bb531deb42fe648f38318537acf7310c01ab2b06ce23efc158b0beb87;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9544b007fe8421ad8a48ca4e895359cf9fc74f3caf2903b898992186d81a74277cc28246e717c70dca60fe9566ea1372b0af2d9fedcba017eda2ffa300c9bd2067608a3a62e13e25;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58c794ffd7113e1b5a6b158fe63f685025adad9226181f5d3b7b2aecc2edb9b184d0f94d69996fdd903371cd42d2a2a00602f08e3f591a329c42cd7e005076598913800e080bbfd3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1bb81b830324efee199ac2e3cbc1104327547357a62624043cbc29df6f7611980657fb16b8c0d374c6878c54b74467fc4f9c863758083f6ac9b2119e42f6c7da32cce486f170783;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6729ba1e137a58efd18d4f3f587524acd4ee916ac2a0377f5d84a902e0253c08c86916b21a446aa5b13822403b3763ba1fbd713ad81948244e8547f94b4110d100e0d8cddb5acd9b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5388bbdf342a7158287e564c9f0ab1d6bd29bea2c9bb01d6cfd60856c1b9d66cf4082e6b211e1042aacf7bb347af8f9f41916187eca9c655fde17af252cee4b4b5236d222411f77;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h371a82dd529ee0d36120b22a15b5b8d5aea64422c6bceab6a240543ad890ce14ee25569d2a49135689dacd5768214fa1685d7f49af273153cb04b561f5b8b96ad147fa1b4f2d8279;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f09f4e602ce6805ac7979ad98b0fde23dffa2cd7724a0c40248c915f61a8bd4680657a688b14bdfbc4abd0d901ca1f1c064d33337ef7363019f4d1c8eb957afea55370b1a781bfe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36fd42833fbff5d95ed3675858be641c3c95e9ab4bd393eaf1cf226d2841b578ff549dbf0be0248cc1fea0819d9f00b2bd1b3f93afd808abb163fd12e841c24ef3cb25739a867069;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd99e76489154b0bb296abecbf9a728ad996ebe46f61ecde1e557bf439a11c97368c7d479bf6632d2660b42deaca6a3ad1e98b728c1cbcd396fd2b1e43ee6d9536aef15cdd6214ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecb509a2bd64d11ddc332cff9d18c86a24b4da46c413e1081fd0165302261679aa36b9d3c236f8543f40c6aba0d2ee0ba8400008eeb5c8ed9cb265b6df5b604c99160d178a7b251b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca311a42416734dc07ec393407fa0247178668686cebdbe561a143677c059145e4c0556ce79db05008ec354b4ed049a743b542419147678808a3b03b083df8edc6ccccaa35223a6c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21628420b15ae67278e49694784fe0b50f6f91a536afa579b7ec88d3061334ffe4d7c3ae23dc52a3803593c0638f823e9580afc4b91ad02b20e9fcc26d816e2fb8ddf39b9752b74c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf71dd74dc292851a98dff7c2445e0a01e18240c569a9b40239f05499b824b057a61d7b0f85c420a500ef89ac223a4b261554214cecc1024fcc4451ddfd0e6f1ee54037c437cf9665;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a56e9083a847495a9c6e01f35cdd2c8dc3eebec081084ebbd9f36fd486dc930427cabc9803b0653bac96db2519b7bfd0dc44a5867bdc74c1ac87bfc64194a0051e91fa5f0d8b73;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf2c21a553fb92b0619bea6efbe949458db51cd4087d94e2a8519dc7906210d02c01315114bb72b039e72be476428dd73c3aa11c3932eebf56505998c452fb2e3f0e04fadf50a60a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b79d29279044c5b01b0bbc466623cf0caf52ca5abf857d0c5260e05ab0c52d46a2d3d5cbec9f209897945e6f965f8a7c59b288b9b13178b33cb2e45e451f89a6928bf9d2ddc5aa5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3c513456be521dbf792f71c0cd8fcdd8682f9952cdcf28fde34062f442e80d1bab2a1dcc73f02f460aba35cbeaa69d530cc50fe2d1d66b2a296e86d5852d7710a278410d3030ed1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h689ccba7c1cf299703558ef29836828ad30bb1c397d20eab1e3bc2becf810abe4120f77263979164c531c0b9584cdb05c5b77342d67eb735f255e7b1afa3f44bcf4b551050f7383e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60c21a071898bb2156d71a186752b1a864c17804cfe083edd045405da4f4540deca3bdebb515a0e86fc8cad1d5a8eee669bd4b5a613897f43e8256f0bc9e4f3a83ca2c088ed747ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23eca55f249d75709d35802b60b7d2e813d16885a151f182341a81277fdf8c4e1a8b48bf4ee843266c447bd30d006df9a4a3f81f4d5cdb01fa3892089ef257c3274c426e77271cbd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4457896e19535709d494f9de44f80e58eff1687c10f8fcc53530f59b9004375e79ccc6986654439aa83bd3f0b9930f86d7d037f6ac1fc67c5ddaf17b166553cc18eb448cf1b99634;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd841c33fc88e34a53ad25bd4f18d0701db7c6214fc51f61d8abe626658a76934d4cf2b4cf5104cb81471bf5686ec310a546169b240ae32dc7f5bfd575a9fff6b6cba748a24e9ce35;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8d6b730f7e1ae723a078a3103624adeab9d59fc10a8c0bd440e5b197d61cf437cb55eb144092f2f36b03a835a0676c75df8915348c6c83cfce2bd0cf0e50a8b308ec80067185e3d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38f4353cf6e0ef17eb9c0f374b29c36c9e86d59c37a3b58346043624eb90f775bdf0dcf35b91c650fc06f69d01660b3ef6fb9e6e282ac1026884e2d26726eed95567ee7636f609da;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h876309bc74188b51c1939aa8e6848cae1de647842b8f5bb9848477994b84c452503292f58bf5cb7404aadfbee8757f81775012639fe22025d90faa631a4757852848f58bffd309e4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73986a034d0a8112d73a13ecf4a0cbb672b2032a9ab679dc86072d7daceb5d2e85a464ed8eae59c63c4882c0a9802a855b280581f84c117ccaa83032c6db40edbafb253069001385;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h873a190ef716a979fa3b17fbf99a80066032ebd1736bcdb10503d4c0d99945f21d1e6d13fee1a4b75928d031111f669934d72b56675683a6c966478df5c5e74807ac882a89f08aab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c1f9a4ea423caedce9fb1efb6449a62e499e83bf3a02cb8f50f534417c1e4c31f75ee35fa6097531a0ccbcb5d3e24bd6ca076288d8f26b5bbb72d348f018c6060a9a6bc0d054087;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88260d926dad858cd4fa2654ebfb018696686260ce10fb3057f704590076fbac015811ccf62b01ae3625a4985c47bed578489a81433d50a66bddd2de372075109023527eb1625019;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcba35902af674a2c97802a9ac2e2f09116409e09afde13b544e487b365c30712ffba9562899978beee3b24523045a5659e707c2aa118d48b27ae4ee7853e351e98686f353be12b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67549b0719683bf88b7678c0b5ce508edfb605b249f32774899197645c774440558252ee3981604e02491d620e3a18d9bd2824d8313e7a9e89b22e618241c1b03a3d0fc8e0eb298f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haaf09bfb3c3e768e5bce952a8cef33bd7c2b5b92dc6c8d28771b6e8017f2f6b87a324b22f6c6c850a341e333ee274e76ee9296fc88a34fabf098e431f8beaf3ee7dc76d7cbb8297d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83d942e3747db9c79e89bad2b0e3ac4647127f2266432e34b3a59851c88a743d0b45d26163af62d7597a0a364741bc34be4cdbc7869817e3ad2b59f900292a6476aad61b9016de41;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26e61f101a8e3f34302ed641a8d052f93fefd15b5802457db559c461020572435bea1e65aa03a8e52fe8bf2396488cfa9cafa3661683fdb211c0f9a93eeb89700bd4b35dedd42655;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc5c23fe47cdfbbf8b76c2c51bfc9b732bb7638542cf1396d04d36e5c1fe8451efc3810a3d79fc9bc3628a357dc94a5445bfb502f3fd93d31457d5f11522e87729fc439725f0ac33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b9e574bf0ad93b50c5583e47ac193fecdcfb68f60a175ad07827849abbade29f474988c4d78ba4be956173250bace005fc6aff7b65619d743bf5934e00bacfca15cc0e0248edf5e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8581357c6e0e8b7b44af03d2fc7c2ee11d3d340ba48bc4ffea6cbbb9f7796a1b42efebfb763b2fabbb802fc5dc95300b88c7474986853aafc035fa90084afba68373db9b3a83d88f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe9a87777b31ca45cfa5479ff026d8a8b2d724ec00ac09abe06c165086638f9cb149955c0bba764854a066ef6fc2594e3c19aee78047019cc55c7f2ec28f6d73c304c16924ec7c26;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1bce15f1924d4567decf2ab8691a694fb28f48d847412a59a0940a658e7d502ad084fbb5bf7fffaea55614b41b582950ae3fcbf36a7247800ba6ddcff5cddbf3d94a6954e3935b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h679d23b8b84ad548d3ea80727e41c1f4fd23eca381f5bb7a392ca9c829119d5a7933672fc9cf9dfa037af9ffb2cf731580a371e648f018519f03dba6d40334a7be6b30936586c750;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23cacb330e9a4d8cc0631bf215f8404896f1d04507eb0e541975a67651a80061b670cf3078c2219f6be582fc2b62e955d527cdd0415dc94ac43b4512341e2921c6acd6e1d48bf03;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6fbd6b54ea82d4773b729b0ef33a6a445b46f42e240439c8bd04aee670a373655d00cb8510e93e73e814b63e499a60a356e86a09a959ee0c0e72331a4e81143d13f3fb157674643a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he044fb1f4f706057bc88261489e3d836df6f2673384c768f407b0372cc19e9bfdae23de0c39eb40821800187562a345fef271719004e963d64f1fea395b9c134cab850ebc5e7d931;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5327d7534f885374dc58dae7a69e98a9bb2376e82f29dbdbaadf35cc7c57792a1d41cf335b3c26f607854fbaf9d7f6cc951f16ac4ea2003df9dc84d22b24860496f4b7dabd627d6c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h337b35c4908886e2d7fe994a45dafae2fafe157b76f7a49e155de9c9e510bb1115f0fbf80edd28bd7710cb72148a26fd99e33a364dfc7aa1df5a12949adb66c8e2a4fa1053b3b832;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59066129cc23ade1315433c486abc518f2b0c025e4952397807219fc8ae89e6a56a5dfbdf5d64ad1de195966805308eff5003c6824dd7b8c7e31d0d911068376620b8147f4c5e894;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6aba8fc26447b3471468672cd95350f394b79bfced24a61b8dad78aa74bb6e5a2f234e79f69a8368e39a46702704695ff8593ff36d0a642a0bc255d39fc8c1a764dd502e7f7fdb4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7545ca2edc9b18fb59d65f0e177af2d7fdfb66241d1baf1e03f78c29a5451ad76a63727883273312c4c3a63bd242fe2b910d9cd38e7e36dcc78a3c9a580c53890052ad552c7e3b81;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb285903a5da305caf8dd5ea0f20ee02ce0a7143a9650b87e473ec1bfc6280fc0bff3e75c33f98611c8cafacf59754312bb380e948a00236baa2127c3dff7dcd6afc8e98722984723;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57ad01f4b717da6bed6d902a2e04128f6ec5f403d50a93f758217f02f05c9994eb25b55eca3e40a50637fd6bcb507f63259e3877772d4f7de0b8b5f542bce1fd0a1b3790909e06aa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0b3172efc24197d5998744b387a6871c3aaf9b8c67f6383c1e2ae48c7a496c888f1b781beda29856079a6da7cddd79754b8725e80e15a2a64104f4482bed666843fdcd89894444;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35175b219393873f422121754541b642147725ef1b2be8a1febd91dbdbbe40cb81bcebbb8ef44a3a0a7c376142a61a1d93c84cc7c402dd14c00296d024ed247c89f1ab93a52ff43b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e26c89557c32bbdff8350f7cec383ae27dc70a95a4a767095727492b1318738e8b2368c4088163f8da94079a17b76bc88336522da20362ca416bbcfdfc0ecdd8e1f138918d1d4b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a3b1f94fbebad529d77a929722ec7a5bc6d7fc5424d961ba08ff9a29631f3aaf221231f5e3756e87d1668d68625f72c7c01c9ecf2933765993c347ce02120e32d9434079854ac90;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0d651f74c4d0c6c9439f68b8556b881c623030f0f5f6bde7cfd1faa49536f261dbfc7448d65ad7e190e70da6d0288b72e1d596ed6f92a51ec4ac4b3f555594c48969f573f4df85c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19a06be5e81b69b7c7213183e981ed03ab963d9e73004e8428d246ad398b95091611395c0cd978685b060c95900e88a8f4a66f8654ba17680a7d30852ce82244cd82e98351006d78;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbefa47084b61dc9ed4e7479e52502adf4a9d8d7ed4a8cd76daf697919e33726605faff07c36b4da5877e0e4171d5bb140a9f94b049dd782ab8d8c60b121019724667b6306dde987;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h347afa9dbdabc5234743cde48ecf0c54167302e4ef61b42539870218ecd016345b9559bb09a675a59851374ff041481264b8c7a846a507e2d46a18aea3fd9c54da85c08e35131b95;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1381dc25b4680dd5bdbe2d723354d4a070f6493aec5d161ce16591243d4d52b8c843a7c799d19a8d48254ed9fbe0c8696247439f99a54a04ea91fc0c406e8982bf31c10cd5c73470;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1be46e6469915f50bd69fbd1e447c6fde71a0ad66705b9ab34cf34b7d10852263eb28496b8fb66dab68c3bbe42b33fcd19facf1fda19f2d6250f70133dcbc28b64ffdc7557c5a84b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e7a46239a7fdf52d4b0b3aeef1fa55d700f8a23ee9b52eaca1675ce9cc55fbca1f6f5f7e3ea00a61d4041d55a93f7dbdaaf499d7fcd2794e6ee36bc0a8d28ff41491731a51b02e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cc772edcffa5ffa87f96b0e3075737f9945dc3142272073fbd30d750ff308f9c486e71e7d8b7e9092791b00a1f3e1c4aaf08c08e95f3a6cfcdfafa82c857c3de8d516b8bc1bc2a0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1f1151600f6f8ef49b74ecb8d2d46640571954bc4728140ba93b3374de721b168c670251e95fbd843ac6885d0e01ffac8d02b013f773f6ca3b9df37eea1fe444a548dca3b991d14;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d0e706864784b2b5d5d966dca594e662de1e1bd3a771a71ed40423196a6669402628447f1e9ac129020a1a703b13f4d72e1f4d0c981ef2509370a7c4ff0da38a66ad2d000b121c9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82c755cf622f619b6f49f84876b1c19604ed67f22a7639cbd3446624602c6c7431fbc690e0c41163f3b8fa0dee14f4844bb86c43e8d8357366b0c453dd8b9bbd984b8d3af27edda1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c50e6a662e7f06361e2db55f86466286687d95fd21c6bb54e1244fdc3e898821202507a61f54cc63f1b48cbbd5c16b93c3ae49fdb0e545f23be73aaf900548b9ecc91857ee1131d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd76b2db0df03e15d1f02a999435a7c3cf849a42ce15ec7465d8c78d6755dba9c9f817076285145111994b7964d5c5f8600a19cd381c849d32cd3535bafe504234491a3148f34d62;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he64d30a7338609da000314d3e66ebca90a37d5907b7c0fe5d647407398c0f9e38220beb9b1b9898f5d7bf45075e2570478392526b3d940c0de346043565dca1456dd1c484d7d2a43;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he13c1a78934bf154ca26ee4cd34ccc6ee6af7eb9a50368bfc07babca43e7aeafd9d4da898741aa33a5005051f0cf18e98abcf032a5ee6c4ceaeb0af36ef4d27904b51cc6195c7b48;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59bc10f064fd6ce355637c19c547769aba9e861c514533f817b259c0fce93d6694fd0fffbab68f846b093ee6c97513a1684f4b2e0f86fb1e717e77ec6a236dfda8189a09d73fec73;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h452cc469976183d80d5cfc95a6e8f70330a2c258f7f3af096b3f1b44b8a065f2d5b8eaedeece6e4e9cb6625857e8e6a0e2ac5233e29ddbe8403f617fa0285ba9026ba40dfd112d76;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8991a6a973ece2d764c26ec214555f8818d8b4d7a7f7bb820617b641098e4b1845ef2a3891a44772740a25e4e54242724ec5286a726cac744e616f8fa58c891892bb49b8eda1c0a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7a0e9aac7fd86a4a9b3c55303285d9ff208040705cf34d124133bfa72bab16b5ac12935f3154982e93f92fdd6dc60a69e2a12911736acae979d01118f2348493f6e43e2332ee1a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd34e7a626bf9e6935faff98e24fbb8124def82fa6dce821f857f32210afde58911b47bb6d67eeb7b9f5cb89cedc6510be3947c33ec863b347a4d7e3a8b360be5ce721366e4e6b2d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5fafcbb9d41f720a739791d40be877843b3b389b3eeacce99eae0e9056ee48dcb26b7e3e366e66cb24591120ae5ff9285f13d763cb0dc4d7273eaeebd3da8a56d382eeac1c8b935;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfff23c8ccc7356379d6f56a0755f25e9b0f5a10af9e6eafb76b976a32f42fb1915693b1f93c440945a0630bc835c6b4d0d9bcc624c66af94948b9f0e14c2282e958715c6f919a066;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c1dcadbe3f04503a700bfb7c045bd68f9b50cb32eedc523077a4833b5391e338a1e43e4acc363d70496d2bba5346dd41188c68e08f30e21e974172fd7e4bd7260729855c8bc9b00;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6e226440484456c0ebe74e98b0028d3653216c53a6d669c0afc9b545092b0520044e5e0a841c53fce7c12f098628154969c60684a1b270badd9cd06ebf36d8a108883834457805f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65374eecc43ee29ca283a8ae8279b20f4df8da3744312dd3a3924412aa864f6ef15975b10f438f231e28e374a87e1b3a66b7ce5a036130be6c6fb96f55f8335174619aad2485dafa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5d7f0db18c04eba841f8e9e80b35032d9979344b2a5a20d3d061a390e5bf2d16fbf8854954f391b6f6e241d28896517f04cc886c7dd6dd40d34ab9d3153fde6a84d4ea6dcd0a13b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedca5c1f44a6bdf45ac0bdb5ab245e05318974ec02b3160d8ddb11ce22205116c68cdbdc848437ffab4906ec8262eb87ee8e8ada5ceddacb9144f0b0042ee2b94c6ca93f1491204a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d048274fd0a94b0bb2d84bc05b4679f6f07cf135c9f5e6661b33f0dad740048f7a4de2f1a7435687c9867481ba10aa16338dad11c26f0c0769367226a5413dc27665138477abee5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1683c6938ebeb99a5cf738bb25b5aa9dcf3985f8b9a01c9f99915ea203edd82439027a13e8b0d71a72be03529d45e847d58fbe4da2e7ec217a91c286fb70e4d3b917a758ac2c5d92;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe8a0af809595f7804e2dfb06fb7543612cc2ca8850276cdccdeb37e1ceda3216cc98c3beaf9e711d1ad446d2385e311e09dece9cf2275a57b7bffe46fc98b9b9acd3849c9061baf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35eca77bd4a30d12c308c24ca9df96677d2555650074a0a4eb262becb7b8d56139b7233b10f342c12a113633889954453630b9650884f21c1275783be3347ff2982bb01f1c2207a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2efb12950ba913b0ebcd0ae97965a9797e417586e4455ae1eb6ae01763a3c4025a17207a9620e0fab2ff9e2593d7453bbf29487666d1a0b75102ddb14900e17cf3493ca56e58976;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h949d89edf4ed2377bc91a5abcf532e90d9d3210d860871d4120208a5b5ff969432d3e122b1bd8cb6d0f954186d535c033ae1fe8f50e6837f745d7b22f18ac4e5c7dbb30c8d594540;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73bf99d889ba8bd3e03f799c675c82daf4245dde98e984ae1079e4a485225842b6bb6293cd416c07c59b9b365681567f786c678c73477e983b3a492d01dda5b51fe409b43701f4a3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d85b168e8cebfdd53aa30aec72b6a6ab7f99a194451cf342e648685ff512d8176cba704796cc8a8e011cbd84e47bddec44d0a6bf2e44d85e3504d7b79a37e8978253f19db7a6f80;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6addc7fbb2860e9e4921d154074e1d85abbda677cde4d42cc6c2aedc76d9d791a740bc75132de6b964d1c76ad4273e3920dee79cd10cfa155e5fc6dda084517c2aed42a8ac8221c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0e541c1288293205e690240cb2b0ad09a350e6b27d03ffc1fe0eb07273feec88800e450bc91afe8170317d923836fadae2066ca19cd945e678610a6a2d20d9d61306e4e5b34508e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h665f011b1408ba6a5b946113e5599fe90d95f3140047bc881771b3ac4f58d75fa9aac5005c92556b8a6a1938194b3ed736d5c28dcf831f9dee2a3cab21c39bea5c3a65d012fe8a0a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he70c6544f85ed7ea4a9c5c140fc1859693a1297ee6fea7d6b2f80af6c59eed720260ebcddd2b1e6f2aa285d73bde0409233f30dc70ad837651f98facd16fe653d5c3aa494b0b854f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha59100ea14cdc8d359d4e1eb42a1828d71a535ac7d21985fdfddf48631f85dd3152ef57b5ee182d91b6489f1427f1346797fdde2cd0f362690dd5b853ce56e6779d0d5aa54ca9b73;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e66cb26f50c4c6e79c45fbf970bce6cab189e7d394adaea0131d346cae26e48486e6faacb346db73a550edc0b145887e0eabb6a97bd41efae272640d2e75dd4a25ba70fc0b6e76d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ba8bdd23dab5321f79ac676234c3d0de3f23af372ca41d58ccb08fb5d7af2f509358f762dafe93f874bb0cec2a377b3ba3301ad6155179e636b0f7e5db62b0e17b07d6c7eb53b1a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1118b98924e2e434824881da93d8e2c1fd8e7646b620dbeee231d1c35cb9d6665ff38720c9286c8a4451b3aa6ef11dd9a17b5c4f1f254537a048b7f5be69820e75ba4e2dabd8b4e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f1549587cea20a8b0ec15167a54b73d46c1d2fbfbc805864ec30bcd2b5d09ac083ac1ad2f752d76507c32b578b289bb68db173654b37a63ce55a23d882fb15d48cd0b7387be48a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab67af0ffd4d1aa7b489cf6f645792ecbab9e863314cd6ac7b6624791d7ee662b2bf97616340fa7064c1f335b3b564f38b429fde342d9a5d6f4b7b330cf36edd4cb327ac5c328096;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h546739b0cc72928e4fd004c196692a6d696f8e2c70a2023051b0cf27cd56c3c85788b052f14c27826c2a4eafb676b70b761e83cbc12ea75d49d4bc516ab2212df6fd71c59f4a7114;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92f0a8c9c179d33f00db4825c280d69b470ac92158fb917f2d08420689f08b5c2e70330c52af872b86c80dded5fa02604ef07fab58013b95eb615d0cae230085ed9afbaa99a7b3b2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c83437c9b46cb4936e4bffe8853882742d23580a4ba199326c724bbabaa8a3f1d7864987c1c9c47729c0ef20783493df9931b0b9479f27a84ad91392378ad11af2a3608c7e7860a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d28ade1acc514512b3a80b40a39149a0e0b8c6c769c6e9ae2bc660bbc5275f0b530271fef6ddb6d1de1d4d83d2e012906805d090112063611c75b0b0ce260dda85d987dacaedbdf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab0b028bec95133e96a80057f9f71dcd1ec55496c76eea3e003e144bea14d9c132e1cbd6c6edf7a6e887bc43c7f0bfbdaec23644c56200e9de600610b6438bc008c64d544aab2f49;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1099b4a6f8f58bb2b4d097cbb460b0c444e9f175e56b073c31149942da131d87d901bfbd37b5033a2e6b7e4b858962b9aea2f09ff62609b9598641768c97f5e94b3c011e37508fa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94d15637fea72881063f66b579a74fe6c6f9bb3f8a80965a4b2586c7fd0ec17efd9b99d827044274f2d8c448d643b08ad7303ed6d0df4920f7bd269b95346b4825e6dd299ca5e39c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc435bb03f28cdf268126f5c13f8e9eb34520e4b7dfa18ea2b09c41fa47aed388f1bb6877649cfc83c4968c640558402b4dab6e08da295e59db67b2e3f4c0d9185d40f98158a5f1ac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8bc053e8b41b2ccb3a2903162d0647c73cb90022f444135aa626a8a3eec1bb14d6105f7751908cfa4cf94b7feed011363fe19bb1faa2026a5d204e4999c9c7643ebf8eb6800a8a8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96ac1f57d51de9cf4b5f694732091c8dc458e32a506be3d3908a87ada1b90eb204dbb0d210ddbdfd9f1fb6f6bcbf8a379d3395ed708cfce244296676c1a31d78192c08188c7495a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d12e32913c9d56f7b8bd73c9f465e8fbb3749ae1860afa748497d32c254c5be1795cdd8db48c12c90bbafbcbdaf8dcbc3f10e6b89cef670425ef4888a9ce20b167ef084a193bc45;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d3e57b876887194e0c10c1cf028b5ac40def96eb8e920240e03e61dac6b2343f5ce95d3b0b2ccce50e4f689f290036b8ecad430736bb1b411edc908d2fac722a372a63835206b18;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6b5195df4972886173abf30644bdc0fff24324d55b953ad513afc96244ac56ce6f1cbdd430eb5a61dd91ebdb627313936757866f349d531e7da261d58ee033c94b0a42cdeb3694e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5742ffd7daa14cb65253b2f5fae91d8cbebe8e6e593336a39c9944f91bb582b4180becc1e8bcfaf993ab70492b266014792123299f750d865b78a8d27e0c549de074a7309ff95b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h779c3e9ae7c47ff16125b3538680fa645bb5a6f031d41e603f075ced5db138119acc127ea550bdc191d6f458493d40975b0982376494fc4b15357a4689d01de02f174e04da2309bc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55fd68f4e49f36f4d341297e27a56125a29e90463f5639c84ec1793afffba3c932117e91b7341b5387eefb3229c88300f4d969e89e747b833afe5fab8195d2aa598f57da9581e3ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc17b5fe81395643aeabf22508ebcb5545c416c083081ed44594182d8936b2fbd31994e806c590079a173465672768bb749a4c65691a6cd0a930180522a7d8fff3a23721f85e7589a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h708d8f243c547d18e266f5eda7636464fadfd9fd73da4fdc8d95ec00ac1a9e1d2b160815d1d5220dc9f2d8e7141226d116e04c89d5795261196ab1cb632d415606a74a6ad50cce53;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35f44b4958d25ca58e3f645ce0595b62b6a4baeb8a623b53f3920702fa281d50561ea158e523a363cb6696954dc75e4e949825e01d9418c9fbd60b84d5fd91fc067f9bd2f1281927;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2a6764218f7d7c00fd6074e19915089fc0b2d0c3825f9ab00c12b46b3a1f1e5e0ad1009160f25539c0d6712bac1fe70cf3366d24cfd42b5660098679761d5947859a2b1e775c1c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf1565a65c9e203b887c9c1f808bfb7270bad086df8a3fcec727486adf86a0b3d5d86912ab3d6c687aa23314c3ddca9c2556ef59178a9772a1dfafd8bea3dc9507d455896b05daa9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h953b09080510f50f080007c169c54d632c81709b4888b5c8c419d99975b3532e48ef3f3bbb2fd471be842dc4c65dc40984894e6d2ec0f954d3524efab5d87d801d2b5aa9ab2bb3dc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ef204c8a755951510830e537528099f2d9ce75608703f712715c09cb654ea019fbcebe59ffa26717fca0d1fd47414039d09db2fd70350c0b8d16495d6454e9a9b5737bcad8f364;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85c3ed01f70d7d02dfca0d073b94d31c80e22808a2144e03a057d5bd6deb45b337fdaef486ad73bceed8a1b72d1a94901fb88e5dfbd195002f0e471577c84d1cfccc21cc49a2fe8f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h699b7f72893bd2617d17dfcad49a7383c34ba42f65043d9f8a118eb397bf038d0c647302879d90837626c0766ed2a3714f9d1ba4dbcac21042c5e3387f38fb1b106cc9c27e985a67;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf50d71c5f53c489254fd29f0200b93e42a9717bd63a48dee788a322bf3aa6fd2fc0fc424c9d884c280e9ac615dcccfec97b5a8af86b0c0dbf040dba0cd6cedb484f0cb46b6b4b300;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7963fce02cdce02d1d81da8ea7b09b8de472fa31acef28479d8a11e72e6d8a2b21775827ec980f39361908acf3c62cc19cb81bee1c606e289343777dae8a7d951d4fcd2e1c24102b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h538d72f503e3af3599420732955ec2808dae3a27c6d58c5de0d13a78c28df86f37a501cdcec441891dc48effc62c5199765327b284e2ca4cba7c28d6e7c8a5b43f1989458934ad44;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haeb2c98161767f177f817809e633b4d584cd5f48abd7b8662c714e942ef7b9326832645bc27580ace9a3b5f5d31686b80112ff62e11ab50cef2e6018f84997a9d42bb2aeef294b26;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h950f31537f7ebfc5b2e5ab4230d0ef7727837bec48138174a16e9fec6cd07b27141b4fe29ff603d810d289b87e1bfd6c9244f3c7c5a6bc64cdcd47b0aecafa591c5fa9083552cb01;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e8f280e04606519f1dda6110b8d2ddcc51cb075e1d67fc8bd273347703e8871f600b29a003139b8d067fceee961a77fb0ce081f01ee9e6fa3a12e2eed9240ba06c997574e2a1e92;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h626dc7432eeb50a312d13a687e9e640f39d90a9c4f4cf3482b8a0a89c53f8e4963496b3f9c1f9848b73e28a1b94816f2fd1a7611515c9e3ba7cd582c538b7201eba063d4e0ec18eb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7e1c1de5643c5a3472796b26b09aadd0263ea30fb7d78dc1155e49dcfca257f91f5b52329253e07b0ab626b15c68406babbe400d5c5f4a24c6c3f4a33caff294e3815e857b9635;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46a11c4581f00c756d52c4903b1a53058418ee6d3459d67df16b049c000328124b65e50581ddc45190798ef3b177c2730766f1c894c15b85e64f212eafef3cfcba63e53e18be120d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb88e4b5dbd2588b019b58d3965aefc0204c48451adb66215f1f6c5f449a6f6e390a0f200ceae3bdcc3a0224bf7af72e10b09b04152440c6c87e244be61d737bb717a566705b02e87;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f3f0b64efc953992f73d40c46145ff85a5db2c84b8024ce5f5ef9b1dfda19c8053d13aeb05a686dd49fc86338fc368045167369c71adaf92cc203a0fae4975f8192a4fa840efc5e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca28bbf586b4a83be4f1e21763a5e8a430954b9bf360c2a17c1be6b1583be8495a9c1400cdeb2de08c4dcc8137575cfbde56c696e6a0209df55d7da1fd0a34a1eba35fa17226c658;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ffa9683e4c8dc49f579e397d00877b7e3c99613606952123cc74b5ded9e99b03db705cf7d3090276222f68356c067e6dff26ace57275a4e0e11e89a8fd462ab3c2d7b7600787a76;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h672f7230e667cffed0c46c1f321f7438df73ef2aaff23907358b45c6a49f2ca6171ced535fde1b0b6ed1f7aafb213c82fc9094163668abed6433c5004ea5bf0ab88610c50a4164ca;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8568f67b17f3c8a088d3a604b1ecae68e4d915d45d6cec97dc207cdfc4b4ffd48e9c810a3d17fb1b1cf349f1248d34c8c9e8932642997b50000e5cabbb23896cd1fefd6e50717a5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7143a5853c7fec85f3c37380fcdb29ae095f2b1552a68fefb7649fe204a33b03079e9ab54cc29ee18cd3b8bd2aa26d2ea3bdc6cfed43a3daff9858b17aa6f0392384a865acc1327e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b0bb40bdffff74d6469f350db16e99bb17cbffb0df2597812495aaf7b35202112f150306a1c87db46b34e1ef7b7bdfa147653216eea4a5edc0e15b729f8571c997912f17582888f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h978b799497e73c2d473531859898609fb342869925f3c2894a03286c1b9f143396bc0fcad105313b09aa1d975a6637c5bf09dd21638169437e92876752ad4134067ba27805468806;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3d2ea542f380ec37e95bad6b0018d83baeb25f7be45c0083d285336f626e42e85febbcb856a656e7c74fc2c4187fb28c157c09535fc234b1048a77dd8eff0af542a6c9d42aa7808;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6dd755eb8826c2cbb67a37570748cbecb227a9a32bcce1c5cbcd884ee277095af167c775bd8093e7d6a525d55105b74a8dfa8b05487ba299e401203c7940154d1cfaf0eb14ac298e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87e85654ce4c7d3d671ec777dd116126a0c29053aacbe92428e914ad10ee51ada0b067d0f212427901149e99aebab8038eda0da05cb8c8019f9839b320d1ccc378f5a90ab85b9928;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36c275ae1ab59edd8796ee18fe338115a7a124702fb2d13b36178272a6567b5178a1a7d8124e4cf6e7f444f3a01b3d87d080daecf3c102510c7d37414c6793d3dcbc30ef048f13a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b1b87fe6b492b1d6a268091d98d99644bc376fc9b0f7ce320f14c280cc2a54821ea64dc6e77daf4592fbbd49fd0d4af4199d4d788f25517d6b54c0ca55e909a0f35f93fca5d379a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h546eb96dfac265780f382c084651e83f34fa676ac12568769c542a2a83f15d5f4d8ca094d0b78b94e53f2a76f3bc8c860d84400e6ab170393ee3be42d45fb7fc417cc3d8c7616c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a3b750de6a4997670f9e0ce4699b2660b95ca34ad1e61239835557b1a53f2ed6a8a6125e9204c5a9c1afd7e07123cf72bcd823068442e80c3652dbef553c95a5070b627a3716750;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e4a729bb055c4030b04fc2989058e05ae5f6e38c821344543f34d272f0eb35ef323b765bb81b076a971887a77e6779be445c8c9ddd4582f60ec02628f5e5dbdb7ccbba2b00308f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73cadd47ac734cb08e50622f9116c52b27173411c3e809920d2d5b5da4b678ed3962fd3098818f99f0d9da8f30d153a9ddb8775269ef860a7aedba4184db4c9b23da77bd28930b4d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92b21dde6f56d924bc58a374427fbbbb786032b6e04833ef0f2068a1ab07810f32bd0791ae0b514d9715073af82e7b0c7828dd46418084618a1bfa09873a3672f1bd97faf3779aba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20f3a83566ca6a947a1ac41b22789e368f062524864a9a7c449f3cb8b4a969d66a873e6d75d17c7ee44636b8b3a50339131cdf52ba4c0c21e25c503e92030fc12986e20ed050a8f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb384bef69fc36c6cffe730e13a81f1549d727efa2582c604281b07de57cf7eaf290ff25ba05ed3b17e0ef77cbe70cae17de48d42e2296bb4ad3d872e0273442a44ecd2f08397d32e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a4a93417b5bf5c3fc7b24e2434bc500aea6169775b0ad1215f9a797fbe7f0f9c5f97d7e35d840deb24477cd7b2d3eacc68ee150d2db04dbe999ba280e238beb64bc7fb529b6fa6f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c5e72be0566c50a969b3bf88a8fa6cf7d3617c0f972f0cb2ee60d7b7b634dad850f2d6c7eff91a7a637dcb84296406893e0080ef2a2a3a3dc3688fe9a3d1e742e3c178ac06c2565;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d09b94f2f8465402a2f706602040be23ab5a67c6ad134c4934b11622bb0642d7d965f0a5ee1830b4994548f27cf5f1fcd7880d37a27dc4bb9afe33c056b8a16027465930b1179a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef3bff46c8bf5fd8c0cc4b4e4d1d64cfd40e04a64221def27cb38c8cbe3259bf3526907d8858b09a1eb165407eecbef7d5e96afb6110413e859fcb6a7f9cd2cf0849555ee57e7f22;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdca43a2272c1a45fd5939a40b86eb6c3d8f4444bbd501116778b4995c313989a4fe26a57a4fe6cefefc9ae4aced1793abe118202b5395896a8d8e55f694f56b6865d252c201b2ae3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54ce88b3063b2f604f949713130ca2e52a1d48684f6191d8221c9fbe5ce9237e027286c2ff6aed948cfaba2f4298fa488f535c45abbf615ae77793729f182ee6c61ae77ba4879221;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecfdc6f9a23f750b3ccd936dcf9809f13fd30325dc08f60d44989ad9ea7388d1304f360bbf5d93f526761bb9ef9037c888381a9fb4f3a78d98fbf6df1fdc516dedf91cc9ff2df89;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc6925aee412404e4176bc048d3821b11b8fb5818a018f5b619f95776f221fac5e23c98102f563a7a9ce76fa989a7ce2946b5ef5e815f5982eb396c6fac9c53284d6a8ff7388087f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c8196a78968616b7ce20ca789edf7353681c49afd067a8184e12e8e5efe282ccfcba0eadfde736c5ea883463685da7e66189f7e51bb80392955003b66d205eda7b06fdc81f46eaf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb73ebf693e25ac30228a79cf1d43c60cd16e6fe4c5e35d196d5196d125ceea585b17f5648301c1c6b9cd8d47b9f70acdabb6b01898bd21436badccd6f1ef231cdfbe864d3ab6b07d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54e355814de78152c5c6431135aff1f748f130ed8755bd69da86f0004dd53358127bf124890f8d5c0a6fb8adf237edc85e772e09e1eae21de4a8b13eacc6343532d0c57b86b038de;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ce30f4feb3ee3aa0fdb6c0e71a8906f2238575e9958b81b6988eeb0c19ef066674c038e755ed31eea3b873316a4a71ac0390fa7f465def974b6969ca5213b61d638b64d47a9eac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1fc9415ac5e0944e12f986a034253433dbfc13b4c62f3a04c00f9e81d371b58ca80bb0021962a2037747d2d1fef65601ed4de67630402800db06139142081dd5066b7dc3eef897d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9305564e76e2c379fb3475e37a72dc692470a8c67bde812446131ba2890ff6c3cf51dc0864ade8b80555762fcd9c7371b1d1547c8cc966c6c39ae622c6a702e154caf7d97c137671;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bb256707be601349a8491a3818d18f9052be8a88fe628aa5284ce4bd53b30b1183275d020391f44b52f4512c9a3552cb499e5ac6538330c5aa62cd1c875a57f6788fdf10b73e946;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86ad719c47debc84e706f7de96ae3c8eb469c3493601bc66add0366a8201d0741005f24b3b71664566180e5817b054b1276ae1d4381d87228888ebf222e34cf3c4c5e39915fab074;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6fceb5d3c8d60d9a6d9f748d12ffc98a37d7d95f2f2e8a6d08ed20fdeceda8cafb5723f26f160dfe3e288d8f354f2971198d297f97356e31d947edd832e9eadd948182666aa4af79;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb577552c2f71c3a06f415b01059564ac206129b5ad47632b87323927793283d0dc8eceef824cf53a5da9f05ee7657818d3de124c4334759b36443a20598b46950e6bb989290a5ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23bffefdd2040f5ac329a71ab587fe5381d33fc1ad5926acdd690e1d695670af8b3bdbebf26098a5c0751a2c323b013d515e3830fa2bbb9d6454b4a0113750ed8c0f725afe0f4d3a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47d1639db246b198cfd83f89d375b0756ad3b78d06095ca51273a495b092912c33ffb1e1e57b510c63d8880c0ad9059b855b082a21099abfcb9f52028f665e7fd9125d48d77669d4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59db5df352a2be8399059606b9eaf8e4785b0a7b8a4fe35ca34748353b99de63054ad4d94943a403124a84170799892d4fb8778cecae96e57a14fa2f2f3e9f0e7b3bd5e37d536d0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf7e2d905ec3e563a43e8492ce8af230ff6a4e4fbcab5e30453a65013f05586ff87293fe6356cb45b45b12ca5fb78b40cea2333bb6246889497cb20cebe8280912c1bdb7f1d92680;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bd6b3d83e3a902837cbb42bc9a205f846784fd66ec6c0c9432d9744181cd0461b2e6ed142be8e3f51a3286c8a1110ef658370af0ece2d77a8b1b38d69bd922585b19d0e1bf9b1d0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb895d384b19a878bead1ed00898d1a223662191ed98718e92f94d596238cb5312d56febe77b934ad70349638a6c0a47b75f2a1de25c3fd10cd05fef04068d7e937745749669b3a7a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4affac5420fb0cd1b4770d4081343b0c4e1c00e03765e0ecae75e1db16b10cd1b716e753aa23979c9ee28bac51bc83f161e228cded670b2a92256e404e47fe5b056451d83dccdc0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61e5ee29356b19b649e46318032a5e670f5952b5b1287eb00416a58db00241eb8365bbd3011bcf418543249a37dec3bceb4663c1d8fc4216402bbe4e5aa69a0a7fad4948537ea1d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbcb169b8b15338b628944e8e20e5ae7827ed619ef72fdae508efd9709cfdc0c8efe9fc6365e20afabe53dd98b28c8438ac4502eab367246ed0a9133509f49af96f7d081bb6c2e22f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8bcdc995aeabf3d986dd2e232fb0112184c54afc53dcd8c627c9e5b7135dc6ad03023b06fc52b11d2ded73c40a24ef7a7b6d03d418f25a0fd020a259fd9a9fe0820e0ae35c1de8c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69c9c0b9aba1b3cd41df5349d822efae814226f75baeae22bdad927587e1f2c87433544d1518531656af2d925713637cd38a3ec1865fb81f2d3c851a2433b612d5d0fbcc7b43ee76;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcfc75b9f4c35e702de47d1fc607bba32b418a9dcf7a100121618b08166f4cf59ba61af81bd4553f073c38e47c057e8c5b4a10ba95c4abec605500701625237ad3704b8362c9d9cbb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c22c61971c73676415a845157f4ec89aabcaafa6a9da77beecf8f6c6967713e9ac3c81820b6729d79a52f11be42a6df3987075007b236568993792ab783b465a3625b910e11e092;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha28eef063d7fa2f786d0e4df9d9f8fbcb7bfcaeb20244ebebdcb0916ca9faf057b417a72fb4a36183f21e0ff3c9035cc210c9d8bcb0cd848ed6c2d77e9610062870e87a5b47f234b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50c6b9c68af3d499f9cbeb1e0bf0611ce4972a4afbbd3a834da542f79247420b385b25d8476a9577fedf1fc7437e75b1b6fb2f5948cf2bcc3a9ae9291a08e5824769b55976e54858;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf37e5a5c0e44e32e68176163c263253cb333c203c556aace2ee532a91962edff8e323ca2d9a4f36967bfa671251b96e70d47412420f80c7106fc16f94d832b1f9be90d8f80293c39;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2eac7a3cfc4bcbddb40533ef0e6a89f684996970fcf0a9134dcdebf59b29bdccd8570fe888c17fac3fd1bbb99ca202f3577e841ea620f44e41a051454fd6f257330c36cf739d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2319d89a1bbf57d3337d0d6de68766de4ef7addf2e74f005265978a0fd6a1ba7359c7f0a8bca36d10ca07cbd4364e90a91b2961da89307bb6b79a590f2ab7c2ec550bc1011073ddb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29c184e326289fdfd224dcc8483481f9297ba2229ffe26e6a1a71f89ff685df31c1e085d44d6294f2ce718cb54ae773f2926f49edee5f0324c4a7cf24d395b43d3ae405712b22798;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29cf0ce0538c0e4545108d4bd462c6df963fc601668ea73c2a891544bf5425e4c4cbda4e9cc80b60dafea3e26dc4eaaffd5b20da50fcd94acbfe13a28c65237cb0ebcccde2dc13ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc8af8b9f5b233c8fa0a21189f377cf2092ae2ba66fbfe998dd8d1cab590072bca1964106df313cec58ae2d96b41e709dda7fb7a950da976c1cdf2e1570ee53af290fa3559def523;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc258fb7053cbd8789a9068b8effb23e0cad237c49dab3f306ddf0023ccbada6dd9c41553443bb8089f2c85a0f77d9cd69fe2aa063980199281ef80e9243d3631faedbe7ed281455;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h39d491ce953852869d8e5ca3eb23c95da3d13e847fb5faa26870b2b1c5de1d52577bbf5713eaae784e92c1f9ffedf4bdd9447246de5b7af4c7b8649e7a1f23f1540f512c20f55035;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha160e9cd0dfafeb15534cf39fd10bb141958c3e4f467a6528cdc21da0af29c18a5dee4ade70e5461f8af618d0ad22463dc89f5a4eaf7521be7903e5b7dea37dae4a99fde2ac3b536;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha55d0d73e4b26adb7a40201bb3426cd5508047d7d785b49bd2afb84f801df301576c9fb70c48fe6aa2c63ae56d6dd1da463de64b4352cd9f8bdb6a7fd888149eef5b23f7b42a498f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdba2661d36c79e71e75215150473917468167ceb38b47c45d7233943504643e4ed8b738c0a101eb995742487e06e53841c9ff8a1dbce6cadea182ee13fe98c9e5b85304c06da3311;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcce32cbeeb5fd4346321c193b2188b3faee334b7ad1253a5749db2b7d4460c3fe093fc988ebcd326354aee7c4bfc325fa5c2aa94f302a9d9a598e0e81d073f91f34272d4a78c3941;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e183634a049a5fc85432e177d82804d15a425d1d29ba64a2064530026be6a5f49b4be5b7e9b7dc863217f813e0a80a0bf6c5d1b7dc89b7b2fdf3ae2ce32641c9876ddd02029239a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h987906b902ed26fe5799e1d51266131dc6377830e30e2a6654e96948fa1c5cfb80e0d186e7dd98d32350a59f8013c79f6f1a4268307282922f53c5330f13577e5fd6b02b7bf55ff2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60d9b8925e3f7306698cdeecfd552045fc117b5c38a0b0ceffbd5730be870d5f3a542fa41aaa3a05ae446443d3b8c58f3f28b04e3ee0398e49f4c91115dd5fb5694c3e93332c600a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31baca198f1d556b957de1495a2d0357f3ad8361693c4217e79f8b991e5b157a5e047d2f180bf07d8545cb06efe7c137d978f1f56c7aa7296cc72320da5dd2c3a413e66f20212675;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c6737e549cb0cc1699447ac4a6f478a42d69253570801a23e12ea6f37223d6e85a93ef5db6f2e89325c4594503af3e292e98568cd2069acff78b7eb5019a114509f0278931e6392;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f4adb1ca77861b0a6a46711d5bdcc7ae7a7e9524ef1de8b004f4cab2a810e4f1e899a7c197083211f2149e52ab8e93e4c7d7ae2ed201486f5e8ed665272e2b72af0fb572db5193a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h650308c54844882e9c56f393abcbaee668e8299e0863e38d660e40214816b68a3462977fb59b3280f756b8a940906219f632c4ac4f9719ddff38081546d15d85aa9070d6141c00d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha67261fa35ed32df3630441069eddb57b385d6c670f971d8c76f8df86c303296e6454ff195dcf987024421ce11a9147b1fa8eb3068b74287308f434367e80e42c1622f0e4e03f5b2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0e011c814180b7793452c27f2ade558ea29d9121ec79669e2c70ba41fc375d162d593680190f09983ea82db1fd6c945b2118dc8d0e88e01eb6ba3f0297998e3a6680f07e8a21e19;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55547b91206bda22a385e98575faf840ae3be797d32b764d5abf68122ce08474bfc7f80cfe1bddc8d0af67a51e7bb7615b88190333a96487e8734bb9c35c11093db6e01105283654;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf84dbd80b0fac823ae43c23edbf0f77edc6a5406b1eb413767919456aedb1c3aa2d7fc2fa87f3b3590f5cb760f2208bb4a315d58f727dfd45beb35ed300ddeaa3f43acb67a78c36;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbdc1c945ca2ce6004eec9b11f21da5c060e26db008bb3caa9b57f93a69ef74eae187fd299fe5ed754b1e8a15ab2e3a16940ffc151acc2a377b77b09290629df092692dac795b1482;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1ab2e7b869b9634b1bf5cc1204833ec71fc33a7084a7b25fe1de4e30816be620290e0724469ddbd5ebeeeaa9555b4a645def3b6e0bbdafb9b25ebd4e5d6ff2930851cd6183caae1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc2628895703a626270bc269b4e47f39439d874fb28dbb002d85853c7be72caeddfe3165a17b3fbe7454129a369d07852d4b99d4100b87f2e2914bfccfcf4fd911f1c96ad3b4d95c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ffb3fd46af458df0d4920a29549166f0eefdd8f4b4631791adddc5d38b76f0cf7d589b7d66b131e78434f96c34f364a5128bea2d0c643d4be6aaaa900b549d8bf2c36e71b14123c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha622f9609af26061a5d449228ac35dd8cb2e50183ee0e0cb681b6db510f1a18a57940dc37e9842c0a9d1807737f1f6c58c2bb70ac9a0af2713465004801bff965440002543e7cf08;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97514d87bc9268deef523e46b4ba27ebdd9635c313e4325f30c212055499f3256a4c7d7bcf6adb6fa8fcda534b4dc6cc11d0a1eabfc348b02d9a5b02cee98bd0950f4e68965339f1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7541a77b9b0b6316e3331a4f034c7975f6c358f4b847fc29afb03a13a10b572b0c7ede42931f78c3a6d79ed865033df5ad56909933e6e8d77f8c809032d3bdc0f50d8bda6134a138;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd98ba9ab7a10fcba4b1927f5a9f234cf638bfbdd70fda28a927d1fe2a108ab7d1b7cb581819ba9f47769edc7672f63b17164219abf6e0ea40ca1216dbe8af96341b516f942375bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c0b8a2787346ad5d5b253dfcb5d138b9cacacf0497ea6a4dbd5616647c7c0321eceb527605211f1184937cc4ada56cda0c94df26baf1c7723e015a9769aaf831a56dba6f9691690;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94c9ee9ffebc3d08ca5386c3c47940a21a2b13b807a2d46b58af9a6481f36f3c8bbe465a4cc8ab4cf961d9b2a311c52987626106ee26a1ff80bff11088cd4980a628b3a5ea37e1f2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2778d966f7d796e13ec0a35bea1ca7cf2c583c6013c425cc6adb6dde5e92754e1538379ed9cc4ba1ccb0f801e092b805c7e8939c3da72dc688b42002ddc51e14c57bcbd920bee7d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12e40a80158ca02f6b27a07cd65271788df1f36120c9b833443f466bd9872fe9256a437818b175a988c5984f36fcaefabfe195913c5b3bf101c578d9a118f034e4700fee9762510e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58886ab764ba5cf2f2d2276fbeb50b5f43babaaf5541d7e781a3460e567ccb0f72895028aa9b97719b01c55264ff311a1f6555afb1a0f4230238b7f89f1df8e0db335a3ea45954ef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heba08b719fdff743601d2551941d5570c9ecff035cf7313f21b56ba64f8ae0f7ffead220b0fd4bfcb9d1bf4a4499fb39e3b2d9f6a9023fe28b09c313ae27c1df385b09ad839326b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b8a4c812c88f9795a609064ddaf31a4d3dfb4fb44bd467a2065f4c594b87357fa6fa86303347cb92bf7a58f7790d8a8a78ea2923caba966dd8c1fd8091590b8ac6f109ad93b16a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3dc17f667e880a3fdde52a6d39ee0fb3f0f0cd48a0efc45c23118138e284b9f988fd1737f4e2be3a84b90c8fa5d0ab1fb4bdc78d8c50d772b59261b3c9d621e3dae4668a1ad93d32;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf94fa504d75ddd1adaf42f6a35bfd625330c44104c605d63f778994d97256c566ff2ac380101ac1def5661a60f701dd6972e89981035e4874b039aa0ca87d031a5ed16578b62f149;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h921cbcdff4c5898e94f855a929c9f37df33d1fd5da343cb5f9be61f10e45a1168578d2a5e6b0020716685a90df22e19fbf30a9838c171917b5224370464b94ce4c2b6cac12dca0d9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2374f394d0c93d51136fa2f09cc0476b080732c2ff8b4bfa174d93aaca34bc8f1162c3d26f5e86aa917b57ff1d372d5bac3e46536e69234b46311f1c7044f4b3269bef649615a57;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0701948eb4f9ce6f1817965aba5d62a2315e222b11204288306ffa7559ff86afca38b148de51225d72bae5892b6467fae0f29408999dbd53b47fffb7ab1cc2ebaef507740f1d8ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h422017209867dec9bd069d87c07ce137e26c1d4c44d65679cda273239ad48415c8273c863b61d1d1c594a1b5f36aab6c419fb18c5b988ee681da81ab68c2342ec99aef7f79b52f3f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9fbb4360ce3d211e4053c6bd724c7d628e4242bd846ee228b7003f011dd2dcc9ca39834d5d38f118188fb56b08881b723c7480c1d574efbbc3eb4e2373fa933ca512319e3f7edbe6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9a925b36953d5a9a53feb557016df089b6c9038926148b00efb8d6f8868dd42b7701965cfda586a1e4cb486564f1a9b785181626ba199eade1e9694a9314ea80e8415be444c1a68;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0ddeb1267cb7cb1b078c592bfcbfcf1bab8770184f1a0ff00ae3a256d468b941c41206434f60d22f9fc0377a68b2e17cef88e38f532e51658709bfbad92a39a88b6b54229c37655;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h194391de045895a3fe76f76c676a9095c447cea3e66f83ae8819d3ab51566315ec0050f6249d3018ceb91354844e277a045e21f3f8aaf98b8a59fb54085749baa62333739003cb31;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79fbf61d417c78e2822fe013d3dd7dbca29ddae95ac5bc6ff7ec2052d52fea8e3b87c04b8833627c3fa43272ceed64cfcbae7db17ffd54e430b94d6032a7a2cb6634f0316146a0a7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38b95639fd7da04e4511d8d9515350bcb5f76874ee8997a91524294bc15462eb854a9eab78e7170ec0c759254e32e621a5bd092dbefed05dc0fa6e8331b3cae9d45240f3484afcee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3dceee4123755c83bbbcf287909cc19f42274698fc9fbf3fc8598721ea3b440a129242c0ebd6ff432e11edaf8ac135d28489e67825370ded09fa6c11185aff19203bc3d887d2c192;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc7291f293f25ff35fd777fd786d4a0ee89bf076e2e790a79ac616c0d57704addbe1f1ded01539411505e3fbab79d9d0179e992e56fb64ac922e4a75a7066a026bc55e43bbdc4f7c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9c9a20d532fbfa15402bf6c44a9993d183cadc01305fdaccc949487b8bcd01ae8ba3585d973185fe245eaf3812287f110a604ec085f49292e4883499386fc07fb2d87fef2429c75;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcba6c1368b42e0e61002eef979d52c3af211504825d8bc5228538c6b5547f030b0f123522fa97ed18e70e197689f2d0e25c5db954336e4e85244ec08f796754ea2d5382ee1bb4c5d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4470ffa7717ea8db74046e100efbcf44600e4610696f7ce551264d2d3994d6c41acb7416f84c44efb00e4f3b6535b13b1a99bc660e57f447e30981611f7a08030644aafa8fca0381;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9a1f7ceea823d8d86c8c4dc1a934eb983747ebb3408567bae6f429a06be73afbc946aed0ec2f891ebce70a309003a826bf4ed3cfb55030f9e5490ca959b2323c5ec1e2bb8e4f596;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7791a38fe9c9b8831a34c2b6e99f97028ac4fe534d89bb94f9eef4f85f7f65369e3e5154d58dbf707a07724dcc0dc5a0081eb883950630d9e99b91cc5597303c47938828e132e1e2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he539489250335e569e0aa04314214b7b4a6415dbdfed8ca81cd7bdb5b83339e66812714021d76ff3bf08c58f11a3fababfce0d40e9dd02d2a6bd7f0430d28229395c597303571062;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f734915bc8b13f1e55803ac5c9c80868d6243748f53e3bb2c5779fb8b53cfe2efba6b180952be11830663692544a45ca66f1b8f024c04d640158a54d0becc04fb3449b40641e7a0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b55da8f311a52c04ebac7d496498ba382b552f200d43334f522e6634c84dd8c0ffdcd926ffe834ae582b8ce86ba561c1a674c501849db6a476849c549a5d128c5d522d764a4f0d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h474b8a1857beb97dc834df3b5d0c680b89f981940e773b5f9ad5a962207f1e5bbe7a246493982c20be27f568ec6a3aecfd93d42c63c7991b7bfa0101688ab4bd23f788df60d1483b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb901796b9f427ceaf86ddffe05a753668376541c462bf04eaafea9c61cd638bbbdef93cc5522177faa01469bb60ecf16f9c381785b24a286abd157758391559c3c2ca007aeb3ba8d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71e20457e93cb46dcff6841b1c710346cd1a22cb265ebeb19d94a94a678597fad4d661ff1ece5c54cce21a897c0d0eaf428ed699e6ec0af48065c5f60be5615e5ad3b5f607b1cb4b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5393d4424156d80107a242ee4d580bd3009f0f8834c193a3f2f0de513b46e77d2d67ad44a8c2848a8551463254ec8c0143f4e544ad4e158778f9d3fe3942b984230bc8ee401fb3c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2519398a0058fe5aff5f0c830a60904b0c8db4087a9166de27fb95666ffda3d720aa10a9771fd92798ea88a2ff74a1fb07c9a82632768dd2f588a02366d091442f921997fea487f4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26cc0650ed825d5b07adab36a9c3c7ec0af193f8055cdbc50d3826ac9a6a81fb7b326502ec98d5c4c3a15f85250c61478b4f4c8bc3b2877f725f2418d8b06bf9d3f15eec2a8cfcdb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc940bb24b079ccad58de8e03f12610da179059317e1577bc74ef7b467ecbc47f5214969cc8c92473032bb9fd888b8e6b4511371ff94a3716ab863ecc49ab5594264bb3ad946c8ecd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26aec03cef3c8bdab8bf370e7d69bec3d4f8439770763dde3487968ac0098c74385c1ac0f8aac6918bb9e8567ed3bb57c240cd6233cf86fa0b145cf1845b3a73325aa62d99590c05;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ee7f3d96316e26789f8cedefbcb11fc416bf662ae6641cc4372e0ffcebb49105470f88102cc6654acdea417c117fe9e4a7bd2f239eb5fdc1e65ebef40c3e3ba4d2f63b3b732ed18;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h17b40e6fc388dd4c64dfabfa38c736c5d36ab94bbb0d41cf5856d5f4ee952ffe1dfe4ba0ede099776689818d7a2d33e51e2e159bf0b5c605ac10e9c1ceede5c21a73e59a09f97304;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c52fbf0459faf7259594d56c0a0108e01e47bfa2ffdd632c2e2ebbf3f2e58c621fdea569e41fb1f6f4e6868a45c19cdeca49f3d07e7a776c089bff1323f97b6dde008a590264963;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9dcc73db095554723b0c2b68bd2194add8522c77fc13f63cd3697737ee1bffaf9fa051e70393fedccf15333f83d01dc39b24d49140bb1cfec57fa2344f4234c3c9427ea7b009ae0d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58417747f456b72a061d9585d2252dd9a19b71304eb01e4a6ced1d05f68cb952d355e2abb4cce7020ff5715684f2a2100e80370d8a1acff327cffd6b1c840c8df6d1f4f16ee55b01;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1742e8e4d0a702e5c8f09fa54b91cc63ce9fe2a65f137777e261009003ce2a6132f8f4773336b8f3bd78de07eec69b9a9578d2d13d011cf7fab22d7cfd1cac13bcb138492ba8c9c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc33a6f70dc8aafaa06bddc555fe16784d3adcab3561d330dbaf6f53ecc5e304216dd9fda06420266896dee03e075b6026ae01b53c2b54888512266c3c5e9642bf16a5d8b2b1290e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0465fe2f4090cf089e27831d7a9577f77f1f298847eee6824eca6dce812bcb254b886f1b97af0a6e88141bf684a715cae7f01ff3f9ccebf7b10698f76ddf4506ada5f901bf2f743;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff9c76e377e4e4e8e16973d9d1f9cb67e4a9f5ac3fbbcfb98d62e86fcea6f5eb2cba79dae0caab85ca826f7ad1ca6ac038fd8bcc0eb307406e07137a44a240cd15adeba082afba64;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc79f0ffff5f0ae80a42b17591dd77d4466514a9438bac39c754c474bc6257ec0f37173548e043204c1eba4dd7641729988f6dd4c7b3f5faca50fd4e8b3c7c8fedd1cb21fdbb2649;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6aa84b4f234be64da7c7d7fa68151262250ab852cf481765fe326907ae7abfb6782a0fb3aaf5a30bbce03a3cf9f7e9badcd5757df3410cb02e32f369d075212bc779a866b28e8870;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h693cd6fce280551351783f3b6ab6a4df130fdf2460cbdc5c25e685fbe60a19731826cfcab65372dc6ccebd6c827707df1bb07836b738545084016bc238c188dbe121fd5d1f320d3d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c16c10e0308d682caef742bc9777505fb2f46f7334356c9a792ac95b2ccf48aed4354cfd58491faadfd7323307163d0b3cea5a1d2047109fdb97ddedd6e9f210179ebe5b947b368;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee6728c26b1049ce354c3f5f3f46ad323041fb19878db5a859f76acd0b6977f48712924c005296fca619b147f0c403e22c5d16d8951d97e09bdea77558bf39a1ce630cfef953f1d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cc2f5eed72e936060681c51296d41a2bade1e7d2a7d013bc7facaf3ba190abddd1751a71b988e51715176a1cb5c3170fb2e64bac8c5170757c727168836f7043f4b9ca967731525;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0453500176674a0d7a06cf7541df63435dcf629b3ac55f696f436504a03337eb2c678df3bbe8936240b7491a57eafdc3f635de38267e5fe4584204a26da270ca38546cafdbb417e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5482061a89e117706b4cffad591b553770c10e9cebbc5b79a0c5b7d601ecbf4b39d0285741ac7e93f593945b83f8d733967cf414226a8d997b48b6b289bf8ebc78452f3a8200c34;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h747b376a5c98ac6a631c92b7747b6331faaaa19345420d4dd831d695400791fd888ad8d4ddd6442e6049de26700a3897293a6c02d1c6ee44b4d6a3deb591ff48c68aa030d2b6dc3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6cc5e8a62e9bbbdc530e45241387b9ec071a83f56e6cde3175258dd1dc19bf966741ed8b35681db60b20fd85c9bf340b2d31477615111007f3191d9272fe83d00707baad73dbfcb7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd30b46cc8e45e3f1d73ceb153c24b2fd77d2f1b6b1f40c370c3cb5fe443cad49fd0562ac8960218a0958f66ba4d5254b4f7dfe031e49a9648da42eb0eaf6682f73994a531cd5a569;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc133efd98d847fc5eec8f1a884d03a6281f03a140014c8e046598c055889e183e6615c716fe05d13039a9b82ae314a721962afd14fa2334014dd749ca1d37e6a8b9725b021a06af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7800a5e56b66a1925fdd86d8a701b5aaae383e2c9d8a139802594dce835b39a5c0a4a11e8e1576f754203ba5651e3c8aadf922adbe1f553681d528cb3831ebe4f63e0e5e1d0fcfb6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h230211d75aa70ef0828a903da498162feb0fa3e2cb694051994ad72868afb31ec219d95a6faf7dbdb12647b7495289b1b1e49d5bc3350664576ff3c0a2e03a3a6f102946f22a99be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd6d1d5a48126e2f6646cad344792131ef7caf6a8814b093d07b2c4441ae6a340ae85361d7bb9bb6ebda9c1b865a815b37504083c6e6596617a6971522392acfda2534583c0f8885;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc50c02285b815b6a171e51ad11ed32e63dee3539e60129fb6e89e4b783420ea590fc369e634846451478b702695cd61a6e07eca9702406c9626c87548f4c27359ba4b6056d7c99a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f66cfda862e10508d4260a8422de474f73cec3b04687476355b1d07b02488c934b89e6f6ed5f00a9145d364bc290474ea0f5fd292cad14d2e63cfb71d970b49aed999ab7223406f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2d4cf943969492445ca9578f84f51c4be28327359b450cc94c96fa389e74578a6775dabbc55761e18404d28ed0a7558ebe0e77a48034fb7b76d47f60d5a915702abc05321aae474;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4c237dbf126442510532377a406ebe6440d12729884f4caeb6eb89d13abab1f41acfcb1de567874a6bc4e35d3689554c31cec3c39261f5dae50da6e670186b5a25506964a6cac4e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcde84f41adf263e024e822a3e0df40d9a98062ffaa9f6b76f080ca8a66bd7018af0842e5b358b013ebf3c260f383137893c05325b0a9b5723265bd411d32e56f3289b3ef0db6e2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54790c59e031be88dca9a52388ed8d8d1727418445c20508eac426b7a8573a55fb7c6eea214969e67b3439d0df20c7db791e5d61cc408e9a43fcd158e89b16b9bb69d54b4d7c9314;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4058752aaa213adf30d5b949c86b120def797117a6a9e1e2ebbb9e14650808062a34218bab7a782e7de6faf379807d2eacb0c79166e04640ee3df3a40a2ee7b29f5ca1aaa07e002;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e06fe69b56e313a4e9df65606f1fec572540e7d69ec60ee5301ecde8026cc3399aea0940641c4c5a11bba70c14d4d52913f9ffba22dfa6a145be0a9ec0bd101bde0e67197a0ee26;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h17a7bf5ce85452e1e2bd119009eb9ebfe76fc572d998db027a363df9a123057ffd731e04ec207d2519fd79acf381a9eb466e91abdb3d7a96406242b1d7aa47ceb94d739dbd4bd463;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcce9ba824f71c8eb23527cb4265826e9f6fe9b0108539d8401b9806ebf4c9507f7f0095543caf62d763f11113b675c7a3473f66a49556f50d2716f4894e2587c2791e7547977ad3f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6ea570782098217ecf1ef9ca1413c3cb661d0a8d54e76fe50917ecda90e855774e1186f775edc38c29aaabc8685ecb9c71bbcd17404a961425dce9ea22f85e4b4eaae269b90a83c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7713aae19ae868fb5193900e46048b3b076c7c603f5fd3cb783b5d61efeb230b1b9fb31e5a6a2e121bfa28846d0e1df9b5aa34c3b310584d77086811390049343fa68d4714f0edb6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cfcb1ae1df40f34c8721a7e147d2749a926d50ac85e5606f814cfb208cb0fbbb9b607e961d548902ea6bb8398c490214554d58c3b46096ca5dd266ee7bd7f5f7cfb9eb937bae2a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8490a5043b9d6e0b76c2921a064f8f2a6d348039c9dcc10613ac0ff96eef1f5b016b285031952f44cc5dab2d313cdf4291cc8a87f758ee6719c635647333c3a87d7a837ded4b9ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h943703a9d3555c478b6cc0a7ed15990ada2af2506cb080597c492390b9743edf193a16fec6234cdff0b85cc900080d3cc7c97f75200f9ace3604705278afd9deb67ba4fae7bc9085;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc45bea48cf432c5657426d03d49265c13bf701e3c885c054ad1fe536be9860fc3e270b37cfd03016941e1771a121c60cfb76bad346fca88796c5b6208064025aa0d39144d3a4ef71;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23400ca31b1cf1da56d35133ea168d600427356c659206b0ce53f225091c2e6e6385c818bd9c39425cf3c49cb01242e7b19c2d6bede30d1faf0bfd223aa6dcfcb4eef4f31d6b55e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5279651db8653d118c9c29f3bfce7f4cee24377f96536176e401df9913722846d75096a48c7bc1524667ddc4859523b7f9c56ed18b10cbbda5c41b587425cc4a4877f0c61f53c1b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfca9744161451205b37475afac0accada5c3da3be45d42b4eb01f1e8958a73ef6edd99ec20935262cdbd08eb1acb4b2a9bbff460405ed52a7aa04c4217480c1329c50b915f56ebd8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41ceffa31469a5b84913951d1aa5ae4ab41e0b70d9163050ac85dfafb22198dcd8fd58b0c1884e7636b11cb250745dfd9cf248313b94500fd682f3596681c182619c17782a5d0714;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8051756224f2927213bc697b4dd9bf31f8b3f8e6b7e313f787f183f5fac6658830bea37699f36ac4b9a5730079e44b0b4b97db81012b5caafaba454f2efedb588b2844444ccc25a5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9bc7546b76354f206f41b55ff0f748e7282e609c98dd9559735b253b5957005da0c7e50b220c97f8e1ecd4f6193b014d143f5fb64f616f1e58c18757e7192ba99da17279fed44c44;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75b2caed9d2ad61b218950cc272a5a29bc26ec322ba540281707793aede201e24f43406b5ff4a26d184bf52825b6132e716287baeeebe059534bec75a958a3a3fb1ec839fab6813d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc993429527d84dda746c3fa3a8e0d498c5bc553567fae3566452927c86eb29d8054e7a35044ec0d8b381fdd6551f5a34943a30640fb4870624b87551570b882ec0f1a673301f3988;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca5cf3dac6a84b42dcf7866b3cd1264f038c9efaac60d479b27c359bb0cd9af10d1d64ac7a3d6b84df11b1cc54d378b140b9bc876ee7e007c7510ae8902086de1623803fddc5c38b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d4fe4c481e29d8367d29e0c4e7d23942860f06a3ec9cad3ff77b595e4a7ef44a8e8dd1706d8814f79831b7eb442e904b1d7fde21a771736f73d697d1516a2bb9d0027eef53aa0aa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50559bd4c1cc2b55604499877cdb03f8a83ee411dabd30511f88fb24cf68f9df491d74df71132ab90571b47a11a129be141e16727055e7ff08dedbfa525533b9a5762a9cb7958885;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf4448b2cda0a7479a6f8e429fe4cabc1fb499e95224e8580bd7b030008f9968f5fa6a96f3054cab5785e63f7ce577f87789d0d48fc6da6f10088b190d9d46a7ef6adb54059a530c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80bbeee12e9ab8697dc69bd1cb3e48414b0507e48dd4a914709be866fea6f29cbe651431bc13615f3e70fb762558f174361226cbdb27ce130a82bf1f459ad98bb6beebd8dd249926;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2df4ae2346d6fed1934a67af281dddbb8ad969bc4ad44900af4a3ee55be95c7d53c359f26759161badb368d69b2bef17228bc01a665adbcc3870ba9330d6179f6c9b9de83ad989df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b0bed38a46461401ac8080dc843ae9e3fc46571449d6c24b02211fc05b3869c4f420ed5d178f3f7fe0bd669e99b81b7f610d4069a5e205f14f6232967382f3a74ffe4f8fc9803c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36f8f8dcac0ef09628a6a9c9c7783d842750a16742013573f3b9ac595838e2b20fdc69bade77a0ce129364da1ed7f508effe3032a292762a114b9c29c889424a1ef66780152e92f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e2297cf935d8f7e101c145398ede5080ff99c1107452c132f7890c2b5793e332bcda05cbfdd7542a93eef9835c3d02f022bddbaf39839f65bfd920e8af521eb1d446134c9bf174c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbac31e9fd2aef0132f54f98dc43d8ef441c08847432cc41051b4772f19dc8753b7a938293fc0e8242cc2afcc605851bb7fea213e9a6abac9f169556cc381ad64b1f7b794efdb750;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54c12e2427c03baf2d6991f0b87c397ffb111214f137265938c5ca9facbe9196ff6e4746ad94f022a5fe67ff43c66214158cdfde2df7f476a9614d76c2359e851427816e1a5c4766;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce1c7f9d2698932307acb443879bca92e7f3b0f23faec4f936bb26385d355602e5241bc54f4f1242c7608dc79c892287a6e54e76bee0b57a516bc29a32276573c36009a6f08ae005;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b9693c4b85aea60c8557bd581c2cf29de6db32f67aeb3ccbd2f784f8ea6677c7d905a827e6044d2f40e07d5cb74b7e3fb4382cf71c7b0b279e98cb517a13b2672f7a472ab0a37db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6823b7ba913f519520d2da6da8cf1d5fac4d48522e0be6b1fb15a241ffd59aec027e7787d2bb6e19d3b6c8360d594be978691db6bd20efee5abf6192899f244a3c16d9ee5670ad87;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5973948fe677dec50e71f6cf9fd9049fbff42a84df7c4f444f126171b41deee293cc9ba691375939d2e33ffc98c11b05f947a5a290daaad615b595188f592cec041401f32380c250;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c2b73380426532a837888dd6b1cc01b982cb304a95e9e86eca209ac8bb315c21d1ad61d7dc2a45396134e35f4de5951b08f264b6eabfef55fe91a3eb2bf9e9a4b0422f6683d4294;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5fced2dca57650e50593e62f9a9bd8e5771dcdacb61a7f1da57ae4db9b33750d63b726d5a995fa4d187c4b4271a214ca5680f13442529d31f304bfa38527ba453c015f1cc579c1b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85d3be5caf60334505c0f8fa95fdf00ccb10c77d66d1983587f6380538e69225a99f6450b22f6ccf0237fef2121bc529283b362a92e6ea8cb5f7fa28e3945969721bc70e42037a69;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8d5a3a8e8af045b5fd61efc95ed14ea9aac77920d438dcb19d3053e4e36a4693ebc5183c97256fbca72a52d34ccd8a948cda39d30a638884b6d40ffe368f0b7721e456f68f7cbdb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he113f3f5b7b0125fd75bb0a4dc67b189b02baead0c6f67b7c5043e7c522f8b71b4ba53fcaa331be6ee1129dd6405aa143ec76b9b72f40573a61a1b168eac21e478276e9df079928a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2600b378555ede6e82db2a304a8a9a783d089dda6b3e6cb49973d4efa1492ec739cdf5902b96aee01f1709f512f9f5b8969a6d00504882988847ed0ccb5ab7927de68da47249e818;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h231d60034c3d1b0e147aaad52da14076b8e7245814304a0fa8199a80375709578f07dd50dee97c9c18651562e48e070a10d9e36db75c4aa9723d24843b83ea1cbeff9fe401364b33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32317de4088406de830487fe54276bd34f084dd8f29692eda6167db5dca5beed389133b632312f1da418d3bb9f5fb1dbc00dba18926e5cd28c3ee8c8a8dfeddcfbe289e0bfa91572;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h769710571ffe7b8fef0b3560ec5941aac327509c1ad599753e82cfd1dc0e78f8e2c00b811f7ad8110112a33556ab6e6ef216ae5f927c455d4f0c81ccd49b43c782ed1317865e750;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30cabf890537423b95b3e6bbd3bc16e993c56ebaa1dbdae5e192557619e24a6cef5658d95c3ca5b691c092a79ea43f34dd3f81d7a332c4cc6f1e95bdb620a8d66f8cc4c612b31914;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7be648a0daac60268feddae79f11cc7f22d7bf38aede440f40b37985ca444cfed4837eb58fbef8132cce6dab32d636e05f3dcfc88b5daea0213d2e8b0c623fe2ed5cbee0c2488d1e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a9d9f2378c18e9879e94468403420c17168f238bc4205b4894aa2fbb9d047b452fd3775d1878446792c9acd471256fdfadb76e0d53fbf41b20e74b74aa3e5d04c61a9babfaa5e46;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb33eb05c76d2b3ae50e36cc0d034b30fe07421f6d830c633ee8df53c7fc537fc008813369ef0be9f192f8ad0d02a1d0591fc8f59e66eeff309da5e871d17ddf3e4c179709feb964;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b260a81a271b966857358675832c80f6d269056da45f0af110ea190345bd023bf7496b9a70bde10c0d276f40546c0c7bf6e7992aa3ed59298f264d1558b76f002d9e8a5f4ffed58;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e0cda92de9927b9aa37474ddef96df2500c2531c576bbc0e1f4f00969697a338b383c3f6390a0b6c38874157801e2205a9c7c3f96a5949c250fdf8e91d927aca213e7978001bd1c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95606676b8ece944d7586b9bb64ff5b894a1accefc854f2e1ef87d179fc027591329edddffd6fe2d8616be191101a6401d41e4fcbdb6a8bdce6432b32261b227778cbbd918e871f2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75cb0ec3e3d28b034be011e7305aa001540545738658c1c428e3106bdbb9a7e152c6d6a13d75f1f04bc31569e9f910904f647d7d4c9215510429bcb3941529a74c9fce83c1520249;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbcf7644e15740bbdb44314a9e135ad1e633a4ac98d4724c82eb03a258f8f44620849ceffe6888c1b2f6e69c3788c864822a996ac65459622d24c6ae7843279d20379492d046ba124;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd0126302d4b09ffd316f33b5a9022bffa95264ab913d594a8f8209cd0f5b72141b472a8c9e427aa6544c613689576b311ec92f470c80bbe0a9618da30e1824965c792cd0acb912c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9d75024d314649923bd2fcf202f76ba8f55dd95d10f9e031ede6e4314547c0e1db8493e7817e363dc201bfbbc64b6c167bf19785fbf1d44fa914e171b78854cef7a7d15f03c3b99;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had6250eba5bcf4e8f7758a763719b799ce67c981f3488864b22ac8da6a152b311277d08398532cf443c7af81c27106ffadeaba8eb04017ff893e3558ba7c95916d8c917f71b30f5c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44967e160e12c659b7b6b625e357a07d3a6e562d6a8f42e30ecfec637bb34c5acec7054c90bc5e58e4b1aa1337c01f07a571e7949c6bb769fc6dd4fe04ed4ce5153adea1695ff3b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8f69202fa94f1e46c9ef09b249a7278c81d1b0bcd99926d118a62eb0773a1d870f3c6b9dfcc5476051d30051f84906b27be0e4ebff25745abfcbdc8eb07ff44bf7f43a7d738460f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71168d6e905954f264a7189f4f8eb84cff50cd11a3424cd0d241cb42fa8175019df3aac4224221c1702443b0a6b87d2b7f0b1334728c0f9f4a9d08ec834fe38928d3a73189f2837f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b6574f211adf3dfc95366c343c6cc1bd6882f2fdc613f2546bc730fe4f11eabb36b08598da4443dc1ee1e163202431a52bd28994e9d1166f2f9f1c854e1bff00e1cce49d942e621;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5365a98282527b98554a4b63bca8c436140e7fcfe859a2c32e81455d5f3681f4c4d5926e8056fa4ed53639d1085ed31677b4cd4186238903f0372008255bc5091af3c6d0e713ea2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9221b25972168e31a7217a9969c0ed0e0d17473bc062a8b31d764c7fc40e24ef93b75e75debfffe3faab8d62baca3240d5e346a45e956f6b2826553481e79e7e6edb2eea27a3444f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5bf8e8df5e8ac1def9da7978cc75e944f576bc926414e997defac2d613a7c73f4fe914d8cb987be502b486572f03a61d6fedd01024d1bd3f8e70b1d19fcf2d56195b476e3103a06;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha82c82c7ee42afc931271418fc3c7fbf40b87bd584162ffbc34ee0f8f0d6d36480be2b22e9559f2d97c2abe1bf425363871dd08d49114bae84b6a9f3ee77fd9149dbfb291e6709d5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h784af8d5b8260c88326a660f14c9046fa5834ba691b65ff2816c73e2dfcd7bf4e7398589fdb356860caca4cd4394d3b454fe87c06756d93a01ed85c173be0872010dcaecd0ef81ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f58e3e0ddcda470ee6f53502f9d58a738b89c0aa977000389dc5458daa7132d533e524325b94d5514d01b954610d32aef9269c101558e708764b01d59c8fbc4ea66aad8d684943e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h460dcccf4ff88f7eda42d92e676a55ebddbacb50ade7b8680a1efc4013c8bd2ab47713bcda99eb378d66361965a2f4d2cafd4c191c2ffa2f292f11127a4e8f5a0f584a0c414c32b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ecc46edb839c8c081eac71c9298169f368ae19c341415c686c7031a040628bdeff562711fa2c782747eca3e4c2045f38e6ed6d0c25f97759b85b7de323e3bfecba159e41e696794;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59b94fdbdff68cc8420515c3600522e5650ae578583009f4c1273c4d7a54fa55683d28dde7489afc93bfec173e06c6e19f8b2f97f8de4fa78d3aab4c5391f3b176ef30d5424c195b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3b238688ae102a1e63e590a13349a66e219b6a823f479e3fc6e2c4acbe407719801ec70acc355beb35173f59f6232986cb4d0be3b9fac49ada5d0679de9808d01e57603e6c3bd3a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9073db74fcbe2eb5b047c118816d71baeb6f9b42184a7d2c31804faf6143aec1cd7d5793e3d5d6bd0fcf69b224400a6bc61a7e434768b3a01ff44350a100c97b4ab4a8088df992f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heeb371db28e0252697768dca90962dbdeb42c73e76a3682c9d26e298211cc9f045d54357da22710b7c1b8f6aa59d7a2b8fb9ce16867ac4383f857cc5c01669db1fde592dd60b3e7c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc872bb7915a006fa9ad06403d4b5a5aa037ea54f19a576e0f1518369f4ec3d7fcb9f3aca330d63a4d099e6728a107d691add4a33b0fc8719ae30a0bee3341ba2d10b91ee6db0ebc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h328fa25ad5a1ae385e96996b6025d71518e30b559b94ae1a2539a24da21d101ec40ea08e79a1b0ea15cb341ce4db6d505fab2b8d1ab682ce82e2001276d1ecfb1d1e0810714eb8cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd20bd971e2ce0b46c86383b98bb30edcc08c6692d52bfa3156a6f4c11757987e0419647caa31e5e8ca208e2b74105262e3fbda729c93fe6199859765bd492d5dabe05880b73bd749;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5923c32213b2c0f566643acffc79ac39bdff9a2e4715c0d508c2c16320f14cc6059ec7fbff47763458f54ae4a98d70466175a8c7f809b933c7b649ff563e6915d00486fb4f0b2012;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha09ec4c8836098136005fb0a6b1c63378d4268adad182d36f15565f198d4c2de50d109f8d9cc737a6ee1debe6317f0ae8d57d0f3a28748ed6b9be8cefc5214e72df9d9d18aa44bf0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8735ac954af3c5552a8e6d9dc6a4fad9a3c8e6b68588552e13e00139820d38e951b9105e33efa0bacc62811b8d045dcee97e8e4c3f1e16cb542de63a3c8f4c204ca56f219a27535;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a2dac6d0e8289e1cd79fd0f5dcb00d0445c024632d71f419ec1aa63591f5d95c9b4c687213f4f516a4451569c0548178d0527444927be210ea2c732478b0c3fade5fcc5e07d248d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ea15af923b20c1b2bceed11430d5cfab91a170ea4fd1962649d56c3edfccab788824fe49f995121274c58b1dcc73316615b26f4baf97bdbfc64fb9a3b87ab424cea3b7d61bf6d27;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h784fb29a8c555a43d2246654b841a36522d48dddbdca195fa2d19b07c063636d2814df9e2bd2220f7de0dd5ab27f9ddbb332661edfea9cbce31644a2c5158812344d5a29d70a5d15;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3397a8c8004d63268de5278225d90e1872d4d35be53cf455fc3fc3f9301bfb40482a6dc539fe452a29883c458b38ee38cc2d2748ec6525fcae71db3af3bd2f9f804278e72e1eb52;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd49cb692356c0bc7d00b793754383d4a85173db2796610109050a130152a1419381c80644343435253c33aebc34f8bac36bf577d04bdae39bcc53b6a431bff5ba3c4e3538ab35f40;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd13c26649c5801c46d1d4a22c61c986b9dcbb586c8593a5020886f270283b1abaf3d1722ce863b4027a08cee403d907146aef82b25fb56f4c2763acf822820017ec1afd35ff1e5f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5abcbb11e2219ae940f79602db4cd246199e253c2fb7e781358f54aa2d49992a795bfd0cb7e943fcfdfebf70809ea0fda913349ed23a1c8d48fdeda0de4668092698bf8ac6c1e87;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea8c5528468fd17b828c44823211a81f8dfa27f15eb98e39e92fa27e1be6c9377614510da3335f4b10b39f8af949f765944104418a48d2d2312f4a2cb5880d36ede76bdffdeeb51b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3c23ed0c0b8d6ee58320a6ba20379a30d0e1222b350f5b39ccde7492cbebff09c41011e76469765cad9a87a3ff6c9104e1aba3301cba4434e394ee80a2e6fcb73c62f28399021d3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8a37f2eb1d4b1b92ed1d1da0944ade3a6e6ed37df4d2208ec198c321960964564487f69873e93d3d8e85bd6aa60dc97f4783e20758b2c42d254fca69e7b017cc9364a64f179f427;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99ca6eee3d1a26eba88b7a8127fdf9b9a092dcca394a227b9907b4c9480758125a1e05e06f604eec21753271d79dd14e67d67fbecc35224b54a8b97c7dc0fe899cc24b7cd84b5a33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a6a7d5e998da716b08f7bbde751b924ddf1076c62e763e9e0c0279b2504029b682c2fa9fa7d508be08384499d24f5f5e2fdb8ff9ce3aec9d75147ea678b015508e4f16b3cf3bdc2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1b38b43649a22148d422e53c272895ee145bc381ad37af424ea7772226facea67b4c7007745301999dd82c0950cbdf0ae71eca7dafce994b491f446aba6a671913449f256707417;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd528197d6942f48097eca8ee1bcc8e57abda0e3af3a1f5bbe48c7a2de2c0910caf36938377238f30d4f113bc077134b872253e4e68d0ccfec3ae48fe240377194e61dbbb86bdd88f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7fca3043ef47377a85e6b2f94280f9e9e7d20ebd88d9b4b7b09e9d7e57e4c201a2956a868b274a39a631ad382b3b4a39734d9e0439996e594427f11f788b2eb7bfa983f4f2ca5fc8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b1474b74a78576bbfc6d4370207c22752c3b8663d3bf2f5acf4c74ba2ba669eb8a451ebdc3a4296a6645aef6218d322196fdeb3ec033a0b6a4a49f6d7f79af6eac31b717cc6aad7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7654ec67b2bc943c1cf30bc7769d1ceff5abb499aa0f9db10a395c21ddcd40e3db99a653ab5102406adf6f74213b831966f813d0cfa22fed3ad3e81d754ad1f7f0139fd5db9ebd0a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7db7d721158564c6fd1da6df0885710b2381e4bb91b8d539c0fcd31288db5db4847b723ba92b78e10f07f41299728f1a5f168c763ed650929af39b6119cf20b5b65f2a36c4392d3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d6dbf87cb76de12e3599a4353341900ad79286262bfd063e8260245f54a03e25879cad1fb34ff1801533d07f970251729c0b86c20978ddab76284b9d6f82029d0c428fa50eed8a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f90f779df821c4d0c7896fa06c6f598ff7192c2cd59fe763f40e00db016a64063a7c18a8e03e17bb135fc069b787c4546888503043d72f78482c56b8577197b387172cf6edbcc51;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8cf65ca5a19ca1b69051e352168684e639905ad37ffee6e3c1e62e40acd01235dcc4fa539a771e79c083322a86ea40b06bf5227825ef26bc0840675f1c99d131862139b978b9e63;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86858480bb90b628e9d9d5442627a4f17125230441a7ce0be9fe90d02b16d52fc231288963e9688fca941a05ec8d6b6d9f654923624a92f8ff8ee3045226a8742efc2ac327bfa1d2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbfc13c8eae2f0844248d6120fd74e53881e26938b2c9c0350421f79decaca85732fd4b6a2e3a4782ad46dc43a218353b0a0587c5b023ee3470e88d52a0e7460c774ca2e8788546c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12ef3b8a7eb2b2cc0e0a01649c2ecf00213aada8b621497dda119e8e67b35188769e0d1e3b130dbb7c92b7ff5bbaeefb1c36192e34e941d05fb4b6bd96e37962cf3dd5d04106b1b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b15457ee82047c8ddbd837cb8081c91f31d506d5f4d0fced72134f54dc1a95b4844a84c47e8882a602e335fd036329fa13148bdeaed1c6798ed8d366eceeb1d7ae56f68f1f29b70;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7454367f8f8dec56695b3782bfc28a6824d9969878600b348a0b852c8a1ae5422ef5403fb3201c596e48053384de374617b5750662879063d05c4ae683dcce951c49e5be83e5de8f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6099e014a7727922d2bbab5e9d343a20da83243193cd6a9327252a1984b98735ca1f9c2d878a97bc995ee7e69481652d7101d9c89e7fb1547ca780d2d4577764491df0531cffdf8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa05a412d80b77a131aa933f9fe0765b5acdc0c76d15b35dc84dd8192caf9d8103c1fab4809020aeb7a27aff3f3b70386836e74c82c43a600f7d854e9e73d705462f4375c0af4d62;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc56329d61e233aa3d278555d0c0bd6d80fa5941ed948cf7d3124a3705ee973e440958567891ed3c036d4ca37c51b67d94ccd047f057e03cebf32480d85810e5a1059759a3a7d0b6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf924f0335a2b5ad9b7ff30e21cb05bfb799a2f3042620bf7bcdc90e626d49b98d29915ab86d908229fc2624fe1179271fec5c91b839038089dd644ffbeb0a7ae0b7ebaa3bb63aee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5428136efdf845c17264af52358bef16c6875448f2260688cb7de038a8c868ce50fa4a93b04b3b276e250fdb0d42cf7425a0a459a3ece1a1f0590dade69476d3a0b1843c3b97e934;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2535ae9bacc4812a0d8c57b5beac8ec17fa27feb25f5e4a73dd23796c4bc812c3c4ca03794c685eeabeeae3540862d9a904fb46601188be74fbf67072c4257c485ac2272ec91eaf4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64f5586d7d43bf1f28f4f748e4c4b690fa2b54f2c37570882c4b55893f2f5dda7ef3aa7081774a70048f61ae544aae9255dcf26fb6acf0df2084a1b0465b81fcb6085db8ed0f3258;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8cb45c194d8e94906af4d169427d26d3d521a8e1302bebb0df03ad4cecacd1f4f03978e3fb04d62a69990433ba302afafde8a1ea0c86f663882de1b08fa44a6d128483229b9dd93;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb010bf24b016956364807175ece27596f11253a54da999d4447081767024771515c2cc676def85e1319662cca910dc903d32a52966942c5c00b802c7a54b457273924f14e19538ec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc304d18788cb11fcbf866e97cda9ffb6dc1f6da1a3ae90173df4cab0dc7b717e0ab66d50b3dc1085e01dbb9a8e74dc8ab2da325832f9776d9a0b709b322b6bde33f45da3de9e4dcf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c9f713521381cb94f908ff89e80742c7168fef9c7f1d94e8718013351eb41683d4347a537f56a8b756a7bace070f256ce768a9949637c9877d90f5831a0e27cc8b18feb4c395fb6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57a8430133cbec235af7195736e1e7ff071577d8afaf7fd4befaf0d14a75ac4566b1b5d8a60ffc8e411dc112e0ddbd725a5461b7e2e401e67ea8c0ce6415f39cdf3bbb296faa3fae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac6809051327ebcd0cb0360de6d2470d7b104160085a5a9d699723adad7a73d4d0a54ec7cd715fcd5d1bc142060f9dbdf7521624c37d200cfb6d253e58f8c79799c027d6187045f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2017c92659f03a099f08f5da9bcb056a1ccec89ec34af003e8e7457404361bff13316c31e2bec8fcf4de5fa51f8ea912d6e0a619c314855347e744c79053f8eca027590d71d91aa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69865cf706d7cfff98a5386f93f6c2ac89db0c9a5fb8c6f7e62c1b2aa421debadc2289ed7c19cded33e1f8b2018f01c4977618c2daeefda9f9f26bfbf8dc61aa0eb0c8d693c85d57;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc88ae916ac5389928359e409774828e873bd9033ebdad173e26cee3db97c1914cb45733cae5ac7898868071b76ee41eceaa44f0993d4442a9428665f5caaabf42214303f6f666280;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d818b873768d7b7efb72c8e85cdb1b88af0be37e8d5f884b5c8d3e47658ceedf06c4993653d0422a94a230e5c80aaf08da1dfdec9cad3da51c82e3321637d2187c16e49fdf92fc6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd65123937b620de74487a149dc9ee43bd9df8a0ab8cf70435b8a4bddd4f9818e7e5b550e5a56d569b6ac5851fe7cc21caca0ae35bae35b54b970c352981dfe4efc0b34af63830002;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44e75be21f1514a10ab0b0fe5e1c53710cba2a9a8c5453cf4b9f93ad16469ac2da66d300843ae1814ecb0e47540bb949747cc713681aa6b09699f0c386f32152ecc1e80c4d144748;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c2699689f0854f580cf6d3d499036bb274b0e05fec52c22dcc441528e3788d06ab12c3f7fcf3f579ff07a911b371f3ed5556a213c3674c74b9891197928d670db8189aa53fcf5b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h712792ffb03cb856d816249c91e082dd55445f065459e542dfcae80b928c94016b767cb8ab8e17d7b58b28b85ae3bcb66ff3c02651c33db448ce66c409f409f1566e3b0d89e59ecf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9129a4b32373aa89aabe143a4d261e619ebd389ce475d989dbef4295f97725da507d01e9d9b80cd258f3494036d1d32b66767c4be53bacd38c0276819fd252681e5c1adada8c8c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3390fd7b402d4d2104f15d964f80ec80921abe2ff28aa10aeafe489efad9b2b81a67cd370e33e10860ffcabc5c0db790be6b5343f31396a24b3525aa67f8ee118be86bb779626b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha754a196822d1b5ccfb1df3269d5879f40feea789653412b12dfe9d57413ad8e173c027bef27d5a3fafe5106b65b0055865058612dc238825ecf702c2f8dd19d9c624fb96e270da8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42966ec0cfd7d148dd5fd44eadedc93e263c4ce98ecdda7d29137bf4159a5fb2f7e218522ae507ff45f5540e7759a5e4879259adbbc2ca7885f477967c8b51649fd14b68adafbeeb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6d3f4ed06292eedb46ba3e90abccc209aa52c9cec01a69e8d8b36d7a1c16f8cdd68927716d50334c79d0ce794bae7777e6cfdbc1c7c359e99f7a12d1f8ee46a157a2815b466ea9e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71c8fa32ab9e3e727a9a904f0868b2423b61e746e8a16ead3dc71c2d12ae34bee79f53b48b77d47bafccb7857b8cc75a6ea725952419e45906ff34fd322c3f56fe57700c6474ff04;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbe909e35cee6de2574cdfe73cee122cb5723d76da75ada34fc64f9b9efb537b4e465c24f653708cf81efa2188e5495eb597bb299d3d8cada4b4230267120e371ee4fe20bb1ddc7c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6dbc9023d4d1c9718a0625f7d6ea4bf6941de24c7b06fe347aecfdb24f881749564fea6e7c1bccf9ad51d8d80ccbf0b80cd59417aba58d69b2e2f81519586002e8402d91137a5d0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fbaa8583a4c2a31a6dba08ccf4219b8061849453e9f18d0609fad1fcd7d189e65ecf18b716edc2f0617a48741c09ab2c1f9111c58215154feab92d1316bdc8583d72b0e26671aee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha345097723cd2abe248bc3007bade69bad905c1f483b79f0df3a76a2def09e8780c90642e005518989a36b526d937588493855538317e4169391a43cb4c4e4e049cf8977346c3b8a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32e5f67239ba85cf7894b71ada882e71090453d13393a6a737394db1854c5a8d8354134a54491c2b47c3af37b3baf96a6e49c752868872725cfcccb21e5ec49c459100affadd89d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6d417e377e6bf2136da1f1592979b378b40e740cf12c51d98e37d4b37fda01dbb6cfa135161d6a4e2bb7acd7a50ee0ec4dc0b059e788c6c21c959fed3a5aa957300d69d6752216c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb819aa0ea5ace6c1b3822ec0a48b4fd6853900b00fe6ead2f9b2d3ef879860106f777689f04367b436683d5de9fc36283f24949ce101802e3a6973565a0c52c195557ed270990ca4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41d67a60e84d004ffb0fd6fc9d538581b0dc1a8dcd207850ef3c9b6838c0c3ad731ca184208cd92e0efce747e5956c983bbb7efb6a78fa09f1632efca1a217815f8f56a02beed47e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16f6d537156fd4cc7cff0e1ef6beea4b7f1996da2400943c8f10df2edaaa3b9880c4287d38afb5ad1746122c054cb153dd14093f6f014bac70826a81b330120daa4754fb509636e3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h17fe7ea541647fb93a597dc2212d2d8fb75a2b379598b355fb09a0494b3794eb11f367db8ed1bb929f0020e8c89547801a81aa84366d4916cd55131d074867e46921d7b9cf3265f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1a44ed16b6237bff024b432c5093524c19c7f10c666d3c2164df3ea98ceae50166fca279215d62c58bec628d38c24c1ff252805a8999ecf8f7e54318d42ccea9ac03046d8b4d5a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h582090946257d49bb44a06df5a6e6000545f51bf808aa5cf15f250288a9e3452fb7dd3342bab5fdb18ba44e7f816fb52255d590448e44db83be5274b713db48e9d08c7ec18762fac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3948d13352383ae65d4a29322d01549794d68a2be954161336b77a73160694d1930b02a38259e52f3ba1874ae3cad8b3d9748e859f2a0084063dc703022d4d8fd7d4be8442618fe1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfca36cc1ccfd205e9d758a0e017413fdc9095752248670aba810752aceaa039d4b4c66022e60e05326da3b7d42984529c7d53d840093f3eb5fcd6c295dcd276a3fb854c93c7920ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3a5f426f7c8713994525fa56160302a399ddf3d8dc126815d4644de69282df4e8ca639b3f4ef1f2c43076f617f997d6fec2c8bbe2883cb9f9b575c07d73a7536a1cf9f1c9470ffc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19e6f71622aef95d5fbaf228cb4de6251462f29a130c1acd15d9f13433f29e92f0e605725dd51da88b9312fb26b250a44f74b2fb8c8bd3f714c3ba6cc796dbecb392844e42181db8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3e42ff3d39527c78b18f6d513d274c773c13eb0c226504631aa81bdaee08a3a548621d874f3b71bbc32d028b0f99f2bc14778c9f387dd47a7558d587f2723cd95a5c02b2581a341;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76117a4e03fcb30d89d508254c3e4ea2ba105d3837b15ef4df6b003f33e0d72cc879214c85446acc51bca4a25d7c7e348084a53870db68d16cf7b24403970c432f0f12c1f19bee5a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h708599efeb667a9c7136c8f729acf94eb80812eb43924582605914c46b66257be1edf6f7913dedb8cbb9cde9910a0e5ffda945674fbc871d6eba2a8b26dd8a9c79e2bed43c8c6a87;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b06279a4fa0f6359f77505b690242a180c1a671d7b84bc693b4c8c446f047945cffb3a56ab34b738a4d5884aa9c1e9c09ff37eb1a04bc0811600b4cbe70f3e4f82be57cff451f7b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdac8bac711451e16e043e14c4313dfcb0eb911334a72053d13ea15bbf2e0c660b8b1928d9c16ba4e595224f358ace656eba1fc2ca1e5110e3ac6cfc2e85c32b8e4fb56e9e85da81;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9d11440ae4e57d3d87d2ac711fd03e1f3d5c4e6b7bd4b57683cf847cc94adbb893e5b89292b149482b1d9ba6bddd016fa3c67fceda29409903639bb1ba28a91456c0b8b1e96cdf1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85c7f0e605c8e58d773a5f335f83deb64edfa6241a59610fc40a190fc48219d1a8bb6f9676110d89ea8dcc3bfe8d6c864dcea422e0152011bb1ddbe6afc959cf83c69577aac8a398;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94225b75133c5ebdb3047b00d0875fdc6e8ab8868530277f7fc733bdc8c8e035173fcc4b3c0d84f1301585d5ff76ba8a467879c998fc0376de999cf25b50baa508325c678887a5c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e46e962b42d219976b65d6ab5e1f1d65f1bcdee970e3c2bb980012beda90b2fe57b201c67ba6029cf09f6abecdff69316e7007f20a3491a7d9968a619323a79ae7e4ed96159d7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5047256f1068a50e712cd0d8b54f014456c183fddd6834f5d941e84ef9c84a31c2bf622428ff5ca08661590a6350a61489403bb67f0705237e3fd1c10f35d00ad06c3e9827a7418f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc84c9c73ebe1ca08ae9e0001fb6d86d69b573593074323ab0c0d57e737332f893bef418c06d8d63182c1a9eead4766a51122f7ae3f0075f802239cb20e78f5c8537c1f1e12d8a64;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6d44fc9e2594ade499fc76318a2107905177b380db2eb68ce4fa944e6054af7caeed452f46334d343ac8a7491aa49b9d601a5ef1b828bda931409d3e4739d081b87fcf72cf8e0a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h810d8e71ac7fa30c39cebe420e5e920cb9263eaa4435e1a03bf7ecd0adf9d3ab02ab84ed29d30b29a17b6df7cacd56a036cc1499c7843023373d79da4b24a2ee8e65f3c7f9ef9ba6;
        #1
        $finish();
    end
endmodule
