module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17);
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    compressor_CLA54_12 compressor_CLA54_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17));
    initial begin
        src0 <= 54'h0;
        src1 <= 54'h0;
        src2 <= 54'h0;
        src3 <= 54'h0;
        src4 <= 54'h0;
        src5 <= 54'h0;
        src6 <= 54'h0;
        src7 <= 54'h0;
        src8 <= 54'h0;
        src9 <= 54'h0;
        src10 <= 54'h0;
        src11 <= 54'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA54_12(
    input [53:0]src0,
    input [53:0]src1,
    input [53:0]src2,
    input [53:0]src3,
    input [53:0]src4,
    input [53:0]src5,
    input [53:0]src6,
    input [53:0]src7,
    input [53:0]src8,
    input [53:0]src9,
    input [53:0]src10,
    input [53:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [17:0] stage1_0;
   wire [17:0] stage1_1;
   wire [17:0] stage1_2;
   wire [17:0] stage1_3;
   wire [25:0] stage1_4;
   wire [29:0] stage1_5;
   wire [18:0] stage1_6;
   wire [17:0] stage1_7;
   wire [26:0] stage1_8;
   wire [25:0] stage1_9;
   wire [19:0] stage1_10;
   wire [24:0] stage1_11;
   wire [16:0] stage1_12;
   wire [6:0] stage1_13;
   wire [7:0] stage2_0;
   wire [8:0] stage2_1;
   wire [5:0] stage2_2;
   wire [7:0] stage2_3;
   wire [11:0] stage2_4;
   wire [7:0] stage2_5;
   wire [12:0] stage2_6;
   wire [10:0] stage2_7;
   wire [7:0] stage2_8;
   wire [11:0] stage2_9;
   wire [10:0] stage2_10;
   wire [7:0] stage2_11;
   wire [12:0] stage2_12;
   wire [6:0] stage2_13;
   wire [2:0] stage2_14;
   wire [0:0] stage2_15;
   wire [3:0] stage3_0;
   wire [6:0] stage3_1;
   wire [5:0] stage3_2;
   wire [1:0] stage3_3;
   wire [5:0] stage3_4;
   wire [2:0] stage3_5;
   wire [3:0] stage3_6;
   wire [5:0] stage3_7;
   wire [4:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [2:0] stage3_14;
   wire [1:0] stage3_15;
   wire [0:0] stage3_16;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc615_5 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28]},
      {stage0_1[0]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc615_5 gpc5 (
      {stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33]},
      {stage0_1[1]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc615_5 gpc6 (
      {stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_1[2]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc615_5 gpc7 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43]},
      {stage0_1[3]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39]},
      {stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35]},
      {stage1_5[5],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45]},
      {stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41]},
      {stage1_5[6],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51]},
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage1_5[7],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc615_5 gpc16 (
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52]},
      {stage0_3[48]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[8],stage1_4[16],stage1_3[16],stage1_2[16]}
   );
   gpc615_5 gpc17 (
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53]},
      {stage0_4[6]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[1],stage1_5[9],stage1_4[17],stage1_3[17]}
   );
   gpc606_5 gpc18 (
      {stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[2],stage1_5[10],stage1_4[18]}
   );
   gpc606_5 gpc19 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[3],stage1_5[11],stage1_4[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[4],stage1_5[12],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[5],stage1_5[13],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[6],stage1_5[14],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[7],stage1_5[15],stage1_4[23]}
   );
   gpc606_5 gpc24 (
      {stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[8],stage1_5[16],stage1_4[24]}
   );
   gpc615_5 gpc25 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_5[6]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[9],stage1_5[17],stage1_4[25]}
   );
   gpc606_5 gpc26 (
      {stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[8],stage1_7[9],stage1_6[10],stage1_5[18]}
   );
   gpc606_5 gpc27 (
      {stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[9],stage1_7[10],stage1_6[11],stage1_5[19]}
   );
   gpc606_5 gpc28 (
      {stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[10],stage1_7[11],stage1_6[12],stage1_5[20]}
   );
   gpc615_5 gpc29 (
      {stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_6[48]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[11],stage1_7[12],stage1_6[13],stage1_5[21]}
   );
   gpc615_5 gpc30 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34]},
      {stage0_6[49]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[12],stage1_7[13],stage1_6[14],stage1_5[22]}
   );
   gpc615_5 gpc31 (
      {stage0_5[35], stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39]},
      {stage0_6[50]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[13],stage1_7[14],stage1_6[15],stage1_5[23]}
   );
   gpc615_5 gpc32 (
      {stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43], stage0_5[44]},
      {stage0_6[51]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[14],stage1_7[15],stage1_6[16],stage1_5[24]}
   );
   gpc615_5 gpc33 (
      {stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48], stage0_5[49]},
      {stage0_6[52]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[15],stage1_7[16],stage1_6[17],stage1_5[25]}
   );
   gpc606_5 gpc34 (
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[0],stage1_9[8],stage1_8[16],stage1_7[17]}
   );
   gpc2135_5 gpc35 (
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4]},
      {stage0_9[6], stage0_9[7], stage0_9[8]},
      {stage0_10[0]},
      {stage0_11[0], stage0_11[1]},
      {stage1_12[0],stage1_11[1],stage1_10[1],stage1_9[9],stage1_8[17]}
   );
   gpc2135_5 gpc36 (
      {stage0_8[5], stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9]},
      {stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_10[1]},
      {stage0_11[2], stage0_11[3]},
      {stage1_12[1],stage1_11[2],stage1_10[2],stage1_9[10],stage1_8[18]}
   );
   gpc1406_5 gpc37 (
      {stage0_8[10], stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage0_11[4]},
      {stage1_12[2],stage1_11[3],stage1_10[3],stage1_9[11],stage1_8[19]}
   );
   gpc606_5 gpc38 (
      {stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[3],stage1_11[4],stage1_10[4],stage1_9[12],stage1_8[20]}
   );
   gpc606_5 gpc39 (
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[4],stage1_11[5],stage1_10[5],stage1_9[13],stage1_8[21]}
   );
   gpc606_5 gpc40 (
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[5],stage1_11[6],stage1_10[6],stage1_9[14],stage1_8[22]}
   );
   gpc615_5 gpc41 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38]},
      {stage0_9[12]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[6],stage1_11[7],stage1_10[7],stage1_9[15],stage1_8[23]}
   );
   gpc615_5 gpc42 (
      {stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_9[13]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[7],stage1_11[8],stage1_10[8],stage1_9[16],stage1_8[24]}
   );
   gpc615_5 gpc43 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_9[14]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[8],stage1_11[9],stage1_10[9],stage1_9[17],stage1_8[25]}
   );
   gpc615_5 gpc44 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_9[15]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[9],stage1_11[10],stage1_10[10],stage1_9[18],stage1_8[26]}
   );
   gpc606_5 gpc45 (
      {stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_11[5], stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10]},
      {stage1_13[0],stage1_12[10],stage1_11[11],stage1_10[11],stage1_9[19]}
   );
   gpc606_5 gpc46 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27]},
      {stage0_11[11], stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16]},
      {stage1_13[1],stage1_12[11],stage1_11[12],stage1_10[12],stage1_9[20]}
   );
   gpc606_5 gpc47 (
      {stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33]},
      {stage0_11[17], stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22]},
      {stage1_13[2],stage1_12[12],stage1_11[13],stage1_10[13],stage1_9[21]}
   );
   gpc615_5 gpc48 (
      {stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38]},
      {stage0_10[48]},
      {stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28]},
      {stage1_13[3],stage1_12[13],stage1_11[14],stage1_10[14],stage1_9[22]}
   );
   gpc615_5 gpc49 (
      {stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_10[49]},
      {stage0_11[29], stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34]},
      {stage1_13[4],stage1_12[14],stage1_11[15],stage1_10[15],stage1_9[23]}
   );
   gpc615_5 gpc50 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48]},
      {stage0_10[50]},
      {stage0_11[35], stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40]},
      {stage1_13[5],stage1_12[15],stage1_11[16],stage1_10[16],stage1_9[24]}
   );
   gpc615_5 gpc51 (
      {stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_10[51]},
      {stage0_11[41], stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46]},
      {stage1_13[6],stage1_12[16],stage1_11[17],stage1_10[17],stage1_9[25]}
   );
   gpc1_1 gpc52 (
      {stage0_0[44]},
      {stage1_0[8]}
   );
   gpc1_1 gpc53 (
      {stage0_0[45]},
      {stage1_0[9]}
   );
   gpc1_1 gpc54 (
      {stage0_0[46]},
      {stage1_0[10]}
   );
   gpc1_1 gpc55 (
      {stage0_0[47]},
      {stage1_0[11]}
   );
   gpc1_1 gpc56 (
      {stage0_0[48]},
      {stage1_0[12]}
   );
   gpc1_1 gpc57 (
      {stage0_0[49]},
      {stage1_0[13]}
   );
   gpc1_1 gpc58 (
      {stage0_0[50]},
      {stage1_0[14]}
   );
   gpc1_1 gpc59 (
      {stage0_0[51]},
      {stage1_0[15]}
   );
   gpc1_1 gpc60 (
      {stage0_0[52]},
      {stage1_0[16]}
   );
   gpc1_1 gpc61 (
      {stage0_0[53]},
      {stage1_0[17]}
   );
   gpc1_1 gpc62 (
      {stage0_1[52]},
      {stage1_1[16]}
   );
   gpc1_1 gpc63 (
      {stage0_1[53]},
      {stage1_1[17]}
   );
   gpc1_1 gpc64 (
      {stage0_2[53]},
      {stage1_2[17]}
   );
   gpc1_1 gpc65 (
      {stage0_5[50]},
      {stage1_5[26]}
   );
   gpc1_1 gpc66 (
      {stage0_5[51]},
      {stage1_5[27]}
   );
   gpc1_1 gpc67 (
      {stage0_5[52]},
      {stage1_5[28]}
   );
   gpc1_1 gpc68 (
      {stage0_5[53]},
      {stage1_5[29]}
   );
   gpc1_1 gpc69 (
      {stage0_6[53]},
      {stage1_6[18]}
   );
   gpc1_1 gpc70 (
      {stage0_10[52]},
      {stage1_10[18]}
   );
   gpc1_1 gpc71 (
      {stage0_10[53]},
      {stage1_10[19]}
   );
   gpc1_1 gpc72 (
      {stage0_11[47]},
      {stage1_11[18]}
   );
   gpc1_1 gpc73 (
      {stage0_11[48]},
      {stage1_11[19]}
   );
   gpc1_1 gpc74 (
      {stage0_11[49]},
      {stage1_11[20]}
   );
   gpc1_1 gpc75 (
      {stage0_11[50]},
      {stage1_11[21]}
   );
   gpc1_1 gpc76 (
      {stage0_11[51]},
      {stage1_11[22]}
   );
   gpc1_1 gpc77 (
      {stage0_11[52]},
      {stage1_11[23]}
   );
   gpc1_1 gpc78 (
      {stage0_11[53]},
      {stage1_11[24]}
   );
   gpc2135_5 gpc79 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc80 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc81 (
      {stage1_0[10], stage1_0[11], stage1_0[12]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[2]},
      {stage1_3[4]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc615_5 gpc82 (
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7]},
      {stage1_3[5]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[3],stage2_3[3],stage2_2[3]}
   );
   gpc615_5 gpc83 (
      {stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage1_3[6]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc615_5 gpc84 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_3[7]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc85 (
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage1_4[18]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[3],stage2_5[3],stage2_4[6],stage2_3[6]}
   );
   gpc615_5 gpc86 (
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage1_4[19]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[4],stage2_5[4],stage2_4[7],stage2_3[7]}
   );
   gpc1163_5 gpc87 (
      {stage1_4[20], stage1_4[21], stage1_4[22]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[2],stage2_6[5],stage2_5[5],stage2_4[8]}
   );
   gpc606_5 gpc88 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6]},
      {stage2_9[0],stage2_8[1],stage2_7[3],stage2_6[6],stage2_5[6]}
   );
   gpc606_5 gpc89 (
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage2_9[1],stage2_8[2],stage2_7[4],stage2_6[7],stage2_5[7]}
   );
   gpc606_5 gpc90 (
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[2],stage2_8[3],stage2_7[5],stage2_6[8]}
   );
   gpc615_5 gpc91 (
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage1_7[13]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[3],stage2_8[4],stage2_7[6],stage2_6[9]}
   );
   gpc615_5 gpc92 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[14]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[4],stage2_8[5],stage2_7[7],stage2_6[10]}
   );
   gpc1163_5 gpc93 (
      {stage1_8[18], stage1_8[19], stage1_8[20]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_10[0]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[0],stage2_10[3],stage2_9[5],stage2_8[6]}
   );
   gpc606_5 gpc94 (
      {stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26]},
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage2_12[1],stage2_11[1],stage2_10[4],stage2_9[6],stage2_8[7]}
   );
   gpc606_5 gpc95 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6]},
      {stage2_13[0],stage2_12[2],stage2_11[2],stage2_10[5],stage2_9[7]}
   );
   gpc606_5 gpc96 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12]},
      {stage2_13[1],stage2_12[3],stage2_11[3],stage2_10[6],stage2_9[8]}
   );
   gpc606_5 gpc97 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage2_13[2],stage2_12[4],stage2_11[4],stage2_10[7],stage2_9[9]}
   );
   gpc606_5 gpc98 (
      {stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[3],stage2_12[5],stage2_11[5],stage2_10[8]}
   );
   gpc606_5 gpc99 (
      {stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[4],stage2_12[6],stage2_11[6],stage2_10[9]}
   );
   gpc606_5 gpc100 (
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[2],stage2_13[5],stage2_12[7],stage2_11[7]}
   );
   gpc1_1 gpc101 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc102 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc103 (
      {stage1_0[15]},
      {stage2_0[5]}
   );
   gpc1_1 gpc104 (
      {stage1_0[16]},
      {stage2_0[6]}
   );
   gpc1_1 gpc105 (
      {stage1_0[17]},
      {stage2_0[7]}
   );
   gpc1_1 gpc106 (
      {stage1_1[12]},
      {stage2_1[3]}
   );
   gpc1_1 gpc107 (
      {stage1_1[13]},
      {stage2_1[4]}
   );
   gpc1_1 gpc108 (
      {stage1_1[14]},
      {stage2_1[5]}
   );
   gpc1_1 gpc109 (
      {stage1_1[15]},
      {stage2_1[6]}
   );
   gpc1_1 gpc110 (
      {stage1_1[16]},
      {stage2_1[7]}
   );
   gpc1_1 gpc111 (
      {stage1_1[17]},
      {stage2_1[8]}
   );
   gpc1_1 gpc112 (
      {stage1_4[23]},
      {stage2_4[9]}
   );
   gpc1_1 gpc113 (
      {stage1_4[24]},
      {stage2_4[10]}
   );
   gpc1_1 gpc114 (
      {stage1_4[25]},
      {stage2_4[11]}
   );
   gpc1_1 gpc115 (
      {stage1_6[17]},
      {stage2_6[11]}
   );
   gpc1_1 gpc116 (
      {stage1_6[18]},
      {stage2_6[12]}
   );
   gpc1_1 gpc117 (
      {stage1_7[15]},
      {stage2_7[8]}
   );
   gpc1_1 gpc118 (
      {stage1_7[16]},
      {stage2_7[9]}
   );
   gpc1_1 gpc119 (
      {stage1_7[17]},
      {stage2_7[10]}
   );
   gpc1_1 gpc120 (
      {stage1_9[24]},
      {stage2_9[10]}
   );
   gpc1_1 gpc121 (
      {stage1_9[25]},
      {stage2_9[11]}
   );
   gpc1_1 gpc122 (
      {stage1_10[19]},
      {stage2_10[10]}
   );
   gpc1_1 gpc123 (
      {stage1_12[12]},
      {stage2_12[8]}
   );
   gpc1_1 gpc124 (
      {stage1_12[13]},
      {stage2_12[9]}
   );
   gpc1_1 gpc125 (
      {stage1_12[14]},
      {stage2_12[10]}
   );
   gpc1_1 gpc126 (
      {stage1_12[15]},
      {stage2_12[11]}
   );
   gpc1_1 gpc127 (
      {stage1_12[16]},
      {stage2_12[12]}
   );
   gpc1_1 gpc128 (
      {stage1_13[6]},
      {stage2_13[6]}
   );
   gpc2135_5 gpc129 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage2_3[0], stage2_3[1]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc130 (
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[1]}
   );
   gpc615_5 gpc131 (
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4]},
      {stage2_5[6]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[2]}
   );
   gpc615_5 gpc132 (
      {stage2_4[5], stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9]},
      {stage2_5[7]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[2],stage3_6[2],stage3_5[2],stage3_4[3]}
   );
   gpc615_5 gpc133 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[3]}
   );
   gpc615_5 gpc134 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[4]}
   );
   gpc606_5 gpc135 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[2],stage3_9[2],stage3_8[4]}
   );
   gpc615_5 gpc136 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10]},
      {stage2_11[0]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[1],stage3_11[3],stage3_10[3]}
   );
   gpc606_5 gpc137 (
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[1],stage3_12[2],stage3_11[4]}
   );
   gpc1325_5 gpc138 (
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10]},
      {stage2_13[6], 1'b0},
      {stage2_14[0], stage2_14[1], stage2_14[2]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[1],stage3_14[2],stage3_13[2],stage3_12[3]}
   );
   gpc1_1 gpc139 (
      {stage2_0[5]},
      {stage3_0[1]}
   );
   gpc1_1 gpc140 (
      {stage2_0[6]},
      {stage3_0[2]}
   );
   gpc1_1 gpc141 (
      {stage2_0[7]},
      {stage3_0[3]}
   );
   gpc1_1 gpc142 (
      {stage2_1[3]},
      {stage3_1[1]}
   );
   gpc1_1 gpc143 (
      {stage2_1[4]},
      {stage3_1[2]}
   );
   gpc1_1 gpc144 (
      {stage2_1[5]},
      {stage3_1[3]}
   );
   gpc1_1 gpc145 (
      {stage2_1[6]},
      {stage3_1[4]}
   );
   gpc1_1 gpc146 (
      {stage2_1[7]},
      {stage3_1[5]}
   );
   gpc1_1 gpc147 (
      {stage2_1[8]},
      {stage3_1[6]}
   );
   gpc1_1 gpc148 (
      {stage2_2[1]},
      {stage3_2[1]}
   );
   gpc1_1 gpc149 (
      {stage2_2[2]},
      {stage3_2[2]}
   );
   gpc1_1 gpc150 (
      {stage2_2[3]},
      {stage3_2[3]}
   );
   gpc1_1 gpc151 (
      {stage2_2[4]},
      {stage3_2[4]}
   );
   gpc1_1 gpc152 (
      {stage2_2[5]},
      {stage3_2[5]}
   );
   gpc1_1 gpc153 (
      {stage2_4[10]},
      {stage3_4[4]}
   );
   gpc1_1 gpc154 (
      {stage2_4[11]},
      {stage3_4[5]}
   );
   gpc1_1 gpc155 (
      {stage2_6[12]},
      {stage3_6[3]}
   );
   gpc1_1 gpc156 (
      {stage2_7[10]},
      {stage3_7[5]}
   );
   gpc1_1 gpc157 (
      {stage2_11[7]},
      {stage3_11[5]}
   );
   gpc1_1 gpc158 (
      {stage2_12[11]},
      {stage3_12[4]}
   );
   gpc1_1 gpc159 (
      {stage2_12[12]},
      {stage3_12[5]}
   );
   gpc1163_5 gpc160 (
      {stage3_0[0], stage3_0[1], stage3_0[2]},
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_2[0]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc161 (
      {stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage3_3[1]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc1343_5 gpc162 (
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[0], stage3_7[1], stage3_7[2]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[1]}
   );
   gpc1343_5 gpc163 (
      {stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc164 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc165 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], stage3_14[2]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc1_1 gpc166 (
      {stage3_0[3]},
      {stage4_0[1]}
   );
   gpc1_1 gpc167 (
      {stage3_1[6]},
      {stage4_1[1]}
   );
   gpc1_1 gpc168 (
      {stage3_15[1]},
      {stage4_15[1]}
   );
   gpc1_1 gpc169 (
      {stage3_16[0]},
      {stage4_16[1]}
   );
endmodule

module testbench();
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor_CLA54_12 compressor_CLA54_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h7d45632c2ad67d26a6db68fa5eae6aea5718385439e36f9c661a568818b27bd765bdf7a92c0de006b384825f5305ffb65554562a27ad86a26ab39a3d8c79527a5cc2315648ddc057c2582a5dca7dd6863e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'he9fb8f7bfedee90e8a1cd98a51d93f9a1a58fb8b82a285d827fa0ef5c1c34c98eeaf597b166259d5ad3ce70049b2762c9a605abf4f27383fe2805a836b5cae6c7a61178b0c3f21956f3ab8ab5fbd6190f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h8d0a1f92f7cc03db0c0e695884ed4f77c48d7986f7286788d4b4a71a22ebdeb894f64d08bd66fb56d00df769a07c94df78ade6616dd6fa2ec078d45ab130b6594ea096baed7e89f4bc2a7fc42775b10f01;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hf41fe9d5333c8bf95d95266aeb346641d0ac9b7a18d134ee693856a9fe0c387f584c70bead468eeadd4f231b06be76800bc9d844d42536f7b2f9a5e4b6d4acf7c4009fbda3595d41385b99b127fae81326;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h69f7bcb5994693cf8d243e97002dce4fb82c4d1429c42db285027599b81bc7c6598c9a0c4b12935c1ee06988d5e4fc7fa2694391e9d63864f5dd1d6e32767570d8c16c4e154ae451cd483d1bdc31e1921a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hcfb03aff5a05ea3a5dceea991696e6bfeded04b409fe03c797293122a953174deb98c78889867060e97ab02947abe704733eff0239707e52426b50d43537ed6688139ad10e08fcb7b11b4413a9598ff12c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h97d9f042890fd1276536f957afdf05050a109a44228b3d485543a4c02e7ce52b7d02b057030a8f51a9af4e9e4108d5718cbd7579e1456fc67b00040a03f83edbac7272f93f9b6fffcbf8a94db81f573a73;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'he931bf23a9a80d7c1c11b31954903d79299f710932f3ce0111baf080df5e828ea6dfa68f8b7d895c9a9b44f9c13c7abf7e16a526e201ee44282881b08bdc530c48bdcef0e8060a844bf09758cbba2c37b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hca305ae11cb2e4dee83185adb6b921968cdab061a9cc00fb9856a9a5c922e7e06b573f239f1b5bd2d78be4e1078d401b6a21facf94954e97d33980efdd94fa715de68e235f77f44e29db5817b0fe413a9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'ha747e9e8215d1b46639850eb83cab4f7cfc8a1ceb189a37ee6e6045ddc226d2033870da8563e9ea98395da4d30ee3f41f6521157f15b6cd4d0a0874cfb1af1d9303e5b7180d066fb8a0adf2fa7056e7528;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hda5192defb5eeca947eb7134534c57e25186c8a85c6e651d0024b003e87764e1a9b9a4d765030da9d463bc419ca253404e13c6bae80daf0048fc9536b089fc29ea8a96c127053247bf6580febb5aec688f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hcd4bace65b84feac78be5372402843d5dcac9a2c3a35bec9c4f31da0444a897e3ef622039fb26f050b364771b704e9f18c3b8677b8fb55a812025ed4b2f15f1a508fd94c7f7b9074905f710becf1520f22;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'ha00353c8bcec643b46fe905ab7f074272d8efb28179c809f64bb3e72e516814ee83a84ae04f2fb8af69ee051085aa7d01c075acf472e20f7c3696fdb015ce1b4bef1eddcc75a9426417e3ee56011dfff17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'heabed49f160df8325e19bcb5a1a10c2bcb6b0477922f205dad08adc9ad163d857fa8df0a1e34e4fff7368d8a57ce64608f4f9b9f80ac406a2bd5b4abc6d4af7e81941de7c6955d8d8f505e105d4390387b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h3ff855d775c941217fed3eb0094c07390e04ada54c84e2fc7dabcd8b5ae81cc3cf0b185f45dcdac2a731d830014752fb9125eb592407b2ffb3b71575dd51554039392410c6135c85e9c21936d0d9eadbfc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h1a9bbdab20073c6865c063d6c103f5a9a299ed9a5ee71aeed4238037d568ad11a500572afe9d3b551646b9bf42fa747d073cbba80e8bf3d9bc8b0b78494599672f636f26408e68df11767e43d59339c239;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h2e01f6b0ac8b6ac3d89052c928036217f08f90148ef77443780a54b82dadb68eaef5a8603694d7cfa153e893ebcd6ae800cffd692b6c6894d808619472c95428b35956ea26e1fdac92c26cb6869cb8d113;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9f428820fcccfcccf46bd19ae540b865a3d8addd52919a013314fde630e244aa1f7d76b9c726773bd2663cdd6efc1c4217bc3b50885bc69d373f1c0f134bc8aa30e475d011376abe0f47955e6da07685ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h51025b2598ff0d67b62120c5bddc43057c8021fda6094f29ab1f95cc2b99ff1719fa7f23af1f602f381786c40b18b3f0d1fc2b5e3b4ca9e08e14191917109f6d4cfe235392c1931a62b3bbf1d8b535f236;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h896ce5bd2977d6b433f9b1e3134c3410d68d1302374f01bda1d4cf3f795c61443f6c4da03927672caaadc67b15fa43218b8d67b105a65a32527df3563ae7b7f38ed03b837ffffbd7100de84bcf5f7f2ba4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h5a3d7de5af77ef075a8d9bf6fd9e8d9d97732e70b9a22584c1807124d8baac192440c524bbd01b62b79933639b24efe90086cd1c3ab9212bd08eadff8fe732de269ba6a11760dab299ab5bea3299132f7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hed206e0c64727fe1f634b98c122e3eb27c6c4a172ebf1b6e5ec262a595980a35703beaf3195972c1593bf3c5a18c792080baba10c2fbc10679df59517ae273e4d0ae7831e7a55d76426600a7e98407e63a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'he4940b24e26d758c19f52df2a0cc4ebea9109147b67ecd3ecad0ddc30e564c1fae2b08e2bf9fb8e76609df973823b199bad9839efeed7193848f2cc577df7c6a51d58f0dd57fa2a46a0479bf3eb99d27f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h6cafee894d8f82765696ce1932ebe086ae0a0fde7cf0d0d0914c4526884fcc45522aef1df9c20cc089ca969aa113240d894bed9540b79fdd18b47556e565ed7f1ca18f7a442b2115d0e2073a86b517f17a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h7834c4f2320a8fded8d857b4caac120fafc81792d64416edead863b5df500956f97fae4eeab77efd8d18818f23edbcb244916a40411b0a05bc0cceea0cd925c38f716d4a48bd782ca77d3d71094eabe8e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb275116400b44961c042c484be8a8749743b158354c51ca66a586e382899bad5e8180ce9d3eec379873d4e2341ea7f53685d9511e8006b5bd1ee471d86929b209aa09b657d693f60ab02807f6b7e969ef6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hd27e7188e1f5f9f85a0e2beddfaba696fe7f2644c7ddb2887da892569908c03b15313d82173a3cac6490446b7a0d6472581ac258af43485dab7458cb8f5229ce7a49d30a7cead188bf50941dda8f778cdb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hfb7a679e40ab2477837826a6792d8ffb8d9aa8f9afeeee27578051fe645e5c5a63ff7dd87212c313076234556327038ddd659f71336358c087efca9da493a26686bd3439f2e34448f3d5df70a6dc2bf5c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hc5f604999d03cb05d3c92bcaa68eedb5d71bbba7a356b3609b6d933ed15ccfad52d2ec2e2d19aeb9831bdb2fe93eef579515ff8f5de49441e20b1cf349f4e83a49dab6ee35d2b6858adb3d8b5fa1e9727a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h6fa0197f7b7ce5422076e0db67e8a87c9221825f06fd2c41e7f78221cfde438996200839c5d952d9fc1ad72888de6366ed626952fd9e3df6d717774bd7aab963d1a5bcf601166e4821599cbc33c060b8c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h111ae2c1b81feff424efd2fcccef47bf26c3c491f6002e0384c09f2c36f65047a0df38792a893ef43fbe9fa8b99e3f04e4919316f30a9487b920f2e23ca0346e04b0c176f60dfce7fd19354d7afa206cc2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hfca7ed60812bd64ba329a8276a104997332dbce8d9ef33a2ebdc86b5bcd798e2ad581567b8e1626172d5279fefb544626879f0746628c2bf6af341e0481c7b28af2afcd4fc79b24a7e4536d79adaf2763f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h2067d0b12c0855fe0d5dd9c3e04bce403878f4aaac5c1de5da0423e18d16e560eaa0ded5b03d74672ec9c248732ee5a07447d4b8cd4cfb6ccc52c210f9086303f322e543832ba1d76733d3a147f97dd254;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hbfb379d9ed28fd3515416367b60332bcc7badf380f20bb2ad2db8dfbf9d86b20c72f52bf2575ca4c688eb458593378c43ce1abbb57d518efd980940f6a99b34baa144e87ec11d6a8080edec7efe2e30a00;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h236ea9e2a766a486db5c2a4f1d207e9640016631d4e553448c71203c9a7c05fa913bf88653b614697323f9aaf7015530040d3faa4b89c10d9059c378fb49fb4d558cf2be3dcaf45fdf0f9150ce7753c929;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hdd6a90bb952c0710272ccc39011939401dcf29ddd05b1992ad685110a56f3c9976a045186c8736ccb105a04806960bd8e1c2b642fcabbf68f87b3e8dab1786e412e386f34fd1007c60af3e27f1de3a7816;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hcedcdc50f66c1e3153169beb14660d6500e9936f38fd57cdb2b7bd26ed1f02e81b87e8d5e2b803af82e9713df3e016b31026b1f3a7e2565ad4079cdd8d5fe27294b67c759259af3fd4eeaac527b1f90ece;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hd20e8a695a261be177bb6d288d9423b7d0a4bf1ff0485c6796509cd17ffed6340ec5a14fb5af36c66e5dcda3c03918104d436e9ca4c8ac65b7e0379b2b9afde5c6ba1e386f5644337e42d86ef3874266a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h275d7f6e88782ec7d28acaa3d594e70475fd3cbff6e199c49317989dd7cded88781fa5ae7292f635ccd29f1f8959e887a75d719c0b017d0dc180f1bbff91a587bc7902ac3c7715767509607ff290bde048;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h5ecc9858994b04b7d9f28322c1dacb295cfcfbb5d9b15a3fc29e4b4cefbc5ccd93ded5942a22966b7d95bf4e16ce4af0f45883e19f82856f92a9b07e3c53752ae4f441ec919ab6890646c4fed3b4de2848;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb6b9f6d096a5feaa5ff6b1a059f43fa6205d43e3f64e9875c47eceb5b4d2972c8cd7f4c3506666483af1303bdb6416ca71ff174553e77904061ec982116edf1b9a118ff1b41bc6c301c7b60ac826e7353a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hd320a227cd577d50b9752767597df82a0cd4d65ba036c1f39a5aed3812ef2d462d7dcce143bd7548cb5d2c08f7e375d9c401bb1649371d7f7dc6efb8a7d92ed281f3aad5b37827233fa93fc422872d30c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hae0375da763849377dcd427f858a5e08e8a5a298e4de6ed7e79a2bdf1e43713227d8d7a909bf2b70d95a7f54bb61fdd14f2e18b44be9ec0cdde655cc38fd8de79db1c56dbbaf1e494e054d4f6a174defbc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9c8a125cc678ce0868186055db5855ad43973876ebc0077a1ae52b93d84b0010f7f4bf02cc7ee4e14df377b6c32ca69c3efa2f2afd9fc97da3bc8a38692a449b5d88de1c1bbaa675d6d440f5fc1ce3e4fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h1f3b7195b5dc968d18ccf57aeef680b3b966f7f417c5fe99a0528e14811263c0653eec765875cbf0fdf7b53ef2f26478588f2266caa5fddb4367bd99320e432afd83c35043448be67dadb136c5ba4acd38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h5c6ddf91441b592c7f43689d7765c3caf0bca24a775a827badb81cba68b4b211628b26d74b68243b7c6d5f8096246791d0ff14925b63c0ccaccf64b58e6199b2f6f8db593ce86a77499028af3f67c97d60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hd5a1cb6cfbff165c6c79ae20d807f3746a354ad6aa8750803c55053537f3e3b8ea7ebd6a88ee81039c020fa3b54b4e717e9a844a6a21cdcce5dc99d99a1b4a0fd353a48b4fa5469c40074c2e9bd26452e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h7e6b19c34856f751e8d5519bb196230adea9b22e11f7f2475fc4d0870f4b54fa065b96b44887afbad0f7f3b9b7cae9bc5f37ffb9b8e614ab780c6c81746864dfc8f0e022ceb2b834d56bafdd72e5d8ac73;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hea65be6a2aa6ec5808204fc468ee8b30a24d92846076c531b12935e47e649c39b6ad89272c3da79f692a28b5344ce8dcd96525c574e8965a7cbf28035926f07f056490044b0653607a196fdb49a6bd2c9a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hdbf42be735a3b5a40dcab7c088c4eff6986e52856724e68cc0e5b650a40d2cdde675a86b25db0db7af15ff84ea3ddb8e6386a79950d3918b39ed9b3969354dfc8a9c6c8bf1e90f399f66bcd26d33cca462;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h456d8290598b776b8020cb1386b271c3a05d663c983e3601999c4169d6fc59369c4c2598d3452dc72c9b2204b2aabbc2c804c731f91857b074da2f0a6abecd0f149fa47590f8aa130778fdea165af713a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hc7f8e51f9ee1e1b276e5652369b49931842ecc5b438b956b3b6918c2383157d4953eecc2cf378b1b7aa8042949c05d68b604a518c4b9bc0be48320d3bcf0fe1ed413fcf891d8943b4fa9da29b09cde9829;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h3f670b5ee18c594dd90ec2399e0c73ba196277c4724f7129718336c5fa3aa5491c222245a73d9a5d1a8cabf79460a3b8291f590a24f3808b352aa163c4e64d087bf58b181ecb990a1b20b4f557a057b3fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h180763bb045023e3d6b0f276cc3923d2828a3e26a70fe77e5f4906f2689f026f23b472f5b88d3a1f1e9d343521fd34044d2882833c9ca41d989f2207d7c795185fcba333f7a8e1fece05dab7a3db086bd8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h87750bf981ac8490c94b9d7eb6f084f24017fd9f04fde1c257e5933467a15e6c8527ab43143058dd4f96ec8e9398f41399bae0165cb063d34fff466c1cb8846a5b62029461c0d5070636f2000d50180f3c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h59ce85c527dbf298a5e408a9503b956f3bbd82fb94a6a574dbe512395bdd826b385222a4017c74f6a59599dfdfbdf8c3d922b28976bb5130acc40277e6cb0bc0cfa370466e8830ff0f760d8b404dd69536;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb3f31e64dcff9797a94a47ec0cd51b1d6eb5e98b75628fac27a326acf36291120d498e099c83201df6f0268f796f8efee61f303461e7bf7642c1614ad6317766a5ec9cc0a60e6ec8a18ce7b740e75dc29f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h4eb0ed8de3dd73a7bf192468e9e0c3a075618b4ea01d4023dfebd2bc33ad0eac74b565d964c39afaf331da8b042d3f9a10dab0c0bf41e5c8e31a33a98dfd8b0d66d8b1e36e11f9567b13608e14c8c25a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hab1d733119e46ec8894ff654d5473de437879ad668a87532fd53bbcb3bed9f48f738794dd2706e41818bde670db6468bdd9b0f8bd974ba3581c35c6f67f3cfc74814e93e61faf71ae8cd10bf135f5bae17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h11e2c68c7b2b75f772de9d9513faccbf0efed3d92e5780aceb6860a07d18da8b2e7d2ac0d98a74c327a38db041df4fd3b13979ef6549ef004f15846d81a695915b2f2b3c4202043fecddddfb6883df1cac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hc6c775a29182de5cfcadef3e62ed025bd8dd5fc545b54bbf8d9a67848fc0d4955a951714204f2c697d31679f01054ae1cc6f8d358d7a3c546c43dac32f98c49b227d198db605b6bc252916aef93f798ec5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h36b64abe1fd94c57750c49e988138956724cf19cd2185fd253b5d0849c788f80445d59ced70089f1f00383545c6612b12c36e456fc52b14188617770ab512bc5eed3a1f8bd3708920aab838bca5b4861e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hbf2f57ac3a09e98f9404133ef04a3876fe073edfca6c964139a0d1ffc2ac0d24d9a6c4e509997b8320ec69aaadf3ba1a41b1a196fd9465619c457e6dedbba00c98d85339e08a7aebb445c2ef6165d961da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9d6a94c20b6313458d3d7f826530cf94f728e701ac2b1e7a03a0571d6d541e092939d776163295b6bcd075280f116ba9bef57c33db4b366c83ad9a1b90059ab141403c42a047d406f8641f4a3c2c0b912b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hf2c69300c48366d83d12802826ac6805fc2d5c599cbeb03460f90b75112da7f1c734785cfcac5b489a7637583dc412193d9d7a4e01acfdd053457f4557ae67a1849a1f76a060c87ffd3bc337423e02413b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hd637cd57d6a39ec8d4d723e9b470ea9d93c2a575e101a75eea36d889f69ef1438937be11bc70359dcb02d4880bf6010d99fe24c0a02ca16623df68ee7b8e9a1d06b074c5e5416ac4b09998470106adbfe1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9ac54184b014abbea196a1c3c487e16457bb756d6392944c3f67170b219740a8371a48248f333434dea55e35e39298bdc613870a1d98106348df33a6476a06c5590f9f98d975ed5eeb6398d416a77391dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h678d5375e99a0f117f2e0219f13dd76e0668706b58593aabfa6bae5051366d8b4a2466f2e81956de2142b998286ebdc5c80ac88c148e6860a5a522ae162a80b4f082a986d32239519f643d166f1974d416;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h1f3384f2115d40896587d37d31fda16b9a4cda1039580038a88f1f900baa57b2b1da860a83d7f2ac4672561b248df431767cbd1a035e2f9246ce00786efd998fa53078b49bfe6803b206ffa7d0d33e3d1c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h19bc6d055c03a3145ada18eb1ab742fef93da6e9a2bd330159c52d4e81c863f556653b274d4c527ca443759003de2d68e3ca434afc887ad5cbdf4db282f0a6d3e7369544869d820e79cfa85b5143c3c76f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h152e0f98f40d3ac1250713607ba9c7f9455244ec4c72dd080871546c45cbd1c99d1e67f7609101d825d66a1257f8937a92ff32ac8375f711f886ea70a37ee5d7540938a5c6473f1061fab6ff6d98813719;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hcf7d9af750b72bdc49b0c804f7eb194ca419e3b0b0884d04a5bf223f5a2484f6aa0eadcc2c4cc806cf3244cebbf7674bad5d4cedcac8261ec4690225e9762337b3605cdb359fa16b4e2f54fa3efffed843;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h15938fe53d8520bcbefa5d71a50f89ae406b02b699350240d7d245a571be87f771066223bbcc3a0e783dcd41738ab7978e92c055563565da904c591d5a0009fda57991cf28cffbc690ceb99adf576e0d78;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h96c8c19a6dd055ef9836d68f3b8dab98e8d05f30061ee9eaa703785605ba6824791dc3bddb09eff989d8f56dbb6803d47e6940b455131007510afa7ac53c22d108cb70f1572d1f5334d93f0d580a04a8be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h62691c9c4056ba91955548a29e7d41fa76c3cd6fd59470324e301573beff5c12d9860f777e989edf294c09276212745cb78e21d2c433b552c2daff1587b5c5680207c8673298e022d52ba34f125df2c8cf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hfcb9d0bf0614f706f26a8e3cf4ca0f76bef2f38d869f9fd878d96da9388009a8ecf826a06d818aa53661608066b1b2a09387b66990a0be341df1f0c0a43c1afbad2da8b7efb0b0fce2e3426b205ade9e73;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h65e3b44a54a420dcc674814eb36eb7e533860b19cbc93af6ed36290cea1caa1badf50a3c9d06890e075ad6def08429094c8b1fd105575cb1114e8fd30554b39d18a43acfca0bbacaf27dca1f2341fba618;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h1da4beb32e1bc15ac585091a9a68e32de9f6e00df0ef3b43116f7aa20d2eaffdc6ae6df4263e820c7100c297eea5a40b4af63c8ec225aef35b8aee524ab986d4a446b1af7249985916159a28d2743098f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9edc7e18024b9682c25344bdcc8978bc925a8f7c0a78cc173f678384857941d131868468acc47abcb1ff3d15058e9cd21e37a1723a8b30fd1cddb1a39d9e262ec610c399be57a3e0967a8bf29e6d9b1c4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'he17133dd392dbcd94a5606b27fbb08f29261235ac9f27189da8c863eff5af12273cf0b86af001b8c998b9eface7ff2d56467f63f1959b248cd870a14386f078f2d4276457a4bdfa8724bf9404a12d867ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'ha9ac0bfa4f8ae0abd6267736ec88708ad2365c8a3dbb995c0f2c656926e80f666d8e0b538715532bc1783721333575dd85372e1cd956247f17fa3de9f9d418290e1ed3ccbf7bdb4c23567614c204cf3379;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h1407fbdfdeee8f7a5c39cec7836af45cadff0d66dd19c1138db5d55122c90ca90fc9f2baccf7a8399ff51fc548f297f13f2d83299ba766fb73da22ac6485f6f6777d5a32fede556b2fc9779f0fbb93544c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h68a367d3f097911c49f0306f9e7372895edab7ec140e147603ee3fcae88c6b20177095b1480455be4be53108c193aaf8c32008b661bae14caa32fbad36261ae776834bd4217f5112142222064dea007173;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9782aaa87be7c2a8d2a2e8c3c0ea29b1b033c1125836ee69bb07fbb21047dc643de787ed809c52272d833cb2c7fad04f2d206d60bc64cec2b81b81bd6e4239a7df969b8f0d2b5f5901de7dec7dee8e87e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h5e0395b3044d997a4c6f7ee515fc78e11a6c562f1c6cced7c8fe0cad74fb6583bb00c1ce0d1c054f58454f7d5e66c44450889fc59ccb325712b4cba5a6d8cacddf3a5def01afb9e2a0c5395e2601f079be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hfc9f73253dbb8d1d345c43aaf227dea6453a26b60e3ae99897d27eabbca8ab49b476baab86026759433ebc8859a83e04409cc8a1bc6756cf411cb236d51d39d457e47db935032edb6153267f88c46de2ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9f963d209ad18ce4dffbcc7660b3e36f4c4159c542f3a85e0c9452ee09114b49236ae041416a230682b8bd9a7e8f7750f0d3630d3ec8f7286373065512950cce32dce3493d47da742b62435f5e5cf06345;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h4db176c2a6bd0acd469cc220205b5b8ca821a1bbf0513fea27f58c5af40d1c516153f58825eac2998be09d197f12cf365295272ccf7a0e9efae26824a891532d0558901c2e8ff534e9b12aa583e374a55c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'ha801066e7045d655f9710802c6cea9c58a5a2fb23c39539a9195da14be5daa348793ebf70fba57f4edebb7dee6d8cbabf8aa47c7a08c1395b0b23ea222cbbcf933b433e6e0269a7073fe571b4b3ed0eba5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hed8e1d2ddac88d2fd3ecaba7d36d4ebf90ca8c157a5da643837019ca0e28d21a49f1379356d9afe52b90393e7b9ca14f6c7f12ca7cb2530c15290d77d04ec0b6c743f7832236ec7c41e213ccf05573593a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h713b7debcc1efc88d035604a2e40c83cfde1ecbff241126e944a01cc7bc9b17983f368509045d5001fb8f8d2729ce104e2bbdf3aa49f96a8139dfe16cc820b45d81a0a351be4a530cf0daf7b488f183bf5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hda6822172f2b74abeb9256094466635e5806162d33524f19d9162fa288f533ffbe0a5eec030e5b7c5738348bcfbe4491627947d49f1614547681d5b0bc4a1f9e56fd25ec6f8ee2cb43bfaff28ab8890094;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h1bc8e399707cab35d5460aab46d8a4bcad6aa93e7c35b190d6517f0fbb6a5b8319b242c73e90ed6606e1cf30a26813560d7b923a58b2c39f522bce9d41c4932efc0fdf0c9b0556182fa9ff19523c9a63e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'he6cd60406cb57bd180de02cb665eb2fe338afea5c832df64c14e963398928410c7cf5e60f0f23902f540cda0f9df8683f5146c45b007d38cb4095d0e784ae71b61ba87efedd7224cdf8572f16add161c2d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h6807f475fbce643774e229b23c3c84100cd0e2f3f63bf10b9458b527a8978a36977192deea12f719b1cf7d7e2dfdb93d99fd4e1cef92a3354f834062710640c50c52186bd4eeeca57f380de2a10bab4d48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h156b2a6cadc1ff5039285a957a2638d5aafa1cace3c1414ed3d81804d998416c97c21cb739c627ce984a8ca0c57a6262cdd1986e9f0b3578ec390c7feb56fd960e5e9cb475bab75aedecd218f002edf1ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h78d06d36f2f76a75c857a97365c548f28af0ab51feda20db612af4f621096ac6269922294aa4eb5e92030c25bbf28aa18a28bce1cd7824c91224665a2a6cbd1808fe5b42249fa4122c1359fdbe1c41778;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h2a5487c19420dbbd0d7599bae14e3a469803e6068f1848fb5647cd26eae9dede7bd225aa5c93ee006d3d90b75f94916e31353efab94c2c887eec5ae83742a11a4c951be9ebd82624a0a93862f75ba4408e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h4fb11be1289a76b8a450c857701518af93947913ca54ce891c4a315d3350e285e154b9761767943a7afa18a30a329331cb59c598075ca79fed0c8a7cb9e0edcd3b8a364913665ea1bf3b33bc8f17a27344;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h143a807e1ef12c1bcb11dd1a2e69dd0789ae3a7204d2d7883623c8b46adae0c51884387d59c7a8915152b72ffa11f224351eada2eabd414b495430f8241f72bbf05c4c5afabae8913083811f883de1db68;
        #1
        $finish();
    end
endmodule
