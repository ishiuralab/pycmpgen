module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69);
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    reg [63:0] src16;
    reg [63:0] src17;
    reg [63:0] src18;
    reg [63:0] src19;
    reg [63:0] src20;
    reg [63:0] src21;
    reg [63:0] src22;
    reg [63:0] src23;
    reg [63:0] src24;
    reg [63:0] src25;
    reg [63:0] src26;
    reg [63:0] src27;
    reg [63:0] src28;
    reg [63:0] src29;
    reg [63:0] src30;
    reg [63:0] src31;
    reg [63:0] src32;
    reg [63:0] src33;
    reg [63:0] src34;
    reg [63:0] src35;
    reg [63:0] src36;
    reg [63:0] src37;
    reg [63:0] src38;
    reg [63:0] src39;
    reg [63:0] src40;
    reg [63:0] src41;
    reg [63:0] src42;
    reg [63:0] src43;
    reg [63:0] src44;
    reg [63:0] src45;
    reg [63:0] src46;
    reg [63:0] src47;
    reg [63:0] src48;
    reg [63:0] src49;
    reg [63:0] src50;
    reg [63:0] src51;
    reg [63:0] src52;
    reg [63:0] src53;
    reg [63:0] src54;
    reg [63:0] src55;
    reg [63:0] src56;
    reg [63:0] src57;
    reg [63:0] src58;
    reg [63:0] src59;
    reg [63:0] src60;
    reg [63:0] src61;
    reg [63:0] src62;
    reg [63:0] src63;
    compressor2_1_64_64 compressor2_1_64_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69));
    initial begin
        src0 <= 64'h0;
        src1 <= 64'h0;
        src2 <= 64'h0;
        src3 <= 64'h0;
        src4 <= 64'h0;
        src5 <= 64'h0;
        src6 <= 64'h0;
        src7 <= 64'h0;
        src8 <= 64'h0;
        src9 <= 64'h0;
        src10 <= 64'h0;
        src11 <= 64'h0;
        src12 <= 64'h0;
        src13 <= 64'h0;
        src14 <= 64'h0;
        src15 <= 64'h0;
        src16 <= 64'h0;
        src17 <= 64'h0;
        src18 <= 64'h0;
        src19 <= 64'h0;
        src20 <= 64'h0;
        src21 <= 64'h0;
        src22 <= 64'h0;
        src23 <= 64'h0;
        src24 <= 64'h0;
        src25 <= 64'h0;
        src26 <= 64'h0;
        src27 <= 64'h0;
        src28 <= 64'h0;
        src29 <= 64'h0;
        src30 <= 64'h0;
        src31 <= 64'h0;
        src32 <= 64'h0;
        src33 <= 64'h0;
        src34 <= 64'h0;
        src35 <= 64'h0;
        src36 <= 64'h0;
        src37 <= 64'h0;
        src38 <= 64'h0;
        src39 <= 64'h0;
        src40 <= 64'h0;
        src41 <= 64'h0;
        src42 <= 64'h0;
        src43 <= 64'h0;
        src44 <= 64'h0;
        src45 <= 64'h0;
        src46 <= 64'h0;
        src47 <= 64'h0;
        src48 <= 64'h0;
        src49 <= 64'h0;
        src50 <= 64'h0;
        src51 <= 64'h0;
        src52 <= 64'h0;
        src53 <= 64'h0;
        src54 <= 64'h0;
        src55 <= 64'h0;
        src56 <= 64'h0;
        src57 <= 64'h0;
        src58 <= 64'h0;
        src59 <= 64'h0;
        src60 <= 64'h0;
        src61 <= 64'h0;
        src62 <= 64'h0;
        src63 <= 64'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor2_1_64_64(
    input [63:0]src0,
    input [63:0]src1,
    input [63:0]src2,
    input [63:0]src3,
    input [63:0]src4,
    input [63:0]src5,
    input [63:0]src6,
    input [63:0]src7,
    input [63:0]src8,
    input [63:0]src9,
    input [63:0]src10,
    input [63:0]src11,
    input [63:0]src12,
    input [63:0]src13,
    input [63:0]src14,
    input [63:0]src15,
    input [63:0]src16,
    input [63:0]src17,
    input [63:0]src18,
    input [63:0]src19,
    input [63:0]src20,
    input [63:0]src21,
    input [63:0]src22,
    input [63:0]src23,
    input [63:0]src24,
    input [63:0]src25,
    input [63:0]src26,
    input [63:0]src27,
    input [63:0]src28,
    input [63:0]src29,
    input [63:0]src30,
    input [63:0]src31,
    input [63:0]src32,
    input [63:0]src33,
    input [63:0]src34,
    input [63:0]src35,
    input [63:0]src36,
    input [63:0]src37,
    input [63:0]src38,
    input [63:0]src39,
    input [63:0]src40,
    input [63:0]src41,
    input [63:0]src42,
    input [63:0]src43,
    input [63:0]src44,
    input [63:0]src45,
    input [63:0]src46,
    input [63:0]src47,
    input [63:0]src48,
    input [63:0]src49,
    input [63:0]src50,
    input [63:0]src51,
    input [63:0]src52,
    input [63:0]src53,
    input [63:0]src54,
    input [63:0]src55,
    input [63:0]src56,
    input [63:0]src57,
    input [63:0]src58,
    input [63:0]src59,
    input [63:0]src60,
    input [63:0]src61,
    input [63:0]src62,
    input [63:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [0:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [0:0] comp_out67;
    wire [1:0] comp_out68;
    wire [0:0] comp_out69;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69)
    );
    rowadder2_1_70 rowadder2_1inst(
        .src0({comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out68[1], 1'h0, comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], 1'h0, 1'h0, comp_out1[1], comp_out0[1]}),
        .dst0({dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [63:0] src0,
      input wire [63:0] src1,
      input wire [63:0] src2,
      input wire [63:0] src3,
      input wire [63:0] src4,
      input wire [63:0] src5,
      input wire [63:0] src6,
      input wire [63:0] src7,
      input wire [63:0] src8,
      input wire [63:0] src9,
      input wire [63:0] src10,
      input wire [63:0] src11,
      input wire [63:0] src12,
      input wire [63:0] src13,
      input wire [63:0] src14,
      input wire [63:0] src15,
      input wire [63:0] src16,
      input wire [63:0] src17,
      input wire [63:0] src18,
      input wire [63:0] src19,
      input wire [63:0] src20,
      input wire [63:0] src21,
      input wire [63:0] src22,
      input wire [63:0] src23,
      input wire [63:0] src24,
      input wire [63:0] src25,
      input wire [63:0] src26,
      input wire [63:0] src27,
      input wire [63:0] src28,
      input wire [63:0] src29,
      input wire [63:0] src30,
      input wire [63:0] src31,
      input wire [63:0] src32,
      input wire [63:0] src33,
      input wire [63:0] src34,
      input wire [63:0] src35,
      input wire [63:0] src36,
      input wire [63:0] src37,
      input wire [63:0] src38,
      input wire [63:0] src39,
      input wire [63:0] src40,
      input wire [63:0] src41,
      input wire [63:0] src42,
      input wire [63:0] src43,
      input wire [63:0] src44,
      input wire [63:0] src45,
      input wire [63:0] src46,
      input wire [63:0] src47,
      input wire [63:0] src48,
      input wire [63:0] src49,
      input wire [63:0] src50,
      input wire [63:0] src51,
      input wire [63:0] src52,
      input wire [63:0] src53,
      input wire [63:0] src54,
      input wire [63:0] src55,
      input wire [63:0] src56,
      input wire [63:0] src57,
      input wire [63:0] src58,
      input wire [63:0] src59,
      input wire [63:0] src60,
      input wire [63:0] src61,
      input wire [63:0] src62,
      input wire [63:0] src63,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [0:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [0:0] dst67,
      output wire [1:0] dst68,
      output wire [0:0] dst69);

   wire [63:0] stage0_0;
   wire [63:0] stage0_1;
   wire [63:0] stage0_2;
   wire [63:0] stage0_3;
   wire [63:0] stage0_4;
   wire [63:0] stage0_5;
   wire [63:0] stage0_6;
   wire [63:0] stage0_7;
   wire [63:0] stage0_8;
   wire [63:0] stage0_9;
   wire [63:0] stage0_10;
   wire [63:0] stage0_11;
   wire [63:0] stage0_12;
   wire [63:0] stage0_13;
   wire [63:0] stage0_14;
   wire [63:0] stage0_15;
   wire [63:0] stage0_16;
   wire [63:0] stage0_17;
   wire [63:0] stage0_18;
   wire [63:0] stage0_19;
   wire [63:0] stage0_20;
   wire [63:0] stage0_21;
   wire [63:0] stage0_22;
   wire [63:0] stage0_23;
   wire [63:0] stage0_24;
   wire [63:0] stage0_25;
   wire [63:0] stage0_26;
   wire [63:0] stage0_27;
   wire [63:0] stage0_28;
   wire [63:0] stage0_29;
   wire [63:0] stage0_30;
   wire [63:0] stage0_31;
   wire [63:0] stage0_32;
   wire [63:0] stage0_33;
   wire [63:0] stage0_34;
   wire [63:0] stage0_35;
   wire [63:0] stage0_36;
   wire [63:0] stage0_37;
   wire [63:0] stage0_38;
   wire [63:0] stage0_39;
   wire [63:0] stage0_40;
   wire [63:0] stage0_41;
   wire [63:0] stage0_42;
   wire [63:0] stage0_43;
   wire [63:0] stage0_44;
   wire [63:0] stage0_45;
   wire [63:0] stage0_46;
   wire [63:0] stage0_47;
   wire [63:0] stage0_48;
   wire [63:0] stage0_49;
   wire [63:0] stage0_50;
   wire [63:0] stage0_51;
   wire [63:0] stage0_52;
   wire [63:0] stage0_53;
   wire [63:0] stage0_54;
   wire [63:0] stage0_55;
   wire [63:0] stage0_56;
   wire [63:0] stage0_57;
   wire [63:0] stage0_58;
   wire [63:0] stage0_59;
   wire [63:0] stage0_60;
   wire [63:0] stage0_61;
   wire [63:0] stage0_62;
   wire [63:0] stage0_63;
   wire [18:0] stage1_0;
   wire [47:0] stage1_1;
   wire [23:0] stage1_2;
   wire [27:0] stage1_3;
   wire [37:0] stage1_4;
   wire [26:0] stage1_5;
   wire [21:0] stage1_6;
   wire [35:0] stage1_7;
   wire [26:0] stage1_8;
   wire [28:0] stage1_9;
   wire [33:0] stage1_10;
   wire [32:0] stage1_11;
   wire [26:0] stage1_12;
   wire [30:0] stage1_13;
   wire [24:0] stage1_14;
   wire [44:0] stage1_15;
   wire [30:0] stage1_16;
   wire [44:0] stage1_17;
   wire [22:0] stage1_18;
   wire [28:0] stage1_19;
   wire [40:0] stage1_20;
   wire [32:0] stage1_21;
   wire [30:0] stage1_22;
   wire [34:0] stage1_23;
   wire [26:0] stage1_24;
   wire [44:0] stage1_25;
   wire [28:0] stage1_26;
   wire [40:0] stage1_27;
   wire [26:0] stage1_28;
   wire [28:0] stage1_29;
   wire [25:0] stage1_30;
   wire [22:0] stage1_31;
   wire [30:0] stage1_32;
   wire [37:0] stage1_33;
   wire [23:0] stage1_34;
   wire [29:0] stage1_35;
   wire [43:0] stage1_36;
   wire [23:0] stage1_37;
   wire [41:0] stage1_38;
   wire [22:0] stage1_39;
   wire [26:0] stage1_40;
   wire [35:0] stage1_41;
   wire [28:0] stage1_42;
   wire [35:0] stage1_43;
   wire [32:0] stage1_44;
   wire [47:0] stage1_45;
   wire [16:0] stage1_46;
   wire [40:0] stage1_47;
   wire [31:0] stage1_48;
   wire [24:0] stage1_49;
   wire [24:0] stage1_50;
   wire [31:0] stage1_51;
   wire [42:0] stage1_52;
   wire [26:0] stage1_53;
   wire [32:0] stage1_54;
   wire [24:0] stage1_55;
   wire [25:0] stage1_56;
   wire [25:0] stage1_57;
   wire [40:0] stage1_58;
   wire [41:0] stage1_59;
   wire [32:0] stage1_60;
   wire [30:0] stage1_61;
   wire [32:0] stage1_62;
   wire [27:0] stage1_63;
   wire [15:0] stage1_64;
   wire [8:0] stage1_65;
   wire [5:0] stage2_0;
   wire [8:0] stage2_1;
   wire [11:0] stage2_2;
   wire [11:0] stage2_3;
   wire [25:0] stage2_4;
   wire [21:0] stage2_5;
   wire [13:0] stage2_6;
   wire [19:0] stage2_7;
   wire [19:0] stage2_8;
   wire [10:0] stage2_9;
   wire [30:0] stage2_10;
   wire [15:0] stage2_11;
   wire [18:0] stage2_12;
   wire [8:0] stage2_13;
   wire [15:0] stage2_14;
   wire [20:0] stage2_15;
   wire [15:0] stage2_16;
   wire [21:0] stage2_17;
   wire [18:0] stage2_18;
   wire [14:0] stage2_19;
   wire [23:0] stage2_20;
   wire [12:0] stage2_21;
   wire [10:0] stage2_22;
   wire [16:0] stage2_23;
   wire [13:0] stage2_24;
   wire [13:0] stage2_25;
   wire [19:0] stage2_26;
   wire [25:0] stage2_27;
   wire [15:0] stage2_28;
   wire [9:0] stage2_29;
   wire [19:0] stage2_30;
   wire [12:0] stage2_31;
   wire [18:0] stage2_32;
   wire [22:0] stage2_33;
   wire [12:0] stage2_34;
   wire [12:0] stage2_35;
   wire [17:0] stage2_36;
   wire [17:0] stage2_37;
   wire [23:0] stage2_38;
   wire [12:0] stage2_39;
   wire [11:0] stage2_40;
   wire [19:0] stage2_41;
   wire [14:0] stage2_42;
   wire [12:0] stage2_43;
   wire [17:0] stage2_44;
   wire [13:0] stage2_45;
   wire [11:0] stage2_46;
   wire [18:0] stage2_47;
   wire [16:0] stage2_48;
   wire [10:0] stage2_49;
   wire [11:0] stage2_50;
   wire [15:0] stage2_51;
   wire [11:0] stage2_52;
   wire [17:0] stage2_53;
   wire [14:0] stage2_54;
   wire [16:0] stage2_55;
   wire [9:0] stage2_56;
   wire [13:0] stage2_57;
   wire [17:0] stage2_58;
   wire [19:0] stage2_59;
   wire [13:0] stage2_60;
   wire [14:0] stage2_61;
   wire [12:0] stage2_62;
   wire [12:0] stage2_63;
   wire [10:0] stage2_64;
   wire [7:0] stage2_65;
   wire [3:0] stage2_66;
   wire [1:0] stage2_67;
   wire [5:0] stage3_0;
   wire [3:0] stage3_1;
   wire [2:0] stage3_2;
   wire [4:0] stage3_3;
   wire [6:0] stage3_4;
   wire [8:0] stage3_5;
   wire [7:0] stage3_6;
   wire [10:0] stage3_7;
   wire [8:0] stage3_8;
   wire [11:0] stage3_9;
   wire [6:0] stage3_10;
   wire [8:0] stage3_11;
   wire [7:0] stage3_12;
   wire [8:0] stage3_13;
   wire [6:0] stage3_14;
   wire [8:0] stage3_15;
   wire [7:0] stage3_16;
   wire [6:0] stage3_17;
   wire [12:0] stage3_18;
   wire [6:0] stage3_19;
   wire [5:0] stage3_20;
   wire [8:0] stage3_21;
   wire [6:0] stage3_22;
   wire [7:0] stage3_23;
   wire [6:0] stage3_24;
   wire [7:0] stage3_25;
   wire [6:0] stage3_26;
   wire [6:0] stage3_27;
   wire [8:0] stage3_28;
   wire [8:0] stage3_29;
   wire [5:0] stage3_30;
   wire [6:0] stage3_31;
   wire [6:0] stage3_32;
   wire [16:0] stage3_33;
   wire [6:0] stage3_34;
   wire [5:0] stage3_35;
   wire [9:0] stage3_36;
   wire [5:0] stage3_37;
   wire [10:0] stage3_38;
   wire [6:0] stage3_39;
   wire [5:0] stage3_40;
   wire [13:0] stage3_41;
   wire [3:0] stage3_42;
   wire [5:0] stage3_43;
   wire [16:0] stage3_44;
   wire [4:0] stage3_45;
   wire [6:0] stage3_46;
   wire [8:0] stage3_47;
   wire [5:0] stage3_48;
   wire [5:0] stage3_49;
   wire [6:0] stage3_50;
   wire [8:0] stage3_51;
   wire [6:0] stage3_52;
   wire [5:0] stage3_53;
   wire [5:0] stage3_54;
   wire [9:0] stage3_55;
   wire [5:0] stage3_56;
   wire [7:0] stage3_57;
   wire [7:0] stage3_58;
   wire [7:0] stage3_59;
   wire [13:0] stage3_60;
   wire [6:0] stage3_61;
   wire [4:0] stage3_62;
   wire [5:0] stage3_63;
   wire [4:0] stage3_64;
   wire [5:0] stage3_65;
   wire [2:0] stage3_66;
   wire [2:0] stage3_67;
   wire [0:0] stage3_68;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [2:0] stage4_2;
   wire [1:0] stage4_3;
   wire [3:0] stage4_4;
   wire [1:0] stage4_5;
   wire [2:0] stage4_6;
   wire [4:0] stage4_7;
   wire [4:0] stage4_8;
   wire [2:0] stage4_9;
   wire [3:0] stage4_10;
   wire [4:0] stage4_11;
   wire [2:0] stage4_12;
   wire [3:0] stage4_13;
   wire [3:0] stage4_14;
   wire [3:0] stage4_15;
   wire [4:0] stage4_16;
   wire [2:0] stage4_17;
   wire [3:0] stage4_18;
   wire [2:0] stage4_19;
   wire [3:0] stage4_20;
   wire [7:0] stage4_21;
   wire [1:0] stage4_22;
   wire [3:0] stage4_23;
   wire [3:0] stage4_24;
   wire [2:0] stage4_25;
   wire [3:0] stage4_26;
   wire [3:0] stage4_27;
   wire [3:0] stage4_28;
   wire [3:0] stage4_29;
   wire [2:0] stage4_30;
   wire [2:0] stage4_31;
   wire [3:0] stage4_32;
   wire [5:0] stage4_33;
   wire [4:0] stage4_34;
   wire [2:0] stage4_35;
   wire [3:0] stage4_36;
   wire [4:0] stage4_37;
   wire [2:0] stage4_38;
   wire [2:0] stage4_39;
   wire [2:0] stage4_40;
   wire [3:0] stage4_41;
   wire [3:0] stage4_42;
   wire [3:0] stage4_43;
   wire [5:0] stage4_44;
   wire [2:0] stage4_45;
   wire [3:0] stage4_46;
   wire [3:0] stage4_47;
   wire [3:0] stage4_48;
   wire [3:0] stage4_49;
   wire [3:0] stage4_50;
   wire [5:0] stage4_51;
   wire [1:0] stage4_52;
   wire [1:0] stage4_53;
   wire [2:0] stage4_54;
   wire [6:0] stage4_55;
   wire [1:0] stage4_56;
   wire [3:0] stage4_57;
   wire [5:0] stage4_58;
   wire [2:0] stage4_59;
   wire [5:0] stage4_60;
   wire [4:0] stage4_61;
   wire [2:0] stage4_62;
   wire [1:0] stage4_63;
   wire [6:0] stage4_64;
   wire [2:0] stage4_65;
   wire [1:0] stage4_66;
   wire [0:0] stage4_67;
   wire [0:0] stage4_68;
   wire [0:0] stage4_69;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [0:0] stage5_2;
   wire [0:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [1:0] stage5_19;
   wire [1:0] stage5_20;
   wire [1:0] stage5_21;
   wire [1:0] stage5_22;
   wire [1:0] stage5_23;
   wire [1:0] stage5_24;
   wire [1:0] stage5_25;
   wire [1:0] stage5_26;
   wire [1:0] stage5_27;
   wire [1:0] stage5_28;
   wire [1:0] stage5_29;
   wire [1:0] stage5_30;
   wire [1:0] stage5_31;
   wire [1:0] stage5_32;
   wire [1:0] stage5_33;
   wire [1:0] stage5_34;
   wire [1:0] stage5_35;
   wire [1:0] stage5_36;
   wire [1:0] stage5_37;
   wire [1:0] stage5_38;
   wire [1:0] stage5_39;
   wire [1:0] stage5_40;
   wire [1:0] stage5_41;
   wire [1:0] stage5_42;
   wire [1:0] stage5_43;
   wire [1:0] stage5_44;
   wire [1:0] stage5_45;
   wire [1:0] stage5_46;
   wire [1:0] stage5_47;
   wire [1:0] stage5_48;
   wire [1:0] stage5_49;
   wire [1:0] stage5_50;
   wire [1:0] stage5_51;
   wire [1:0] stage5_52;
   wire [1:0] stage5_53;
   wire [1:0] stage5_54;
   wire [1:0] stage5_55;
   wire [1:0] stage5_56;
   wire [1:0] stage5_57;
   wire [1:0] stage5_58;
   wire [1:0] stage5_59;
   wire [1:0] stage5_60;
   wire [1:0] stage5_61;
   wire [1:0] stage5_62;
   wire [1:0] stage5_63;
   wire [1:0] stage5_64;
   wire [1:0] stage5_65;
   wire [1:0] stage5_66;
   wire [0:0] stage5_67;
   wire [1:0] stage5_68;
   wire [0:0] stage5_69;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;
   assign dst22 = stage5_22;
   assign dst23 = stage5_23;
   assign dst24 = stage5_24;
   assign dst25 = stage5_25;
   assign dst26 = stage5_26;
   assign dst27 = stage5_27;
   assign dst28 = stage5_28;
   assign dst29 = stage5_29;
   assign dst30 = stage5_30;
   assign dst31 = stage5_31;
   assign dst32 = stage5_32;
   assign dst33 = stage5_33;
   assign dst34 = stage5_34;
   assign dst35 = stage5_35;
   assign dst36 = stage5_36;
   assign dst37 = stage5_37;
   assign dst38 = stage5_38;
   assign dst39 = stage5_39;
   assign dst40 = stage5_40;
   assign dst41 = stage5_41;
   assign dst42 = stage5_42;
   assign dst43 = stage5_43;
   assign dst44 = stage5_44;
   assign dst45 = stage5_45;
   assign dst46 = stage5_46;
   assign dst47 = stage5_47;
   assign dst48 = stage5_48;
   assign dst49 = stage5_49;
   assign dst50 = stage5_50;
   assign dst51 = stage5_51;
   assign dst52 = stage5_52;
   assign dst53 = stage5_53;
   assign dst54 = stage5_54;
   assign dst55 = stage5_55;
   assign dst56 = stage5_56;
   assign dst57 = stage5_57;
   assign dst58 = stage5_58;
   assign dst59 = stage5_59;
   assign dst60 = stage5_60;
   assign dst61 = stage5_61;
   assign dst62 = stage5_62;
   assign dst63 = stage5_63;
   assign dst64 = stage5_64;
   assign dst65 = stage5_65;
   assign dst66 = stage5_66;
   assign dst67 = stage5_67;
   assign dst68 = stage5_68;
   assign dst69 = stage5_69;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc615_5 gpc14 (
      {stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34]},
      {stage0_4[0]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[0],stage1_5[5],stage1_4[14],stage1_3[14]}
   );
   gpc615_5 gpc15 (
      {stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39]},
      {stage0_4[1]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[1],stage1_5[6],stage1_4[15],stage1_3[15]}
   );
   gpc615_5 gpc16 (
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage0_4[2]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[2],stage1_5[7],stage1_4[16],stage1_3[16]}
   );
   gpc615_5 gpc17 (
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage0_4[3]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[3],stage1_5[8],stage1_4[17],stage1_3[17]}
   );
   gpc615_5 gpc18 (
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage0_4[4]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[4],stage1_5[9],stage1_4[18],stage1_3[18]}
   );
   gpc606_5 gpc19 (
      {stage0_4[5], stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[5],stage1_6[5],stage1_5[10],stage1_4[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[6],stage1_6[6],stage1_5[11],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[17], stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[7],stage1_6[7],stage1_5[12],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[8],stage1_6[8],stage1_5[13],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[9],stage1_6[9],stage1_5[14],stage1_4[23]}
   );
   gpc606_5 gpc24 (
      {stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[10],stage1_6[10],stage1_5[15],stage1_4[24]}
   );
   gpc606_5 gpc25 (
      {stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[11],stage1_6[11],stage1_5[16],stage1_4[25]}
   );
   gpc606_5 gpc26 (
      {stage0_4[47], stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[12],stage1_6[12],stage1_5[17],stage1_4[26]}
   );
   gpc606_5 gpc27 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[8],stage1_7[13],stage1_6[13],stage1_5[18]}
   );
   gpc606_5 gpc28 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[9],stage1_7[14],stage1_6[14],stage1_5[19]}
   );
   gpc606_5 gpc29 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[10],stage1_7[15],stage1_6[15],stage1_5[20]}
   );
   gpc606_5 gpc30 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[11],stage1_7[16],stage1_6[16],stage1_5[21]}
   );
   gpc606_5 gpc31 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[12],stage1_7[17],stage1_6[17],stage1_5[22]}
   );
   gpc615_5 gpc32 (
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52]},
      {stage0_7[30]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[5],stage1_8[13],stage1_7[18],stage1_6[18]}
   );
   gpc615_5 gpc33 (
      {stage0_6[53], stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57]},
      {stage0_7[31]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[6],stage1_8[14],stage1_7[19],stage1_6[19]}
   );
   gpc615_5 gpc34 (
      {stage0_6[58], stage0_6[59], stage0_6[60], stage0_6[61], stage0_6[62]},
      {stage0_7[32]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[7],stage1_8[15],stage1_7[20],stage1_6[20]}
   );
   gpc615_5 gpc35 (
      {stage0_7[33], stage0_7[34], stage0_7[35], stage0_7[36], stage0_7[37]},
      {stage0_8[18]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[8],stage1_8[16],stage1_7[21]}
   );
   gpc615_5 gpc36 (
      {stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41], stage0_7[42]},
      {stage0_8[19]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[4],stage1_9[9],stage1_8[17],stage1_7[22]}
   );
   gpc615_5 gpc37 (
      {stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage0_8[20]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[5],stage1_9[10],stage1_8[18],stage1_7[23]}
   );
   gpc615_5 gpc38 (
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52]},
      {stage0_8[21]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[6],stage1_9[11],stage1_8[19],stage1_7[24]}
   );
   gpc606_5 gpc39 (
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[4],stage1_10[7],stage1_9[12],stage1_8[20]}
   );
   gpc606_5 gpc40 (
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[5],stage1_10[8],stage1_9[13],stage1_8[21]}
   );
   gpc606_5 gpc41 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[6],stage1_10[9],stage1_9[14],stage1_8[22]}
   );
   gpc606_5 gpc42 (
      {stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[7],stage1_10[10],stage1_9[15],stage1_8[23]}
   );
   gpc606_5 gpc43 (
      {stage0_8[46], stage0_8[47], stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[8],stage1_10[11],stage1_9[16],stage1_8[24]}
   );
   gpc606_5 gpc44 (
      {stage0_8[52], stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[9],stage1_10[12],stage1_9[17],stage1_8[25]}
   );
   gpc606_5 gpc45 (
      {stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[10],stage1_10[13],stage1_9[18],stage1_8[26]}
   );
   gpc606_5 gpc46 (
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[7],stage1_11[11],stage1_10[14],stage1_9[19]}
   );
   gpc606_5 gpc47 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[8],stage1_11[12],stage1_10[15],stage1_9[20]}
   );
   gpc606_5 gpc48 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[9],stage1_11[13],stage1_10[16],stage1_9[21]}
   );
   gpc606_5 gpc49 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[10],stage1_11[14],stage1_10[17],stage1_9[22]}
   );
   gpc606_5 gpc50 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[11],stage1_11[15],stage1_10[18],stage1_9[23]}
   );
   gpc606_5 gpc51 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[12],stage1_11[16],stage1_10[19],stage1_9[24]}
   );
   gpc615_5 gpc52 (
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46]},
      {stage0_11[36]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[6],stage1_12[13],stage1_11[17],stage1_10[20]}
   );
   gpc615_5 gpc53 (
      {stage0_10[47], stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51]},
      {stage0_11[37]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[7],stage1_12[14],stage1_11[18],stage1_10[21]}
   );
   gpc615_5 gpc54 (
      {stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41], stage0_11[42]},
      {stage0_12[12]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[2],stage1_13[8],stage1_12[15],stage1_11[19]}
   );
   gpc615_5 gpc55 (
      {stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage0_12[13]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[3],stage1_13[9],stage1_12[16],stage1_11[20]}
   );
   gpc615_5 gpc56 (
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52]},
      {stage0_12[14]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[4],stage1_13[10],stage1_12[17],stage1_11[21]}
   );
   gpc606_5 gpc57 (
      {stage0_12[15], stage0_12[16], stage0_12[17], stage0_12[18], stage0_12[19], stage0_12[20]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[3],stage1_14[5],stage1_13[11],stage1_12[18]}
   );
   gpc606_5 gpc58 (
      {stage0_12[21], stage0_12[22], stage0_12[23], stage0_12[24], stage0_12[25], stage0_12[26]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[4],stage1_14[6],stage1_13[12],stage1_12[19]}
   );
   gpc606_5 gpc59 (
      {stage0_12[27], stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31], stage0_12[32]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[5],stage1_14[7],stage1_13[13],stage1_12[20]}
   );
   gpc606_5 gpc60 (
      {stage0_12[33], stage0_12[34], stage0_12[35], stage0_12[36], stage0_12[37], stage0_12[38]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[6],stage1_14[8],stage1_13[14],stage1_12[21]}
   );
   gpc606_5 gpc61 (
      {stage0_12[39], stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43], stage0_12[44]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[7],stage1_14[9],stage1_13[15],stage1_12[22]}
   );
   gpc606_5 gpc62 (
      {stage0_12[45], stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49], stage0_12[50]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[8],stage1_14[10],stage1_13[16],stage1_12[23]}
   );
   gpc606_5 gpc63 (
      {stage0_12[51], stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55], stage0_12[56]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[9],stage1_14[11],stage1_13[17],stage1_12[24]}
   );
   gpc606_5 gpc64 (
      {stage0_12[57], stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61], stage0_12[62]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[10],stage1_14[12],stage1_13[18],stage1_12[25]}
   );
   gpc2135_5 gpc65 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22]},
      {stage0_14[48], stage0_14[49], stage0_14[50]},
      {stage0_15[0]},
      {stage0_16[0], stage0_16[1]},
      {stage1_17[0],stage1_16[8],stage1_15[11],stage1_14[13],stage1_13[19]}
   );
   gpc606_5 gpc66 (
      {stage0_13[23], stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28]},
      {stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5], stage0_15[6]},
      {stage1_17[1],stage1_16[9],stage1_15[12],stage1_14[14],stage1_13[20]}
   );
   gpc606_5 gpc67 (
      {stage0_13[29], stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34]},
      {stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11], stage0_15[12]},
      {stage1_17[2],stage1_16[10],stage1_15[13],stage1_14[15],stage1_13[21]}
   );
   gpc606_5 gpc68 (
      {stage0_13[35], stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40]},
      {stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17], stage0_15[18]},
      {stage1_17[3],stage1_16[11],stage1_15[14],stage1_14[16],stage1_13[22]}
   );
   gpc606_5 gpc69 (
      {stage0_13[41], stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46]},
      {stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24]},
      {stage1_17[4],stage1_16[12],stage1_15[15],stage1_14[17],stage1_13[23]}
   );
   gpc606_5 gpc70 (
      {stage0_13[47], stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52]},
      {stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29], stage0_15[30]},
      {stage1_17[5],stage1_16[13],stage1_15[16],stage1_14[18],stage1_13[24]}
   );
   gpc606_5 gpc71 (
      {stage0_13[53], stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58]},
      {stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35], stage0_15[36]},
      {stage1_17[6],stage1_16[14],stage1_15[17],stage1_14[19],stage1_13[25]}
   );
   gpc615_5 gpc72 (
      {stage0_14[51], stage0_14[52], stage0_14[53], stage0_14[54], stage0_14[55]},
      {stage0_15[37]},
      {stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5], stage0_16[6], stage0_16[7]},
      {stage1_18[0],stage1_17[7],stage1_16[15],stage1_15[18],stage1_14[20]}
   );
   gpc615_5 gpc73 (
      {stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59], stage0_14[60]},
      {stage0_15[38]},
      {stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11], stage0_16[12], stage0_16[13]},
      {stage1_18[1],stage1_17[8],stage1_16[16],stage1_15[19],stage1_14[21]}
   );
   gpc606_5 gpc74 (
      {stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17], stage0_16[18], stage0_16[19]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[0],stage1_18[2],stage1_17[9],stage1_16[17]}
   );
   gpc606_5 gpc75 (
      {stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23], stage0_16[24], stage0_16[25]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[1],stage1_18[3],stage1_17[10],stage1_16[18]}
   );
   gpc606_5 gpc76 (
      {stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29], stage0_16[30], stage0_16[31]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[2],stage1_18[4],stage1_17[11],stage1_16[19]}
   );
   gpc606_5 gpc77 (
      {stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35], stage0_16[36], stage0_16[37]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[3],stage1_18[5],stage1_17[12],stage1_16[20]}
   );
   gpc615_5 gpc78 (
      {stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42]},
      {stage0_17[0]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[4],stage1_18[6],stage1_17[13],stage1_16[21]}
   );
   gpc615_5 gpc79 (
      {stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage0_17[1]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[5],stage1_18[7],stage1_17[14],stage1_16[22]}
   );
   gpc615_5 gpc80 (
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52]},
      {stage0_17[2]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[6],stage1_18[8],stage1_17[15],stage1_16[23]}
   );
   gpc615_5 gpc81 (
      {stage0_16[53], stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57]},
      {stage0_17[3]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[7],stage1_18[9],stage1_17[16],stage1_16[24]}
   );
   gpc606_5 gpc82 (
      {stage0_17[4], stage0_17[5], stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[8],stage1_19[8],stage1_18[10],stage1_17[17]}
   );
   gpc606_5 gpc83 (
      {stage0_17[10], stage0_17[11], stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[9],stage1_19[9],stage1_18[11],stage1_17[18]}
   );
   gpc606_5 gpc84 (
      {stage0_17[16], stage0_17[17], stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[10],stage1_19[10],stage1_18[12],stage1_17[19]}
   );
   gpc606_5 gpc85 (
      {stage0_17[22], stage0_17[23], stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[11],stage1_19[11],stage1_18[13],stage1_17[20]}
   );
   gpc606_5 gpc86 (
      {stage0_17[28], stage0_17[29], stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[12],stage1_19[12],stage1_18[14],stage1_17[21]}
   );
   gpc606_5 gpc87 (
      {stage0_17[34], stage0_17[35], stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[13],stage1_19[13],stage1_18[15],stage1_17[22]}
   );
   gpc623_5 gpc88 (
      {stage0_17[40], stage0_17[41], stage0_17[42]},
      {stage0_18[48], stage0_18[49]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[14],stage1_19[14],stage1_18[16],stage1_17[23]}
   );
   gpc615_5 gpc89 (
      {stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53], stage0_18[54]},
      {stage0_19[42]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[7],stage1_20[15],stage1_19[15],stage1_18[17]}
   );
   gpc615_5 gpc90 (
      {stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage0_19[43]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[8],stage1_20[16],stage1_19[16],stage1_18[18]}
   );
   gpc615_5 gpc91 (
      {stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47], stage0_19[48]},
      {stage0_20[12]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[2],stage1_21[9],stage1_20[17],stage1_19[17]}
   );
   gpc615_5 gpc92 (
      {stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage0_20[13]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[3],stage1_21[10],stage1_20[18],stage1_19[18]}
   );
   gpc615_5 gpc93 (
      {stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17], stage0_20[18]},
      {stage0_21[12]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[2],stage1_22[4],stage1_21[11],stage1_20[19]}
   );
   gpc615_5 gpc94 (
      {stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage0_21[13]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[3],stage1_22[5],stage1_21[12],stage1_20[20]}
   );
   gpc615_5 gpc95 (
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28]},
      {stage0_21[14]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[4],stage1_22[6],stage1_21[13],stage1_20[21]}
   );
   gpc615_5 gpc96 (
      {stage0_20[29], stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33]},
      {stage0_21[15]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[5],stage1_22[7],stage1_21[14],stage1_20[22]}
   );
   gpc615_5 gpc97 (
      {stage0_20[34], stage0_20[35], stage0_20[36], stage0_20[37], stage0_20[38]},
      {stage0_21[16]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[6],stage1_22[8],stage1_21[15],stage1_20[23]}
   );
   gpc615_5 gpc98 (
      {stage0_20[39], stage0_20[40], stage0_20[41], stage0_20[42], stage0_20[43]},
      {stage0_21[17]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[7],stage1_22[9],stage1_21[16],stage1_20[24]}
   );
   gpc615_5 gpc99 (
      {stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47], stage0_20[48]},
      {stage0_21[18]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[8],stage1_22[10],stage1_21[17],stage1_20[25]}
   );
   gpc606_5 gpc100 (
      {stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[7],stage1_23[9],stage1_22[11],stage1_21[18]}
   );
   gpc606_5 gpc101 (
      {stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[8],stage1_23[10],stage1_22[12],stage1_21[19]}
   );
   gpc606_5 gpc102 (
      {stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35], stage0_21[36]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[9],stage1_23[11],stage1_22[13],stage1_21[20]}
   );
   gpc606_5 gpc103 (
      {stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[10],stage1_23[12],stage1_22[14],stage1_21[21]}
   );
   gpc606_5 gpc104 (
      {stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47], stage0_21[48]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[11],stage1_23[13],stage1_22[15],stage1_21[22]}
   );
   gpc606_5 gpc105 (
      {stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53], stage0_21[54]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[12],stage1_23[14],stage1_22[16],stage1_21[23]}
   );
   gpc615_5 gpc106 (
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46]},
      {stage0_23[36]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[6],stage1_24[13],stage1_23[15],stage1_22[17]}
   );
   gpc615_5 gpc107 (
      {stage0_22[47], stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51]},
      {stage0_23[37]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[7],stage1_24[14],stage1_23[16],stage1_22[18]}
   );
   gpc615_5 gpc108 (
      {stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41], stage0_23[42]},
      {stage0_24[12]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[2],stage1_25[8],stage1_24[15],stage1_23[17]}
   );
   gpc615_5 gpc109 (
      {stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage0_24[13]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[3],stage1_25[9],stage1_24[16],stage1_23[18]}
   );
   gpc606_5 gpc110 (
      {stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17], stage0_24[18], stage0_24[19]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[2],stage1_26[4],stage1_25[10],stage1_24[17]}
   );
   gpc606_5 gpc111 (
      {stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23], stage0_24[24], stage0_24[25]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[3],stage1_26[5],stage1_25[11],stage1_24[18]}
   );
   gpc606_5 gpc112 (
      {stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29], stage0_24[30], stage0_24[31]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[4],stage1_26[6],stage1_25[12],stage1_24[19]}
   );
   gpc606_5 gpc113 (
      {stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35], stage0_24[36], stage0_24[37]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[5],stage1_26[7],stage1_25[13],stage1_24[20]}
   );
   gpc606_5 gpc114 (
      {stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41], stage0_24[42], stage0_24[43]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[6],stage1_26[8],stage1_25[14],stage1_24[21]}
   );
   gpc606_5 gpc115 (
      {stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47], stage0_24[48], stage0_24[49]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[7],stage1_26[9],stage1_25[15],stage1_24[22]}
   );
   gpc606_5 gpc116 (
      {stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53], stage0_24[54], stage0_24[55]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[8],stage1_26[10],stage1_25[16],stage1_24[23]}
   );
   gpc606_5 gpc117 (
      {stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59], stage0_24[60], stage0_24[61]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[9],stage1_26[11],stage1_25[17],stage1_24[24]}
   );
   gpc606_5 gpc118 (
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[8],stage1_27[10],stage1_26[12],stage1_25[18]}
   );
   gpc606_5 gpc119 (
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[9],stage1_27[11],stage1_26[13],stage1_25[19]}
   );
   gpc606_5 gpc120 (
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[10],stage1_27[12],stage1_26[14],stage1_25[20]}
   );
   gpc606_5 gpc121 (
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[11],stage1_27[13],stage1_26[15],stage1_25[21]}
   );
   gpc606_5 gpc122 (
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[12],stage1_27[14],stage1_26[16],stage1_25[22]}
   );
   gpc615_5 gpc123 (
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52]},
      {stage0_27[30]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[5],stage1_28[13],stage1_27[15],stage1_26[17]}
   );
   gpc615_5 gpc124 (
      {stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage0_28[6]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[1],stage1_29[6],stage1_28[14],stage1_27[16]}
   );
   gpc615_5 gpc125 (
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40]},
      {stage0_28[7]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[2],stage1_29[7],stage1_28[15],stage1_27[17]}
   );
   gpc606_5 gpc126 (
      {stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11], stage0_28[12], stage0_28[13]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[2],stage1_30[3],stage1_29[8],stage1_28[16]}
   );
   gpc606_5 gpc127 (
      {stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17], stage0_28[18], stage0_28[19]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[3],stage1_30[4],stage1_29[9],stage1_28[17]}
   );
   gpc606_5 gpc128 (
      {stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23], stage0_28[24], stage0_28[25]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[4],stage1_30[5],stage1_29[10],stage1_28[18]}
   );
   gpc606_5 gpc129 (
      {stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29], stage0_28[30], stage0_28[31]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[5],stage1_30[6],stage1_29[11],stage1_28[19]}
   );
   gpc606_5 gpc130 (
      {stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35], stage0_28[36], stage0_28[37]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[6],stage1_30[7],stage1_29[12],stage1_28[20]}
   );
   gpc606_5 gpc131 (
      {stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41], stage0_28[42], stage0_28[43]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[7],stage1_30[8],stage1_29[13],stage1_28[21]}
   );
   gpc606_5 gpc132 (
      {stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47], stage0_28[48], stage0_28[49]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[8],stage1_30[9],stage1_29[14],stage1_28[22]}
   );
   gpc606_5 gpc133 (
      {stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53], stage0_28[54], stage0_28[55]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[9],stage1_30[10],stage1_29[15],stage1_28[23]}
   );
   gpc606_5 gpc134 (
      {stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59], stage0_28[60], stage0_28[61]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[10],stage1_30[11],stage1_29[16],stage1_28[24]}
   );
   gpc606_5 gpc135 (
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[9],stage1_31[11],stage1_30[12],stage1_29[17]}
   );
   gpc606_5 gpc136 (
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[10],stage1_31[12],stage1_30[13],stage1_29[18]}
   );
   gpc606_5 gpc137 (
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[11],stage1_31[13],stage1_30[14],stage1_29[19]}
   );
   gpc606_5 gpc138 (
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[12],stage1_31[14],stage1_30[15],stage1_29[20]}
   );
   gpc606_5 gpc139 (
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[13],stage1_31[15],stage1_30[16],stage1_29[21]}
   );
   gpc606_5 gpc140 (
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[14],stage1_31[16],stage1_30[17],stage1_29[22]}
   );
   gpc606_5 gpc141 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[15],stage1_31[17],stage1_30[18],stage1_29[23]}
   );
   gpc606_5 gpc142 (
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[16],stage1_31[18],stage1_30[19],stage1_29[24]}
   );
   gpc615_5 gpc143 (
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58]},
      {stage0_31[48]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[8],stage1_32[17],stage1_31[19],stage1_30[20]}
   );
   gpc615_5 gpc144 (
      {stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage0_32[6]},
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage1_35[0],stage1_34[1],stage1_33[9],stage1_32[18],stage1_31[20]}
   );
   gpc615_5 gpc145 (
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58]},
      {stage0_32[7]},
      {stage0_33[6], stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11]},
      {stage1_35[1],stage1_34[2],stage1_33[10],stage1_32[19],stage1_31[21]}
   );
   gpc615_5 gpc146 (
      {stage0_31[59], stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63]},
      {stage0_32[8]},
      {stage0_33[12], stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17]},
      {stage1_35[2],stage1_34[3],stage1_33[11],stage1_32[20],stage1_31[22]}
   );
   gpc606_5 gpc147 (
      {stage0_32[9], stage0_32[10], stage0_32[11], stage0_32[12], stage0_32[13], stage0_32[14]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[3],stage1_34[4],stage1_33[12],stage1_32[21]}
   );
   gpc606_5 gpc148 (
      {stage0_32[15], stage0_32[16], stage0_32[17], stage0_32[18], stage0_32[19], stage0_32[20]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[4],stage1_34[5],stage1_33[13],stage1_32[22]}
   );
   gpc606_5 gpc149 (
      {stage0_32[21], stage0_32[22], stage0_32[23], stage0_32[24], stage0_32[25], stage0_32[26]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[5],stage1_34[6],stage1_33[14],stage1_32[23]}
   );
   gpc606_5 gpc150 (
      {stage0_32[27], stage0_32[28], stage0_32[29], stage0_32[30], stage0_32[31], stage0_32[32]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[6],stage1_34[7],stage1_33[15],stage1_32[24]}
   );
   gpc606_5 gpc151 (
      {stage0_32[33], stage0_32[34], stage0_32[35], stage0_32[36], stage0_32[37], stage0_32[38]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[7],stage1_34[8],stage1_33[16],stage1_32[25]}
   );
   gpc606_5 gpc152 (
      {stage0_32[39], stage0_32[40], stage0_32[41], stage0_32[42], stage0_32[43], stage0_32[44]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[8],stage1_34[9],stage1_33[17],stage1_32[26]}
   );
   gpc606_5 gpc153 (
      {stage0_32[45], stage0_32[46], stage0_32[47], stage0_32[48], stage0_32[49], stage0_32[50]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[9],stage1_34[10],stage1_33[18],stage1_32[27]}
   );
   gpc606_5 gpc154 (
      {stage0_32[51], stage0_32[52], stage0_32[53], stage0_32[54], stage0_32[55], stage0_32[56]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[10],stage1_34[11],stage1_33[19],stage1_32[28]}
   );
   gpc606_5 gpc155 (
      {stage0_32[57], stage0_32[58], stage0_32[59], stage0_32[60], stage0_32[61], stage0_32[62]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[11],stage1_34[12],stage1_33[20],stage1_32[29]}
   );
   gpc606_5 gpc156 (
      {stage0_33[18], stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[9],stage1_35[12],stage1_34[13],stage1_33[21]}
   );
   gpc606_5 gpc157 (
      {stage0_33[24], stage0_33[25], stage0_33[26], stage0_33[27], stage0_33[28], stage0_33[29]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[10],stage1_35[13],stage1_34[14],stage1_33[22]}
   );
   gpc606_5 gpc158 (
      {stage0_33[30], stage0_33[31], stage0_33[32], stage0_33[33], stage0_33[34], stage0_33[35]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[11],stage1_35[14],stage1_34[15],stage1_33[23]}
   );
   gpc606_5 gpc159 (
      {stage0_33[36], stage0_33[37], stage0_33[38], stage0_33[39], stage0_33[40], stage0_33[41]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[12],stage1_35[15],stage1_34[16],stage1_33[24]}
   );
   gpc606_5 gpc160 (
      {stage0_33[42], stage0_33[43], stage0_33[44], stage0_33[45], stage0_33[46], stage0_33[47]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[13],stage1_35[16],stage1_34[17],stage1_33[25]}
   );
   gpc615_5 gpc161 (
      {stage0_33[48], stage0_33[49], stage0_33[50], stage0_33[51], stage0_33[52]},
      {stage0_34[54]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[14],stage1_35[17],stage1_34[18],stage1_33[26]}
   );
   gpc615_5 gpc162 (
      {stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage0_35[36]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[6],stage1_36[15],stage1_35[18],stage1_34[19]}
   );
   gpc615_5 gpc163 (
      {stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage0_36[6]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[1],stage1_37[7],stage1_36[16],stage1_35[19]}
   );
   gpc615_5 gpc164 (
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46]},
      {stage0_36[7]},
      {stage0_37[6], stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11]},
      {stage1_39[1],stage1_38[2],stage1_37[8],stage1_36[17],stage1_35[20]}
   );
   gpc615_5 gpc165 (
      {stage0_35[47], stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51]},
      {stage0_36[8]},
      {stage0_37[12], stage0_37[13], stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17]},
      {stage1_39[2],stage1_38[3],stage1_37[9],stage1_36[18],stage1_35[21]}
   );
   gpc615_5 gpc166 (
      {stage0_35[52], stage0_35[53], stage0_35[54], stage0_35[55], stage0_35[56]},
      {stage0_36[9]},
      {stage0_37[18], stage0_37[19], stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23]},
      {stage1_39[3],stage1_38[4],stage1_37[10],stage1_36[19],stage1_35[22]}
   );
   gpc606_5 gpc167 (
      {stage0_36[10], stage0_36[11], stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[4],stage1_38[5],stage1_37[11],stage1_36[20]}
   );
   gpc606_5 gpc168 (
      {stage0_36[16], stage0_36[17], stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[5],stage1_38[6],stage1_37[12],stage1_36[21]}
   );
   gpc606_5 gpc169 (
      {stage0_36[22], stage0_36[23], stage0_36[24], stage0_36[25], stage0_36[26], stage0_36[27]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[6],stage1_38[7],stage1_37[13],stage1_36[22]}
   );
   gpc606_5 gpc170 (
      {stage0_36[28], stage0_36[29], stage0_36[30], stage0_36[31], stage0_36[32], stage0_36[33]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[7],stage1_38[8],stage1_37[14],stage1_36[23]}
   );
   gpc606_5 gpc171 (
      {stage0_36[34], stage0_36[35], stage0_36[36], stage0_36[37], stage0_36[38], stage0_36[39]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[8],stage1_38[9],stage1_37[15],stage1_36[24]}
   );
   gpc606_5 gpc172 (
      {stage0_36[40], stage0_36[41], stage0_36[42], stage0_36[43], stage0_36[44], stage0_36[45]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[9],stage1_38[10],stage1_37[16],stage1_36[25]}
   );
   gpc606_5 gpc173 (
      {stage0_37[24], stage0_37[25], stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[6],stage1_39[10],stage1_38[11],stage1_37[17]}
   );
   gpc606_5 gpc174 (
      {stage0_37[30], stage0_37[31], stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[7],stage1_39[11],stage1_38[12],stage1_37[18]}
   );
   gpc606_5 gpc175 (
      {stage0_37[36], stage0_37[37], stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[8],stage1_39[12],stage1_38[13],stage1_37[19]}
   );
   gpc606_5 gpc176 (
      {stage0_37[42], stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[9],stage1_39[13],stage1_38[14],stage1_37[20]}
   );
   gpc606_5 gpc177 (
      {stage0_37[48], stage0_37[49], stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[10],stage1_39[14],stage1_38[15],stage1_37[21]}
   );
   gpc606_5 gpc178 (
      {stage0_37[54], stage0_37[55], stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[11],stage1_39[15],stage1_38[16],stage1_37[22]}
   );
   gpc606_5 gpc179 (
      {stage0_37[60], stage0_37[61], stage0_37[62], stage0_37[63], 1'b0, 1'b0},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[12],stage1_39[16],stage1_38[17],stage1_37[23]}
   );
   gpc615_5 gpc180 (
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40]},
      {stage0_39[42]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[7],stage1_40[13],stage1_39[17],stage1_38[18]}
   );
   gpc615_5 gpc181 (
      {stage0_39[43], stage0_39[44], stage0_39[45], stage0_39[46], stage0_39[47]},
      {stage0_40[6]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[1],stage1_41[8],stage1_40[14],stage1_39[18]}
   );
   gpc615_5 gpc182 (
      {stage0_39[48], stage0_39[49], stage0_39[50], stage0_39[51], stage0_39[52]},
      {stage0_40[7]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[2],stage1_41[9],stage1_40[15],stage1_39[19]}
   );
   gpc615_5 gpc183 (
      {stage0_39[53], stage0_39[54], stage0_39[55], stage0_39[56], stage0_39[57]},
      {stage0_40[8]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[3],stage1_41[10],stage1_40[16],stage1_39[20]}
   );
   gpc615_5 gpc184 (
      {stage0_39[58], stage0_39[59], stage0_39[60], stage0_39[61], stage0_39[62]},
      {stage0_40[9]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[4],stage1_41[11],stage1_40[17],stage1_39[21]}
   );
   gpc606_5 gpc185 (
      {stage0_40[10], stage0_40[11], stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[4],stage1_42[5],stage1_41[12],stage1_40[18]}
   );
   gpc606_5 gpc186 (
      {stage0_40[16], stage0_40[17], stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[5],stage1_42[6],stage1_41[13],stage1_40[19]}
   );
   gpc606_5 gpc187 (
      {stage0_40[22], stage0_40[23], stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[6],stage1_42[7],stage1_41[14],stage1_40[20]}
   );
   gpc606_5 gpc188 (
      {stage0_40[28], stage0_40[29], stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[7],stage1_42[8],stage1_41[15],stage1_40[21]}
   );
   gpc606_5 gpc189 (
      {stage0_40[34], stage0_40[35], stage0_40[36], stage0_40[37], stage0_40[38], stage0_40[39]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[8],stage1_42[9],stage1_41[16],stage1_40[22]}
   );
   gpc606_5 gpc190 (
      {stage0_40[40], stage0_40[41], stage0_40[42], stage0_40[43], stage0_40[44], stage0_40[45]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[9],stage1_42[10],stage1_41[17],stage1_40[23]}
   );
   gpc606_5 gpc191 (
      {stage0_40[46], stage0_40[47], stage0_40[48], stage0_40[49], stage0_40[50], stage0_40[51]},
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage1_44[6],stage1_43[10],stage1_42[11],stage1_41[18],stage1_40[24]}
   );
   gpc606_5 gpc192 (
      {stage0_40[52], stage0_40[53], stage0_40[54], stage0_40[55], stage0_40[56], stage0_40[57]},
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage1_44[7],stage1_43[11],stage1_42[12],stage1_41[19],stage1_40[25]}
   );
   gpc606_5 gpc193 (
      {stage0_40[58], stage0_40[59], stage0_40[60], stage0_40[61], stage0_40[62], stage0_40[63]},
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage1_44[8],stage1_43[12],stage1_42[13],stage1_41[20],stage1_40[26]}
   );
   gpc606_5 gpc194 (
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[9],stage1_43[13],stage1_42[14],stage1_41[21]}
   );
   gpc606_5 gpc195 (
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[10],stage1_43[14],stage1_42[15],stage1_41[22]}
   );
   gpc606_5 gpc196 (
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[11],stage1_43[15],stage1_42[16],stage1_41[23]}
   );
   gpc606_5 gpc197 (
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage0_43[18], stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23]},
      {stage1_45[3],stage1_44[12],stage1_43[16],stage1_42[17],stage1_41[24]}
   );
   gpc606_5 gpc198 (
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage0_43[24], stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage1_45[4],stage1_44[13],stage1_43[17],stage1_42[18],stage1_41[25]}
   );
   gpc615_5 gpc199 (
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34]},
      {stage0_44[0]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[0],stage1_45[5],stage1_44[14],stage1_43[18]}
   );
   gpc615_5 gpc200 (
      {stage0_43[35], stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39]},
      {stage0_44[1]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[1],stage1_45[6],stage1_44[15],stage1_43[19]}
   );
   gpc615_5 gpc201 (
      {stage0_43[40], stage0_43[41], stage0_43[42], stage0_43[43], stage0_43[44]},
      {stage0_44[2]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[2],stage1_45[7],stage1_44[16],stage1_43[20]}
   );
   gpc615_5 gpc202 (
      {stage0_43[45], stage0_43[46], stage0_43[47], stage0_43[48], stage0_43[49]},
      {stage0_44[3]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[3],stage1_45[8],stage1_44[17],stage1_43[21]}
   );
   gpc606_5 gpc203 (
      {stage0_44[4], stage0_44[5], stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[4],stage1_46[4],stage1_45[9],stage1_44[18]}
   );
   gpc606_5 gpc204 (
      {stage0_44[10], stage0_44[11], stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[5],stage1_46[5],stage1_45[10],stage1_44[19]}
   );
   gpc606_5 gpc205 (
      {stage0_44[16], stage0_44[17], stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[6],stage1_46[6],stage1_45[11],stage1_44[20]}
   );
   gpc606_5 gpc206 (
      {stage0_44[22], stage0_44[23], stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[7],stage1_46[7],stage1_45[12],stage1_44[21]}
   );
   gpc606_5 gpc207 (
      {stage0_44[28], stage0_44[29], stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[8],stage1_46[8],stage1_45[13],stage1_44[22]}
   );
   gpc606_5 gpc208 (
      {stage0_44[34], stage0_44[35], stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[9],stage1_46[9],stage1_45[14],stage1_44[23]}
   );
   gpc606_5 gpc209 (
      {stage0_44[40], stage0_44[41], stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[10],stage1_46[10],stage1_45[15],stage1_44[24]}
   );
   gpc606_5 gpc210 (
      {stage0_44[46], stage0_44[47], stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[11],stage1_46[11],stage1_45[16],stage1_44[25]}
   );
   gpc606_5 gpc211 (
      {stage0_44[52], stage0_44[53], stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[12],stage1_46[12],stage1_45[17],stage1_44[26]}
   );
   gpc606_5 gpc212 (
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[9],stage1_47[13],stage1_46[13],stage1_45[18]}
   );
   gpc606_5 gpc213 (
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[10],stage1_47[14],stage1_46[14],stage1_45[19]}
   );
   gpc615_5 gpc214 (
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58]},
      {stage0_47[12]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[2],stage1_48[11],stage1_47[15],stage1_46[15]}
   );
   gpc615_5 gpc215 (
      {stage0_46[59], stage0_46[60], stage0_46[61], stage0_46[62], stage0_46[63]},
      {stage0_47[13]},
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage1_50[1],stage1_49[3],stage1_48[12],stage1_47[16],stage1_46[16]}
   );
   gpc606_5 gpc216 (
      {stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17], stage0_47[18], stage0_47[19]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[2],stage1_49[4],stage1_48[13],stage1_47[17]}
   );
   gpc606_5 gpc217 (
      {stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23], stage0_47[24], stage0_47[25]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[3],stage1_49[5],stage1_48[14],stage1_47[18]}
   );
   gpc615_5 gpc218 (
      {stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29], stage0_47[30]},
      {stage0_48[12]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[4],stage1_49[6],stage1_48[15],stage1_47[19]}
   );
   gpc615_5 gpc219 (
      {stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage0_48[13]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[5],stage1_49[7],stage1_48[16],stage1_47[20]}
   );
   gpc615_5 gpc220 (
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40]},
      {stage0_48[14]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[6],stage1_49[8],stage1_48[17],stage1_47[21]}
   );
   gpc615_5 gpc221 (
      {stage0_47[41], stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45]},
      {stage0_48[15]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[7],stage1_49[9],stage1_48[18],stage1_47[22]}
   );
   gpc606_5 gpc222 (
      {stage0_48[16], stage0_48[17], stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[6],stage1_50[8],stage1_49[10],stage1_48[19]}
   );
   gpc606_5 gpc223 (
      {stage0_48[22], stage0_48[23], stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[7],stage1_50[9],stage1_49[11],stage1_48[20]}
   );
   gpc606_5 gpc224 (
      {stage0_48[28], stage0_48[29], stage0_48[30], stage0_48[31], stage0_48[32], stage0_48[33]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[8],stage1_50[10],stage1_49[12],stage1_48[21]}
   );
   gpc606_5 gpc225 (
      {stage0_48[34], stage0_48[35], stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[9],stage1_50[11],stage1_49[13],stage1_48[22]}
   );
   gpc606_5 gpc226 (
      {stage0_48[40], stage0_48[41], stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[10],stage1_50[12],stage1_49[14],stage1_48[23]}
   );
   gpc606_5 gpc227 (
      {stage0_48[46], stage0_48[47], stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[11],stage1_50[13],stage1_49[15],stage1_48[24]}
   );
   gpc606_5 gpc228 (
      {stage0_48[52], stage0_48[53], stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[12],stage1_50[14],stage1_49[16],stage1_48[25]}
   );
   gpc606_5 gpc229 (
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[7],stage1_51[13],stage1_50[15],stage1_49[17]}
   );
   gpc606_5 gpc230 (
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46], stage0_49[47]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[8],stage1_51[14],stage1_50[16],stage1_49[18]}
   );
   gpc606_5 gpc231 (
      {stage0_49[48], stage0_49[49], stage0_49[50], stage0_49[51], stage0_49[52], stage0_49[53]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[9],stage1_51[15],stage1_50[17],stage1_49[19]}
   );
   gpc606_5 gpc232 (
      {stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58], stage0_49[59]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[10],stage1_51[16],stage1_50[18],stage1_49[20]}
   );
   gpc615_5 gpc233 (
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46]},
      {stage0_51[24]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[4],stage1_52[11],stage1_51[17],stage1_50[19]}
   );
   gpc615_5 gpc234 (
      {stage0_50[47], stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51]},
      {stage0_51[25]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[5],stage1_52[12],stage1_51[18],stage1_50[20]}
   );
   gpc615_5 gpc235 (
      {stage0_50[52], stage0_50[53], stage0_50[54], stage0_50[55], stage0_50[56]},
      {stage0_51[26]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[6],stage1_52[13],stage1_51[19],stage1_50[21]}
   );
   gpc615_5 gpc236 (
      {stage0_50[57], stage0_50[58], stage0_50[59], stage0_50[60], stage0_50[61]},
      {stage0_51[27]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[7],stage1_52[14],stage1_51[20],stage1_50[22]}
   );
   gpc606_5 gpc237 (
      {stage0_51[28], stage0_51[29], stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[4],stage1_53[8],stage1_52[15],stage1_51[21]}
   );
   gpc615_5 gpc238 (
      {stage0_51[34], stage0_51[35], stage0_51[36], stage0_51[37], stage0_51[38]},
      {stage0_52[24]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[5],stage1_53[9],stage1_52[16],stage1_51[22]}
   );
   gpc615_5 gpc239 (
      {stage0_51[39], stage0_51[40], stage0_51[41], stage0_51[42], stage0_51[43]},
      {stage0_52[25]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[6],stage1_53[10],stage1_52[17],stage1_51[23]}
   );
   gpc615_5 gpc240 (
      {stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47], stage0_51[48]},
      {stage0_52[26]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[7],stage1_53[11],stage1_52[18],stage1_51[24]}
   );
   gpc615_5 gpc241 (
      {stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage0_52[27]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[8],stage1_53[12],stage1_52[19],stage1_51[25]}
   );
   gpc615_5 gpc242 (
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58]},
      {stage0_52[28]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[9],stage1_53[13],stage1_52[20],stage1_51[26]}
   );
   gpc606_5 gpc243 (
      {stage0_52[29], stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[6],stage1_54[10],stage1_53[14],stage1_52[21]}
   );
   gpc615_5 gpc244 (
      {stage0_52[35], stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39]},
      {stage0_53[36]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[7],stage1_54[11],stage1_53[15],stage1_52[22]}
   );
   gpc615_5 gpc245 (
      {stage0_52[40], stage0_52[41], stage0_52[42], stage0_52[43], stage0_52[44]},
      {stage0_53[37]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[8],stage1_54[12],stage1_53[16],stage1_52[23]}
   );
   gpc615_5 gpc246 (
      {stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41], stage0_53[42]},
      {stage0_54[18]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[3],stage1_55[9],stage1_54[13],stage1_53[17]}
   );
   gpc615_5 gpc247 (
      {stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage0_54[19]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[4],stage1_55[10],stage1_54[14],stage1_53[18]}
   );
   gpc615_5 gpc248 (
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52]},
      {stage0_54[20]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[5],stage1_55[11],stage1_54[15],stage1_53[19]}
   );
   gpc615_5 gpc249 (
      {stage0_53[53], stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57]},
      {stage0_54[21]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[6],stage1_55[12],stage1_54[16],stage1_53[20]}
   );
   gpc606_5 gpc250 (
      {stage0_54[22], stage0_54[23], stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27]},
      {stage0_56[0], stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5]},
      {stage1_58[0],stage1_57[4],stage1_56[7],stage1_55[13],stage1_54[17]}
   );
   gpc606_5 gpc251 (
      {stage0_54[28], stage0_54[29], stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33]},
      {stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11]},
      {stage1_58[1],stage1_57[5],stage1_56[8],stage1_55[14],stage1_54[18]}
   );
   gpc615_5 gpc252 (
      {stage0_54[34], stage0_54[35], stage0_54[36], stage0_54[37], stage0_54[38]},
      {stage0_55[24]},
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage1_58[2],stage1_57[6],stage1_56[9],stage1_55[15],stage1_54[19]}
   );
   gpc615_5 gpc253 (
      {stage0_54[39], stage0_54[40], stage0_54[41], stage0_54[42], stage0_54[43]},
      {stage0_55[25]},
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23]},
      {stage1_58[3],stage1_57[7],stage1_56[10],stage1_55[16],stage1_54[20]}
   );
   gpc615_5 gpc254 (
      {stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47], stage0_54[48]},
      {stage0_55[26]},
      {stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29]},
      {stage1_58[4],stage1_57[8],stage1_56[11],stage1_55[17],stage1_54[21]}
   );
   gpc615_5 gpc255 (
      {stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage0_55[27]},
      {stage0_56[30], stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35]},
      {stage1_58[5],stage1_57[9],stage1_56[12],stage1_55[18],stage1_54[22]}
   );
   gpc606_5 gpc256 (
      {stage0_55[28], stage0_55[29], stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[6],stage1_57[10],stage1_56[13],stage1_55[19]}
   );
   gpc606_5 gpc257 (
      {stage0_55[34], stage0_55[35], stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[7],stage1_57[11],stage1_56[14],stage1_55[20]}
   );
   gpc606_5 gpc258 (
      {stage0_55[40], stage0_55[41], stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[8],stage1_57[12],stage1_56[15],stage1_55[21]}
   );
   gpc606_5 gpc259 (
      {stage0_55[46], stage0_55[47], stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[9],stage1_57[13],stage1_56[16],stage1_55[22]}
   );
   gpc606_5 gpc260 (
      {stage0_55[52], stage0_55[53], stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57]},
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage1_59[4],stage1_58[10],stage1_57[14],stage1_56[17],stage1_55[23]}
   );
   gpc606_5 gpc261 (
      {stage0_55[58], stage0_55[59], stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63]},
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage1_59[5],stage1_58[11],stage1_57[15],stage1_56[18],stage1_55[24]}
   );
   gpc606_5 gpc262 (
      {stage0_56[36], stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[6],stage1_58[12],stage1_57[16],stage1_56[19]}
   );
   gpc615_5 gpc263 (
      {stage0_56[42], stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46]},
      {stage0_57[36]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[7],stage1_58[13],stage1_57[17],stage1_56[20]}
   );
   gpc615_5 gpc264 (
      {stage0_56[47], stage0_56[48], stage0_56[49], stage0_56[50], stage0_56[51]},
      {stage0_57[37]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[8],stage1_58[14],stage1_57[18],stage1_56[21]}
   );
   gpc615_5 gpc265 (
      {stage0_56[52], stage0_56[53], stage0_56[54], stage0_56[55], stage0_56[56]},
      {stage0_57[38]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[9],stage1_58[15],stage1_57[19],stage1_56[22]}
   );
   gpc615_5 gpc266 (
      {stage0_56[57], stage0_56[58], stage0_56[59], stage0_56[60], stage0_56[61]},
      {stage0_57[39]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[10],stage1_58[16],stage1_57[20],stage1_56[23]}
   );
   gpc615_5 gpc267 (
      {stage0_57[40], stage0_57[41], stage0_57[42], stage0_57[43], stage0_57[44]},
      {stage0_58[30]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[5],stage1_59[11],stage1_58[17],stage1_57[21]}
   );
   gpc615_5 gpc268 (
      {stage0_57[45], stage0_57[46], stage0_57[47], stage0_57[48], stage0_57[49]},
      {stage0_58[31]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[6],stage1_59[12],stage1_58[18],stage1_57[22]}
   );
   gpc615_5 gpc269 (
      {stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53], stage0_57[54]},
      {stage0_58[32]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[7],stage1_59[13],stage1_58[19],stage1_57[23]}
   );
   gpc615_5 gpc270 (
      {stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage0_58[33]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[8],stage1_59[14],stage1_58[20],stage1_57[24]}
   );
   gpc615_5 gpc271 (
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], 1'b0},
      {stage0_58[34]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[9],stage1_59[15],stage1_58[21],stage1_57[25]}
   );
   gpc1406_5 gpc272 (
      {stage0_58[35], stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3]},
      {stage0_61[0]},
      {stage1_62[0],stage1_61[5],stage1_60[10],stage1_59[16],stage1_58[22]}
   );
   gpc606_5 gpc273 (
      {stage0_58[41], stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46]},
      {stage0_60[4], stage0_60[5], stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9]},
      {stage1_62[1],stage1_61[6],stage1_60[11],stage1_59[17],stage1_58[23]}
   );
   gpc606_5 gpc274 (
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage0_61[1], stage0_61[2], stage0_61[3], stage0_61[4], stage0_61[5], stage0_61[6]},
      {stage1_63[0],stage1_62[2],stage1_61[7],stage1_60[12],stage1_59[18]}
   );
   gpc606_5 gpc275 (
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage0_61[7], stage0_61[8], stage0_61[9], stage0_61[10], stage0_61[11], stage0_61[12]},
      {stage1_63[1],stage1_62[3],stage1_61[8],stage1_60[13],stage1_59[19]}
   );
   gpc606_5 gpc276 (
      {stage0_60[10], stage0_60[11], stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[2],stage1_62[4],stage1_61[9],stage1_60[14]}
   );
   gpc606_5 gpc277 (
      {stage0_60[16], stage0_60[17], stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[3],stage1_62[5],stage1_61[10],stage1_60[15]}
   );
   gpc606_5 gpc278 (
      {stage0_60[22], stage0_60[23], stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[4],stage1_62[6],stage1_61[11],stage1_60[16]}
   );
   gpc606_5 gpc279 (
      {stage0_60[28], stage0_60[29], stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[5],stage1_62[7],stage1_61[12],stage1_60[17]}
   );
   gpc606_5 gpc280 (
      {stage0_60[34], stage0_60[35], stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[6],stage1_62[8],stage1_61[13],stage1_60[18]}
   );
   gpc606_5 gpc281 (
      {stage0_60[40], stage0_60[41], stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[7],stage1_62[9],stage1_61[14],stage1_60[19]}
   );
   gpc606_5 gpc282 (
      {stage0_60[46], stage0_60[47], stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[8],stage1_62[10],stage1_61[15],stage1_60[20]}
   );
   gpc615_5 gpc283 (
      {stage0_61[13], stage0_61[14], stage0_61[15], stage0_61[16], stage0_61[17]},
      {stage0_62[42]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[7],stage1_63[9],stage1_62[11],stage1_61[16]}
   );
   gpc615_5 gpc284 (
      {stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21], stage0_61[22]},
      {stage0_62[43]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[8],stage1_63[10],stage1_62[12],stage1_61[17]}
   );
   gpc615_5 gpc285 (
      {stage0_61[23], stage0_61[24], stage0_61[25], stage0_61[26], stage0_61[27]},
      {stage0_62[44]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[9],stage1_63[11],stage1_62[13],stage1_61[18]}
   );
   gpc615_5 gpc286 (
      {stage0_61[28], stage0_61[29], stage0_61[30], stage0_61[31], stage0_61[32]},
      {stage0_62[45]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[10],stage1_63[12],stage1_62[14],stage1_61[19]}
   );
   gpc615_5 gpc287 (
      {stage0_61[33], stage0_61[34], stage0_61[35], stage0_61[36], stage0_61[37]},
      {stage0_62[46]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[11],stage1_63[13],stage1_62[15],stage1_61[20]}
   );
   gpc615_5 gpc288 (
      {stage0_61[38], stage0_61[39], stage0_61[40], stage0_61[41], stage0_61[42]},
      {stage0_62[47]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[12],stage1_63[14],stage1_62[16],stage1_61[21]}
   );
   gpc615_5 gpc289 (
      {stage0_61[43], stage0_61[44], stage0_61[45], stage0_61[46], stage0_61[47]},
      {stage0_62[48]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[13],stage1_63[15],stage1_62[17],stage1_61[22]}
   );
   gpc615_5 gpc290 (
      {stage0_61[48], stage0_61[49], stage0_61[50], stage0_61[51], stage0_61[52]},
      {stage0_62[49]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[14],stage1_63[16],stage1_62[18],stage1_61[23]}
   );
   gpc615_5 gpc291 (
      {stage0_61[53], stage0_61[54], stage0_61[55], stage0_61[56], stage0_61[57]},
      {stage0_62[50]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[15],stage1_63[17],stage1_62[19],stage1_61[24]}
   );
   gpc1_1 gpc292 (
      {stage0_0[54]},
      {stage1_0[9]}
   );
   gpc1_1 gpc293 (
      {stage0_0[55]},
      {stage1_0[10]}
   );
   gpc1_1 gpc294 (
      {stage0_0[56]},
      {stage1_0[11]}
   );
   gpc1_1 gpc295 (
      {stage0_0[57]},
      {stage1_0[12]}
   );
   gpc1_1 gpc296 (
      {stage0_0[58]},
      {stage1_0[13]}
   );
   gpc1_1 gpc297 (
      {stage0_0[59]},
      {stage1_0[14]}
   );
   gpc1_1 gpc298 (
      {stage0_0[60]},
      {stage1_0[15]}
   );
   gpc1_1 gpc299 (
      {stage0_0[61]},
      {stage1_0[16]}
   );
   gpc1_1 gpc300 (
      {stage0_0[62]},
      {stage1_0[17]}
   );
   gpc1_1 gpc301 (
      {stage0_0[63]},
      {stage1_0[18]}
   );
   gpc1_1 gpc302 (
      {stage0_1[30]},
      {stage1_1[14]}
   );
   gpc1_1 gpc303 (
      {stage0_1[31]},
      {stage1_1[15]}
   );
   gpc1_1 gpc304 (
      {stage0_1[32]},
      {stage1_1[16]}
   );
   gpc1_1 gpc305 (
      {stage0_1[33]},
      {stage1_1[17]}
   );
   gpc1_1 gpc306 (
      {stage0_1[34]},
      {stage1_1[18]}
   );
   gpc1_1 gpc307 (
      {stage0_1[35]},
      {stage1_1[19]}
   );
   gpc1_1 gpc308 (
      {stage0_1[36]},
      {stage1_1[20]}
   );
   gpc1_1 gpc309 (
      {stage0_1[37]},
      {stage1_1[21]}
   );
   gpc1_1 gpc310 (
      {stage0_1[38]},
      {stage1_1[22]}
   );
   gpc1_1 gpc311 (
      {stage0_1[39]},
      {stage1_1[23]}
   );
   gpc1_1 gpc312 (
      {stage0_1[40]},
      {stage1_1[24]}
   );
   gpc1_1 gpc313 (
      {stage0_1[41]},
      {stage1_1[25]}
   );
   gpc1_1 gpc314 (
      {stage0_1[42]},
      {stage1_1[26]}
   );
   gpc1_1 gpc315 (
      {stage0_1[43]},
      {stage1_1[27]}
   );
   gpc1_1 gpc316 (
      {stage0_1[44]},
      {stage1_1[28]}
   );
   gpc1_1 gpc317 (
      {stage0_1[45]},
      {stage1_1[29]}
   );
   gpc1_1 gpc318 (
      {stage0_1[46]},
      {stage1_1[30]}
   );
   gpc1_1 gpc319 (
      {stage0_1[47]},
      {stage1_1[31]}
   );
   gpc1_1 gpc320 (
      {stage0_1[48]},
      {stage1_1[32]}
   );
   gpc1_1 gpc321 (
      {stage0_1[49]},
      {stage1_1[33]}
   );
   gpc1_1 gpc322 (
      {stage0_1[50]},
      {stage1_1[34]}
   );
   gpc1_1 gpc323 (
      {stage0_1[51]},
      {stage1_1[35]}
   );
   gpc1_1 gpc324 (
      {stage0_1[52]},
      {stage1_1[36]}
   );
   gpc1_1 gpc325 (
      {stage0_1[53]},
      {stage1_1[37]}
   );
   gpc1_1 gpc326 (
      {stage0_1[54]},
      {stage1_1[38]}
   );
   gpc1_1 gpc327 (
      {stage0_1[55]},
      {stage1_1[39]}
   );
   gpc1_1 gpc328 (
      {stage0_1[56]},
      {stage1_1[40]}
   );
   gpc1_1 gpc329 (
      {stage0_1[57]},
      {stage1_1[41]}
   );
   gpc1_1 gpc330 (
      {stage0_1[58]},
      {stage1_1[42]}
   );
   gpc1_1 gpc331 (
      {stage0_1[59]},
      {stage1_1[43]}
   );
   gpc1_1 gpc332 (
      {stage0_1[60]},
      {stage1_1[44]}
   );
   gpc1_1 gpc333 (
      {stage0_1[61]},
      {stage1_1[45]}
   );
   gpc1_1 gpc334 (
      {stage0_1[62]},
      {stage1_1[46]}
   );
   gpc1_1 gpc335 (
      {stage0_1[63]},
      {stage1_1[47]}
   );
   gpc1_1 gpc336 (
      {stage0_2[54]},
      {stage1_2[14]}
   );
   gpc1_1 gpc337 (
      {stage0_2[55]},
      {stage1_2[15]}
   );
   gpc1_1 gpc338 (
      {stage0_2[56]},
      {stage1_2[16]}
   );
   gpc1_1 gpc339 (
      {stage0_2[57]},
      {stage1_2[17]}
   );
   gpc1_1 gpc340 (
      {stage0_2[58]},
      {stage1_2[18]}
   );
   gpc1_1 gpc341 (
      {stage0_2[59]},
      {stage1_2[19]}
   );
   gpc1_1 gpc342 (
      {stage0_2[60]},
      {stage1_2[20]}
   );
   gpc1_1 gpc343 (
      {stage0_2[61]},
      {stage1_2[21]}
   );
   gpc1_1 gpc344 (
      {stage0_2[62]},
      {stage1_2[22]}
   );
   gpc1_1 gpc345 (
      {stage0_2[63]},
      {stage1_2[23]}
   );
   gpc1_1 gpc346 (
      {stage0_3[55]},
      {stage1_3[19]}
   );
   gpc1_1 gpc347 (
      {stage0_3[56]},
      {stage1_3[20]}
   );
   gpc1_1 gpc348 (
      {stage0_3[57]},
      {stage1_3[21]}
   );
   gpc1_1 gpc349 (
      {stage0_3[58]},
      {stage1_3[22]}
   );
   gpc1_1 gpc350 (
      {stage0_3[59]},
      {stage1_3[23]}
   );
   gpc1_1 gpc351 (
      {stage0_3[60]},
      {stage1_3[24]}
   );
   gpc1_1 gpc352 (
      {stage0_3[61]},
      {stage1_3[25]}
   );
   gpc1_1 gpc353 (
      {stage0_3[62]},
      {stage1_3[26]}
   );
   gpc1_1 gpc354 (
      {stage0_3[63]},
      {stage1_3[27]}
   );
   gpc1_1 gpc355 (
      {stage0_4[53]},
      {stage1_4[27]}
   );
   gpc1_1 gpc356 (
      {stage0_4[54]},
      {stage1_4[28]}
   );
   gpc1_1 gpc357 (
      {stage0_4[55]},
      {stage1_4[29]}
   );
   gpc1_1 gpc358 (
      {stage0_4[56]},
      {stage1_4[30]}
   );
   gpc1_1 gpc359 (
      {stage0_4[57]},
      {stage1_4[31]}
   );
   gpc1_1 gpc360 (
      {stage0_4[58]},
      {stage1_4[32]}
   );
   gpc1_1 gpc361 (
      {stage0_4[59]},
      {stage1_4[33]}
   );
   gpc1_1 gpc362 (
      {stage0_4[60]},
      {stage1_4[34]}
   );
   gpc1_1 gpc363 (
      {stage0_4[61]},
      {stage1_4[35]}
   );
   gpc1_1 gpc364 (
      {stage0_4[62]},
      {stage1_4[36]}
   );
   gpc1_1 gpc365 (
      {stage0_4[63]},
      {stage1_4[37]}
   );
   gpc1_1 gpc366 (
      {stage0_5[60]},
      {stage1_5[23]}
   );
   gpc1_1 gpc367 (
      {stage0_5[61]},
      {stage1_5[24]}
   );
   gpc1_1 gpc368 (
      {stage0_5[62]},
      {stage1_5[25]}
   );
   gpc1_1 gpc369 (
      {stage0_5[63]},
      {stage1_5[26]}
   );
   gpc1_1 gpc370 (
      {stage0_6[63]},
      {stage1_6[21]}
   );
   gpc1_1 gpc371 (
      {stage0_7[53]},
      {stage1_7[25]}
   );
   gpc1_1 gpc372 (
      {stage0_7[54]},
      {stage1_7[26]}
   );
   gpc1_1 gpc373 (
      {stage0_7[55]},
      {stage1_7[27]}
   );
   gpc1_1 gpc374 (
      {stage0_7[56]},
      {stage1_7[28]}
   );
   gpc1_1 gpc375 (
      {stage0_7[57]},
      {stage1_7[29]}
   );
   gpc1_1 gpc376 (
      {stage0_7[58]},
      {stage1_7[30]}
   );
   gpc1_1 gpc377 (
      {stage0_7[59]},
      {stage1_7[31]}
   );
   gpc1_1 gpc378 (
      {stage0_7[60]},
      {stage1_7[32]}
   );
   gpc1_1 gpc379 (
      {stage0_7[61]},
      {stage1_7[33]}
   );
   gpc1_1 gpc380 (
      {stage0_7[62]},
      {stage1_7[34]}
   );
   gpc1_1 gpc381 (
      {stage0_7[63]},
      {stage1_7[35]}
   );
   gpc1_1 gpc382 (
      {stage0_9[60]},
      {stage1_9[25]}
   );
   gpc1_1 gpc383 (
      {stage0_9[61]},
      {stage1_9[26]}
   );
   gpc1_1 gpc384 (
      {stage0_9[62]},
      {stage1_9[27]}
   );
   gpc1_1 gpc385 (
      {stage0_9[63]},
      {stage1_9[28]}
   );
   gpc1_1 gpc386 (
      {stage0_10[52]},
      {stage1_10[22]}
   );
   gpc1_1 gpc387 (
      {stage0_10[53]},
      {stage1_10[23]}
   );
   gpc1_1 gpc388 (
      {stage0_10[54]},
      {stage1_10[24]}
   );
   gpc1_1 gpc389 (
      {stage0_10[55]},
      {stage1_10[25]}
   );
   gpc1_1 gpc390 (
      {stage0_10[56]},
      {stage1_10[26]}
   );
   gpc1_1 gpc391 (
      {stage0_10[57]},
      {stage1_10[27]}
   );
   gpc1_1 gpc392 (
      {stage0_10[58]},
      {stage1_10[28]}
   );
   gpc1_1 gpc393 (
      {stage0_10[59]},
      {stage1_10[29]}
   );
   gpc1_1 gpc394 (
      {stage0_10[60]},
      {stage1_10[30]}
   );
   gpc1_1 gpc395 (
      {stage0_10[61]},
      {stage1_10[31]}
   );
   gpc1_1 gpc396 (
      {stage0_10[62]},
      {stage1_10[32]}
   );
   gpc1_1 gpc397 (
      {stage0_10[63]},
      {stage1_10[33]}
   );
   gpc1_1 gpc398 (
      {stage0_11[53]},
      {stage1_11[22]}
   );
   gpc1_1 gpc399 (
      {stage0_11[54]},
      {stage1_11[23]}
   );
   gpc1_1 gpc400 (
      {stage0_11[55]},
      {stage1_11[24]}
   );
   gpc1_1 gpc401 (
      {stage0_11[56]},
      {stage1_11[25]}
   );
   gpc1_1 gpc402 (
      {stage0_11[57]},
      {stage1_11[26]}
   );
   gpc1_1 gpc403 (
      {stage0_11[58]},
      {stage1_11[27]}
   );
   gpc1_1 gpc404 (
      {stage0_11[59]},
      {stage1_11[28]}
   );
   gpc1_1 gpc405 (
      {stage0_11[60]},
      {stage1_11[29]}
   );
   gpc1_1 gpc406 (
      {stage0_11[61]},
      {stage1_11[30]}
   );
   gpc1_1 gpc407 (
      {stage0_11[62]},
      {stage1_11[31]}
   );
   gpc1_1 gpc408 (
      {stage0_11[63]},
      {stage1_11[32]}
   );
   gpc1_1 gpc409 (
      {stage0_12[63]},
      {stage1_12[26]}
   );
   gpc1_1 gpc410 (
      {stage0_13[59]},
      {stage1_13[26]}
   );
   gpc1_1 gpc411 (
      {stage0_13[60]},
      {stage1_13[27]}
   );
   gpc1_1 gpc412 (
      {stage0_13[61]},
      {stage1_13[28]}
   );
   gpc1_1 gpc413 (
      {stage0_13[62]},
      {stage1_13[29]}
   );
   gpc1_1 gpc414 (
      {stage0_13[63]},
      {stage1_13[30]}
   );
   gpc1_1 gpc415 (
      {stage0_14[61]},
      {stage1_14[22]}
   );
   gpc1_1 gpc416 (
      {stage0_14[62]},
      {stage1_14[23]}
   );
   gpc1_1 gpc417 (
      {stage0_14[63]},
      {stage1_14[24]}
   );
   gpc1_1 gpc418 (
      {stage0_15[39]},
      {stage1_15[20]}
   );
   gpc1_1 gpc419 (
      {stage0_15[40]},
      {stage1_15[21]}
   );
   gpc1_1 gpc420 (
      {stage0_15[41]},
      {stage1_15[22]}
   );
   gpc1_1 gpc421 (
      {stage0_15[42]},
      {stage1_15[23]}
   );
   gpc1_1 gpc422 (
      {stage0_15[43]},
      {stage1_15[24]}
   );
   gpc1_1 gpc423 (
      {stage0_15[44]},
      {stage1_15[25]}
   );
   gpc1_1 gpc424 (
      {stage0_15[45]},
      {stage1_15[26]}
   );
   gpc1_1 gpc425 (
      {stage0_15[46]},
      {stage1_15[27]}
   );
   gpc1_1 gpc426 (
      {stage0_15[47]},
      {stage1_15[28]}
   );
   gpc1_1 gpc427 (
      {stage0_15[48]},
      {stage1_15[29]}
   );
   gpc1_1 gpc428 (
      {stage0_15[49]},
      {stage1_15[30]}
   );
   gpc1_1 gpc429 (
      {stage0_15[50]},
      {stage1_15[31]}
   );
   gpc1_1 gpc430 (
      {stage0_15[51]},
      {stage1_15[32]}
   );
   gpc1_1 gpc431 (
      {stage0_15[52]},
      {stage1_15[33]}
   );
   gpc1_1 gpc432 (
      {stage0_15[53]},
      {stage1_15[34]}
   );
   gpc1_1 gpc433 (
      {stage0_15[54]},
      {stage1_15[35]}
   );
   gpc1_1 gpc434 (
      {stage0_15[55]},
      {stage1_15[36]}
   );
   gpc1_1 gpc435 (
      {stage0_15[56]},
      {stage1_15[37]}
   );
   gpc1_1 gpc436 (
      {stage0_15[57]},
      {stage1_15[38]}
   );
   gpc1_1 gpc437 (
      {stage0_15[58]},
      {stage1_15[39]}
   );
   gpc1_1 gpc438 (
      {stage0_15[59]},
      {stage1_15[40]}
   );
   gpc1_1 gpc439 (
      {stage0_15[60]},
      {stage1_15[41]}
   );
   gpc1_1 gpc440 (
      {stage0_15[61]},
      {stage1_15[42]}
   );
   gpc1_1 gpc441 (
      {stage0_15[62]},
      {stage1_15[43]}
   );
   gpc1_1 gpc442 (
      {stage0_15[63]},
      {stage1_15[44]}
   );
   gpc1_1 gpc443 (
      {stage0_16[58]},
      {stage1_16[25]}
   );
   gpc1_1 gpc444 (
      {stage0_16[59]},
      {stage1_16[26]}
   );
   gpc1_1 gpc445 (
      {stage0_16[60]},
      {stage1_16[27]}
   );
   gpc1_1 gpc446 (
      {stage0_16[61]},
      {stage1_16[28]}
   );
   gpc1_1 gpc447 (
      {stage0_16[62]},
      {stage1_16[29]}
   );
   gpc1_1 gpc448 (
      {stage0_16[63]},
      {stage1_16[30]}
   );
   gpc1_1 gpc449 (
      {stage0_17[43]},
      {stage1_17[24]}
   );
   gpc1_1 gpc450 (
      {stage0_17[44]},
      {stage1_17[25]}
   );
   gpc1_1 gpc451 (
      {stage0_17[45]},
      {stage1_17[26]}
   );
   gpc1_1 gpc452 (
      {stage0_17[46]},
      {stage1_17[27]}
   );
   gpc1_1 gpc453 (
      {stage0_17[47]},
      {stage1_17[28]}
   );
   gpc1_1 gpc454 (
      {stage0_17[48]},
      {stage1_17[29]}
   );
   gpc1_1 gpc455 (
      {stage0_17[49]},
      {stage1_17[30]}
   );
   gpc1_1 gpc456 (
      {stage0_17[50]},
      {stage1_17[31]}
   );
   gpc1_1 gpc457 (
      {stage0_17[51]},
      {stage1_17[32]}
   );
   gpc1_1 gpc458 (
      {stage0_17[52]},
      {stage1_17[33]}
   );
   gpc1_1 gpc459 (
      {stage0_17[53]},
      {stage1_17[34]}
   );
   gpc1_1 gpc460 (
      {stage0_17[54]},
      {stage1_17[35]}
   );
   gpc1_1 gpc461 (
      {stage0_17[55]},
      {stage1_17[36]}
   );
   gpc1_1 gpc462 (
      {stage0_17[56]},
      {stage1_17[37]}
   );
   gpc1_1 gpc463 (
      {stage0_17[57]},
      {stage1_17[38]}
   );
   gpc1_1 gpc464 (
      {stage0_17[58]},
      {stage1_17[39]}
   );
   gpc1_1 gpc465 (
      {stage0_17[59]},
      {stage1_17[40]}
   );
   gpc1_1 gpc466 (
      {stage0_17[60]},
      {stage1_17[41]}
   );
   gpc1_1 gpc467 (
      {stage0_17[61]},
      {stage1_17[42]}
   );
   gpc1_1 gpc468 (
      {stage0_17[62]},
      {stage1_17[43]}
   );
   gpc1_1 gpc469 (
      {stage0_17[63]},
      {stage1_17[44]}
   );
   gpc1_1 gpc470 (
      {stage0_18[60]},
      {stage1_18[19]}
   );
   gpc1_1 gpc471 (
      {stage0_18[61]},
      {stage1_18[20]}
   );
   gpc1_1 gpc472 (
      {stage0_18[62]},
      {stage1_18[21]}
   );
   gpc1_1 gpc473 (
      {stage0_18[63]},
      {stage1_18[22]}
   );
   gpc1_1 gpc474 (
      {stage0_19[54]},
      {stage1_19[19]}
   );
   gpc1_1 gpc475 (
      {stage0_19[55]},
      {stage1_19[20]}
   );
   gpc1_1 gpc476 (
      {stage0_19[56]},
      {stage1_19[21]}
   );
   gpc1_1 gpc477 (
      {stage0_19[57]},
      {stage1_19[22]}
   );
   gpc1_1 gpc478 (
      {stage0_19[58]},
      {stage1_19[23]}
   );
   gpc1_1 gpc479 (
      {stage0_19[59]},
      {stage1_19[24]}
   );
   gpc1_1 gpc480 (
      {stage0_19[60]},
      {stage1_19[25]}
   );
   gpc1_1 gpc481 (
      {stage0_19[61]},
      {stage1_19[26]}
   );
   gpc1_1 gpc482 (
      {stage0_19[62]},
      {stage1_19[27]}
   );
   gpc1_1 gpc483 (
      {stage0_19[63]},
      {stage1_19[28]}
   );
   gpc1_1 gpc484 (
      {stage0_20[49]},
      {stage1_20[26]}
   );
   gpc1_1 gpc485 (
      {stage0_20[50]},
      {stage1_20[27]}
   );
   gpc1_1 gpc486 (
      {stage0_20[51]},
      {stage1_20[28]}
   );
   gpc1_1 gpc487 (
      {stage0_20[52]},
      {stage1_20[29]}
   );
   gpc1_1 gpc488 (
      {stage0_20[53]},
      {stage1_20[30]}
   );
   gpc1_1 gpc489 (
      {stage0_20[54]},
      {stage1_20[31]}
   );
   gpc1_1 gpc490 (
      {stage0_20[55]},
      {stage1_20[32]}
   );
   gpc1_1 gpc491 (
      {stage0_20[56]},
      {stage1_20[33]}
   );
   gpc1_1 gpc492 (
      {stage0_20[57]},
      {stage1_20[34]}
   );
   gpc1_1 gpc493 (
      {stage0_20[58]},
      {stage1_20[35]}
   );
   gpc1_1 gpc494 (
      {stage0_20[59]},
      {stage1_20[36]}
   );
   gpc1_1 gpc495 (
      {stage0_20[60]},
      {stage1_20[37]}
   );
   gpc1_1 gpc496 (
      {stage0_20[61]},
      {stage1_20[38]}
   );
   gpc1_1 gpc497 (
      {stage0_20[62]},
      {stage1_20[39]}
   );
   gpc1_1 gpc498 (
      {stage0_20[63]},
      {stage1_20[40]}
   );
   gpc1_1 gpc499 (
      {stage0_21[55]},
      {stage1_21[24]}
   );
   gpc1_1 gpc500 (
      {stage0_21[56]},
      {stage1_21[25]}
   );
   gpc1_1 gpc501 (
      {stage0_21[57]},
      {stage1_21[26]}
   );
   gpc1_1 gpc502 (
      {stage0_21[58]},
      {stage1_21[27]}
   );
   gpc1_1 gpc503 (
      {stage0_21[59]},
      {stage1_21[28]}
   );
   gpc1_1 gpc504 (
      {stage0_21[60]},
      {stage1_21[29]}
   );
   gpc1_1 gpc505 (
      {stage0_21[61]},
      {stage1_21[30]}
   );
   gpc1_1 gpc506 (
      {stage0_21[62]},
      {stage1_21[31]}
   );
   gpc1_1 gpc507 (
      {stage0_21[63]},
      {stage1_21[32]}
   );
   gpc1_1 gpc508 (
      {stage0_22[52]},
      {stage1_22[19]}
   );
   gpc1_1 gpc509 (
      {stage0_22[53]},
      {stage1_22[20]}
   );
   gpc1_1 gpc510 (
      {stage0_22[54]},
      {stage1_22[21]}
   );
   gpc1_1 gpc511 (
      {stage0_22[55]},
      {stage1_22[22]}
   );
   gpc1_1 gpc512 (
      {stage0_22[56]},
      {stage1_22[23]}
   );
   gpc1_1 gpc513 (
      {stage0_22[57]},
      {stage1_22[24]}
   );
   gpc1_1 gpc514 (
      {stage0_22[58]},
      {stage1_22[25]}
   );
   gpc1_1 gpc515 (
      {stage0_22[59]},
      {stage1_22[26]}
   );
   gpc1_1 gpc516 (
      {stage0_22[60]},
      {stage1_22[27]}
   );
   gpc1_1 gpc517 (
      {stage0_22[61]},
      {stage1_22[28]}
   );
   gpc1_1 gpc518 (
      {stage0_22[62]},
      {stage1_22[29]}
   );
   gpc1_1 gpc519 (
      {stage0_22[63]},
      {stage1_22[30]}
   );
   gpc1_1 gpc520 (
      {stage0_23[48]},
      {stage1_23[19]}
   );
   gpc1_1 gpc521 (
      {stage0_23[49]},
      {stage1_23[20]}
   );
   gpc1_1 gpc522 (
      {stage0_23[50]},
      {stage1_23[21]}
   );
   gpc1_1 gpc523 (
      {stage0_23[51]},
      {stage1_23[22]}
   );
   gpc1_1 gpc524 (
      {stage0_23[52]},
      {stage1_23[23]}
   );
   gpc1_1 gpc525 (
      {stage0_23[53]},
      {stage1_23[24]}
   );
   gpc1_1 gpc526 (
      {stage0_23[54]},
      {stage1_23[25]}
   );
   gpc1_1 gpc527 (
      {stage0_23[55]},
      {stage1_23[26]}
   );
   gpc1_1 gpc528 (
      {stage0_23[56]},
      {stage1_23[27]}
   );
   gpc1_1 gpc529 (
      {stage0_23[57]},
      {stage1_23[28]}
   );
   gpc1_1 gpc530 (
      {stage0_23[58]},
      {stage1_23[29]}
   );
   gpc1_1 gpc531 (
      {stage0_23[59]},
      {stage1_23[30]}
   );
   gpc1_1 gpc532 (
      {stage0_23[60]},
      {stage1_23[31]}
   );
   gpc1_1 gpc533 (
      {stage0_23[61]},
      {stage1_23[32]}
   );
   gpc1_1 gpc534 (
      {stage0_23[62]},
      {stage1_23[33]}
   );
   gpc1_1 gpc535 (
      {stage0_23[63]},
      {stage1_23[34]}
   );
   gpc1_1 gpc536 (
      {stage0_24[62]},
      {stage1_24[25]}
   );
   gpc1_1 gpc537 (
      {stage0_24[63]},
      {stage1_24[26]}
   );
   gpc1_1 gpc538 (
      {stage0_25[42]},
      {stage1_25[23]}
   );
   gpc1_1 gpc539 (
      {stage0_25[43]},
      {stage1_25[24]}
   );
   gpc1_1 gpc540 (
      {stage0_25[44]},
      {stage1_25[25]}
   );
   gpc1_1 gpc541 (
      {stage0_25[45]},
      {stage1_25[26]}
   );
   gpc1_1 gpc542 (
      {stage0_25[46]},
      {stage1_25[27]}
   );
   gpc1_1 gpc543 (
      {stage0_25[47]},
      {stage1_25[28]}
   );
   gpc1_1 gpc544 (
      {stage0_25[48]},
      {stage1_25[29]}
   );
   gpc1_1 gpc545 (
      {stage0_25[49]},
      {stage1_25[30]}
   );
   gpc1_1 gpc546 (
      {stage0_25[50]},
      {stage1_25[31]}
   );
   gpc1_1 gpc547 (
      {stage0_25[51]},
      {stage1_25[32]}
   );
   gpc1_1 gpc548 (
      {stage0_25[52]},
      {stage1_25[33]}
   );
   gpc1_1 gpc549 (
      {stage0_25[53]},
      {stage1_25[34]}
   );
   gpc1_1 gpc550 (
      {stage0_25[54]},
      {stage1_25[35]}
   );
   gpc1_1 gpc551 (
      {stage0_25[55]},
      {stage1_25[36]}
   );
   gpc1_1 gpc552 (
      {stage0_25[56]},
      {stage1_25[37]}
   );
   gpc1_1 gpc553 (
      {stage0_25[57]},
      {stage1_25[38]}
   );
   gpc1_1 gpc554 (
      {stage0_25[58]},
      {stage1_25[39]}
   );
   gpc1_1 gpc555 (
      {stage0_25[59]},
      {stage1_25[40]}
   );
   gpc1_1 gpc556 (
      {stage0_25[60]},
      {stage1_25[41]}
   );
   gpc1_1 gpc557 (
      {stage0_25[61]},
      {stage1_25[42]}
   );
   gpc1_1 gpc558 (
      {stage0_25[62]},
      {stage1_25[43]}
   );
   gpc1_1 gpc559 (
      {stage0_25[63]},
      {stage1_25[44]}
   );
   gpc1_1 gpc560 (
      {stage0_26[53]},
      {stage1_26[18]}
   );
   gpc1_1 gpc561 (
      {stage0_26[54]},
      {stage1_26[19]}
   );
   gpc1_1 gpc562 (
      {stage0_26[55]},
      {stage1_26[20]}
   );
   gpc1_1 gpc563 (
      {stage0_26[56]},
      {stage1_26[21]}
   );
   gpc1_1 gpc564 (
      {stage0_26[57]},
      {stage1_26[22]}
   );
   gpc1_1 gpc565 (
      {stage0_26[58]},
      {stage1_26[23]}
   );
   gpc1_1 gpc566 (
      {stage0_26[59]},
      {stage1_26[24]}
   );
   gpc1_1 gpc567 (
      {stage0_26[60]},
      {stage1_26[25]}
   );
   gpc1_1 gpc568 (
      {stage0_26[61]},
      {stage1_26[26]}
   );
   gpc1_1 gpc569 (
      {stage0_26[62]},
      {stage1_26[27]}
   );
   gpc1_1 gpc570 (
      {stage0_26[63]},
      {stage1_26[28]}
   );
   gpc1_1 gpc571 (
      {stage0_27[41]},
      {stage1_27[18]}
   );
   gpc1_1 gpc572 (
      {stage0_27[42]},
      {stage1_27[19]}
   );
   gpc1_1 gpc573 (
      {stage0_27[43]},
      {stage1_27[20]}
   );
   gpc1_1 gpc574 (
      {stage0_27[44]},
      {stage1_27[21]}
   );
   gpc1_1 gpc575 (
      {stage0_27[45]},
      {stage1_27[22]}
   );
   gpc1_1 gpc576 (
      {stage0_27[46]},
      {stage1_27[23]}
   );
   gpc1_1 gpc577 (
      {stage0_27[47]},
      {stage1_27[24]}
   );
   gpc1_1 gpc578 (
      {stage0_27[48]},
      {stage1_27[25]}
   );
   gpc1_1 gpc579 (
      {stage0_27[49]},
      {stage1_27[26]}
   );
   gpc1_1 gpc580 (
      {stage0_27[50]},
      {stage1_27[27]}
   );
   gpc1_1 gpc581 (
      {stage0_27[51]},
      {stage1_27[28]}
   );
   gpc1_1 gpc582 (
      {stage0_27[52]},
      {stage1_27[29]}
   );
   gpc1_1 gpc583 (
      {stage0_27[53]},
      {stage1_27[30]}
   );
   gpc1_1 gpc584 (
      {stage0_27[54]},
      {stage1_27[31]}
   );
   gpc1_1 gpc585 (
      {stage0_27[55]},
      {stage1_27[32]}
   );
   gpc1_1 gpc586 (
      {stage0_27[56]},
      {stage1_27[33]}
   );
   gpc1_1 gpc587 (
      {stage0_27[57]},
      {stage1_27[34]}
   );
   gpc1_1 gpc588 (
      {stage0_27[58]},
      {stage1_27[35]}
   );
   gpc1_1 gpc589 (
      {stage0_27[59]},
      {stage1_27[36]}
   );
   gpc1_1 gpc590 (
      {stage0_27[60]},
      {stage1_27[37]}
   );
   gpc1_1 gpc591 (
      {stage0_27[61]},
      {stage1_27[38]}
   );
   gpc1_1 gpc592 (
      {stage0_27[62]},
      {stage1_27[39]}
   );
   gpc1_1 gpc593 (
      {stage0_27[63]},
      {stage1_27[40]}
   );
   gpc1_1 gpc594 (
      {stage0_28[62]},
      {stage1_28[25]}
   );
   gpc1_1 gpc595 (
      {stage0_28[63]},
      {stage1_28[26]}
   );
   gpc1_1 gpc596 (
      {stage0_29[60]},
      {stage1_29[25]}
   );
   gpc1_1 gpc597 (
      {stage0_29[61]},
      {stage1_29[26]}
   );
   gpc1_1 gpc598 (
      {stage0_29[62]},
      {stage1_29[27]}
   );
   gpc1_1 gpc599 (
      {stage0_29[63]},
      {stage1_29[28]}
   );
   gpc1_1 gpc600 (
      {stage0_30[59]},
      {stage1_30[21]}
   );
   gpc1_1 gpc601 (
      {stage0_30[60]},
      {stage1_30[22]}
   );
   gpc1_1 gpc602 (
      {stage0_30[61]},
      {stage1_30[23]}
   );
   gpc1_1 gpc603 (
      {stage0_30[62]},
      {stage1_30[24]}
   );
   gpc1_1 gpc604 (
      {stage0_30[63]},
      {stage1_30[25]}
   );
   gpc1_1 gpc605 (
      {stage0_32[63]},
      {stage1_32[30]}
   );
   gpc1_1 gpc606 (
      {stage0_33[53]},
      {stage1_33[27]}
   );
   gpc1_1 gpc607 (
      {stage0_33[54]},
      {stage1_33[28]}
   );
   gpc1_1 gpc608 (
      {stage0_33[55]},
      {stage1_33[29]}
   );
   gpc1_1 gpc609 (
      {stage0_33[56]},
      {stage1_33[30]}
   );
   gpc1_1 gpc610 (
      {stage0_33[57]},
      {stage1_33[31]}
   );
   gpc1_1 gpc611 (
      {stage0_33[58]},
      {stage1_33[32]}
   );
   gpc1_1 gpc612 (
      {stage0_33[59]},
      {stage1_33[33]}
   );
   gpc1_1 gpc613 (
      {stage0_33[60]},
      {stage1_33[34]}
   );
   gpc1_1 gpc614 (
      {stage0_33[61]},
      {stage1_33[35]}
   );
   gpc1_1 gpc615 (
      {stage0_33[62]},
      {stage1_33[36]}
   );
   gpc1_1 gpc616 (
      {stage0_33[63]},
      {stage1_33[37]}
   );
   gpc1_1 gpc617 (
      {stage0_34[60]},
      {stage1_34[20]}
   );
   gpc1_1 gpc618 (
      {stage0_34[61]},
      {stage1_34[21]}
   );
   gpc1_1 gpc619 (
      {stage0_34[62]},
      {stage1_34[22]}
   );
   gpc1_1 gpc620 (
      {stage0_34[63]},
      {stage1_34[23]}
   );
   gpc1_1 gpc621 (
      {stage0_35[57]},
      {stage1_35[23]}
   );
   gpc1_1 gpc622 (
      {stage0_35[58]},
      {stage1_35[24]}
   );
   gpc1_1 gpc623 (
      {stage0_35[59]},
      {stage1_35[25]}
   );
   gpc1_1 gpc624 (
      {stage0_35[60]},
      {stage1_35[26]}
   );
   gpc1_1 gpc625 (
      {stage0_35[61]},
      {stage1_35[27]}
   );
   gpc1_1 gpc626 (
      {stage0_35[62]},
      {stage1_35[28]}
   );
   gpc1_1 gpc627 (
      {stage0_35[63]},
      {stage1_35[29]}
   );
   gpc1_1 gpc628 (
      {stage0_36[46]},
      {stage1_36[26]}
   );
   gpc1_1 gpc629 (
      {stage0_36[47]},
      {stage1_36[27]}
   );
   gpc1_1 gpc630 (
      {stage0_36[48]},
      {stage1_36[28]}
   );
   gpc1_1 gpc631 (
      {stage0_36[49]},
      {stage1_36[29]}
   );
   gpc1_1 gpc632 (
      {stage0_36[50]},
      {stage1_36[30]}
   );
   gpc1_1 gpc633 (
      {stage0_36[51]},
      {stage1_36[31]}
   );
   gpc1_1 gpc634 (
      {stage0_36[52]},
      {stage1_36[32]}
   );
   gpc1_1 gpc635 (
      {stage0_36[53]},
      {stage1_36[33]}
   );
   gpc1_1 gpc636 (
      {stage0_36[54]},
      {stage1_36[34]}
   );
   gpc1_1 gpc637 (
      {stage0_36[55]},
      {stage1_36[35]}
   );
   gpc1_1 gpc638 (
      {stage0_36[56]},
      {stage1_36[36]}
   );
   gpc1_1 gpc639 (
      {stage0_36[57]},
      {stage1_36[37]}
   );
   gpc1_1 gpc640 (
      {stage0_36[58]},
      {stage1_36[38]}
   );
   gpc1_1 gpc641 (
      {stage0_36[59]},
      {stage1_36[39]}
   );
   gpc1_1 gpc642 (
      {stage0_36[60]},
      {stage1_36[40]}
   );
   gpc1_1 gpc643 (
      {stage0_36[61]},
      {stage1_36[41]}
   );
   gpc1_1 gpc644 (
      {stage0_36[62]},
      {stage1_36[42]}
   );
   gpc1_1 gpc645 (
      {stage0_36[63]},
      {stage1_36[43]}
   );
   gpc1_1 gpc646 (
      {stage0_38[41]},
      {stage1_38[19]}
   );
   gpc1_1 gpc647 (
      {stage0_38[42]},
      {stage1_38[20]}
   );
   gpc1_1 gpc648 (
      {stage0_38[43]},
      {stage1_38[21]}
   );
   gpc1_1 gpc649 (
      {stage0_38[44]},
      {stage1_38[22]}
   );
   gpc1_1 gpc650 (
      {stage0_38[45]},
      {stage1_38[23]}
   );
   gpc1_1 gpc651 (
      {stage0_38[46]},
      {stage1_38[24]}
   );
   gpc1_1 gpc652 (
      {stage0_38[47]},
      {stage1_38[25]}
   );
   gpc1_1 gpc653 (
      {stage0_38[48]},
      {stage1_38[26]}
   );
   gpc1_1 gpc654 (
      {stage0_38[49]},
      {stage1_38[27]}
   );
   gpc1_1 gpc655 (
      {stage0_38[50]},
      {stage1_38[28]}
   );
   gpc1_1 gpc656 (
      {stage0_38[51]},
      {stage1_38[29]}
   );
   gpc1_1 gpc657 (
      {stage0_38[52]},
      {stage1_38[30]}
   );
   gpc1_1 gpc658 (
      {stage0_38[53]},
      {stage1_38[31]}
   );
   gpc1_1 gpc659 (
      {stage0_38[54]},
      {stage1_38[32]}
   );
   gpc1_1 gpc660 (
      {stage0_38[55]},
      {stage1_38[33]}
   );
   gpc1_1 gpc661 (
      {stage0_38[56]},
      {stage1_38[34]}
   );
   gpc1_1 gpc662 (
      {stage0_38[57]},
      {stage1_38[35]}
   );
   gpc1_1 gpc663 (
      {stage0_38[58]},
      {stage1_38[36]}
   );
   gpc1_1 gpc664 (
      {stage0_38[59]},
      {stage1_38[37]}
   );
   gpc1_1 gpc665 (
      {stage0_38[60]},
      {stage1_38[38]}
   );
   gpc1_1 gpc666 (
      {stage0_38[61]},
      {stage1_38[39]}
   );
   gpc1_1 gpc667 (
      {stage0_38[62]},
      {stage1_38[40]}
   );
   gpc1_1 gpc668 (
      {stage0_38[63]},
      {stage1_38[41]}
   );
   gpc1_1 gpc669 (
      {stage0_39[63]},
      {stage1_39[22]}
   );
   gpc1_1 gpc670 (
      {stage0_41[54]},
      {stage1_41[26]}
   );
   gpc1_1 gpc671 (
      {stage0_41[55]},
      {stage1_41[27]}
   );
   gpc1_1 gpc672 (
      {stage0_41[56]},
      {stage1_41[28]}
   );
   gpc1_1 gpc673 (
      {stage0_41[57]},
      {stage1_41[29]}
   );
   gpc1_1 gpc674 (
      {stage0_41[58]},
      {stage1_41[30]}
   );
   gpc1_1 gpc675 (
      {stage0_41[59]},
      {stage1_41[31]}
   );
   gpc1_1 gpc676 (
      {stage0_41[60]},
      {stage1_41[32]}
   );
   gpc1_1 gpc677 (
      {stage0_41[61]},
      {stage1_41[33]}
   );
   gpc1_1 gpc678 (
      {stage0_41[62]},
      {stage1_41[34]}
   );
   gpc1_1 gpc679 (
      {stage0_41[63]},
      {stage1_41[35]}
   );
   gpc1_1 gpc680 (
      {stage0_42[54]},
      {stage1_42[19]}
   );
   gpc1_1 gpc681 (
      {stage0_42[55]},
      {stage1_42[20]}
   );
   gpc1_1 gpc682 (
      {stage0_42[56]},
      {stage1_42[21]}
   );
   gpc1_1 gpc683 (
      {stage0_42[57]},
      {stage1_42[22]}
   );
   gpc1_1 gpc684 (
      {stage0_42[58]},
      {stage1_42[23]}
   );
   gpc1_1 gpc685 (
      {stage0_42[59]},
      {stage1_42[24]}
   );
   gpc1_1 gpc686 (
      {stage0_42[60]},
      {stage1_42[25]}
   );
   gpc1_1 gpc687 (
      {stage0_42[61]},
      {stage1_42[26]}
   );
   gpc1_1 gpc688 (
      {stage0_42[62]},
      {stage1_42[27]}
   );
   gpc1_1 gpc689 (
      {stage0_42[63]},
      {stage1_42[28]}
   );
   gpc1_1 gpc690 (
      {stage0_43[50]},
      {stage1_43[22]}
   );
   gpc1_1 gpc691 (
      {stage0_43[51]},
      {stage1_43[23]}
   );
   gpc1_1 gpc692 (
      {stage0_43[52]},
      {stage1_43[24]}
   );
   gpc1_1 gpc693 (
      {stage0_43[53]},
      {stage1_43[25]}
   );
   gpc1_1 gpc694 (
      {stage0_43[54]},
      {stage1_43[26]}
   );
   gpc1_1 gpc695 (
      {stage0_43[55]},
      {stage1_43[27]}
   );
   gpc1_1 gpc696 (
      {stage0_43[56]},
      {stage1_43[28]}
   );
   gpc1_1 gpc697 (
      {stage0_43[57]},
      {stage1_43[29]}
   );
   gpc1_1 gpc698 (
      {stage0_43[58]},
      {stage1_43[30]}
   );
   gpc1_1 gpc699 (
      {stage0_43[59]},
      {stage1_43[31]}
   );
   gpc1_1 gpc700 (
      {stage0_43[60]},
      {stage1_43[32]}
   );
   gpc1_1 gpc701 (
      {stage0_43[61]},
      {stage1_43[33]}
   );
   gpc1_1 gpc702 (
      {stage0_43[62]},
      {stage1_43[34]}
   );
   gpc1_1 gpc703 (
      {stage0_43[63]},
      {stage1_43[35]}
   );
   gpc1_1 gpc704 (
      {stage0_44[58]},
      {stage1_44[27]}
   );
   gpc1_1 gpc705 (
      {stage0_44[59]},
      {stage1_44[28]}
   );
   gpc1_1 gpc706 (
      {stage0_44[60]},
      {stage1_44[29]}
   );
   gpc1_1 gpc707 (
      {stage0_44[61]},
      {stage1_44[30]}
   );
   gpc1_1 gpc708 (
      {stage0_44[62]},
      {stage1_44[31]}
   );
   gpc1_1 gpc709 (
      {stage0_44[63]},
      {stage1_44[32]}
   );
   gpc1_1 gpc710 (
      {stage0_45[36]},
      {stage1_45[20]}
   );
   gpc1_1 gpc711 (
      {stage0_45[37]},
      {stage1_45[21]}
   );
   gpc1_1 gpc712 (
      {stage0_45[38]},
      {stage1_45[22]}
   );
   gpc1_1 gpc713 (
      {stage0_45[39]},
      {stage1_45[23]}
   );
   gpc1_1 gpc714 (
      {stage0_45[40]},
      {stage1_45[24]}
   );
   gpc1_1 gpc715 (
      {stage0_45[41]},
      {stage1_45[25]}
   );
   gpc1_1 gpc716 (
      {stage0_45[42]},
      {stage1_45[26]}
   );
   gpc1_1 gpc717 (
      {stage0_45[43]},
      {stage1_45[27]}
   );
   gpc1_1 gpc718 (
      {stage0_45[44]},
      {stage1_45[28]}
   );
   gpc1_1 gpc719 (
      {stage0_45[45]},
      {stage1_45[29]}
   );
   gpc1_1 gpc720 (
      {stage0_45[46]},
      {stage1_45[30]}
   );
   gpc1_1 gpc721 (
      {stage0_45[47]},
      {stage1_45[31]}
   );
   gpc1_1 gpc722 (
      {stage0_45[48]},
      {stage1_45[32]}
   );
   gpc1_1 gpc723 (
      {stage0_45[49]},
      {stage1_45[33]}
   );
   gpc1_1 gpc724 (
      {stage0_45[50]},
      {stage1_45[34]}
   );
   gpc1_1 gpc725 (
      {stage0_45[51]},
      {stage1_45[35]}
   );
   gpc1_1 gpc726 (
      {stage0_45[52]},
      {stage1_45[36]}
   );
   gpc1_1 gpc727 (
      {stage0_45[53]},
      {stage1_45[37]}
   );
   gpc1_1 gpc728 (
      {stage0_45[54]},
      {stage1_45[38]}
   );
   gpc1_1 gpc729 (
      {stage0_45[55]},
      {stage1_45[39]}
   );
   gpc1_1 gpc730 (
      {stage0_45[56]},
      {stage1_45[40]}
   );
   gpc1_1 gpc731 (
      {stage0_45[57]},
      {stage1_45[41]}
   );
   gpc1_1 gpc732 (
      {stage0_45[58]},
      {stage1_45[42]}
   );
   gpc1_1 gpc733 (
      {stage0_45[59]},
      {stage1_45[43]}
   );
   gpc1_1 gpc734 (
      {stage0_45[60]},
      {stage1_45[44]}
   );
   gpc1_1 gpc735 (
      {stage0_45[61]},
      {stage1_45[45]}
   );
   gpc1_1 gpc736 (
      {stage0_45[62]},
      {stage1_45[46]}
   );
   gpc1_1 gpc737 (
      {stage0_45[63]},
      {stage1_45[47]}
   );
   gpc1_1 gpc738 (
      {stage0_47[46]},
      {stage1_47[23]}
   );
   gpc1_1 gpc739 (
      {stage0_47[47]},
      {stage1_47[24]}
   );
   gpc1_1 gpc740 (
      {stage0_47[48]},
      {stage1_47[25]}
   );
   gpc1_1 gpc741 (
      {stage0_47[49]},
      {stage1_47[26]}
   );
   gpc1_1 gpc742 (
      {stage0_47[50]},
      {stage1_47[27]}
   );
   gpc1_1 gpc743 (
      {stage0_47[51]},
      {stage1_47[28]}
   );
   gpc1_1 gpc744 (
      {stage0_47[52]},
      {stage1_47[29]}
   );
   gpc1_1 gpc745 (
      {stage0_47[53]},
      {stage1_47[30]}
   );
   gpc1_1 gpc746 (
      {stage0_47[54]},
      {stage1_47[31]}
   );
   gpc1_1 gpc747 (
      {stage0_47[55]},
      {stage1_47[32]}
   );
   gpc1_1 gpc748 (
      {stage0_47[56]},
      {stage1_47[33]}
   );
   gpc1_1 gpc749 (
      {stage0_47[57]},
      {stage1_47[34]}
   );
   gpc1_1 gpc750 (
      {stage0_47[58]},
      {stage1_47[35]}
   );
   gpc1_1 gpc751 (
      {stage0_47[59]},
      {stage1_47[36]}
   );
   gpc1_1 gpc752 (
      {stage0_47[60]},
      {stage1_47[37]}
   );
   gpc1_1 gpc753 (
      {stage0_47[61]},
      {stage1_47[38]}
   );
   gpc1_1 gpc754 (
      {stage0_47[62]},
      {stage1_47[39]}
   );
   gpc1_1 gpc755 (
      {stage0_47[63]},
      {stage1_47[40]}
   );
   gpc1_1 gpc756 (
      {stage0_48[58]},
      {stage1_48[26]}
   );
   gpc1_1 gpc757 (
      {stage0_48[59]},
      {stage1_48[27]}
   );
   gpc1_1 gpc758 (
      {stage0_48[60]},
      {stage1_48[28]}
   );
   gpc1_1 gpc759 (
      {stage0_48[61]},
      {stage1_48[29]}
   );
   gpc1_1 gpc760 (
      {stage0_48[62]},
      {stage1_48[30]}
   );
   gpc1_1 gpc761 (
      {stage0_48[63]},
      {stage1_48[31]}
   );
   gpc1_1 gpc762 (
      {stage0_49[60]},
      {stage1_49[21]}
   );
   gpc1_1 gpc763 (
      {stage0_49[61]},
      {stage1_49[22]}
   );
   gpc1_1 gpc764 (
      {stage0_49[62]},
      {stage1_49[23]}
   );
   gpc1_1 gpc765 (
      {stage0_49[63]},
      {stage1_49[24]}
   );
   gpc1_1 gpc766 (
      {stage0_50[62]},
      {stage1_50[23]}
   );
   gpc1_1 gpc767 (
      {stage0_50[63]},
      {stage1_50[24]}
   );
   gpc1_1 gpc768 (
      {stage0_51[59]},
      {stage1_51[27]}
   );
   gpc1_1 gpc769 (
      {stage0_51[60]},
      {stage1_51[28]}
   );
   gpc1_1 gpc770 (
      {stage0_51[61]},
      {stage1_51[29]}
   );
   gpc1_1 gpc771 (
      {stage0_51[62]},
      {stage1_51[30]}
   );
   gpc1_1 gpc772 (
      {stage0_51[63]},
      {stage1_51[31]}
   );
   gpc1_1 gpc773 (
      {stage0_52[45]},
      {stage1_52[24]}
   );
   gpc1_1 gpc774 (
      {stage0_52[46]},
      {stage1_52[25]}
   );
   gpc1_1 gpc775 (
      {stage0_52[47]},
      {stage1_52[26]}
   );
   gpc1_1 gpc776 (
      {stage0_52[48]},
      {stage1_52[27]}
   );
   gpc1_1 gpc777 (
      {stage0_52[49]},
      {stage1_52[28]}
   );
   gpc1_1 gpc778 (
      {stage0_52[50]},
      {stage1_52[29]}
   );
   gpc1_1 gpc779 (
      {stage0_52[51]},
      {stage1_52[30]}
   );
   gpc1_1 gpc780 (
      {stage0_52[52]},
      {stage1_52[31]}
   );
   gpc1_1 gpc781 (
      {stage0_52[53]},
      {stage1_52[32]}
   );
   gpc1_1 gpc782 (
      {stage0_52[54]},
      {stage1_52[33]}
   );
   gpc1_1 gpc783 (
      {stage0_52[55]},
      {stage1_52[34]}
   );
   gpc1_1 gpc784 (
      {stage0_52[56]},
      {stage1_52[35]}
   );
   gpc1_1 gpc785 (
      {stage0_52[57]},
      {stage1_52[36]}
   );
   gpc1_1 gpc786 (
      {stage0_52[58]},
      {stage1_52[37]}
   );
   gpc1_1 gpc787 (
      {stage0_52[59]},
      {stage1_52[38]}
   );
   gpc1_1 gpc788 (
      {stage0_52[60]},
      {stage1_52[39]}
   );
   gpc1_1 gpc789 (
      {stage0_52[61]},
      {stage1_52[40]}
   );
   gpc1_1 gpc790 (
      {stage0_52[62]},
      {stage1_52[41]}
   );
   gpc1_1 gpc791 (
      {stage0_52[63]},
      {stage1_52[42]}
   );
   gpc1_1 gpc792 (
      {stage0_53[58]},
      {stage1_53[21]}
   );
   gpc1_1 gpc793 (
      {stage0_53[59]},
      {stage1_53[22]}
   );
   gpc1_1 gpc794 (
      {stage0_53[60]},
      {stage1_53[23]}
   );
   gpc1_1 gpc795 (
      {stage0_53[61]},
      {stage1_53[24]}
   );
   gpc1_1 gpc796 (
      {stage0_53[62]},
      {stage1_53[25]}
   );
   gpc1_1 gpc797 (
      {stage0_53[63]},
      {stage1_53[26]}
   );
   gpc1_1 gpc798 (
      {stage0_54[54]},
      {stage1_54[23]}
   );
   gpc1_1 gpc799 (
      {stage0_54[55]},
      {stage1_54[24]}
   );
   gpc1_1 gpc800 (
      {stage0_54[56]},
      {stage1_54[25]}
   );
   gpc1_1 gpc801 (
      {stage0_54[57]},
      {stage1_54[26]}
   );
   gpc1_1 gpc802 (
      {stage0_54[58]},
      {stage1_54[27]}
   );
   gpc1_1 gpc803 (
      {stage0_54[59]},
      {stage1_54[28]}
   );
   gpc1_1 gpc804 (
      {stage0_54[60]},
      {stage1_54[29]}
   );
   gpc1_1 gpc805 (
      {stage0_54[61]},
      {stage1_54[30]}
   );
   gpc1_1 gpc806 (
      {stage0_54[62]},
      {stage1_54[31]}
   );
   gpc1_1 gpc807 (
      {stage0_54[63]},
      {stage1_54[32]}
   );
   gpc1_1 gpc808 (
      {stage0_56[62]},
      {stage1_56[24]}
   );
   gpc1_1 gpc809 (
      {stage0_56[63]},
      {stage1_56[25]}
   );
   gpc1_1 gpc810 (
      {stage0_58[47]},
      {stage1_58[24]}
   );
   gpc1_1 gpc811 (
      {stage0_58[48]},
      {stage1_58[25]}
   );
   gpc1_1 gpc812 (
      {stage0_58[49]},
      {stage1_58[26]}
   );
   gpc1_1 gpc813 (
      {stage0_58[50]},
      {stage1_58[27]}
   );
   gpc1_1 gpc814 (
      {stage0_58[51]},
      {stage1_58[28]}
   );
   gpc1_1 gpc815 (
      {stage0_58[52]},
      {stage1_58[29]}
   );
   gpc1_1 gpc816 (
      {stage0_58[53]},
      {stage1_58[30]}
   );
   gpc1_1 gpc817 (
      {stage0_58[54]},
      {stage1_58[31]}
   );
   gpc1_1 gpc818 (
      {stage0_58[55]},
      {stage1_58[32]}
   );
   gpc1_1 gpc819 (
      {stage0_58[56]},
      {stage1_58[33]}
   );
   gpc1_1 gpc820 (
      {stage0_58[57]},
      {stage1_58[34]}
   );
   gpc1_1 gpc821 (
      {stage0_58[58]},
      {stage1_58[35]}
   );
   gpc1_1 gpc822 (
      {stage0_58[59]},
      {stage1_58[36]}
   );
   gpc1_1 gpc823 (
      {stage0_58[60]},
      {stage1_58[37]}
   );
   gpc1_1 gpc824 (
      {stage0_58[61]},
      {stage1_58[38]}
   );
   gpc1_1 gpc825 (
      {stage0_58[62]},
      {stage1_58[39]}
   );
   gpc1_1 gpc826 (
      {stage0_58[63]},
      {stage1_58[40]}
   );
   gpc1_1 gpc827 (
      {stage0_59[42]},
      {stage1_59[20]}
   );
   gpc1_1 gpc828 (
      {stage0_59[43]},
      {stage1_59[21]}
   );
   gpc1_1 gpc829 (
      {stage0_59[44]},
      {stage1_59[22]}
   );
   gpc1_1 gpc830 (
      {stage0_59[45]},
      {stage1_59[23]}
   );
   gpc1_1 gpc831 (
      {stage0_59[46]},
      {stage1_59[24]}
   );
   gpc1_1 gpc832 (
      {stage0_59[47]},
      {stage1_59[25]}
   );
   gpc1_1 gpc833 (
      {stage0_59[48]},
      {stage1_59[26]}
   );
   gpc1_1 gpc834 (
      {stage0_59[49]},
      {stage1_59[27]}
   );
   gpc1_1 gpc835 (
      {stage0_59[50]},
      {stage1_59[28]}
   );
   gpc1_1 gpc836 (
      {stage0_59[51]},
      {stage1_59[29]}
   );
   gpc1_1 gpc837 (
      {stage0_59[52]},
      {stage1_59[30]}
   );
   gpc1_1 gpc838 (
      {stage0_59[53]},
      {stage1_59[31]}
   );
   gpc1_1 gpc839 (
      {stage0_59[54]},
      {stage1_59[32]}
   );
   gpc1_1 gpc840 (
      {stage0_59[55]},
      {stage1_59[33]}
   );
   gpc1_1 gpc841 (
      {stage0_59[56]},
      {stage1_59[34]}
   );
   gpc1_1 gpc842 (
      {stage0_59[57]},
      {stage1_59[35]}
   );
   gpc1_1 gpc843 (
      {stage0_59[58]},
      {stage1_59[36]}
   );
   gpc1_1 gpc844 (
      {stage0_59[59]},
      {stage1_59[37]}
   );
   gpc1_1 gpc845 (
      {stage0_59[60]},
      {stage1_59[38]}
   );
   gpc1_1 gpc846 (
      {stage0_59[61]},
      {stage1_59[39]}
   );
   gpc1_1 gpc847 (
      {stage0_59[62]},
      {stage1_59[40]}
   );
   gpc1_1 gpc848 (
      {stage0_59[63]},
      {stage1_59[41]}
   );
   gpc1_1 gpc849 (
      {stage0_60[52]},
      {stage1_60[21]}
   );
   gpc1_1 gpc850 (
      {stage0_60[53]},
      {stage1_60[22]}
   );
   gpc1_1 gpc851 (
      {stage0_60[54]},
      {stage1_60[23]}
   );
   gpc1_1 gpc852 (
      {stage0_60[55]},
      {stage1_60[24]}
   );
   gpc1_1 gpc853 (
      {stage0_60[56]},
      {stage1_60[25]}
   );
   gpc1_1 gpc854 (
      {stage0_60[57]},
      {stage1_60[26]}
   );
   gpc1_1 gpc855 (
      {stage0_60[58]},
      {stage1_60[27]}
   );
   gpc1_1 gpc856 (
      {stage0_60[59]},
      {stage1_60[28]}
   );
   gpc1_1 gpc857 (
      {stage0_60[60]},
      {stage1_60[29]}
   );
   gpc1_1 gpc858 (
      {stage0_60[61]},
      {stage1_60[30]}
   );
   gpc1_1 gpc859 (
      {stage0_60[62]},
      {stage1_60[31]}
   );
   gpc1_1 gpc860 (
      {stage0_60[63]},
      {stage1_60[32]}
   );
   gpc1_1 gpc861 (
      {stage0_61[58]},
      {stage1_61[25]}
   );
   gpc1_1 gpc862 (
      {stage0_61[59]},
      {stage1_61[26]}
   );
   gpc1_1 gpc863 (
      {stage0_61[60]},
      {stage1_61[27]}
   );
   gpc1_1 gpc864 (
      {stage0_61[61]},
      {stage1_61[28]}
   );
   gpc1_1 gpc865 (
      {stage0_61[62]},
      {stage1_61[29]}
   );
   gpc1_1 gpc866 (
      {stage0_61[63]},
      {stage1_61[30]}
   );
   gpc1_1 gpc867 (
      {stage0_62[51]},
      {stage1_62[20]}
   );
   gpc1_1 gpc868 (
      {stage0_62[52]},
      {stage1_62[21]}
   );
   gpc1_1 gpc869 (
      {stage0_62[53]},
      {stage1_62[22]}
   );
   gpc1_1 gpc870 (
      {stage0_62[54]},
      {stage1_62[23]}
   );
   gpc1_1 gpc871 (
      {stage0_62[55]},
      {stage1_62[24]}
   );
   gpc1_1 gpc872 (
      {stage0_62[56]},
      {stage1_62[25]}
   );
   gpc1_1 gpc873 (
      {stage0_62[57]},
      {stage1_62[26]}
   );
   gpc1_1 gpc874 (
      {stage0_62[58]},
      {stage1_62[27]}
   );
   gpc1_1 gpc875 (
      {stage0_62[59]},
      {stage1_62[28]}
   );
   gpc1_1 gpc876 (
      {stage0_62[60]},
      {stage1_62[29]}
   );
   gpc1_1 gpc877 (
      {stage0_62[61]},
      {stage1_62[30]}
   );
   gpc1_1 gpc878 (
      {stage0_62[62]},
      {stage1_62[31]}
   );
   gpc1_1 gpc879 (
      {stage0_62[63]},
      {stage1_62[32]}
   );
   gpc1_1 gpc880 (
      {stage0_63[54]},
      {stage1_63[18]}
   );
   gpc1_1 gpc881 (
      {stage0_63[55]},
      {stage1_63[19]}
   );
   gpc1_1 gpc882 (
      {stage0_63[56]},
      {stage1_63[20]}
   );
   gpc1_1 gpc883 (
      {stage0_63[57]},
      {stage1_63[21]}
   );
   gpc1_1 gpc884 (
      {stage0_63[58]},
      {stage1_63[22]}
   );
   gpc1_1 gpc885 (
      {stage0_63[59]},
      {stage1_63[23]}
   );
   gpc1_1 gpc886 (
      {stage0_63[60]},
      {stage1_63[24]}
   );
   gpc1_1 gpc887 (
      {stage0_63[61]},
      {stage1_63[25]}
   );
   gpc1_1 gpc888 (
      {stage0_63[62]},
      {stage1_63[26]}
   );
   gpc1_1 gpc889 (
      {stage0_63[63]},
      {stage1_63[27]}
   );
   gpc1163_5 gpc890 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc891 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc892 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc893 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc894 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc895 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], 1'b0, 1'b0},
      {stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc606_5 gpc896 (
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_3[5], stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10]},
      {stage2_5[0],stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6]}
   );
   gpc606_5 gpc897 (
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage2_5[1],stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7]}
   );
   gpc606_5 gpc898 (
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22]},
      {stage2_5[2],stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8]}
   );
   gpc606_5 gpc899 (
      {stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[3],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc606_5 gpc900 (
      {stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[4],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc615_5 gpc901 (
      {stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage1_4[12]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[2],stage2_5[5],stage2_4[11],stage2_3[11]}
   );
   gpc1163_5 gpc902 (
      {stage1_4[13], stage1_4[14], stage1_4[15]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[1],stage2_6[3],stage2_5[6],stage2_4[12]}
   );
   gpc606_5 gpc903 (
      {stage1_4[16], stage1_4[17], stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[2],stage2_6[4],stage2_5[7],stage2_4[13]}
   );
   gpc1325_5 gpc904 (
      {stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage1_5[12], stage1_5[13]},
      {stage1_6[7], stage1_6[8], stage1_6[9]},
      {stage1_7[1]},
      {stage2_8[2],stage2_7[3],stage2_6[5],stage2_5[8],stage2_4[14]}
   );
   gpc615_5 gpc905 (
      {stage1_6[10], stage1_6[11], stage1_6[12], stage1_6[13], stage1_6[14]},
      {stage1_7[2]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[3],stage2_7[4],stage2_6[6]}
   );
   gpc117_4 gpc906 (
      {stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9]},
      {stage1_8[6]},
      {stage1_9[0]},
      {stage2_10[1],stage2_9[1],stage2_8[4],stage2_7[5]}
   );
   gpc615_5 gpc907 (
      {stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13], stage1_7[14]},
      {stage1_8[7]},
      {stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5], stage1_9[6]},
      {stage2_11[0],stage2_10[2],stage2_9[2],stage2_8[5],stage2_7[6]}
   );
   gpc615_5 gpc908 (
      {stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18], stage1_7[19]},
      {stage1_8[8]},
      {stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11], stage1_9[12]},
      {stage2_11[1],stage2_10[3],stage2_9[3],stage2_8[6],stage2_7[7]}
   );
   gpc615_5 gpc909 (
      {stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24]},
      {stage1_8[9]},
      {stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17], stage1_9[18]},
      {stage2_11[2],stage2_10[4],stage2_9[4],stage2_8[7],stage2_7[8]}
   );
   gpc606_5 gpc910 (
      {stage1_8[10], stage1_8[11], stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[3],stage2_10[5],stage2_9[5],stage2_8[8]}
   );
   gpc606_5 gpc911 (
      {stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23], stage1_9[24]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[1],stage2_11[4],stage2_10[6],stage2_9[6]}
   );
   gpc615_5 gpc912 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10]},
      {stage1_11[6]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[2],stage2_11[5],stage2_10[7]}
   );
   gpc615_5 gpc913 (
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[1],stage2_13[2],stage2_12[3],stage2_11[6]}
   );
   gpc615_5 gpc914 (
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16]},
      {stage1_12[7]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[2],stage2_13[3],stage2_12[4],stage2_11[7]}
   );
   gpc615_5 gpc915 (
      {stage1_11[17], stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21]},
      {stage1_12[8]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[3],stage2_13[4],stage2_12[5],stage2_11[8]}
   );
   gpc615_5 gpc916 (
      {stage1_11[22], stage1_11[23], stage1_11[24], stage1_11[25], stage1_11[26]},
      {stage1_12[9]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[4],stage2_13[5],stage2_12[6],stage2_11[9]}
   );
   gpc606_5 gpc917 (
      {stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[4],stage2_14[5],stage2_13[6],stage2_12[7]}
   );
   gpc615_5 gpc918 (
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28]},
      {stage1_14[6]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[1],stage2_15[5],stage2_14[6],stage2_13[7]}
   );
   gpc615_5 gpc919 (
      {stage1_13[29], stage1_13[30], 1'b0, 1'b0, 1'b0},
      {stage1_14[7]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[2],stage2_15[6],stage2_14[7],stage2_13[8]}
   );
   gpc606_5 gpc920 (
      {stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12], stage1_14[13]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[2],stage2_16[3],stage2_15[7],stage2_14[8]}
   );
   gpc615_5 gpc921 (
      {stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18]},
      {stage1_15[12]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[3],stage2_16[4],stage2_15[8],stage2_14[9]}
   );
   gpc615_5 gpc922 (
      {stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_16[12]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[4],stage2_16[5],stage2_15[9]}
   );
   gpc615_5 gpc923 (
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22]},
      {stage1_16[13]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[3],stage2_17[5],stage2_16[6],stage2_15[10]}
   );
   gpc615_5 gpc924 (
      {stage1_15[23], stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27]},
      {stage1_16[14]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[4],stage2_17[6],stage2_16[7],stage2_15[11]}
   );
   gpc615_5 gpc925 (
      {stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31], stage1_15[32]},
      {stage1_16[15]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[5],stage2_17[7],stage2_16[8],stage2_15[12]}
   );
   gpc615_5 gpc926 (
      {stage1_15[33], stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37]},
      {stage1_16[16]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[6],stage2_17[8],stage2_16[9],stage2_15[13]}
   );
   gpc615_5 gpc927 (
      {stage1_16[17], stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21]},
      {stage1_17[30]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[5],stage2_18[7],stage2_17[9],stage2_16[10]}
   );
   gpc615_5 gpc928 (
      {stage1_16[22], stage1_16[23], stage1_16[24], stage1_16[25], stage1_16[26]},
      {stage1_17[31]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[6],stage2_18[8],stage2_17[10],stage2_16[11]}
   );
   gpc623_5 gpc929 (
      {stage1_17[32], stage1_17[33], stage1_17[34]},
      {stage1_18[12], stage1_18[13]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[7],stage2_18[9],stage2_17[11]}
   );
   gpc615_5 gpc930 (
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10]},
      {stage1_20[0]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[0],stage2_21[1],stage2_20[3],stage2_19[8]}
   );
   gpc615_5 gpc931 (
      {stage1_19[11], stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15]},
      {stage1_20[1]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[1],stage2_21[2],stage2_20[4],stage2_19[9]}
   );
   gpc615_5 gpc932 (
      {stage1_19[16], stage1_19[17], stage1_19[18], stage1_19[19], stage1_19[20]},
      {stage1_20[2]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[2],stage2_21[3],stage2_20[5],stage2_19[10]}
   );
   gpc615_5 gpc933 (
      {stage1_19[21], stage1_19[22], stage1_19[23], stage1_19[24], stage1_19[25]},
      {stage1_20[3]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[3],stage2_21[4],stage2_20[6],stage2_19[11]}
   );
   gpc606_5 gpc934 (
      {stage1_20[4], stage1_20[5], stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[4],stage2_22[4],stage2_21[5],stage2_20[7]}
   );
   gpc606_5 gpc935 (
      {stage1_20[10], stage1_20[11], stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[5],stage2_22[5],stage2_21[6],stage2_20[8]}
   );
   gpc606_5 gpc936 (
      {stage1_20[16], stage1_20[17], stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[6],stage2_22[6],stage2_21[7],stage2_20[9]}
   );
   gpc606_5 gpc937 (
      {stage1_20[22], stage1_20[23], stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[7],stage2_22[7],stage2_21[8],stage2_20[10]}
   );
   gpc606_5 gpc938 (
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[4],stage2_23[8],stage2_22[8],stage2_21[9]}
   );
   gpc1415_5 gpc939 (
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28]},
      {stage1_23[6]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3]},
      {stage1_25[0]},
      {stage2_26[0],stage2_25[1],stage2_24[5],stage2_23[9],stage2_22[9]}
   );
   gpc623_5 gpc940 (
      {stage1_22[29], stage1_22[30], 1'b0},
      {stage1_23[7], stage1_23[8]},
      {stage1_24[4], stage1_24[5], stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9]},
      {stage2_26[1],stage2_25[2],stage2_24[6],stage2_23[10],stage2_22[10]}
   );
   gpc615_5 gpc941 (
      {stage1_23[9], stage1_23[10], stage1_23[11], stage1_23[12], stage1_23[13]},
      {stage1_24[10]},
      {stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5], stage1_25[6]},
      {stage2_27[0],stage2_26[2],stage2_25[3],stage2_24[7],stage2_23[11]}
   );
   gpc615_5 gpc942 (
      {stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17], stage1_23[18]},
      {stage1_24[11]},
      {stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11], stage1_25[12]},
      {stage2_27[1],stage2_26[3],stage2_25[4],stage2_24[8],stage2_23[12]}
   );
   gpc615_5 gpc943 (
      {stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage1_24[12]},
      {stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17], stage1_25[18]},
      {stage2_27[2],stage2_26[4],stage2_25[5],stage2_24[9],stage2_23[13]}
   );
   gpc615_5 gpc944 (
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28]},
      {stage1_24[13]},
      {stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23], stage1_25[24]},
      {stage2_27[3],stage2_26[5],stage2_25[6],stage2_24[10],stage2_23[14]}
   );
   gpc615_5 gpc945 (
      {stage1_23[29], stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33]},
      {stage1_24[14]},
      {stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29], stage1_25[30]},
      {stage2_27[4],stage2_26[6],stage2_25[7],stage2_24[11],stage2_23[15]}
   );
   gpc606_5 gpc946 (
      {stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18], stage1_24[19], stage1_24[20]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[5],stage2_26[7],stage2_25[8],stage2_24[12]}
   );
   gpc606_5 gpc947 (
      {stage1_24[21], stage1_24[22], stage1_24[23], stage1_24[24], stage1_24[25], stage1_24[26]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[6],stage2_26[8],stage2_25[9],stage2_24[13]}
   );
   gpc606_5 gpc948 (
      {stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35], stage1_25[36]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[2],stage2_27[7],stage2_26[9],stage2_25[10]}
   );
   gpc606_5 gpc949 (
      {stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41], stage1_25[42]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[3],stage2_27[8],stage2_26[10],stage2_25[11]}
   );
   gpc615_5 gpc950 (
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16]},
      {stage1_27[12]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[2],stage2_28[4],stage2_27[9],stage2_26[11]}
   );
   gpc615_5 gpc951 (
      {stage1_26[17], stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21]},
      {stage1_27[13]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[3],stage2_28[5],stage2_27[10],stage2_26[12]}
   );
   gpc615_5 gpc952 (
      {stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17], stage1_27[18]},
      {stage1_28[12]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[2],stage2_29[4],stage2_28[6],stage2_27[11]}
   );
   gpc615_5 gpc953 (
      {stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage1_28[13]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[3],stage2_29[5],stage2_28[7],stage2_27[12]}
   );
   gpc615_5 gpc954 (
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28]},
      {stage1_28[14]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[4],stage2_29[6],stage2_28[8],stage2_27[13]}
   );
   gpc606_5 gpc955 (
      {stage1_28[15], stage1_28[16], stage1_28[17], stage1_28[18], stage1_28[19], stage1_28[20]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[3],stage2_30[5],stage2_29[7],stage2_28[9]}
   );
   gpc606_5 gpc956 (
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[1],stage2_31[4],stage2_30[6],stage2_29[8]}
   );
   gpc606_5 gpc957 (
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], 1'b0},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[2],stage2_31[5],stage2_30[7],stage2_29[9]}
   );
   gpc615_5 gpc958 (
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10]},
      {stage1_31[12]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[2],stage2_32[3],stage2_31[6],stage2_30[8]}
   );
   gpc615_5 gpc959 (
      {stage1_30[11], stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15]},
      {stage1_31[13]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[3],stage2_32[4],stage2_31[7],stage2_30[9]}
   );
   gpc615_5 gpc960 (
      {stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17], stage1_31[18]},
      {stage1_32[12]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[2],stage2_33[4],stage2_32[5],stage2_31[8]}
   );
   gpc606_5 gpc961 (
      {stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17], stage1_32[18]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[1],stage2_34[3],stage2_33[5],stage2_32[6]}
   );
   gpc606_5 gpc962 (
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[1],stage2_35[2],stage2_34[4],stage2_33[6]}
   );
   gpc606_5 gpc963 (
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[2],stage2_35[3],stage2_34[5],stage2_33[7]}
   );
   gpc606_5 gpc964 (
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[3],stage2_35[4],stage2_34[6],stage2_33[8]}
   );
   gpc615_5 gpc965 (
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10]},
      {stage1_35[18]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[3],stage2_36[4],stage2_35[5],stage2_34[7]}
   );
   gpc615_5 gpc966 (
      {stage1_34[11], stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15]},
      {stage1_35[19]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[4],stage2_36[5],stage2_35[6],stage2_34[8]}
   );
   gpc615_5 gpc967 (
      {stage1_34[16], stage1_34[17], stage1_34[18], stage1_34[19], stage1_34[20]},
      {stage1_35[20]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[5],stage2_36[6],stage2_35[7],stage2_34[9]}
   );
   gpc615_5 gpc968 (
      {stage1_35[21], stage1_35[22], stage1_35[23], stage1_35[24], stage1_35[25]},
      {stage1_36[18]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[3],stage2_37[6],stage2_36[7],stage2_35[8]}
   );
   gpc606_5 gpc969 (
      {stage1_36[19], stage1_36[20], stage1_36[21], stage1_36[22], stage1_36[23], stage1_36[24]},
      {stage1_38[0], stage1_38[1], stage1_38[2], stage1_38[3], stage1_38[4], stage1_38[5]},
      {stage2_40[0],stage2_39[1],stage2_38[4],stage2_37[7],stage2_36[8]}
   );
   gpc606_5 gpc970 (
      {stage1_36[25], stage1_36[26], stage1_36[27], stage1_36[28], stage1_36[29], stage1_36[30]},
      {stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10], stage1_38[11]},
      {stage2_40[1],stage2_39[2],stage2_38[5],stage2_37[8],stage2_36[9]}
   );
   gpc606_5 gpc971 (
      {stage1_36[31], stage1_36[32], stage1_36[33], stage1_36[34], stage1_36[35], stage1_36[36]},
      {stage1_38[12], stage1_38[13], stage1_38[14], stage1_38[15], stage1_38[16], stage1_38[17]},
      {stage2_40[2],stage2_39[3],stage2_38[6],stage2_37[9],stage2_36[10]}
   );
   gpc606_5 gpc972 (
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage2_41[0],stage2_40[3],stage2_39[4],stage2_38[7],stage2_37[10]}
   );
   gpc606_5 gpc973 (
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage1_39[6], stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11]},
      {stage2_41[1],stage2_40[4],stage2_39[5],stage2_38[8],stage2_37[11]}
   );
   gpc1406_5 gpc974 (
      {stage1_38[18], stage1_38[19], stage1_38[20], stage1_38[21], stage1_38[22], stage1_38[23]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3]},
      {stage1_41[0]},
      {stage2_42[0],stage2_41[2],stage2_40[5],stage2_39[6],stage2_38[9]}
   );
   gpc1325_5 gpc975 (
      {stage1_38[24], stage1_38[25], stage1_38[26], stage1_38[27], stage1_38[28]},
      {stage1_39[12], stage1_39[13]},
      {stage1_40[4], stage1_40[5], stage1_40[6]},
      {stage1_41[1]},
      {stage2_42[1],stage2_41[3],stage2_40[6],stage2_39[7],stage2_38[10]}
   );
   gpc615_5 gpc976 (
      {stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17], stage1_39[18]},
      {stage1_40[7]},
      {stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5], stage1_41[6], stage1_41[7]},
      {stage2_43[0],stage2_42[2],stage2_41[4],stage2_40[7],stage2_39[8]}
   );
   gpc606_5 gpc977 (
      {stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11], stage1_40[12], stage1_40[13]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[1],stage2_42[3],stage2_41[5],stage2_40[8]}
   );
   gpc606_5 gpc978 (
      {stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17], stage1_40[18], stage1_40[19]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[2],stage2_42[4],stage2_41[6],stage2_40[9]}
   );
   gpc606_5 gpc979 (
      {stage1_40[20], stage1_40[21], stage1_40[22], stage1_40[23], stage1_40[24], stage1_40[25]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[3],stage2_42[5],stage2_41[7],stage2_40[10]}
   );
   gpc7_3 gpc980 (
      {stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11], stage1_41[12], stage1_41[13], stage1_41[14]},
      {stage2_43[4],stage2_42[6],stage2_41[8]}
   );
   gpc606_5 gpc981 (
      {stage1_41[15], stage1_41[16], stage1_41[17], stage1_41[18], stage1_41[19], stage1_41[20]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[3],stage2_43[5],stage2_42[7],stage2_41[9]}
   );
   gpc606_5 gpc982 (
      {stage1_41[21], stage1_41[22], stage1_41[23], stage1_41[24], stage1_41[25], stage1_41[26]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[4],stage2_43[6],stage2_42[8],stage2_41[10]}
   );
   gpc606_5 gpc983 (
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage2_46[0],stage2_45[2],stage2_44[5],stage2_43[7],stage2_42[9]}
   );
   gpc615_5 gpc984 (
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16]},
      {stage1_44[6]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[1],stage2_45[3],stage2_44[6],stage2_43[8]}
   );
   gpc615_5 gpc985 (
      {stage1_43[17], stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21]},
      {stage1_44[7]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[2],stage2_45[4],stage2_44[7],stage2_43[9]}
   );
   gpc615_5 gpc986 (
      {stage1_43[22], stage1_43[23], stage1_43[24], stage1_43[25], stage1_43[26]},
      {stage1_44[8]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[3],stage2_45[5],stage2_44[8],stage2_43[10]}
   );
   gpc615_5 gpc987 (
      {stage1_43[27], stage1_43[28], stage1_43[29], stage1_43[30], stage1_43[31]},
      {stage1_44[9]},
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage2_47[3],stage2_46[4],stage2_45[6],stage2_44[9],stage2_43[11]}
   );
   gpc615_5 gpc988 (
      {stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35], 1'b0},
      {stage1_44[10]},
      {stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27], stage1_45[28], stage1_45[29]},
      {stage2_47[4],stage2_46[5],stage2_45[7],stage2_44[10],stage2_43[12]}
   );
   gpc606_5 gpc989 (
      {stage1_44[11], stage1_44[12], stage1_44[13], stage1_44[14], stage1_44[15], stage1_44[16]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[5],stage2_46[6],stage2_45[8],stage2_44[11]}
   );
   gpc606_5 gpc990 (
      {stage1_44[17], stage1_44[18], stage1_44[19], stage1_44[20], stage1_44[21], stage1_44[22]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[6],stage2_46[7],stage2_45[9],stage2_44[12]}
   );
   gpc606_5 gpc991 (
      {stage1_44[23], stage1_44[24], stage1_44[25], stage1_44[26], stage1_44[27], stage1_44[28]},
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16], 1'b0},
      {stage2_48[2],stage2_47[7],stage2_46[8],stage2_45[10],stage2_44[13]}
   );
   gpc606_5 gpc992 (
      {stage1_45[30], stage1_45[31], stage1_45[32], stage1_45[33], stage1_45[34], stage1_45[35]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[3],stage2_47[8],stage2_46[9],stage2_45[11]}
   );
   gpc606_5 gpc993 (
      {stage1_45[36], stage1_45[37], stage1_45[38], stage1_45[39], stage1_45[40], stage1_45[41]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[4],stage2_47[9],stage2_46[10],stage2_45[12]}
   );
   gpc606_5 gpc994 (
      {stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45], stage1_45[46], stage1_45[47]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[5],stage2_47[10],stage2_46[11],stage2_45[13]}
   );
   gpc606_5 gpc995 (
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[0],stage2_49[3],stage2_48[6],stage2_47[11]}
   );
   gpc606_5 gpc996 (
      {stage1_47[24], stage1_47[25], stage1_47[26], stage1_47[27], stage1_47[28], stage1_47[29]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[1],stage2_49[4],stage2_48[7],stage2_47[12]}
   );
   gpc606_5 gpc997 (
      {stage1_47[30], stage1_47[31], stage1_47[32], stage1_47[33], stage1_47[34], stage1_47[35]},
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage2_51[2],stage2_50[2],stage2_49[5],stage2_48[8],stage2_47[13]}
   );
   gpc117_4 gpc998 (
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5], stage1_48[6]},
      {stage1_49[18]},
      {stage1_50[0]},
      {stage2_51[3],stage2_50[3],stage2_49[6],stage2_48[9]}
   );
   gpc117_4 gpc999 (
      {stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11], stage1_48[12], stage1_48[13]},
      {stage1_49[19]},
      {stage1_50[1]},
      {stage2_51[4],stage2_50[4],stage2_49[7],stage2_48[10]}
   );
   gpc117_4 gpc1000 (
      {stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17], stage1_48[18], stage1_48[19], stage1_48[20]},
      {stage1_49[20]},
      {stage1_50[2]},
      {stage2_51[5],stage2_50[5],stage2_49[8],stage2_48[11]}
   );
   gpc207_4 gpc1001 (
      {stage1_48[21], stage1_48[22], stage1_48[23], stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27]},
      {stage1_50[3], stage1_50[4]},
      {stage2_51[6],stage2_50[6],stage2_49[9],stage2_48[12]}
   );
   gpc606_5 gpc1002 (
      {stage1_49[21], stage1_49[22], stage1_49[23], stage1_49[24], 1'b0, 1'b0},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[0],stage2_51[7],stage2_50[7],stage2_49[10]}
   );
   gpc615_5 gpc1003 (
      {stage1_50[5], stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9]},
      {stage1_51[6]},
      {stage1_52[0], stage1_52[1], stage1_52[2], stage1_52[3], stage1_52[4], stage1_52[5]},
      {stage2_54[0],stage2_53[1],stage2_52[1],stage2_51[8],stage2_50[8]}
   );
   gpc615_5 gpc1004 (
      {stage1_50[10], stage1_50[11], stage1_50[12], stage1_50[13], stage1_50[14]},
      {stage1_51[7]},
      {stage1_52[6], stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10], stage1_52[11]},
      {stage2_54[1],stage2_53[2],stage2_52[2],stage2_51[9],stage2_50[9]}
   );
   gpc615_5 gpc1005 (
      {stage1_50[15], stage1_50[16], stage1_50[17], stage1_50[18], stage1_50[19]},
      {stage1_51[8]},
      {stage1_52[12], stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16], stage1_52[17]},
      {stage2_54[2],stage2_53[3],stage2_52[3],stage2_51[10],stage2_50[10]}
   );
   gpc615_5 gpc1006 (
      {stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23], stage1_50[24]},
      {stage1_51[9]},
      {stage1_52[18], stage1_52[19], stage1_52[20], stage1_52[21], stage1_52[22], stage1_52[23]},
      {stage2_54[3],stage2_53[4],stage2_52[4],stage2_51[11],stage2_50[11]}
   );
   gpc2116_5 gpc1007 (
      {stage1_51[10], stage1_51[11], stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15]},
      {stage1_52[24]},
      {stage1_53[0]},
      {stage1_54[0], stage1_54[1]},
      {stage2_55[0],stage2_54[4],stage2_53[5],stage2_52[5],stage2_51[12]}
   );
   gpc2116_5 gpc1008 (
      {stage1_51[16], stage1_51[17], stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21]},
      {stage1_52[25]},
      {stage1_53[1]},
      {stage1_54[2], stage1_54[3]},
      {stage2_55[1],stage2_54[5],stage2_53[6],stage2_52[6],stage2_51[13]}
   );
   gpc615_5 gpc1009 (
      {stage1_51[22], stage1_51[23], stage1_51[24], stage1_51[25], stage1_51[26]},
      {stage1_52[26]},
      {stage1_53[2], stage1_53[3], stage1_53[4], stage1_53[5], stage1_53[6], stage1_53[7]},
      {stage2_55[2],stage2_54[6],stage2_53[7],stage2_52[7],stage2_51[14]}
   );
   gpc615_5 gpc1010 (
      {stage1_51[27], stage1_51[28], stage1_51[29], stage1_51[30], stage1_51[31]},
      {stage1_52[27]},
      {stage1_53[8], stage1_53[9], stage1_53[10], stage1_53[11], stage1_53[12], stage1_53[13]},
      {stage2_55[3],stage2_54[7],stage2_53[8],stage2_52[8],stage2_51[15]}
   );
   gpc615_5 gpc1011 (
      {stage1_52[28], stage1_52[29], stage1_52[30], stage1_52[31], stage1_52[32]},
      {stage1_53[14]},
      {stage1_54[4], stage1_54[5], stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9]},
      {stage2_56[0],stage2_55[4],stage2_54[8],stage2_53[9],stage2_52[9]}
   );
   gpc615_5 gpc1012 (
      {stage1_52[33], stage1_52[34], stage1_52[35], stage1_52[36], stage1_52[37]},
      {stage1_53[15]},
      {stage1_54[10], stage1_54[11], stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15]},
      {stage2_56[1],stage2_55[5],stage2_54[9],stage2_53[10],stage2_52[10]}
   );
   gpc615_5 gpc1013 (
      {stage1_52[38], stage1_52[39], stage1_52[40], stage1_52[41], stage1_52[42]},
      {stage1_53[16]},
      {stage1_54[16], stage1_54[17], stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21]},
      {stage2_56[2],stage2_55[6],stage2_54[10],stage2_53[11],stage2_52[11]}
   );
   gpc615_5 gpc1014 (
      {stage1_53[17], stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21]},
      {stage1_54[22]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[3],stage2_55[7],stage2_54[11],stage2_53[12]}
   );
   gpc1163_5 gpc1015 (
      {stage1_54[23], stage1_54[24], stage1_54[25]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage1_56[0]},
      {stage1_57[0]},
      {stage2_58[0],stage2_57[1],stage2_56[4],stage2_55[8],stage2_54[12]}
   );
   gpc1163_5 gpc1016 (
      {stage1_54[26], stage1_54[27], stage1_54[28]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage1_56[1]},
      {stage1_57[1]},
      {stage2_58[1],stage2_57[2],stage2_56[5],stage2_55[9],stage2_54[13]}
   );
   gpc615_5 gpc1017 (
      {stage1_54[29], stage1_54[30], stage1_54[31], stage1_54[32], 1'b0},
      {stage1_55[18]},
      {stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5], stage1_56[6], stage1_56[7]},
      {stage2_58[2],stage2_57[3],stage2_56[6],stage2_55[10],stage2_54[14]}
   );
   gpc606_5 gpc1018 (
      {stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11], stage1_56[12], stage1_56[13]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[0],stage2_58[3],stage2_57[4],stage2_56[7]}
   );
   gpc606_5 gpc1019 (
      {stage1_56[14], stage1_56[15], stage1_56[16], stage1_56[17], stage1_56[18], stage1_56[19]},
      {stage1_58[6], stage1_58[7], stage1_58[8], stage1_58[9], stage1_58[10], stage1_58[11]},
      {stage2_60[1],stage2_59[1],stage2_58[4],stage2_57[5],stage2_56[8]}
   );
   gpc606_5 gpc1020 (
      {stage1_56[20], stage1_56[21], stage1_56[22], stage1_56[23], stage1_56[24], stage1_56[25]},
      {stage1_58[12], stage1_58[13], stage1_58[14], stage1_58[15], stage1_58[16], stage1_58[17]},
      {stage2_60[2],stage2_59[2],stage2_58[5],stage2_57[6],stage2_56[9]}
   );
   gpc606_5 gpc1021 (
      {stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5], stage1_57[6], stage1_57[7]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[3],stage2_59[3],stage2_58[6],stage2_57[7]}
   );
   gpc615_5 gpc1022 (
      {stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11], stage1_57[12]},
      {stage1_58[18]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[4],stage2_59[4],stage2_58[7],stage2_57[8]}
   );
   gpc615_5 gpc1023 (
      {stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16], stage1_57[17]},
      {stage1_58[19]},
      {stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17]},
      {stage2_61[2],stage2_60[5],stage2_59[5],stage2_58[8],stage2_57[9]}
   );
   gpc615_5 gpc1024 (
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22]},
      {stage1_58[20]},
      {stage1_59[18], stage1_59[19], stage1_59[20], stage1_59[21], stage1_59[22], stage1_59[23]},
      {stage2_61[3],stage2_60[6],stage2_59[6],stage2_58[9],stage2_57[10]}
   );
   gpc615_5 gpc1025 (
      {stage1_58[21], stage1_58[22], stage1_58[23], stage1_58[24], stage1_58[25]},
      {stage1_59[24]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[4],stage2_60[7],stage2_59[7],stage2_58[10]}
   );
   gpc615_5 gpc1026 (
      {stage1_58[26], stage1_58[27], stage1_58[28], stage1_58[29], stage1_58[30]},
      {stage1_59[25]},
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage2_62[1],stage2_61[5],stage2_60[8],stage2_59[8],stage2_58[11]}
   );
   gpc615_5 gpc1027 (
      {stage1_58[31], stage1_58[32], stage1_58[33], stage1_58[34], stage1_58[35]},
      {stage1_59[26]},
      {stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage2_62[2],stage2_61[6],stage2_60[9],stage2_59[9],stage2_58[12]}
   );
   gpc606_5 gpc1028 (
      {stage1_59[27], stage1_59[28], stage1_59[29], stage1_59[30], stage1_59[31], stage1_59[32]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[3],stage2_61[7],stage2_60[10],stage2_59[10]}
   );
   gpc615_5 gpc1029 (
      {stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21], stage1_60[22]},
      {stage1_61[6]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage2_64[0],stage2_63[1],stage2_62[4],stage2_61[8],stage2_60[11]}
   );
   gpc615_5 gpc1030 (
      {stage1_60[23], stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27]},
      {stage1_61[7]},
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11]},
      {stage2_64[1],stage2_63[2],stage2_62[5],stage2_61[9],stage2_60[12]}
   );
   gpc615_5 gpc1031 (
      {stage1_60[28], stage1_60[29], stage1_60[30], stage1_60[31], stage1_60[32]},
      {stage1_61[8]},
      {stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17]},
      {stage2_64[2],stage2_63[3],stage2_62[6],stage2_61[10],stage2_60[13]}
   );
   gpc2135_5 gpc1032 (
      {stage1_61[9], stage1_61[10], stage1_61[11], stage1_61[12], stage1_61[13]},
      {stage1_62[18], stage1_62[19], stage1_62[20]},
      {stage1_63[0]},
      {stage1_64[0], stage1_64[1]},
      {stage2_65[0],stage2_64[3],stage2_63[4],stage2_62[7],stage2_61[11]}
   );
   gpc2135_5 gpc1033 (
      {stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17], stage1_61[18]},
      {stage1_62[21], stage1_62[22], stage1_62[23]},
      {stage1_63[1]},
      {stage1_64[2], stage1_64[3]},
      {stage2_65[1],stage2_64[4],stage2_63[5],stage2_62[8],stage2_61[12]}
   );
   gpc606_5 gpc1034 (
      {stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23], stage1_61[24]},
      {stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5], stage1_63[6], stage1_63[7]},
      {stage2_65[2],stage2_64[5],stage2_63[6],stage2_62[9],stage2_61[13]}
   );
   gpc606_5 gpc1035 (
      {stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29], stage1_61[30]},
      {stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11], stage1_63[12], stage1_63[13]},
      {stage2_65[3],stage2_64[6],stage2_63[7],stage2_62[10],stage2_61[14]}
   );
   gpc606_5 gpc1036 (
      {stage1_62[24], stage1_62[25], stage1_62[26], stage1_62[27], stage1_62[28], stage1_62[29]},
      {stage1_64[4], stage1_64[5], stage1_64[6], stage1_64[7], stage1_64[8], stage1_64[9]},
      {stage2_66[0],stage2_65[4],stage2_64[7],stage2_63[8],stage2_62[11]}
   );
   gpc615_5 gpc1037 (
      {stage1_62[30], stage1_62[31], stage1_62[32], 1'b0, 1'b0},
      {stage1_63[14]},
      {stage1_64[10], stage1_64[11], stage1_64[12], stage1_64[13], stage1_64[14], stage1_64[15]},
      {stage2_66[1],stage2_65[5],stage2_64[8],stage2_63[9],stage2_62[12]}
   );
   gpc606_5 gpc1038 (
      {stage1_63[15], stage1_63[16], stage1_63[17], stage1_63[18], stage1_63[19], stage1_63[20]},
      {stage1_65[0], stage1_65[1], stage1_65[2], stage1_65[3], stage1_65[4], stage1_65[5]},
      {stage2_67[0],stage2_66[2],stage2_65[6],stage2_64[9],stage2_63[10]}
   );
   gpc606_5 gpc1039 (
      {stage1_63[21], stage1_63[22], stage1_63[23], stage1_63[24], stage1_63[25], stage1_63[26]},
      {stage1_65[6], stage1_65[7], stage1_65[8], 1'b0, 1'b0, 1'b0},
      {stage2_67[1],stage2_66[3],stage2_65[7],stage2_64[10],stage2_63[11]}
   );
   gpc1_1 gpc1040 (
      {stage1_2[23]},
      {stage2_2[11]}
   );
   gpc1_1 gpc1041 (
      {stage1_4[27]},
      {stage2_4[15]}
   );
   gpc1_1 gpc1042 (
      {stage1_4[28]},
      {stage2_4[16]}
   );
   gpc1_1 gpc1043 (
      {stage1_4[29]},
      {stage2_4[17]}
   );
   gpc1_1 gpc1044 (
      {stage1_4[30]},
      {stage2_4[18]}
   );
   gpc1_1 gpc1045 (
      {stage1_4[31]},
      {stage2_4[19]}
   );
   gpc1_1 gpc1046 (
      {stage1_4[32]},
      {stage2_4[20]}
   );
   gpc1_1 gpc1047 (
      {stage1_4[33]},
      {stage2_4[21]}
   );
   gpc1_1 gpc1048 (
      {stage1_4[34]},
      {stage2_4[22]}
   );
   gpc1_1 gpc1049 (
      {stage1_4[35]},
      {stage2_4[23]}
   );
   gpc1_1 gpc1050 (
      {stage1_4[36]},
      {stage2_4[24]}
   );
   gpc1_1 gpc1051 (
      {stage1_4[37]},
      {stage2_4[25]}
   );
   gpc1_1 gpc1052 (
      {stage1_5[14]},
      {stage2_5[9]}
   );
   gpc1_1 gpc1053 (
      {stage1_5[15]},
      {stage2_5[10]}
   );
   gpc1_1 gpc1054 (
      {stage1_5[16]},
      {stage2_5[11]}
   );
   gpc1_1 gpc1055 (
      {stage1_5[17]},
      {stage2_5[12]}
   );
   gpc1_1 gpc1056 (
      {stage1_5[18]},
      {stage2_5[13]}
   );
   gpc1_1 gpc1057 (
      {stage1_5[19]},
      {stage2_5[14]}
   );
   gpc1_1 gpc1058 (
      {stage1_5[20]},
      {stage2_5[15]}
   );
   gpc1_1 gpc1059 (
      {stage1_5[21]},
      {stage2_5[16]}
   );
   gpc1_1 gpc1060 (
      {stage1_5[22]},
      {stage2_5[17]}
   );
   gpc1_1 gpc1061 (
      {stage1_5[23]},
      {stage2_5[18]}
   );
   gpc1_1 gpc1062 (
      {stage1_5[24]},
      {stage2_5[19]}
   );
   gpc1_1 gpc1063 (
      {stage1_5[25]},
      {stage2_5[20]}
   );
   gpc1_1 gpc1064 (
      {stage1_5[26]},
      {stage2_5[21]}
   );
   gpc1_1 gpc1065 (
      {stage1_6[15]},
      {stage2_6[7]}
   );
   gpc1_1 gpc1066 (
      {stage1_6[16]},
      {stage2_6[8]}
   );
   gpc1_1 gpc1067 (
      {stage1_6[17]},
      {stage2_6[9]}
   );
   gpc1_1 gpc1068 (
      {stage1_6[18]},
      {stage2_6[10]}
   );
   gpc1_1 gpc1069 (
      {stage1_6[19]},
      {stage2_6[11]}
   );
   gpc1_1 gpc1070 (
      {stage1_6[20]},
      {stage2_6[12]}
   );
   gpc1_1 gpc1071 (
      {stage1_6[21]},
      {stage2_6[13]}
   );
   gpc1_1 gpc1072 (
      {stage1_7[25]},
      {stage2_7[9]}
   );
   gpc1_1 gpc1073 (
      {stage1_7[26]},
      {stage2_7[10]}
   );
   gpc1_1 gpc1074 (
      {stage1_7[27]},
      {stage2_7[11]}
   );
   gpc1_1 gpc1075 (
      {stage1_7[28]},
      {stage2_7[12]}
   );
   gpc1_1 gpc1076 (
      {stage1_7[29]},
      {stage2_7[13]}
   );
   gpc1_1 gpc1077 (
      {stage1_7[30]},
      {stage2_7[14]}
   );
   gpc1_1 gpc1078 (
      {stage1_7[31]},
      {stage2_7[15]}
   );
   gpc1_1 gpc1079 (
      {stage1_7[32]},
      {stage2_7[16]}
   );
   gpc1_1 gpc1080 (
      {stage1_7[33]},
      {stage2_7[17]}
   );
   gpc1_1 gpc1081 (
      {stage1_7[34]},
      {stage2_7[18]}
   );
   gpc1_1 gpc1082 (
      {stage1_7[35]},
      {stage2_7[19]}
   );
   gpc1_1 gpc1083 (
      {stage1_8[16]},
      {stage2_8[9]}
   );
   gpc1_1 gpc1084 (
      {stage1_8[17]},
      {stage2_8[10]}
   );
   gpc1_1 gpc1085 (
      {stage1_8[18]},
      {stage2_8[11]}
   );
   gpc1_1 gpc1086 (
      {stage1_8[19]},
      {stage2_8[12]}
   );
   gpc1_1 gpc1087 (
      {stage1_8[20]},
      {stage2_8[13]}
   );
   gpc1_1 gpc1088 (
      {stage1_8[21]},
      {stage2_8[14]}
   );
   gpc1_1 gpc1089 (
      {stage1_8[22]},
      {stage2_8[15]}
   );
   gpc1_1 gpc1090 (
      {stage1_8[23]},
      {stage2_8[16]}
   );
   gpc1_1 gpc1091 (
      {stage1_8[24]},
      {stage2_8[17]}
   );
   gpc1_1 gpc1092 (
      {stage1_8[25]},
      {stage2_8[18]}
   );
   gpc1_1 gpc1093 (
      {stage1_8[26]},
      {stage2_8[19]}
   );
   gpc1_1 gpc1094 (
      {stage1_9[25]},
      {stage2_9[7]}
   );
   gpc1_1 gpc1095 (
      {stage1_9[26]},
      {stage2_9[8]}
   );
   gpc1_1 gpc1096 (
      {stage1_9[27]},
      {stage2_9[9]}
   );
   gpc1_1 gpc1097 (
      {stage1_9[28]},
      {stage2_9[10]}
   );
   gpc1_1 gpc1098 (
      {stage1_10[11]},
      {stage2_10[8]}
   );
   gpc1_1 gpc1099 (
      {stage1_10[12]},
      {stage2_10[9]}
   );
   gpc1_1 gpc1100 (
      {stage1_10[13]},
      {stage2_10[10]}
   );
   gpc1_1 gpc1101 (
      {stage1_10[14]},
      {stage2_10[11]}
   );
   gpc1_1 gpc1102 (
      {stage1_10[15]},
      {stage2_10[12]}
   );
   gpc1_1 gpc1103 (
      {stage1_10[16]},
      {stage2_10[13]}
   );
   gpc1_1 gpc1104 (
      {stage1_10[17]},
      {stage2_10[14]}
   );
   gpc1_1 gpc1105 (
      {stage1_10[18]},
      {stage2_10[15]}
   );
   gpc1_1 gpc1106 (
      {stage1_10[19]},
      {stage2_10[16]}
   );
   gpc1_1 gpc1107 (
      {stage1_10[20]},
      {stage2_10[17]}
   );
   gpc1_1 gpc1108 (
      {stage1_10[21]},
      {stage2_10[18]}
   );
   gpc1_1 gpc1109 (
      {stage1_10[22]},
      {stage2_10[19]}
   );
   gpc1_1 gpc1110 (
      {stage1_10[23]},
      {stage2_10[20]}
   );
   gpc1_1 gpc1111 (
      {stage1_10[24]},
      {stage2_10[21]}
   );
   gpc1_1 gpc1112 (
      {stage1_10[25]},
      {stage2_10[22]}
   );
   gpc1_1 gpc1113 (
      {stage1_10[26]},
      {stage2_10[23]}
   );
   gpc1_1 gpc1114 (
      {stage1_10[27]},
      {stage2_10[24]}
   );
   gpc1_1 gpc1115 (
      {stage1_10[28]},
      {stage2_10[25]}
   );
   gpc1_1 gpc1116 (
      {stage1_10[29]},
      {stage2_10[26]}
   );
   gpc1_1 gpc1117 (
      {stage1_10[30]},
      {stage2_10[27]}
   );
   gpc1_1 gpc1118 (
      {stage1_10[31]},
      {stage2_10[28]}
   );
   gpc1_1 gpc1119 (
      {stage1_10[32]},
      {stage2_10[29]}
   );
   gpc1_1 gpc1120 (
      {stage1_10[33]},
      {stage2_10[30]}
   );
   gpc1_1 gpc1121 (
      {stage1_11[27]},
      {stage2_11[10]}
   );
   gpc1_1 gpc1122 (
      {stage1_11[28]},
      {stage2_11[11]}
   );
   gpc1_1 gpc1123 (
      {stage1_11[29]},
      {stage2_11[12]}
   );
   gpc1_1 gpc1124 (
      {stage1_11[30]},
      {stage2_11[13]}
   );
   gpc1_1 gpc1125 (
      {stage1_11[31]},
      {stage2_11[14]}
   );
   gpc1_1 gpc1126 (
      {stage1_11[32]},
      {stage2_11[15]}
   );
   gpc1_1 gpc1127 (
      {stage1_12[16]},
      {stage2_12[8]}
   );
   gpc1_1 gpc1128 (
      {stage1_12[17]},
      {stage2_12[9]}
   );
   gpc1_1 gpc1129 (
      {stage1_12[18]},
      {stage2_12[10]}
   );
   gpc1_1 gpc1130 (
      {stage1_12[19]},
      {stage2_12[11]}
   );
   gpc1_1 gpc1131 (
      {stage1_12[20]},
      {stage2_12[12]}
   );
   gpc1_1 gpc1132 (
      {stage1_12[21]},
      {stage2_12[13]}
   );
   gpc1_1 gpc1133 (
      {stage1_12[22]},
      {stage2_12[14]}
   );
   gpc1_1 gpc1134 (
      {stage1_12[23]},
      {stage2_12[15]}
   );
   gpc1_1 gpc1135 (
      {stage1_12[24]},
      {stage2_12[16]}
   );
   gpc1_1 gpc1136 (
      {stage1_12[25]},
      {stage2_12[17]}
   );
   gpc1_1 gpc1137 (
      {stage1_12[26]},
      {stage2_12[18]}
   );
   gpc1_1 gpc1138 (
      {stage1_14[19]},
      {stage2_14[10]}
   );
   gpc1_1 gpc1139 (
      {stage1_14[20]},
      {stage2_14[11]}
   );
   gpc1_1 gpc1140 (
      {stage1_14[21]},
      {stage2_14[12]}
   );
   gpc1_1 gpc1141 (
      {stage1_14[22]},
      {stage2_14[13]}
   );
   gpc1_1 gpc1142 (
      {stage1_14[23]},
      {stage2_14[14]}
   );
   gpc1_1 gpc1143 (
      {stage1_14[24]},
      {stage2_14[15]}
   );
   gpc1_1 gpc1144 (
      {stage1_15[38]},
      {stage2_15[14]}
   );
   gpc1_1 gpc1145 (
      {stage1_15[39]},
      {stage2_15[15]}
   );
   gpc1_1 gpc1146 (
      {stage1_15[40]},
      {stage2_15[16]}
   );
   gpc1_1 gpc1147 (
      {stage1_15[41]},
      {stage2_15[17]}
   );
   gpc1_1 gpc1148 (
      {stage1_15[42]},
      {stage2_15[18]}
   );
   gpc1_1 gpc1149 (
      {stage1_15[43]},
      {stage2_15[19]}
   );
   gpc1_1 gpc1150 (
      {stage1_15[44]},
      {stage2_15[20]}
   );
   gpc1_1 gpc1151 (
      {stage1_16[27]},
      {stage2_16[12]}
   );
   gpc1_1 gpc1152 (
      {stage1_16[28]},
      {stage2_16[13]}
   );
   gpc1_1 gpc1153 (
      {stage1_16[29]},
      {stage2_16[14]}
   );
   gpc1_1 gpc1154 (
      {stage1_16[30]},
      {stage2_16[15]}
   );
   gpc1_1 gpc1155 (
      {stage1_17[35]},
      {stage2_17[12]}
   );
   gpc1_1 gpc1156 (
      {stage1_17[36]},
      {stage2_17[13]}
   );
   gpc1_1 gpc1157 (
      {stage1_17[37]},
      {stage2_17[14]}
   );
   gpc1_1 gpc1158 (
      {stage1_17[38]},
      {stage2_17[15]}
   );
   gpc1_1 gpc1159 (
      {stage1_17[39]},
      {stage2_17[16]}
   );
   gpc1_1 gpc1160 (
      {stage1_17[40]},
      {stage2_17[17]}
   );
   gpc1_1 gpc1161 (
      {stage1_17[41]},
      {stage2_17[18]}
   );
   gpc1_1 gpc1162 (
      {stage1_17[42]},
      {stage2_17[19]}
   );
   gpc1_1 gpc1163 (
      {stage1_17[43]},
      {stage2_17[20]}
   );
   gpc1_1 gpc1164 (
      {stage1_17[44]},
      {stage2_17[21]}
   );
   gpc1_1 gpc1165 (
      {stage1_18[14]},
      {stage2_18[10]}
   );
   gpc1_1 gpc1166 (
      {stage1_18[15]},
      {stage2_18[11]}
   );
   gpc1_1 gpc1167 (
      {stage1_18[16]},
      {stage2_18[12]}
   );
   gpc1_1 gpc1168 (
      {stage1_18[17]},
      {stage2_18[13]}
   );
   gpc1_1 gpc1169 (
      {stage1_18[18]},
      {stage2_18[14]}
   );
   gpc1_1 gpc1170 (
      {stage1_18[19]},
      {stage2_18[15]}
   );
   gpc1_1 gpc1171 (
      {stage1_18[20]},
      {stage2_18[16]}
   );
   gpc1_1 gpc1172 (
      {stage1_18[21]},
      {stage2_18[17]}
   );
   gpc1_1 gpc1173 (
      {stage1_18[22]},
      {stage2_18[18]}
   );
   gpc1_1 gpc1174 (
      {stage1_19[26]},
      {stage2_19[12]}
   );
   gpc1_1 gpc1175 (
      {stage1_19[27]},
      {stage2_19[13]}
   );
   gpc1_1 gpc1176 (
      {stage1_19[28]},
      {stage2_19[14]}
   );
   gpc1_1 gpc1177 (
      {stage1_20[28]},
      {stage2_20[11]}
   );
   gpc1_1 gpc1178 (
      {stage1_20[29]},
      {stage2_20[12]}
   );
   gpc1_1 gpc1179 (
      {stage1_20[30]},
      {stage2_20[13]}
   );
   gpc1_1 gpc1180 (
      {stage1_20[31]},
      {stage2_20[14]}
   );
   gpc1_1 gpc1181 (
      {stage1_20[32]},
      {stage2_20[15]}
   );
   gpc1_1 gpc1182 (
      {stage1_20[33]},
      {stage2_20[16]}
   );
   gpc1_1 gpc1183 (
      {stage1_20[34]},
      {stage2_20[17]}
   );
   gpc1_1 gpc1184 (
      {stage1_20[35]},
      {stage2_20[18]}
   );
   gpc1_1 gpc1185 (
      {stage1_20[36]},
      {stage2_20[19]}
   );
   gpc1_1 gpc1186 (
      {stage1_20[37]},
      {stage2_20[20]}
   );
   gpc1_1 gpc1187 (
      {stage1_20[38]},
      {stage2_20[21]}
   );
   gpc1_1 gpc1188 (
      {stage1_20[39]},
      {stage2_20[22]}
   );
   gpc1_1 gpc1189 (
      {stage1_20[40]},
      {stage2_20[23]}
   );
   gpc1_1 gpc1190 (
      {stage1_21[30]},
      {stage2_21[10]}
   );
   gpc1_1 gpc1191 (
      {stage1_21[31]},
      {stage2_21[11]}
   );
   gpc1_1 gpc1192 (
      {stage1_21[32]},
      {stage2_21[12]}
   );
   gpc1_1 gpc1193 (
      {stage1_23[34]},
      {stage2_23[16]}
   );
   gpc1_1 gpc1194 (
      {stage1_25[43]},
      {stage2_25[12]}
   );
   gpc1_1 gpc1195 (
      {stage1_25[44]},
      {stage2_25[13]}
   );
   gpc1_1 gpc1196 (
      {stage1_26[22]},
      {stage2_26[13]}
   );
   gpc1_1 gpc1197 (
      {stage1_26[23]},
      {stage2_26[14]}
   );
   gpc1_1 gpc1198 (
      {stage1_26[24]},
      {stage2_26[15]}
   );
   gpc1_1 gpc1199 (
      {stage1_26[25]},
      {stage2_26[16]}
   );
   gpc1_1 gpc1200 (
      {stage1_26[26]},
      {stage2_26[17]}
   );
   gpc1_1 gpc1201 (
      {stage1_26[27]},
      {stage2_26[18]}
   );
   gpc1_1 gpc1202 (
      {stage1_26[28]},
      {stage2_26[19]}
   );
   gpc1_1 gpc1203 (
      {stage1_27[29]},
      {stage2_27[14]}
   );
   gpc1_1 gpc1204 (
      {stage1_27[30]},
      {stage2_27[15]}
   );
   gpc1_1 gpc1205 (
      {stage1_27[31]},
      {stage2_27[16]}
   );
   gpc1_1 gpc1206 (
      {stage1_27[32]},
      {stage2_27[17]}
   );
   gpc1_1 gpc1207 (
      {stage1_27[33]},
      {stage2_27[18]}
   );
   gpc1_1 gpc1208 (
      {stage1_27[34]},
      {stage2_27[19]}
   );
   gpc1_1 gpc1209 (
      {stage1_27[35]},
      {stage2_27[20]}
   );
   gpc1_1 gpc1210 (
      {stage1_27[36]},
      {stage2_27[21]}
   );
   gpc1_1 gpc1211 (
      {stage1_27[37]},
      {stage2_27[22]}
   );
   gpc1_1 gpc1212 (
      {stage1_27[38]},
      {stage2_27[23]}
   );
   gpc1_1 gpc1213 (
      {stage1_27[39]},
      {stage2_27[24]}
   );
   gpc1_1 gpc1214 (
      {stage1_27[40]},
      {stage2_27[25]}
   );
   gpc1_1 gpc1215 (
      {stage1_28[21]},
      {stage2_28[10]}
   );
   gpc1_1 gpc1216 (
      {stage1_28[22]},
      {stage2_28[11]}
   );
   gpc1_1 gpc1217 (
      {stage1_28[23]},
      {stage2_28[12]}
   );
   gpc1_1 gpc1218 (
      {stage1_28[24]},
      {stage2_28[13]}
   );
   gpc1_1 gpc1219 (
      {stage1_28[25]},
      {stage2_28[14]}
   );
   gpc1_1 gpc1220 (
      {stage1_28[26]},
      {stage2_28[15]}
   );
   gpc1_1 gpc1221 (
      {stage1_30[16]},
      {stage2_30[10]}
   );
   gpc1_1 gpc1222 (
      {stage1_30[17]},
      {stage2_30[11]}
   );
   gpc1_1 gpc1223 (
      {stage1_30[18]},
      {stage2_30[12]}
   );
   gpc1_1 gpc1224 (
      {stage1_30[19]},
      {stage2_30[13]}
   );
   gpc1_1 gpc1225 (
      {stage1_30[20]},
      {stage2_30[14]}
   );
   gpc1_1 gpc1226 (
      {stage1_30[21]},
      {stage2_30[15]}
   );
   gpc1_1 gpc1227 (
      {stage1_30[22]},
      {stage2_30[16]}
   );
   gpc1_1 gpc1228 (
      {stage1_30[23]},
      {stage2_30[17]}
   );
   gpc1_1 gpc1229 (
      {stage1_30[24]},
      {stage2_30[18]}
   );
   gpc1_1 gpc1230 (
      {stage1_30[25]},
      {stage2_30[19]}
   );
   gpc1_1 gpc1231 (
      {stage1_31[19]},
      {stage2_31[9]}
   );
   gpc1_1 gpc1232 (
      {stage1_31[20]},
      {stage2_31[10]}
   );
   gpc1_1 gpc1233 (
      {stage1_31[21]},
      {stage2_31[11]}
   );
   gpc1_1 gpc1234 (
      {stage1_31[22]},
      {stage2_31[12]}
   );
   gpc1_1 gpc1235 (
      {stage1_32[19]},
      {stage2_32[7]}
   );
   gpc1_1 gpc1236 (
      {stage1_32[20]},
      {stage2_32[8]}
   );
   gpc1_1 gpc1237 (
      {stage1_32[21]},
      {stage2_32[9]}
   );
   gpc1_1 gpc1238 (
      {stage1_32[22]},
      {stage2_32[10]}
   );
   gpc1_1 gpc1239 (
      {stage1_32[23]},
      {stage2_32[11]}
   );
   gpc1_1 gpc1240 (
      {stage1_32[24]},
      {stage2_32[12]}
   );
   gpc1_1 gpc1241 (
      {stage1_32[25]},
      {stage2_32[13]}
   );
   gpc1_1 gpc1242 (
      {stage1_32[26]},
      {stage2_32[14]}
   );
   gpc1_1 gpc1243 (
      {stage1_32[27]},
      {stage2_32[15]}
   );
   gpc1_1 gpc1244 (
      {stage1_32[28]},
      {stage2_32[16]}
   );
   gpc1_1 gpc1245 (
      {stage1_32[29]},
      {stage2_32[17]}
   );
   gpc1_1 gpc1246 (
      {stage1_32[30]},
      {stage2_32[18]}
   );
   gpc1_1 gpc1247 (
      {stage1_33[24]},
      {stage2_33[9]}
   );
   gpc1_1 gpc1248 (
      {stage1_33[25]},
      {stage2_33[10]}
   );
   gpc1_1 gpc1249 (
      {stage1_33[26]},
      {stage2_33[11]}
   );
   gpc1_1 gpc1250 (
      {stage1_33[27]},
      {stage2_33[12]}
   );
   gpc1_1 gpc1251 (
      {stage1_33[28]},
      {stage2_33[13]}
   );
   gpc1_1 gpc1252 (
      {stage1_33[29]},
      {stage2_33[14]}
   );
   gpc1_1 gpc1253 (
      {stage1_33[30]},
      {stage2_33[15]}
   );
   gpc1_1 gpc1254 (
      {stage1_33[31]},
      {stage2_33[16]}
   );
   gpc1_1 gpc1255 (
      {stage1_33[32]},
      {stage2_33[17]}
   );
   gpc1_1 gpc1256 (
      {stage1_33[33]},
      {stage2_33[18]}
   );
   gpc1_1 gpc1257 (
      {stage1_33[34]},
      {stage2_33[19]}
   );
   gpc1_1 gpc1258 (
      {stage1_33[35]},
      {stage2_33[20]}
   );
   gpc1_1 gpc1259 (
      {stage1_33[36]},
      {stage2_33[21]}
   );
   gpc1_1 gpc1260 (
      {stage1_33[37]},
      {stage2_33[22]}
   );
   gpc1_1 gpc1261 (
      {stage1_34[21]},
      {stage2_34[10]}
   );
   gpc1_1 gpc1262 (
      {stage1_34[22]},
      {stage2_34[11]}
   );
   gpc1_1 gpc1263 (
      {stage1_34[23]},
      {stage2_34[12]}
   );
   gpc1_1 gpc1264 (
      {stage1_35[26]},
      {stage2_35[9]}
   );
   gpc1_1 gpc1265 (
      {stage1_35[27]},
      {stage2_35[10]}
   );
   gpc1_1 gpc1266 (
      {stage1_35[28]},
      {stage2_35[11]}
   );
   gpc1_1 gpc1267 (
      {stage1_35[29]},
      {stage2_35[12]}
   );
   gpc1_1 gpc1268 (
      {stage1_36[37]},
      {stage2_36[11]}
   );
   gpc1_1 gpc1269 (
      {stage1_36[38]},
      {stage2_36[12]}
   );
   gpc1_1 gpc1270 (
      {stage1_36[39]},
      {stage2_36[13]}
   );
   gpc1_1 gpc1271 (
      {stage1_36[40]},
      {stage2_36[14]}
   );
   gpc1_1 gpc1272 (
      {stage1_36[41]},
      {stage2_36[15]}
   );
   gpc1_1 gpc1273 (
      {stage1_36[42]},
      {stage2_36[16]}
   );
   gpc1_1 gpc1274 (
      {stage1_36[43]},
      {stage2_36[17]}
   );
   gpc1_1 gpc1275 (
      {stage1_37[18]},
      {stage2_37[12]}
   );
   gpc1_1 gpc1276 (
      {stage1_37[19]},
      {stage2_37[13]}
   );
   gpc1_1 gpc1277 (
      {stage1_37[20]},
      {stage2_37[14]}
   );
   gpc1_1 gpc1278 (
      {stage1_37[21]},
      {stage2_37[15]}
   );
   gpc1_1 gpc1279 (
      {stage1_37[22]},
      {stage2_37[16]}
   );
   gpc1_1 gpc1280 (
      {stage1_37[23]},
      {stage2_37[17]}
   );
   gpc1_1 gpc1281 (
      {stage1_38[29]},
      {stage2_38[11]}
   );
   gpc1_1 gpc1282 (
      {stage1_38[30]},
      {stage2_38[12]}
   );
   gpc1_1 gpc1283 (
      {stage1_38[31]},
      {stage2_38[13]}
   );
   gpc1_1 gpc1284 (
      {stage1_38[32]},
      {stage2_38[14]}
   );
   gpc1_1 gpc1285 (
      {stage1_38[33]},
      {stage2_38[15]}
   );
   gpc1_1 gpc1286 (
      {stage1_38[34]},
      {stage2_38[16]}
   );
   gpc1_1 gpc1287 (
      {stage1_38[35]},
      {stage2_38[17]}
   );
   gpc1_1 gpc1288 (
      {stage1_38[36]},
      {stage2_38[18]}
   );
   gpc1_1 gpc1289 (
      {stage1_38[37]},
      {stage2_38[19]}
   );
   gpc1_1 gpc1290 (
      {stage1_38[38]},
      {stage2_38[20]}
   );
   gpc1_1 gpc1291 (
      {stage1_38[39]},
      {stage2_38[21]}
   );
   gpc1_1 gpc1292 (
      {stage1_38[40]},
      {stage2_38[22]}
   );
   gpc1_1 gpc1293 (
      {stage1_38[41]},
      {stage2_38[23]}
   );
   gpc1_1 gpc1294 (
      {stage1_39[19]},
      {stage2_39[9]}
   );
   gpc1_1 gpc1295 (
      {stage1_39[20]},
      {stage2_39[10]}
   );
   gpc1_1 gpc1296 (
      {stage1_39[21]},
      {stage2_39[11]}
   );
   gpc1_1 gpc1297 (
      {stage1_39[22]},
      {stage2_39[12]}
   );
   gpc1_1 gpc1298 (
      {stage1_40[26]},
      {stage2_40[11]}
   );
   gpc1_1 gpc1299 (
      {stage1_41[27]},
      {stage2_41[11]}
   );
   gpc1_1 gpc1300 (
      {stage1_41[28]},
      {stage2_41[12]}
   );
   gpc1_1 gpc1301 (
      {stage1_41[29]},
      {stage2_41[13]}
   );
   gpc1_1 gpc1302 (
      {stage1_41[30]},
      {stage2_41[14]}
   );
   gpc1_1 gpc1303 (
      {stage1_41[31]},
      {stage2_41[15]}
   );
   gpc1_1 gpc1304 (
      {stage1_41[32]},
      {stage2_41[16]}
   );
   gpc1_1 gpc1305 (
      {stage1_41[33]},
      {stage2_41[17]}
   );
   gpc1_1 gpc1306 (
      {stage1_41[34]},
      {stage2_41[18]}
   );
   gpc1_1 gpc1307 (
      {stage1_41[35]},
      {stage2_41[19]}
   );
   gpc1_1 gpc1308 (
      {stage1_42[24]},
      {stage2_42[10]}
   );
   gpc1_1 gpc1309 (
      {stage1_42[25]},
      {stage2_42[11]}
   );
   gpc1_1 gpc1310 (
      {stage1_42[26]},
      {stage2_42[12]}
   );
   gpc1_1 gpc1311 (
      {stage1_42[27]},
      {stage2_42[13]}
   );
   gpc1_1 gpc1312 (
      {stage1_42[28]},
      {stage2_42[14]}
   );
   gpc1_1 gpc1313 (
      {stage1_44[29]},
      {stage2_44[14]}
   );
   gpc1_1 gpc1314 (
      {stage1_44[30]},
      {stage2_44[15]}
   );
   gpc1_1 gpc1315 (
      {stage1_44[31]},
      {stage2_44[16]}
   );
   gpc1_1 gpc1316 (
      {stage1_44[32]},
      {stage2_44[17]}
   );
   gpc1_1 gpc1317 (
      {stage1_47[36]},
      {stage2_47[14]}
   );
   gpc1_1 gpc1318 (
      {stage1_47[37]},
      {stage2_47[15]}
   );
   gpc1_1 gpc1319 (
      {stage1_47[38]},
      {stage2_47[16]}
   );
   gpc1_1 gpc1320 (
      {stage1_47[39]},
      {stage2_47[17]}
   );
   gpc1_1 gpc1321 (
      {stage1_47[40]},
      {stage2_47[18]}
   );
   gpc1_1 gpc1322 (
      {stage1_48[28]},
      {stage2_48[13]}
   );
   gpc1_1 gpc1323 (
      {stage1_48[29]},
      {stage2_48[14]}
   );
   gpc1_1 gpc1324 (
      {stage1_48[30]},
      {stage2_48[15]}
   );
   gpc1_1 gpc1325 (
      {stage1_48[31]},
      {stage2_48[16]}
   );
   gpc1_1 gpc1326 (
      {stage1_53[22]},
      {stage2_53[13]}
   );
   gpc1_1 gpc1327 (
      {stage1_53[23]},
      {stage2_53[14]}
   );
   gpc1_1 gpc1328 (
      {stage1_53[24]},
      {stage2_53[15]}
   );
   gpc1_1 gpc1329 (
      {stage1_53[25]},
      {stage2_53[16]}
   );
   gpc1_1 gpc1330 (
      {stage1_53[26]},
      {stage2_53[17]}
   );
   gpc1_1 gpc1331 (
      {stage1_55[19]},
      {stage2_55[11]}
   );
   gpc1_1 gpc1332 (
      {stage1_55[20]},
      {stage2_55[12]}
   );
   gpc1_1 gpc1333 (
      {stage1_55[21]},
      {stage2_55[13]}
   );
   gpc1_1 gpc1334 (
      {stage1_55[22]},
      {stage2_55[14]}
   );
   gpc1_1 gpc1335 (
      {stage1_55[23]},
      {stage2_55[15]}
   );
   gpc1_1 gpc1336 (
      {stage1_55[24]},
      {stage2_55[16]}
   );
   gpc1_1 gpc1337 (
      {stage1_57[23]},
      {stage2_57[11]}
   );
   gpc1_1 gpc1338 (
      {stage1_57[24]},
      {stage2_57[12]}
   );
   gpc1_1 gpc1339 (
      {stage1_57[25]},
      {stage2_57[13]}
   );
   gpc1_1 gpc1340 (
      {stage1_58[36]},
      {stage2_58[13]}
   );
   gpc1_1 gpc1341 (
      {stage1_58[37]},
      {stage2_58[14]}
   );
   gpc1_1 gpc1342 (
      {stage1_58[38]},
      {stage2_58[15]}
   );
   gpc1_1 gpc1343 (
      {stage1_58[39]},
      {stage2_58[16]}
   );
   gpc1_1 gpc1344 (
      {stage1_58[40]},
      {stage2_58[17]}
   );
   gpc1_1 gpc1345 (
      {stage1_59[33]},
      {stage2_59[11]}
   );
   gpc1_1 gpc1346 (
      {stage1_59[34]},
      {stage2_59[12]}
   );
   gpc1_1 gpc1347 (
      {stage1_59[35]},
      {stage2_59[13]}
   );
   gpc1_1 gpc1348 (
      {stage1_59[36]},
      {stage2_59[14]}
   );
   gpc1_1 gpc1349 (
      {stage1_59[37]},
      {stage2_59[15]}
   );
   gpc1_1 gpc1350 (
      {stage1_59[38]},
      {stage2_59[16]}
   );
   gpc1_1 gpc1351 (
      {stage1_59[39]},
      {stage2_59[17]}
   );
   gpc1_1 gpc1352 (
      {stage1_59[40]},
      {stage2_59[18]}
   );
   gpc1_1 gpc1353 (
      {stage1_59[41]},
      {stage2_59[19]}
   );
   gpc1_1 gpc1354 (
      {stage1_63[27]},
      {stage2_63[12]}
   );
   gpc606_5 gpc1355 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc606_5 gpc1356 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc606_5 gpc1357 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[2],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc615_5 gpc1358 (
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[12]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[2],stage3_5[3],stage3_4[3],stage3_3[3]}
   );
   gpc606_5 gpc1359 (
      {stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[3],stage3_5[4],stage3_4[4]}
   );
   gpc606_5 gpc1360 (
      {stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[2],stage3_6[4],stage3_5[5],stage3_4[5]}
   );
   gpc606_5 gpc1361 (
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[2],stage3_7[3],stage3_6[5],stage3_5[6]}
   );
   gpc606_5 gpc1362 (
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[3],stage3_7[4],stage3_6[6],stage3_5[7]}
   );
   gpc1325_5 gpc1363 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], 1'b0},
      {stage2_6[12], stage2_6[13]},
      {stage2_7[12], stage2_7[13], stage2_7[14]},
      {stage2_8[0]},
      {stage3_9[2],stage3_8[4],stage3_7[5],stage3_6[7],stage3_5[8]}
   );
   gpc606_5 gpc1364 (
      {stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[0],stage3_9[3],stage3_8[5]}
   );
   gpc606_5 gpc1365 (
      {stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11], stage2_8[12]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[1],stage3_10[1],stage3_9[4],stage3_8[6]}
   );
   gpc606_5 gpc1366 (
      {stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17], stage2_8[18]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[2],stage3_10[2],stage3_9[5],stage3_8[7]}
   );
   gpc606_5 gpc1367 (
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[3],stage3_11[3],stage3_10[3],stage3_9[6]}
   );
   gpc1163_5 gpc1368 (
      {stage2_10[18], stage2_10[19], stage2_10[20]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[0]},
      {stage2_13[0]},
      {stage3_14[0],stage3_13[1],stage3_12[4],stage3_11[4],stage3_10[4]}
   );
   gpc615_5 gpc1369 (
      {stage2_10[21], stage2_10[22], stage2_10[23], stage2_10[24], stage2_10[25]},
      {stage2_11[12]},
      {stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6]},
      {stage3_14[1],stage3_13[2],stage3_12[5],stage3_11[5],stage3_10[5]}
   );
   gpc615_5 gpc1370 (
      {stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29], stage2_10[30]},
      {stage2_11[13]},
      {stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12]},
      {stage3_14[2],stage3_13[3],stage3_12[6],stage3_11[6],stage3_10[6]}
   );
   gpc606_5 gpc1371 (
      {stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[0],stage3_14[3],stage3_13[4],stage3_12[7]}
   );
   gpc615_5 gpc1372 (
      {stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage2_14[6]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[1],stage3_15[1],stage3_14[4],stage3_13[5]}
   );
   gpc615_5 gpc1373 (
      {stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_15[6]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[1],stage3_16[2],stage3_15[2],stage3_14[5]}
   );
   gpc615_5 gpc1374 (
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], 1'b0},
      {stage2_15[7]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[2],stage3_16[3],stage3_15[3],stage3_14[6]}
   );
   gpc615_5 gpc1375 (
      {stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11], stage2_15[12]},
      {stage2_16[12]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[2],stage3_17[3],stage3_16[4],stage3_15[4]}
   );
   gpc615_5 gpc1376 (
      {stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage2_16[13]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[3],stage3_17[4],stage3_16[5],stage3_15[5]}
   );
   gpc606_5 gpc1377 (
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[0],stage3_19[2],stage3_18[4],stage3_17[5]}
   );
   gpc606_5 gpc1378 (
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], 1'b0, 1'b0},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[1],stage3_19[3],stage3_18[5],stage3_17[6]}
   );
   gpc615_5 gpc1379 (
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4]},
      {stage2_19[12]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[2],stage3_20[2],stage3_19[4],stage3_18[6]}
   );
   gpc615_5 gpc1380 (
      {stage2_18[5], stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9]},
      {stage2_19[13]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[3],stage3_20[3],stage3_19[5],stage3_18[7]}
   );
   gpc615_5 gpc1381 (
      {stage2_18[10], stage2_18[11], stage2_18[12], stage2_18[13], stage2_18[14]},
      {stage2_19[14]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[4],stage3_20[4],stage3_19[6],stage3_18[8]}
   );
   gpc606_5 gpc1382 (
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[0],stage3_22[3],stage3_21[5],stage3_20[5]}
   );
   gpc606_5 gpc1383 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[1],stage3_23[1],stage3_22[4],stage3_21[6]}
   );
   gpc606_5 gpc1384 (
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[2],stage3_23[2],stage3_22[5],stage3_21[7]}
   );
   gpc615_5 gpc1385 (
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10]},
      {stage2_23[12]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[2],stage3_24[3],stage3_23[3],stage3_22[6]}
   );
   gpc606_5 gpc1386 (
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[0],stage3_26[1],stage3_25[3],stage3_24[4]}
   );
   gpc606_5 gpc1387 (
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[2],stage3_25[4]}
   );
   gpc606_5 gpc1388 (
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[2],stage3_27[2],stage3_26[3],stage3_25[5]}
   );
   gpc135_4 gpc1389 (
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10]},
      {stage2_27[12], stage2_27[13], stage2_27[14]},
      {stage2_28[0]},
      {stage3_29[2],stage3_28[3],stage3_27[3],stage3_26[4]}
   );
   gpc135_4 gpc1390 (
      {stage2_26[11], stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15]},
      {stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage2_28[1]},
      {stage3_29[3],stage3_28[4],stage3_27[4],stage3_26[5]}
   );
   gpc135_4 gpc1391 (
      {stage2_26[16], stage2_26[17], stage2_26[18], stage2_26[19], 1'b0},
      {stage2_27[18], stage2_27[19], stage2_27[20]},
      {stage2_28[2]},
      {stage3_29[4],stage3_28[5],stage3_27[5],stage3_26[6]}
   );
   gpc615_5 gpc1392 (
      {stage2_27[21], stage2_27[22], stage2_27[23], stage2_27[24], stage2_27[25]},
      {stage2_28[3]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[0],stage3_29[5],stage3_28[6],stage3_27[6]}
   );
   gpc606_5 gpc1393 (
      {stage2_28[4], stage2_28[5], stage2_28[6], stage2_28[7], stage2_28[8], stage2_28[9]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[1],stage3_30[1],stage3_29[6],stage3_28[7]}
   );
   gpc606_5 gpc1394 (
      {stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[2],stage3_30[2],stage3_29[7],stage3_28[8]}
   );
   gpc606_5 gpc1395 (
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], 1'b0, 1'b0},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[2],stage3_31[3],stage3_30[3],stage3_29[8]}
   );
   gpc615_5 gpc1396 (
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16]},
      {stage2_31[6]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[1],stage3_32[3],stage3_31[4],stage3_30[4]}
   );
   gpc615_5 gpc1397 (
      {stage2_30[17], stage2_30[18], stage2_30[19], 1'b0, 1'b0},
      {stage2_31[7]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[2],stage3_32[4],stage3_31[5],stage3_30[5]}
   );
   gpc615_5 gpc1398 (
      {stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11], stage2_31[12]},
      {stage2_32[12]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[2],stage3_33[3],stage3_32[5],stage3_31[6]}
   );
   gpc606_5 gpc1399 (
      {stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17], stage2_32[18]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[1],stage3_34[3],stage3_33[4],stage3_32[6]}
   );
   gpc606_5 gpc1400 (
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[1],stage3_35[2],stage3_34[4],stage3_33[5]}
   );
   gpc615_5 gpc1401 (
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10]},
      {stage2_35[6]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[1],stage3_36[2],stage3_35[3],stage3_34[5]}
   );
   gpc615_5 gpc1402 (
      {stage2_34[11], stage2_34[12], 1'b0, 1'b0, 1'b0},
      {stage2_35[7]},
      {stage2_36[6], stage2_36[7], stage2_36[8], stage2_36[9], stage2_36[10], stage2_36[11]},
      {stage3_38[1],stage3_37[2],stage3_36[3],stage3_35[4],stage3_34[6]}
   );
   gpc615_5 gpc1403 (
      {stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11], stage2_35[12]},
      {stage2_36[12]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[2],stage3_37[3],stage3_36[4],stage3_35[5]}
   );
   gpc606_5 gpc1404 (
      {stage2_37[6], stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5]},
      {stage3_41[0],stage3_40[0],stage3_39[1],stage3_38[3],stage3_37[4]}
   );
   gpc606_5 gpc1405 (
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage2_39[6], stage2_39[7], stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11]},
      {stage3_41[1],stage3_40[1],stage3_39[2],stage3_38[4],stage3_37[5]}
   );
   gpc207_4 gpc1406 (
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5], stage2_38[6]},
      {stage2_40[0], stage2_40[1]},
      {stage3_41[2],stage3_40[2],stage3_39[3],stage3_38[5]}
   );
   gpc207_4 gpc1407 (
      {stage2_38[7], stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11], stage2_38[12], stage2_38[13]},
      {stage2_40[2], stage2_40[3]},
      {stage3_41[3],stage3_40[3],stage3_39[4],stage3_38[6]}
   );
   gpc207_4 gpc1408 (
      {stage2_38[14], stage2_38[15], stage2_38[16], stage2_38[17], stage2_38[18], stage2_38[19], stage2_38[20]},
      {stage2_40[4], stage2_40[5]},
      {stage3_41[4],stage3_40[4],stage3_39[5],stage3_38[7]}
   );
   gpc606_5 gpc1409 (
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[0],stage3_42[0],stage3_41[5],stage3_40[5]}
   );
   gpc135_4 gpc1410 (
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4]},
      {stage2_42[6], stage2_42[7], stage2_42[8]},
      {stage2_43[0]},
      {stage3_44[1],stage3_43[1],stage3_42[1],stage3_41[6]}
   );
   gpc135_4 gpc1411 (
      {stage2_41[5], stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9]},
      {stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage2_43[1]},
      {stage3_44[2],stage3_43[2],stage3_42[2],stage3_41[7]}
   );
   gpc135_4 gpc1412 (
      {stage2_41[10], stage2_41[11], stage2_41[12], stage2_41[13], stage2_41[14]},
      {stage2_42[12], stage2_42[13], stage2_42[14]},
      {stage2_43[2]},
      {stage3_44[3],stage3_43[3],stage3_42[3],stage3_41[8]}
   );
   gpc615_5 gpc1413 (
      {stage2_43[3], stage2_43[4], stage2_43[5], stage2_43[6], stage2_43[7]},
      {stage2_44[0]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[0],stage3_45[0],stage3_44[4],stage3_43[4]}
   );
   gpc615_5 gpc1414 (
      {stage2_43[8], stage2_43[9], stage2_43[10], stage2_43[11], stage2_43[12]},
      {stage2_44[1]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[1],stage3_45[1],stage3_44[5],stage3_43[5]}
   );
   gpc606_5 gpc1415 (
      {stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5], stage2_44[6], stage2_44[7]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[2],stage3_46[2],stage3_45[2],stage3_44[6]}
   );
   gpc1163_5 gpc1416 (
      {stage2_46[6], stage2_46[7], stage2_46[8]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage2_48[0]},
      {stage2_49[0]},
      {stage3_50[0],stage3_49[0],stage3_48[1],stage3_47[3],stage3_46[3]}
   );
   gpc1325_5 gpc1417 (
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10]},
      {stage2_48[1], stage2_48[2]},
      {stage2_49[1], stage2_49[2], stage2_49[3]},
      {stage2_50[0]},
      {stage3_51[0],stage3_50[1],stage3_49[1],stage3_48[2],stage3_47[4]}
   );
   gpc1325_5 gpc1418 (
      {stage2_47[11], stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15]},
      {stage2_48[3], stage2_48[4]},
      {stage2_49[4], stage2_49[5], stage2_49[6]},
      {stage2_50[1]},
      {stage3_51[1],stage3_50[2],stage3_49[2],stage3_48[3],stage3_47[5]}
   );
   gpc1406_5 gpc1419 (
      {stage2_48[5], stage2_48[6], stage2_48[7], stage2_48[8], stage2_48[9], stage2_48[10]},
      {stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage2_51[0]},
      {stage3_52[0],stage3_51[2],stage3_50[3],stage3_49[3],stage3_48[4]}
   );
   gpc1406_5 gpc1420 (
      {stage2_48[11], stage2_48[12], stage2_48[13], stage2_48[14], stage2_48[15], stage2_48[16]},
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9]},
      {stage2_51[1]},
      {stage3_52[1],stage3_51[3],stage3_50[4],stage3_49[4],stage3_48[5]}
   );
   gpc615_5 gpc1421 (
      {stage2_49[7], stage2_49[8], stage2_49[9], stage2_49[10], 1'b0},
      {stage2_50[10]},
      {stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5], stage2_51[6], stage2_51[7]},
      {stage3_53[0],stage3_52[2],stage3_51[4],stage3_50[5],stage3_49[5]}
   );
   gpc615_5 gpc1422 (
      {stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11], stage2_51[12]},
      {stage2_52[0]},
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage3_55[0],stage3_54[0],stage3_53[1],stage3_52[3],stage3_51[5]}
   );
   gpc615_5 gpc1423 (
      {stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5]},
      {stage2_53[6]},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage3_56[0],stage3_55[1],stage3_54[1],stage3_53[2],stage3_52[4]}
   );
   gpc615_5 gpc1424 (
      {stage2_52[6], stage2_52[7], stage2_52[8], stage2_52[9], stage2_52[10]},
      {stage2_53[7]},
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage3_56[1],stage3_55[2],stage3_54[2],stage3_53[3],stage3_52[5]}
   );
   gpc615_5 gpc1425 (
      {stage2_53[8], stage2_53[9], stage2_53[10], stage2_53[11], stage2_53[12]},
      {stage2_54[12]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[2],stage3_55[3],stage3_54[3],stage3_53[4]}
   );
   gpc615_5 gpc1426 (
      {stage2_53[13], stage2_53[14], stage2_53[15], stage2_53[16], stage2_53[17]},
      {stage2_54[13]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[3],stage3_55[4],stage3_54[4],stage3_53[5]}
   );
   gpc615_5 gpc1427 (
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4]},
      {stage2_57[0]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[0],stage3_58[0],stage3_57[2],stage3_56[4]}
   );
   gpc615_5 gpc1428 (
      {stage2_56[5], stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9]},
      {stage2_57[1]},
      {stage2_58[6], stage2_58[7], stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage3_60[1],stage3_59[1],stage3_58[1],stage3_57[3],stage3_56[5]}
   );
   gpc615_5 gpc1429 (
      {stage2_57[2], stage2_57[3], stage2_57[4], stage2_57[5], stage2_57[6]},
      {stage2_58[12]},
      {stage2_59[0], stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5]},
      {stage3_61[0],stage3_60[2],stage3_59[2],stage3_58[2],stage3_57[4]}
   );
   gpc615_5 gpc1430 (
      {stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10], stage2_57[11]},
      {stage2_58[13]},
      {stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11]},
      {stage3_61[1],stage3_60[3],stage3_59[3],stage3_58[3],stage3_57[5]}
   );
   gpc615_5 gpc1431 (
      {stage2_59[12], stage2_59[13], stage2_59[14], stage2_59[15], stage2_59[16]},
      {stage2_60[0]},
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage3_63[0],stage3_62[0],stage3_61[2],stage3_60[4],stage3_59[4]}
   );
   gpc615_5 gpc1432 (
      {stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5]},
      {stage2_61[6]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[1],stage3_62[1],stage3_61[3],stage3_60[5]}
   );
   gpc606_5 gpc1433 (
      {stage2_61[7], stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11], stage2_61[12]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[1],stage3_63[2],stage3_62[2],stage3_61[4]}
   );
   gpc606_5 gpc1434 (
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[1],stage3_64[2],stage3_63[3],stage3_62[3]}
   );
   gpc606_5 gpc1435 (
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11]},
      {stage2_65[0], stage2_65[1], stage2_65[2], stage2_65[3], stage2_65[4], stage2_65[5]},
      {stage3_67[0],stage3_66[1],stage3_65[2],stage3_64[3],stage3_63[4]}
   );
   gpc1406_5 gpc1436 (
      {stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9], stage2_64[10], 1'b0},
      {stage2_66[0], stage2_66[1], stage2_66[2], stage2_66[3]},
      {stage2_67[0]},
      {stage3_68[0],stage3_67[1],stage3_66[2],stage3_65[3],stage3_64[4]}
   );
   gpc1_1 gpc1437 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc1438 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc1439 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc1440 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc1441 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc1442 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc1443 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc1444 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc1445 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc1446 (
      {stage2_3[11]},
      {stage3_3[4]}
   );
   gpc1_1 gpc1447 (
      {stage2_4[25]},
      {stage3_4[6]}
   );
   gpc1_1 gpc1448 (
      {stage2_7[15]},
      {stage3_7[6]}
   );
   gpc1_1 gpc1449 (
      {stage2_7[16]},
      {stage3_7[7]}
   );
   gpc1_1 gpc1450 (
      {stage2_7[17]},
      {stage3_7[8]}
   );
   gpc1_1 gpc1451 (
      {stage2_7[18]},
      {stage3_7[9]}
   );
   gpc1_1 gpc1452 (
      {stage2_7[19]},
      {stage3_7[10]}
   );
   gpc1_1 gpc1453 (
      {stage2_8[19]},
      {stage3_8[8]}
   );
   gpc1_1 gpc1454 (
      {stage2_9[6]},
      {stage3_9[7]}
   );
   gpc1_1 gpc1455 (
      {stage2_9[7]},
      {stage3_9[8]}
   );
   gpc1_1 gpc1456 (
      {stage2_9[8]},
      {stage3_9[9]}
   );
   gpc1_1 gpc1457 (
      {stage2_9[9]},
      {stage3_9[10]}
   );
   gpc1_1 gpc1458 (
      {stage2_9[10]},
      {stage3_9[11]}
   );
   gpc1_1 gpc1459 (
      {stage2_11[14]},
      {stage3_11[7]}
   );
   gpc1_1 gpc1460 (
      {stage2_11[15]},
      {stage3_11[8]}
   );
   gpc1_1 gpc1461 (
      {stage2_13[6]},
      {stage3_13[6]}
   );
   gpc1_1 gpc1462 (
      {stage2_13[7]},
      {stage3_13[7]}
   );
   gpc1_1 gpc1463 (
      {stage2_13[8]},
      {stage3_13[8]}
   );
   gpc1_1 gpc1464 (
      {stage2_15[18]},
      {stage3_15[6]}
   );
   gpc1_1 gpc1465 (
      {stage2_15[19]},
      {stage3_15[7]}
   );
   gpc1_1 gpc1466 (
      {stage2_15[20]},
      {stage3_15[8]}
   );
   gpc1_1 gpc1467 (
      {stage2_16[14]},
      {stage3_16[6]}
   );
   gpc1_1 gpc1468 (
      {stage2_16[15]},
      {stage3_16[7]}
   );
   gpc1_1 gpc1469 (
      {stage2_18[15]},
      {stage3_18[9]}
   );
   gpc1_1 gpc1470 (
      {stage2_18[16]},
      {stage3_18[10]}
   );
   gpc1_1 gpc1471 (
      {stage2_18[17]},
      {stage3_18[11]}
   );
   gpc1_1 gpc1472 (
      {stage2_18[18]},
      {stage3_18[12]}
   );
   gpc1_1 gpc1473 (
      {stage2_21[12]},
      {stage3_21[8]}
   );
   gpc1_1 gpc1474 (
      {stage2_23[13]},
      {stage3_23[4]}
   );
   gpc1_1 gpc1475 (
      {stage2_23[14]},
      {stage3_23[5]}
   );
   gpc1_1 gpc1476 (
      {stage2_23[15]},
      {stage3_23[6]}
   );
   gpc1_1 gpc1477 (
      {stage2_23[16]},
      {stage3_23[7]}
   );
   gpc1_1 gpc1478 (
      {stage2_24[12]},
      {stage3_24[5]}
   );
   gpc1_1 gpc1479 (
      {stage2_24[13]},
      {stage3_24[6]}
   );
   gpc1_1 gpc1480 (
      {stage2_25[12]},
      {stage3_25[6]}
   );
   gpc1_1 gpc1481 (
      {stage2_25[13]},
      {stage3_25[7]}
   );
   gpc1_1 gpc1482 (
      {stage2_33[12]},
      {stage3_33[6]}
   );
   gpc1_1 gpc1483 (
      {stage2_33[13]},
      {stage3_33[7]}
   );
   gpc1_1 gpc1484 (
      {stage2_33[14]},
      {stage3_33[8]}
   );
   gpc1_1 gpc1485 (
      {stage2_33[15]},
      {stage3_33[9]}
   );
   gpc1_1 gpc1486 (
      {stage2_33[16]},
      {stage3_33[10]}
   );
   gpc1_1 gpc1487 (
      {stage2_33[17]},
      {stage3_33[11]}
   );
   gpc1_1 gpc1488 (
      {stage2_33[18]},
      {stage3_33[12]}
   );
   gpc1_1 gpc1489 (
      {stage2_33[19]},
      {stage3_33[13]}
   );
   gpc1_1 gpc1490 (
      {stage2_33[20]},
      {stage3_33[14]}
   );
   gpc1_1 gpc1491 (
      {stage2_33[21]},
      {stage3_33[15]}
   );
   gpc1_1 gpc1492 (
      {stage2_33[22]},
      {stage3_33[16]}
   );
   gpc1_1 gpc1493 (
      {stage2_36[13]},
      {stage3_36[5]}
   );
   gpc1_1 gpc1494 (
      {stage2_36[14]},
      {stage3_36[6]}
   );
   gpc1_1 gpc1495 (
      {stage2_36[15]},
      {stage3_36[7]}
   );
   gpc1_1 gpc1496 (
      {stage2_36[16]},
      {stage3_36[8]}
   );
   gpc1_1 gpc1497 (
      {stage2_36[17]},
      {stage3_36[9]}
   );
   gpc1_1 gpc1498 (
      {stage2_38[21]},
      {stage3_38[8]}
   );
   gpc1_1 gpc1499 (
      {stage2_38[22]},
      {stage3_38[9]}
   );
   gpc1_1 gpc1500 (
      {stage2_38[23]},
      {stage3_38[10]}
   );
   gpc1_1 gpc1501 (
      {stage2_39[12]},
      {stage3_39[6]}
   );
   gpc1_1 gpc1502 (
      {stage2_41[15]},
      {stage3_41[9]}
   );
   gpc1_1 gpc1503 (
      {stage2_41[16]},
      {stage3_41[10]}
   );
   gpc1_1 gpc1504 (
      {stage2_41[17]},
      {stage3_41[11]}
   );
   gpc1_1 gpc1505 (
      {stage2_41[18]},
      {stage3_41[12]}
   );
   gpc1_1 gpc1506 (
      {stage2_41[19]},
      {stage3_41[13]}
   );
   gpc1_1 gpc1507 (
      {stage2_44[8]},
      {stage3_44[7]}
   );
   gpc1_1 gpc1508 (
      {stage2_44[9]},
      {stage3_44[8]}
   );
   gpc1_1 gpc1509 (
      {stage2_44[10]},
      {stage3_44[9]}
   );
   gpc1_1 gpc1510 (
      {stage2_44[11]},
      {stage3_44[10]}
   );
   gpc1_1 gpc1511 (
      {stage2_44[12]},
      {stage3_44[11]}
   );
   gpc1_1 gpc1512 (
      {stage2_44[13]},
      {stage3_44[12]}
   );
   gpc1_1 gpc1513 (
      {stage2_44[14]},
      {stage3_44[13]}
   );
   gpc1_1 gpc1514 (
      {stage2_44[15]},
      {stage3_44[14]}
   );
   gpc1_1 gpc1515 (
      {stage2_44[16]},
      {stage3_44[15]}
   );
   gpc1_1 gpc1516 (
      {stage2_44[17]},
      {stage3_44[16]}
   );
   gpc1_1 gpc1517 (
      {stage2_45[12]},
      {stage3_45[3]}
   );
   gpc1_1 gpc1518 (
      {stage2_45[13]},
      {stage3_45[4]}
   );
   gpc1_1 gpc1519 (
      {stage2_46[9]},
      {stage3_46[4]}
   );
   gpc1_1 gpc1520 (
      {stage2_46[10]},
      {stage3_46[5]}
   );
   gpc1_1 gpc1521 (
      {stage2_46[11]},
      {stage3_46[6]}
   );
   gpc1_1 gpc1522 (
      {stage2_47[16]},
      {stage3_47[6]}
   );
   gpc1_1 gpc1523 (
      {stage2_47[17]},
      {stage3_47[7]}
   );
   gpc1_1 gpc1524 (
      {stage2_47[18]},
      {stage3_47[8]}
   );
   gpc1_1 gpc1525 (
      {stage2_50[11]},
      {stage3_50[6]}
   );
   gpc1_1 gpc1526 (
      {stage2_51[13]},
      {stage3_51[6]}
   );
   gpc1_1 gpc1527 (
      {stage2_51[14]},
      {stage3_51[7]}
   );
   gpc1_1 gpc1528 (
      {stage2_51[15]},
      {stage3_51[8]}
   );
   gpc1_1 gpc1529 (
      {stage2_52[11]},
      {stage3_52[6]}
   );
   gpc1_1 gpc1530 (
      {stage2_54[14]},
      {stage3_54[5]}
   );
   gpc1_1 gpc1531 (
      {stage2_55[12]},
      {stage3_55[5]}
   );
   gpc1_1 gpc1532 (
      {stage2_55[13]},
      {stage3_55[6]}
   );
   gpc1_1 gpc1533 (
      {stage2_55[14]},
      {stage3_55[7]}
   );
   gpc1_1 gpc1534 (
      {stage2_55[15]},
      {stage3_55[8]}
   );
   gpc1_1 gpc1535 (
      {stage2_55[16]},
      {stage3_55[9]}
   );
   gpc1_1 gpc1536 (
      {stage2_57[12]},
      {stage3_57[6]}
   );
   gpc1_1 gpc1537 (
      {stage2_57[13]},
      {stage3_57[7]}
   );
   gpc1_1 gpc1538 (
      {stage2_58[14]},
      {stage3_58[4]}
   );
   gpc1_1 gpc1539 (
      {stage2_58[15]},
      {stage3_58[5]}
   );
   gpc1_1 gpc1540 (
      {stage2_58[16]},
      {stage3_58[6]}
   );
   gpc1_1 gpc1541 (
      {stage2_58[17]},
      {stage3_58[7]}
   );
   gpc1_1 gpc1542 (
      {stage2_59[17]},
      {stage3_59[5]}
   );
   gpc1_1 gpc1543 (
      {stage2_59[18]},
      {stage3_59[6]}
   );
   gpc1_1 gpc1544 (
      {stage2_59[19]},
      {stage3_59[7]}
   );
   gpc1_1 gpc1545 (
      {stage2_60[6]},
      {stage3_60[6]}
   );
   gpc1_1 gpc1546 (
      {stage2_60[7]},
      {stage3_60[7]}
   );
   gpc1_1 gpc1547 (
      {stage2_60[8]},
      {stage3_60[8]}
   );
   gpc1_1 gpc1548 (
      {stage2_60[9]},
      {stage3_60[9]}
   );
   gpc1_1 gpc1549 (
      {stage2_60[10]},
      {stage3_60[10]}
   );
   gpc1_1 gpc1550 (
      {stage2_60[11]},
      {stage3_60[11]}
   );
   gpc1_1 gpc1551 (
      {stage2_60[12]},
      {stage3_60[12]}
   );
   gpc1_1 gpc1552 (
      {stage2_60[13]},
      {stage3_60[13]}
   );
   gpc1_1 gpc1553 (
      {stage2_61[13]},
      {stage3_61[5]}
   );
   gpc1_1 gpc1554 (
      {stage2_61[14]},
      {stage3_61[6]}
   );
   gpc1_1 gpc1555 (
      {stage2_62[12]},
      {stage3_62[4]}
   );
   gpc1_1 gpc1556 (
      {stage2_63[12]},
      {stage3_63[5]}
   );
   gpc1_1 gpc1557 (
      {stage2_65[6]},
      {stage3_65[4]}
   );
   gpc1_1 gpc1558 (
      {stage2_65[7]},
      {stage3_65[5]}
   );
   gpc1_1 gpc1559 (
      {stage2_67[1]},
      {stage3_67[2]}
   );
   gpc135_4 gpc1560 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4]},
      {stage3_1[0], stage3_1[1], stage3_1[2]},
      {stage3_2[0]},
      {stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc1325_5 gpc1561 (
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4]},
      {stage3_4[0], stage3_4[1]},
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[0]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[1]}
   );
   gpc1163_5 gpc1562 (
      {stage3_4[2], stage3_4[3], stage3_4[4]},
      {stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6], stage3_5[7], stage3_5[8]},
      {stage3_6[1]},
      {stage3_7[0]},
      {stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1],stage4_4[1]}
   );
   gpc606_5 gpc1563 (
      {stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5], stage3_6[6], stage3_6[7]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[2],stage4_6[2]}
   );
   gpc615_5 gpc1564 (
      {stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[3]}
   );
   gpc615_5 gpc1565 (
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10]},
      {stage3_8[7]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[2],stage4_9[2],stage4_8[3],stage4_7[4]}
   );
   gpc207_4 gpc1566 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage3_12[0], stage3_12[1]},
      {stage4_13[0],stage4_12[0],stage4_11[2],stage4_10[3]}
   );
   gpc135_4 gpc1567 (
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4]},
      {stage3_12[2], stage3_12[3], stage3_12[4]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[1],stage4_12[1],stage4_11[3]}
   );
   gpc135_4 gpc1568 (
      {stage3_11[5], stage3_11[6], stage3_11[7], stage3_11[8], 1'b0},
      {stage3_12[5], stage3_12[6], stage3_12[7]},
      {stage3_13[1]},
      {stage4_14[1],stage4_13[2],stage4_12[2],stage4_11[4]}
   );
   gpc117_4 gpc1569 (
      {stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7], stage3_13[8]},
      {stage3_14[0]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[2],stage4_13[3]}
   );
   gpc7_3 gpc1570 (
      {stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6], 1'b0},
      {stage4_16[1],stage4_15[1],stage4_14[3]}
   );
   gpc117_4 gpc1571 (
      {stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5], stage3_15[6], stage3_15[7]},
      {stage3_16[0]},
      {stage3_17[0]},
      {stage4_18[0],stage4_17[0],stage4_16[2],stage4_15[2]}
   );
   gpc606_5 gpc1572 (
      {stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5], stage3_16[6]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[1],stage4_16[3]}
   );
   gpc606_5 gpc1573 (
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[1],stage4_19[1],stage4_18[2],stage4_17[2]}
   );
   gpc117_4 gpc1574 (
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12]},
      {stage3_19[6]},
      {stage3_20[0]},
      {stage4_21[1],stage4_20[2],stage4_19[2],stage4_18[3]}
   );
   gpc606_5 gpc1575 (
      {stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5], 1'b0},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[0],stage4_22[0],stage4_21[2],stage4_20[3]}
   );
   gpc215_4 gpc1576 (
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4]},
      {stage3_22[6]},
      {stage3_23[0], stage3_23[1]},
      {stage4_24[1],stage4_23[1],stage4_22[1],stage4_21[3]}
   );
   gpc615_5 gpc1577 (
      {stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5], stage3_23[6]},
      {stage3_24[0]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[0],stage4_25[0],stage4_24[2],stage4_23[2]}
   );
   gpc606_5 gpc1578 (
      {stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5], stage3_24[6]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage4_28[0],stage4_27[1],stage4_26[1],stage4_25[1],stage4_24[3]}
   );
   gpc606_5 gpc1579 (
      {stage3_25[6], stage3_25[7], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[1],stage4_27[2],stage4_26[2],stage4_25[2]}
   );
   gpc2135_5 gpc1580 (
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4]},
      {stage3_29[0], stage3_29[1], stage3_29[2]},
      {stage3_30[0]},
      {stage3_31[0], stage3_31[1]},
      {stage4_32[0],stage4_31[0],stage4_30[0],stage4_29[1],stage4_28[2]}
   );
   gpc2135_5 gpc1581 (
      {stage3_28[5], stage3_28[6], stage3_28[7], stage3_28[8], 1'b0},
      {stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage3_30[1]},
      {stage3_31[2], stage3_31[3]},
      {stage4_32[1],stage4_31[1],stage4_30[1],stage4_29[2],stage4_28[3]}
   );
   gpc1343_5 gpc1582 (
      {stage3_29[6], stage3_29[7], stage3_29[8]},
      {stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[4], stage3_31[5], stage3_31[6]},
      {stage3_32[0]},
      {stage4_33[0],stage4_32[2],stage4_31[2],stage4_30[2],stage4_29[3]}
   );
   gpc7_3 gpc1583 (
      {stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5], stage3_32[6], 1'b0},
      {stage4_34[0],stage4_33[1],stage4_32[3]}
   );
   gpc2135_5 gpc1584 (
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4]},
      {stage3_34[0], stage3_34[1], stage3_34[2]},
      {stage3_35[0]},
      {stage3_36[0], stage3_36[1]},
      {stage4_37[0],stage4_36[0],stage4_35[0],stage4_34[1],stage4_33[2]}
   );
   gpc2135_5 gpc1585 (
      {stage3_33[5], stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9]},
      {stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage3_35[1]},
      {stage3_36[2], stage3_36[3]},
      {stage4_37[1],stage4_36[1],stage4_35[1],stage4_34[2],stage4_33[3]}
   );
   gpc606_5 gpc1586 (
      {stage3_33[10], stage3_33[11], stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15]},
      {stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5], 1'b0, 1'b0},
      {stage4_37[2],stage4_36[2],stage4_35[2],stage4_34[3],stage4_33[4]}
   );
   gpc606_5 gpc1587 (
      {stage3_36[4], stage3_36[5], stage3_36[6], stage3_36[7], stage3_36[8], stage3_36[9]},
      {stage3_38[0], stage3_38[1], stage3_38[2], stage3_38[3], stage3_38[4], stage3_38[5]},
      {stage4_40[0],stage4_39[0],stage4_38[0],stage4_37[3],stage4_36[3]}
   );
   gpc606_5 gpc1588 (
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[1],stage4_39[1],stage4_38[1],stage4_37[4]}
   );
   gpc615_5 gpc1589 (
      {stage3_38[6], stage3_38[7], stage3_38[8], stage3_38[9], stage3_38[10]},
      {stage3_39[6]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[1],stage4_40[2],stage4_39[2],stage4_38[2]}
   );
   gpc207_4 gpc1590 (
      {stage3_41[0], stage3_41[1], stage3_41[2], stage3_41[3], stage3_41[4], stage3_41[5], stage3_41[6]},
      {stage3_43[0], stage3_43[1]},
      {stage4_44[0],stage4_43[0],stage4_42[1],stage4_41[2]}
   );
   gpc207_4 gpc1591 (
      {stage3_41[7], stage3_41[8], stage3_41[9], stage3_41[10], stage3_41[11], stage3_41[12], stage3_41[13]},
      {stage3_43[2], stage3_43[3]},
      {stage4_44[1],stage4_43[1],stage4_42[2],stage4_41[3]}
   );
   gpc615_5 gpc1592 (
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], 1'b0},
      {stage3_43[4]},
      {stage3_44[0], stage3_44[1], stage3_44[2], stage3_44[3], stage3_44[4], stage3_44[5]},
      {stage4_46[0],stage4_45[0],stage4_44[2],stage4_43[2],stage4_42[3]}
   );
   gpc2135_5 gpc1593 (
      {stage3_44[6], stage3_44[7], stage3_44[8], stage3_44[9], stage3_44[10]},
      {stage3_45[0], stage3_45[1], stage3_45[2]},
      {stage3_46[0]},
      {stage3_47[0], stage3_47[1]},
      {stage4_48[0],stage4_47[0],stage4_46[1],stage4_45[1],stage4_44[3]}
   );
   gpc2135_5 gpc1594 (
      {stage3_44[11], stage3_44[12], stage3_44[13], stage3_44[14], stage3_44[15]},
      {stage3_45[3], stage3_45[4], 1'b0},
      {stage3_46[1]},
      {stage3_47[2], stage3_47[3]},
      {stage4_48[1],stage4_47[1],stage4_46[2],stage4_45[2],stage4_44[4]}
   );
   gpc615_5 gpc1595 (
      {stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5], stage3_46[6]},
      {stage3_47[4]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[0],stage4_48[2],stage4_47[2],stage4_46[3]}
   );
   gpc1406_5 gpc1596 (
      {stage3_47[5], stage3_47[6], stage3_47[7], stage3_47[8], 1'b0, 1'b0},
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3]},
      {stage3_50[0]},
      {stage4_51[0],stage4_50[1],stage4_49[1],stage4_48[3],stage4_47[3]}
   );
   gpc615_5 gpc1597 (
      {stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5]},
      {stage3_51[0]},
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5]},
      {stage4_54[0],stage4_53[0],stage4_52[0],stage4_51[1],stage4_50[2]}
   );
   gpc615_5 gpc1598 (
      {stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5]},
      {stage3_52[6]},
      {stage3_53[0], stage3_53[1], stage3_53[2], stage3_53[3], stage3_53[4], stage3_53[5]},
      {stage4_55[0],stage4_54[1],stage4_53[1],stage4_52[1],stage4_51[2]}
   );
   gpc606_5 gpc1599 (
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage3_56[0], stage3_56[1], stage3_56[2], stage3_56[3], stage3_56[4], stage3_56[5]},
      {stage4_58[0],stage4_57[0],stage4_56[0],stage4_55[1],stage4_54[2]}
   );
   gpc606_5 gpc1600 (
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3], stage3_55[4], stage3_55[5]},
      {stage3_57[0], stage3_57[1], stage3_57[2], stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage4_59[0],stage4_58[1],stage4_57[1],stage4_56[1],stage4_55[2]}
   );
   gpc615_5 gpc1601 (
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4]},
      {stage3_59[0]},
      {stage3_60[0], stage3_60[1], stage3_60[2], stage3_60[3], stage3_60[4], stage3_60[5]},
      {stage4_62[0],stage4_61[0],stage4_60[0],stage4_59[1],stage4_58[2]}
   );
   gpc7_3 gpc1602 (
      {stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5], stage3_59[6], stage3_59[7]},
      {stage4_61[1],stage4_60[1],stage4_59[2]}
   );
   gpc615_5 gpc1603 (
      {stage3_60[6], stage3_60[7], stage3_60[8], stage3_60[9], stage3_60[10]},
      {stage3_61[0]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], 1'b0},
      {stage4_64[0],stage4_63[0],stage4_62[1],stage4_61[2],stage4_60[2]}
   );
   gpc615_5 gpc1604 (
      {stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5]},
      {1'b0},
      {stage3_63[0], stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5]},
      {stage4_65[0],stage4_64[1],stage4_63[1],stage4_62[2],stage4_61[3]}
   );
   gpc1325_5 gpc1605 (
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4]},
      {stage3_66[0], stage3_66[1]},
      {stage3_67[0], stage3_67[1], stage3_67[2]},
      {stage3_68[0]},
      {stage4_69[0],stage4_68[0],stage4_67[0],stage4_66[0],stage4_65[1]}
   );
   gpc1_1 gpc1606 (
      {stage3_0[5]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1607 (
      {stage3_1[3]},
      {stage4_1[1]}
   );
   gpc1_1 gpc1608 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc1609 (
      {stage3_2[2]},
      {stage4_2[2]}
   );
   gpc1_1 gpc1610 (
      {stage3_4[5]},
      {stage4_4[2]}
   );
   gpc1_1 gpc1611 (
      {stage3_4[6]},
      {stage4_4[3]}
   );
   gpc1_1 gpc1612 (
      {stage3_8[8]},
      {stage4_8[4]}
   );
   gpc1_1 gpc1613 (
      {stage3_15[8]},
      {stage4_15[3]}
   );
   gpc1_1 gpc1614 (
      {stage3_16[7]},
      {stage4_16[4]}
   );
   gpc1_1 gpc1615 (
      {stage3_21[5]},
      {stage4_21[4]}
   );
   gpc1_1 gpc1616 (
      {stage3_21[6]},
      {stage4_21[5]}
   );
   gpc1_1 gpc1617 (
      {stage3_21[7]},
      {stage4_21[6]}
   );
   gpc1_1 gpc1618 (
      {stage3_21[8]},
      {stage4_21[7]}
   );
   gpc1_1 gpc1619 (
      {stage3_23[7]},
      {stage4_23[3]}
   );
   gpc1_1 gpc1620 (
      {stage3_26[6]},
      {stage4_26[3]}
   );
   gpc1_1 gpc1621 (
      {stage3_27[6]},
      {stage4_27[3]}
   );
   gpc1_1 gpc1622 (
      {stage3_33[16]},
      {stage4_33[5]}
   );
   gpc1_1 gpc1623 (
      {stage3_34[6]},
      {stage4_34[4]}
   );
   gpc1_1 gpc1624 (
      {stage3_43[5]},
      {stage4_43[3]}
   );
   gpc1_1 gpc1625 (
      {stage3_44[16]},
      {stage4_44[5]}
   );
   gpc1_1 gpc1626 (
      {stage3_49[4]},
      {stage4_49[2]}
   );
   gpc1_1 gpc1627 (
      {stage3_49[5]},
      {stage4_49[3]}
   );
   gpc1_1 gpc1628 (
      {stage3_50[6]},
      {stage4_50[3]}
   );
   gpc1_1 gpc1629 (
      {stage3_51[6]},
      {stage4_51[3]}
   );
   gpc1_1 gpc1630 (
      {stage3_51[7]},
      {stage4_51[4]}
   );
   gpc1_1 gpc1631 (
      {stage3_51[8]},
      {stage4_51[5]}
   );
   gpc1_1 gpc1632 (
      {stage3_55[6]},
      {stage4_55[3]}
   );
   gpc1_1 gpc1633 (
      {stage3_55[7]},
      {stage4_55[4]}
   );
   gpc1_1 gpc1634 (
      {stage3_55[8]},
      {stage4_55[5]}
   );
   gpc1_1 gpc1635 (
      {stage3_55[9]},
      {stage4_55[6]}
   );
   gpc1_1 gpc1636 (
      {stage3_57[6]},
      {stage4_57[2]}
   );
   gpc1_1 gpc1637 (
      {stage3_57[7]},
      {stage4_57[3]}
   );
   gpc1_1 gpc1638 (
      {stage3_58[5]},
      {stage4_58[3]}
   );
   gpc1_1 gpc1639 (
      {stage3_58[6]},
      {stage4_58[4]}
   );
   gpc1_1 gpc1640 (
      {stage3_58[7]},
      {stage4_58[5]}
   );
   gpc1_1 gpc1641 (
      {stage3_60[11]},
      {stage4_60[3]}
   );
   gpc1_1 gpc1642 (
      {stage3_60[12]},
      {stage4_60[4]}
   );
   gpc1_1 gpc1643 (
      {stage3_60[13]},
      {stage4_60[5]}
   );
   gpc1_1 gpc1644 (
      {stage3_61[6]},
      {stage4_61[4]}
   );
   gpc1_1 gpc1645 (
      {stage3_64[0]},
      {stage4_64[2]}
   );
   gpc1_1 gpc1646 (
      {stage3_64[1]},
      {stage4_64[3]}
   );
   gpc1_1 gpc1647 (
      {stage3_64[2]},
      {stage4_64[4]}
   );
   gpc1_1 gpc1648 (
      {stage3_64[3]},
      {stage4_64[5]}
   );
   gpc1_1 gpc1649 (
      {stage3_64[4]},
      {stage4_64[6]}
   );
   gpc1_1 gpc1650 (
      {stage3_65[5]},
      {stage4_65[2]}
   );
   gpc1_1 gpc1651 (
      {stage3_66[2]},
      {stage4_66[1]}
   );
   gpc1343_5 gpc1652 (
      {stage4_2[0], stage4_2[1], stage4_2[2]},
      {stage4_3[0], stage4_3[1], 1'b0, 1'b0},
      {stage4_4[0], stage4_4[1], stage4_4[2]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0]}
   );
   gpc623_5 gpc1653 (
      {stage4_6[0], stage4_6[1], stage4_6[2]},
      {stage4_7[0], stage4_7[1]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], 1'b0},
      {stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[1]}
   );
   gpc3_2 gpc1654 (
      {stage4_7[2], stage4_7[3], stage4_7[4]},
      {stage5_8[1],stage5_7[1]}
   );
   gpc1343_5 gpc1655 (
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[1]}
   );
   gpc1423_5 gpc1656 (
      {stage4_11[3], stage4_11[4], 1'b0},
      {stage4_12[1], stage4_12[2]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3]},
      {stage4_14[0]},
      {stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1]}
   );
   gpc1343_5 gpc1657 (
      {stage4_14[1], stage4_14[2], stage4_14[3]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3]},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[1]}
   );
   gpc1423_5 gpc1658 (
      {stage4_16[3], stage4_16[4], 1'b0},
      {stage4_17[1], stage4_17[2]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3]},
      {stage4_19[0]},
      {stage5_20[0],stage5_19[0],stage5_18[1],stage5_17[1],stage5_16[1]}
   );
   gpc1343_5 gpc1659 (
      {stage4_19[1], stage4_19[2], 1'b0},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3]},
      {stage4_21[0], stage4_21[1], stage4_21[2]},
      {stage4_22[0]},
      {stage5_23[0],stage5_22[0],stage5_21[0],stage5_20[1],stage5_19[1]}
   );
   gpc615_5 gpc1660 (
      {stage4_21[3], stage4_21[4], stage4_21[5], stage4_21[6], stage4_21[7]},
      {stage4_22[1]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], 1'b0, 1'b0},
      {stage5_25[0],stage5_24[0],stage5_23[1],stage5_22[1],stage5_21[1]}
   );
   gpc135_4 gpc1661 (
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], 1'b0},
      {stage4_25[0], stage4_25[1], stage4_25[2]},
      {stage4_26[0]},
      {stage5_27[0],stage5_26[0],stage5_25[1],stage5_24[1]}
   );
   gpc1343_5 gpc1662 (
      {stage4_26[1], stage4_26[2], stage4_26[3]},
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3]},
      {stage4_28[0], stage4_28[1], stage4_28[2]},
      {stage4_29[0]},
      {stage5_30[0],stage5_29[0],stage5_28[0],stage5_27[1],stage5_26[1]}
   );
   gpc135_4 gpc1663 (
      {stage4_29[1], stage4_29[2], stage4_29[3], 1'b0, 1'b0},
      {stage4_30[0], stage4_30[1], stage4_30[2]},
      {stage4_31[0]},
      {stage5_32[0],stage5_31[0],stage5_30[1],stage5_29[1]}
   );
   gpc1343_5 gpc1664 (
      {stage4_31[1], stage4_31[2], 1'b0},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3]},
      {stage4_33[0], stage4_33[1], stage4_33[2]},
      {stage4_34[0]},
      {stage5_35[0],stage5_34[0],stage5_33[0],stage5_32[1],stage5_31[1]}
   );
   gpc1343_5 gpc1665 (
      {stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4]},
      {stage4_35[0], stage4_35[1], stage4_35[2]},
      {stage4_36[0]},
      {stage5_37[0],stage5_36[0],stage5_35[1],stage5_34[1],stage5_33[1]}
   );
   gpc1163_5 gpc1666 (
      {stage4_36[1], stage4_36[2], stage4_36[3]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], 1'b0},
      {stage4_38[0]},
      {stage4_39[0]},
      {stage5_40[0],stage5_39[0],stage5_38[0],stage5_37[1],stage5_36[1]}
   );
   gpc1423_5 gpc1667 (
      {stage4_38[1], stage4_38[2], 1'b0},
      {stage4_39[1], stage4_39[2]},
      {stage4_40[0], stage4_40[1], stage4_40[2], 1'b0},
      {stage4_41[0]},
      {stage5_42[0],stage5_41[0],stage5_40[1],stage5_39[1],stage5_38[1]}
   );
   gpc1343_5 gpc1668 (
      {stage4_41[1], stage4_41[2], stage4_41[3]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3]},
      {stage4_43[0], stage4_43[1], stage4_43[2]},
      {stage4_44[0]},
      {stage5_45[0],stage5_44[0],stage5_43[0],stage5_42[1],stage5_41[1]}
   );
   gpc135_4 gpc1669 (
      {stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage4_45[0], stage4_45[1], stage4_45[2]},
      {stage4_46[0]},
      {stage5_47[0],stage5_46[0],stage5_45[1],stage5_44[1]}
   );
   gpc1343_5 gpc1670 (
      {stage4_46[1], stage4_46[2], stage4_46[3]},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3]},
      {stage4_48[0], stage4_48[1], stage4_48[2]},
      {stage4_49[0]},
      {stage5_50[0],stage5_49[0],stage5_48[0],stage5_47[1],stage5_46[1]}
   );
   gpc1163_5 gpc1671 (
      {stage4_49[1], stage4_49[2], stage4_49[3]},
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3], 1'b0, 1'b0},
      {stage4_51[0]},
      {stage4_52[0]},
      {stage5_53[0],stage5_52[0],stage5_51[0],stage5_50[1],stage5_49[1]}
   );
   gpc215_4 gpc1672 (
      {stage4_51[1], stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5]},
      {stage4_52[1]},
      {stage4_53[0], stage4_53[1]},
      {stage5_54[0],stage5_53[1],stage5_52[1],stage5_51[1]}
   );
   gpc3_2 gpc1673 (
      {stage4_54[0], stage4_54[1], stage4_54[2]},
      {stage5_55[0],stage5_54[1]}
   );
   gpc7_3 gpc1674 (
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5], stage4_55[6]},
      {stage5_57[0],stage5_56[0],stage5_55[1]}
   );
   gpc1343_5 gpc1675 (
      {stage4_56[0], stage4_56[1], 1'b0},
      {stage4_57[0], stage4_57[1], stage4_57[2], stage4_57[3]},
      {stage4_58[0], stage4_58[1], stage4_58[2]},
      {stage4_59[0]},
      {stage5_60[0],stage5_59[0],stage5_58[0],stage5_57[1],stage5_56[1]}
   );
   gpc623_5 gpc1676 (
      {stage4_58[3], stage4_58[4], stage4_58[5]},
      {stage4_59[1], stage4_59[2]},
      {stage4_60[0], stage4_60[1], stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5]},
      {stage5_62[0],stage5_61[0],stage5_60[1],stage5_59[1],stage5_58[1]}
   );
   gpc2135_5 gpc1677 (
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4]},
      {stage4_62[0], stage4_62[1], stage4_62[2]},
      {stage4_63[0]},
      {stage4_64[0], stage4_64[1]},
      {stage5_65[0],stage5_64[0],stage5_63[0],stage5_62[1],stage5_61[1]}
   );
   gpc2135_5 gpc1678 (
      {stage4_64[2], stage4_64[3], stage4_64[4], stage4_64[5], stage4_64[6]},
      {stage4_65[0], stage4_65[1], stage4_65[2]},
      {stage4_66[0]},
      {stage4_67[0], 1'b0},
      {stage5_68[0],stage5_67[0],stage5_66[0],stage5_65[1],stage5_64[1]}
   );
   gpc1_1 gpc1679 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1680 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1681 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc1682 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1683 (
      {stage4_4[3]},
      {stage5_4[1]}
   );
   gpc1_1 gpc1684 (
      {stage4_5[1]},
      {stage5_5[1]}
   );
   gpc1_1 gpc1685 (
      {stage4_28[3]},
      {stage5_28[1]}
   );
   gpc1_1 gpc1686 (
      {stage4_43[3]},
      {stage5_43[1]}
   );
   gpc1_1 gpc1687 (
      {stage4_48[3]},
      {stage5_48[1]}
   );
   gpc1_1 gpc1688 (
      {stage4_63[1]},
      {stage5_63[1]}
   );
   gpc1_1 gpc1689 (
      {stage4_66[1]},
      {stage5_66[1]}
   );
   gpc1_1 gpc1690 (
      {stage4_68[0]},
      {stage5_68[1]}
   );
   gpc1_1 gpc1691 (
      {stage4_69[0]},
      {stage5_69[0]}
   );
endmodule
module rowadder2_1_70(input [69:0] src0, input [69:0] src1, output [70:0] dst0);
    wire [69:0] gene;
    wire [69:0] prop;
    wire [71:0] out;
    wire [71:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_24_gene (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(gene[24])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_24_prop (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(prop[24])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_25_gene (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(gene[25])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_25_prop (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(prop[25])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_26_gene (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(gene[26])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_26_prop (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(prop[26])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_27_gene (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(gene[27])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_27_prop (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(prop[27])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_28_gene (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(gene[28])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_28_prop (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(prop[28])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_29_gene (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(gene[29])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_29_prop (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(prop[29])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_30_gene (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(gene[30])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_30_prop (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(prop[30])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_31_gene (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(gene[31])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_31_prop (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(prop[31])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_32_gene (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(gene[32])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_32_prop (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(prop[32])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_33_gene (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(gene[33])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_33_prop (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(prop[33])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_34_gene (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(gene[34])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_34_prop (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(prop[34])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_35_gene (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(gene[35])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_35_prop (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(prop[35])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_36_gene (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(gene[36])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_36_prop (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(prop[36])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_37_gene (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(gene[37])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_37_prop (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(prop[37])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_38_gene (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(gene[38])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_38_prop (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(prop[38])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_39_gene (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(gene[39])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_39_prop (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(prop[39])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_40_gene (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(gene[40])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_40_prop (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(prop[40])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_41_gene (
        .I0(src0[41]),
        .I1(src1[41]),
        .O(gene[41])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_41_prop (
        .I0(src0[41]),
        .I1(src1[41]),
        .O(prop[41])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_42_gene (
        .I0(src0[42]),
        .I1(src1[42]),
        .O(gene[42])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_42_prop (
        .I0(src0[42]),
        .I1(src1[42]),
        .O(prop[42])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_43_gene (
        .I0(src0[43]),
        .I1(src1[43]),
        .O(gene[43])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_43_prop (
        .I0(src0[43]),
        .I1(src1[43]),
        .O(prop[43])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_44_gene (
        .I0(src0[44]),
        .I1(src1[44]),
        .O(gene[44])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_44_prop (
        .I0(src0[44]),
        .I1(src1[44]),
        .O(prop[44])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_45_gene (
        .I0(src0[45]),
        .I1(src1[45]),
        .O(gene[45])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_45_prop (
        .I0(src0[45]),
        .I1(src1[45]),
        .O(prop[45])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_46_gene (
        .I0(src0[46]),
        .I1(src1[46]),
        .O(gene[46])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_46_prop (
        .I0(src0[46]),
        .I1(src1[46]),
        .O(prop[46])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_47_gene (
        .I0(src0[47]),
        .I1(src1[47]),
        .O(gene[47])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_47_prop (
        .I0(src0[47]),
        .I1(src1[47]),
        .O(prop[47])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_48_gene (
        .I0(src0[48]),
        .I1(src1[48]),
        .O(gene[48])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_48_prop (
        .I0(src0[48]),
        .I1(src1[48]),
        .O(prop[48])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_49_gene (
        .I0(src0[49]),
        .I1(src1[49]),
        .O(gene[49])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_49_prop (
        .I0(src0[49]),
        .I1(src1[49]),
        .O(prop[49])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_50_gene (
        .I0(src0[50]),
        .I1(src1[50]),
        .O(gene[50])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_50_prop (
        .I0(src0[50]),
        .I1(src1[50]),
        .O(prop[50])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_51_gene (
        .I0(src0[51]),
        .I1(src1[51]),
        .O(gene[51])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_51_prop (
        .I0(src0[51]),
        .I1(src1[51]),
        .O(prop[51])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_52_gene (
        .I0(src0[52]),
        .I1(src1[52]),
        .O(gene[52])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_52_prop (
        .I0(src0[52]),
        .I1(src1[52]),
        .O(prop[52])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_53_gene (
        .I0(src0[53]),
        .I1(src1[53]),
        .O(gene[53])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_53_prop (
        .I0(src0[53]),
        .I1(src1[53]),
        .O(prop[53])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_54_gene (
        .I0(src0[54]),
        .I1(src1[54]),
        .O(gene[54])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_54_prop (
        .I0(src0[54]),
        .I1(src1[54]),
        .O(prop[54])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_55_gene (
        .I0(src0[55]),
        .I1(src1[55]),
        .O(gene[55])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_55_prop (
        .I0(src0[55]),
        .I1(src1[55]),
        .O(prop[55])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_56_gene (
        .I0(src0[56]),
        .I1(src1[56]),
        .O(gene[56])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_56_prop (
        .I0(src0[56]),
        .I1(src1[56]),
        .O(prop[56])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_57_gene (
        .I0(src0[57]),
        .I1(src1[57]),
        .O(gene[57])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_57_prop (
        .I0(src0[57]),
        .I1(src1[57]),
        .O(prop[57])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_58_gene (
        .I0(src0[58]),
        .I1(src1[58]),
        .O(gene[58])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_58_prop (
        .I0(src0[58]),
        .I1(src1[58]),
        .O(prop[58])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_59_gene (
        .I0(src0[59]),
        .I1(src1[59]),
        .O(gene[59])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_59_prop (
        .I0(src0[59]),
        .I1(src1[59]),
        .O(prop[59])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_60_gene (
        .I0(src0[60]),
        .I1(src1[60]),
        .O(gene[60])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_60_prop (
        .I0(src0[60]),
        .I1(src1[60]),
        .O(prop[60])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_61_gene (
        .I0(src0[61]),
        .I1(src1[61]),
        .O(gene[61])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_61_prop (
        .I0(src0[61]),
        .I1(src1[61]),
        .O(prop[61])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_62_gene (
        .I0(src0[62]),
        .I1(src1[62]),
        .O(gene[62])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_62_prop (
        .I0(src0[62]),
        .I1(src1[62]),
        .O(prop[62])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_63_gene (
        .I0(src0[63]),
        .I1(src1[63]),
        .O(gene[63])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_63_prop (
        .I0(src0[63]),
        .I1(src1[63]),
        .O(prop[63])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_64_gene (
        .I0(src0[64]),
        .I1(src1[64]),
        .O(gene[64])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_64_prop (
        .I0(src0[64]),
        .I1(src1[64]),
        .O(prop[64])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_65_gene (
        .I0(src0[65]),
        .I1(src1[65]),
        .O(gene[65])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_65_prop (
        .I0(src0[65]),
        .I1(src1[65]),
        .O(prop[65])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_66_gene (
        .I0(src0[66]),
        .I1(src1[66]),
        .O(gene[66])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_66_prop (
        .I0(src0[66]),
        .I1(src1[66]),
        .O(prop[66])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_67_gene (
        .I0(src0[67]),
        .I1(src1[67]),
        .O(gene[67])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_67_prop (
        .I0(src0[67]),
        .I1(src1[67]),
        .O(prop[67])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_68_gene (
        .I0(src0[68]),
        .I1(src1[68]),
        .O(gene[68])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_68_prop (
        .I0(src0[68]),
        .I1(src1[68]),
        .O(prop[68])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_69_gene (
        .I0(src0[69]),
        .I1(src1[69]),
        .O(gene[69])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_69_prop (
        .I0(src0[69]),
        .I1(src1[69]),
        .O(prop[69])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_27_24 (
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CI(carryout[23]),
        .CYINIT(1'h0),
        .DI(gene[27:24]),
        .S(prop[27:24])
    );
    CARRY4 carry4_31_28 (
        .CO(carryout[31:28]),
        .O(out[31:28]),
        .CI(carryout[27]),
        .CYINIT(1'h0),
        .DI(gene[31:28]),
        .S(prop[31:28])
    );
    CARRY4 carry4_35_32 (
        .CO(carryout[35:32]),
        .O(out[35:32]),
        .CI(carryout[31]),
        .CYINIT(1'h0),
        .DI(gene[35:32]),
        .S(prop[35:32])
    );
    CARRY4 carry4_39_36 (
        .CO(carryout[39:36]),
        .O(out[39:36]),
        .CI(carryout[35]),
        .CYINIT(1'h0),
        .DI(gene[39:36]),
        .S(prop[39:36])
    );
    CARRY4 carry4_43_40 (
        .CO(carryout[43:40]),
        .O(out[43:40]),
        .CI(carryout[39]),
        .CYINIT(1'h0),
        .DI(gene[43:40]),
        .S(prop[43:40])
    );
    CARRY4 carry4_47_44 (
        .CO(carryout[47:44]),
        .O(out[47:44]),
        .CI(carryout[43]),
        .CYINIT(1'h0),
        .DI(gene[47:44]),
        .S(prop[47:44])
    );
    CARRY4 carry4_51_48 (
        .CO(carryout[51:48]),
        .O(out[51:48]),
        .CI(carryout[47]),
        .CYINIT(1'h0),
        .DI(gene[51:48]),
        .S(prop[51:48])
    );
    CARRY4 carry4_55_52 (
        .CO(carryout[55:52]),
        .O(out[55:52]),
        .CI(carryout[51]),
        .CYINIT(1'h0),
        .DI(gene[55:52]),
        .S(prop[55:52])
    );
    CARRY4 carry4_59_56 (
        .CO(carryout[59:56]),
        .O(out[59:56]),
        .CI(carryout[55]),
        .CYINIT(1'h0),
        .DI(gene[59:56]),
        .S(prop[59:56])
    );
    CARRY4 carry4_63_60 (
        .CO(carryout[63:60]),
        .O(out[63:60]),
        .CI(carryout[59]),
        .CYINIT(1'h0),
        .DI(gene[63:60]),
        .S(prop[63:60])
    );
    CARRY4 carry4_67_64 (
        .CO(carryout[67:64]),
        .O(out[67:64]),
        .CI(carryout[63]),
        .CYINIT(1'h0),
        .DI(gene[67:64]),
        .S(prop[67:64])
    );
    CARRY4 carry4_71_68 (
        .CO(carryout[71:68]),
        .O(out[71:68]),
        .CI(carryout[67]),
        .CYINIT(1'h0),
        .DI({2'h0, gene[69:68]}),
        .S({2'h0, prop[69:68]})
    );
    assign dst0 = {carryout[69], out[69:0]};
endmodule


module testbench();
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    reg [63:0] src16;
    reg [63:0] src17;
    reg [63:0] src18;
    reg [63:0] src19;
    reg [63:0] src20;
    reg [63:0] src21;
    reg [63:0] src22;
    reg [63:0] src23;
    reg [63:0] src24;
    reg [63:0] src25;
    reg [63:0] src26;
    reg [63:0] src27;
    reg [63:0] src28;
    reg [63:0] src29;
    reg [63:0] src30;
    reg [63:0] src31;
    reg [63:0] src32;
    reg [63:0] src33;
    reg [63:0] src34;
    reg [63:0] src35;
    reg [63:0] src36;
    reg [63:0] src37;
    reg [63:0] src38;
    reg [63:0] src39;
    reg [63:0] src40;
    reg [63:0] src41;
    reg [63:0] src42;
    reg [63:0] src43;
    reg [63:0] src44;
    reg [63:0] src45;
    reg [63:0] src46;
    reg [63:0] src47;
    reg [63:0] src48;
    reg [63:0] src49;
    reg [63:0] src50;
    reg [63:0] src51;
    reg [63:0] src52;
    reg [63:0] src53;
    reg [63:0] src54;
    reg [63:0] src55;
    reg [63:0] src56;
    reg [63:0] src57;
    reg [63:0] src58;
    reg [63:0] src59;
    reg [63:0] src60;
    reg [63:0] src61;
    reg [63:0] src62;
    reg [63:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [69:0] srcsum;
    wire [69:0] dstsum;
    wire test;
    compressor2_1_64_64 compressor2_1_64_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc8f276a24e25518b48fffcd47b51803a8d8fc18b3ffd991830917e2ab2a07b0bcfaae8bd4c025234f1171c331aa1a5a10cdffbd15cc36399c995196dd0c8a0e0555e9f0ab1a0499fbf80acba4b31141b5cc081ed3292939398a4fafa46a12a4e5264942894878c973567cdbda2126d76b3779f7e7304a5f7242f2572867eda59fa3dbf7bcd70e34d3e8125a534659a44096d359489da5207d7dc9cf12b2adf12373dbc099272c98003ee0c6555a9682da57557e7f547882c19166c41c1ecc29b42c1471509475b637eb75be7b4a0cdf265529d48c586a59606318ffcd95dfcea889993dc9e52417d88e598695ec0cf788c497fc4c835f882f0b4b48352c122e009e1e7e2b6fc62fdb70f52be4345692f49c54ed972b48b2e553e2c4c6503c1eaee27428c2ebb332a039599a1db14592358b802f543dd542122d06d4e151a3afe710983f32bb8ca4df03ee276d7d4be58571cd35c10869d015fe3502038e07c8c044fddb7aa9fdf428ff7e16e4223f426fe1470f239f32ba62d48cc2d29fd33e0204bd39ff98e9d70f5d64082fe749cb3b549524b1c18c41c0347b16154ba1246f9a62b5b428f71270beac44bacc480b4aeb333a52af315cd1b164b26f68e19d4322cd1f492323025141223bd1618c974fe98068d300037b36450f8b20a2460cc92eefefb5ace44c8329cfe57ba76dd6cb403c2790361809eff6f43c2ccb21dc1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h87e4bc0a8a64cc438628061bd2d6f5f18a0ffaedf72e1a62cb72cd569c2eee15b20fd2172cadbf38e92d5c57ec9fdf5155de06d5ff0379f10e915231ea7bd466e638e98a7c68dceebe205cadee4b12096ede9a2785a6f1b579905a0bec40d1d261485d7b62fa7ffa5620d784f314b0de9570cce2114814c2eba122a90521da8c8bf2e05bdf8fc9b4e2a9993cfa612b6185b00025df74745ef5d24edc9b689a016e509984f56e05f5d602050b8d57948b4e7ad2e6b412371834e8705368d1c5052c697d274751527ca5868561ec2ec67fd5d77952802dca6f5161709357547a6864ab86271abadd13e88101f8e13f0c458fd3bd242f63ea1eda5fe45124ae7764a755991a60b3bfcca079096db900806050cfa8846d426477650330512736b3273a8d6585ca8984dbb3a91686465ead509ce264269e22e6b38e91e8a1391e7788f960e2bddfef2236bbaa0499c07d56c28358d5a2e55578e863ad9bdb01561372167870e971508df8082b0359aace1315dbc8fb7397f7e75adc309a8933b6408cd3884313e2cf834bececceb59abd8f844f3308e49ab68b9dd12bed0ed623311d4b49b5ca78d5cd7bc5e779b3380ac03eb73ccf43cb82612ebd88e208af7337f7951a61c11d4a94ecea2631021bf51cdd7a3860b455672e9346835d98736904125d2f8893fa33641d273d7349f5f5a3cf0683c43f62b475616418096df77b83cb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h73ac18eb8575d0797c3d3b424b9f34a4dc94b3cfcd2e039cdd65fd5099cd5b4860fed3b5b63d0eef4f16c7d0b07863bc7fa2ae1adac65793533e8ad6b7b5f461e41a261fd669bafe1c28b756f047d4e9da7d4358010947861ed6e29254c1ac6c390c62a796062276b46a1db42395ab576d88634a6f0d6469ba60d409000ca3dcef8ca63d1a45a2c810ff124ca1e3e8d5d839ade5a6918944ebe87f2124ee0657598f6c0ac2d8cbf47b482c83cee132363eccf081a6f8ff3c315956908efc1b00804f258e9360c0d06d60f59cc855d9bba3df8599065949d2a09ba643da308107f07ed18d17328c2f979562f2570b4b3a5734d024dcdf041fb35542c79096ea3a54325b0a91c4e388828d3c090a8f8dc247dc52f88fd57bbd046e3350d7fe62e62910497ce06f13d43190ad43d96fd2fa7447ba75ec7ca172a5bcea611f980ea8ca69b201aac219bddcbbebe5917f9605a47dc342f74a83dc74add683bd6037a7e87b2d1afacc3770c3fa75ff7b48d03d6b38566cc99466aa01223370d216313d0e8576cb25f80d50bb795fe753e9bc1c7593ae373007a76b726cf2f616a3b807ef66d52947b08c17b14517c7d29650288e039808868f370f5cee3e53ed7513e54e51aa562b10bdf7329b202b273965c0e723b2b4b947bd559c51eedee0e6e34c18fd5a58ec17295b3e7538334637aea14048afa148899783bbfc1939555b4d16;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb7d38d9b684376fdc5f10a47e0fd447c93be6b428d0d3a7eebbcdfa45f5974e6a28c23cca842b4bd205b8d88887e70e83968046a265ce8a0f5f067c6c52428249e79003854dbe52b440ddc2ae51a7f92f8ce55f398fde3ddab6971725e5da4484bd8caed0d539fc67898bda822a98af17ce590782c73304d69221e6d97280afbdcbaf44120f10a63ffa493174af199540c4eaa5a4be2c14751cad0bda444e7de95f9f4f618641d737f3152981b27ca0a1ef2a80cb3497e9b4afdd5e0d47f7e71ed8fe9bc1f6fb043bca95b01ece237713b99cb366ac47d28052f2d012be3f7bf341d72b3747715f708f264e19ff79de69e9ce92cf7a5add1b1f4a661d528fdfd9401848ecd4c74ac26d2704a1da66ca7be3ce477adeffe2f049914caa1e36e554ae4d24a724941ad1738b74a419fd698bfcb004731b652dd7eb7be82217f020d94693bb092fd14f3bae8c7244255f4ba35450b552e42bbe99f0bebbd263a6b9cd81475c99d652f02fe501a3b9ac72f56aa7b9c9448c7bab2d771777793ec6d4944e3db4f3a8ac1367ee42c6beee6957b307d3147a9090c1207c99dce2e4d117719c1a5a48ece4d058ef6e193c6a2fed6d168c2ca3a1324d1fbb5242fe24070faf1a6cb622aa0a0878612083e5fac86460f327f8ceec99b06c67005a65999ad57861b04727ba652d98522e4dab5035bf2f70d47d9a7d12ce7371a39c7820b0f09;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hec98f3745ee3ab644c2a146f528f0663a35e12da63110eb76b99a2534a8f3d0170e42fd1d7f2ef5e6b6f711335359d4f4a44ec6b741de56739e97ad71552ab9c0212f227f38296c9b4b1d742d024e481ced1c026f29bf5519f3d763a7177204093222cdf917152855f142b9712ba207af5087835ae28efcc95fd2b8fab91062525ab4dc0a5c9391250151eccc4137733f41b383296d3539ab58885180acaee7bd407a7415e2d51d96ed74f5e974d11c7e02834ee1a333952916e0791c9c682ec5c2b3ce4baee2cffb9cf63a015e452d8d19566baedae1cd44008096244a711e323704c1bb92bdaa386ee80eed2180c8d761b8821eabf6436b1b5b5de5b4cd4df1ed722ac36f509c49593867aaabffa218fa04d5350296599009d9f39ebe374b7f9520b34e14609252f692eb1f155b0c1d0d1ae365e1e8739102ec193a013094cd5d817a0d8271ec5c43eb38b5f722f8a92aefecd04bc825d056f8f6f79b23a1923f8e421cbb89057905c49463ec2136f818aeea22bb3a5e91df7e08fa2351b5d2d0b24ba034134ef27d5d96abffede2de4d50fef110507c511199dfd3015ed75ece0acf2649be94054ae13d396f1f50b4bdb52d339cd147419cb7437cfd0be90c6223d04baac7c57704ef66805a89314ce13a9c230decf0946837def4d3d087b580bfe0fe9c73658001dfe59f726bc760f06e586a60e9302db1d191eac17e75;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4ff2616649094c3d4879c24bdf377dd905c9d721f658eb73e4414df21ad2be463b99c8c529016c909053e7e1e3869e1d075b496f027f88ec7b28c10c8f72ace3749f9aee78d993549ff137344e44cf01b977a7a6f641db6f9834a6b41677dffbff3197a1e53791bd449347beed5f936b085d12e66bb6aa6e58017c2ed46ebef400c0dad3604bcc922de2166a82243535ea70ce2bf698c6d87c74152f66b50e3835cc16453f905a779a8d509ccda9b17dfb4211596805d0131080579977028d8d6efa8ba53af9a15aed7ab19cb25e6b1f6237610f06f2c6f637ea03ff72f80e4ebec5d321d41b957dbbf6190b18b03d25ab32404922d0463cc8bb8d5e1761262910181edc5dda15e7b8e74c24e8574e1b090b4240381b9c58bf7d774e01711800bc9ab705430eab640d90953d34489bd9f01e19a2d8608bd94291f50cfad219bc5f1949b280f6ce93d802146898e96289de2a88f082bb0203c09fd18e8843231d561ff11425cfe5f77f577655bf69624b6eba7b5ef7b5d2040aa2e3454aee8100680c0c8305363710ce95e92d7a5e0c7b9f8c7675877a8c5cc040010ff72df3d768426ed6dda4f68a1e9133a8c3cb2790e34cebfb0fc5c28d8a066fa809d03d08c4a32044fbeb777e5ca3d58717f83e20c7c643435c5ac5192fca0e58727a2be7935a37ca1e749e67274b10e8b111559fe37ef8b7eacdff1271f3170b6867bd00;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'heb6fd35543cdbfdb74ed3bb25c87f61705535d5ec9c08544e929ac9c20d58b992dc95db0e26a620f72d992558738a19e6a45920bf172419afa6db3580ca0b8fba88cab53da921e63138afcc0a4d591598cf59ab7fc22c29fb1f816f7e83e64d66533d2d6e1ea5bca74a1f313ae5e5bf4f6f135e0746172f5f16d1f99f5e58fa7f7bf55cbf74b427d4fea0d9a889e8ce675ffa6cc3fcca6ffef7c117f4cec4dda8e4bbc6c68c8707725f11cb16d873658a4cfdc6522f73dcb6b1f956c975af7ce10babdc7257397aa823b0277fb67a8240e949afd745cba9385e66b64aee960bf8a723df661e85dc3745a1c0ac470d19bf3cb67a42525557dd6db45609dabfec23663fe1395b4fd605a2c8b4af84de3a2a82832f6183f3d0c0c795e0584812a0c7a50ea01f45a72c6af29723bc35acd3117de2a4f350493ad0a5cde8e5da499cedaae71f956689fd7c445cc9822e02870dd540bcce9d5c95e94dcce0a747f24547171c368b54c7570a79eb3fa1758585eee0054e6886e1fb69851564ef0dd22329de4fe2e828b1082e4a6eab2f861f14d2a657a0e9dff1feb557f045798ca2a41467069da7f76a56231fe4e1fafb1aa931137855bff694394d51dca8be6a73923cac98c40cd274f2a9fa0193be87da8581ca508c4f8444ffeb528668dcd68f7295d2131a2f5574479dbffb34c5dcdf88ba17e64ca49ccb1d8e175c367dda5a945;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h772dde7bba3ad67be7788d576d8ad90f2a95bcd691e3e4f937b54bb85b87e8cf9a8f4d55e0846b98374936575043d865874ea3093e5ab9ca72afa624e67116b89ff7ba1b3e6f7c3da59e4f8285ef5e30ac97ae76c8d0c94b196fd7f40ff5fdf17df20ed921676b7d27c4c6f864365b60ee65e13fb422d42d73617bf03fc5a069b63d25e893b0e397133dece179105f155bc9755262a0fb88879858190c09888e754ec91276665059f36a2c239b7b3435a87b47450999d6c315bd2338156cbbaba310e50d353dd5c9d80aecc7d5c5b05af0b53fa1917a650f411d83a0ee1e44f24f6f1b94055487d3e15cb999de4ace9879c2d773ba1c7be2ce19099c86cf1ca28d537a1870342185d4ee756be1531a83b2d713d6ac98fdb130feae716b603aea57433809f585cb81a2d0462c150652d2993540d7a79afc67e573399e5fecc7ae0c206e992ea105d54de43748f76a609ebb89c96896b2d363a72f06c06c36af113af9df315b6253a33060f563f4160cb0a6cf533801abfaeadb1a469e519ff1fa38a67b2fb03e4f71cc0f3428f655263133025bdd8008ecb0f6504424d9b89e942ff6802b406a923c3266a63557435e14606e5d084595f8f5671812ce75d53f8338be0a3c27c5294b10a22a2c31fde467eb8ab515d5db435ba1761ca40db3de926b422f9aaea0031df860a93c7e80f7ee1fadf9583bdb1f971e20bd677afb087b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hadbd2a3cdf54d8aca24a177876819fc6c0bf0b21d2604dd41b3f9d926de271c9e17a2fd42f4455cc4baa1f3ef780be25afb147183562b669224de9b400a6e08ed6c326d0f66d78fe1163f4762e625087ebf1b9c9cb80714baf25d981affc47ec76731a4a8ab8303f28b56b4e4990e67612343d67e0e96d0284ccc2d2584503e03c05d542b15dc363e074dd5fcfec86058cd4212665c0bf977e4ccf2df75a98b89de47c750f5f1d1fbc75a4127a3687164494a6535ab57fe7cfd48c966a428a25586cc773c13f378deb8e12a7428a040b640c3311c890b0a86011901fd3b71b3bd3ee28fd138b5d3a88f7b39dd28e18a563e8040845e66d6075c21081c3e8a5f4c60057a3c6a25a25983f22e3ea988af86b3b4ebdfb05ba3bceb207e21e565d790d2f79ec15b2368e50735d9185e13eecc9ad9c01c9698f11687e8382db3d925d5c62398ad18fb46eb04de0905eaa28e93c066f9a75048e58aa4022b052e28a52784118c4a5736b980898e312639622cea4786a774552fbf4a1c4c0d12f237b22e3e2474f0f1b4e0e11f85dd8d4501f85a44262d112384e9f734450fc114b0fe599e8ef4f57fdde5db9b66adcaaae185930293a07bf72c672843d6903764e4ea0445325c9a301185a55c5cc11ea783e6c17f90c82763b266aae1eb614f46756d6c135688f2c45f691a8ed366cea3eb2b72191af9c0432dfaa1124890a4026b1c8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h95c214e0bf2e80511fa5e38f19bdc298ae70123d8bee1ffcafb9642ab3dc39b510f1b86e2140315d46e593caf00274c468e50ccc313121c3176bc491d3a55f2376b29a796a703d64e1c0fd506df791847b78901278c1a406fb287bc554867a5e46f4d080adadd610a91152555b906f39b364236bf406297087283be11f16965470118d027cb110923c996557cfc3a8334534cfafba6c97d85b487b581b81f3272044e3ccfefa9b3aa13e7c07d3ac8dc7224cf2d3b56763659fd2e5a63dfa7ae0e35511f78c9e9cdc367a33a4c68cec71c014a2a45a93db3c16cf8e0e1d57dcb0065028b96e74660375ccfdcc5fc13820de5ec72bf11e95e5d164dbda8d89450cf824bae40f03da6cec1b2dd3872276a80dd485c9893ff79f6880fd6177b6b2177196f10d5ced4406c08afe88fc65b42ebb600976a4fd3a10e89f8bd6f076c8604f3bad33be488893f77059bc0b60d3596a160d2510168f13bc6469815fb1cfe257a20720a531c64c0c175a8e6a220f243794f08812aea79f1f705e1cec88a334455786f8f91df0fb24f570787ded2eb85c4f8e194e803723676c5e9a726cbadc5a04e955c24f25db206a89fd05c1fffc6f4576c490c3c534bd3f09937ed3702ed7373a396366de603c048b7419de9b00347ad2671c03f85f339f46f202602a30ff2ab7f5c3fef9f26622b03ff437a48edcdeb0f8cb2475d6f757d3ab3924437e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcff0c3554b962741bc616830cdcff00c88e5fa20d745b6c89a7f6fb8ff215bf4ae56b4fa1bc13b4cebfd713f7e19960c30cb63f613b6363b0f34d62b5828aa91954f7638cab00ae79f22a132e67d3b585b86b9ca4a73796f6932e567c2fc95d05cf035f80f02822d8072d1543cb5dfdf2f247d509e59d9fb52c72a80f6755455df7e329d4790d91640edcdf45d6a7b16b3d6998293babe070bbe1d6587f1a76601735673aa3028e23be0e409b52a72c623139b2c730edc65f8736faf3ff34e5dd66020c0dc60b84735a650a0a43d367b4a21bbdb45aabfde8c77c877a6c80c7c0dfb0f3820b6a0c6faba63b2e869c656167b54090ae4c5e678306d35967c96fee77c936886a0d2b67f1ea9c787c92d8d27a23d7766bfd99724422d9d5d31254a17ea6473f8a57eb5f41c8a3ec185c2bc38b4915cd37917ce1e61298e53a8e891db7bf76608c2f404c0668c92ccd61744465f43f4f549169b1f170ba2f1ef471e999b340d1372303525df1723b1e3ffd2c889731dde438c87fcf2f6f8774eea310ef8da25ab968a706c9449c0ec4fed283683d5bad3c91d0bada4f016c2a919208e3295ac38eb25e699b0e5d4edd6ed9ffd7966f32d0f93cdb7893b11b475e4652bb95354d51e8c5f908bc5e6bc47fd36f6571d76cd9bc772e9951026d6cacbbcfc873205bf2b032955b66f599c410ed4558784dee2c86f027caf1a8b4cdcc091;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8ee07a52cb7de267a8cc96e2a774730392bcf9d4d18de71395822915954ba4bdd337114725da1929479fc225a44731d5c21cce690d17a3e257729ce9e15f4d1da2cd903fc67e24d69f179420b3cf3258c14051484d470d633d9a23620b38f0985cfedf37a960db2fe68ca152adeb116cda878befe39bd258b73bcc4bb4f9ed5965330eea0c9798b0b15298776ad27f1b59e4a72258965e0d5600bbdbe5921702da6de2083eba7022b049f30cea14c6e7474d98915030f79cd21e423922ba3171b3082027192e62cf210e8ee3ea5c14e179714f1e03963ea2d72da3f37ca4d72d51e0738096ebfb7f270877e415e0948aec6a5d55d4de43ca187536c95e10fd150e68adbf2113b3fdd7813b266708fdb8e3a1ff2c5f13497d8638d2e91333863b7391ed462ab524785371749fcbf00089f8d3cc89dab323c337021d3e154e6393cc45d4a83fa18ac9461dad2e2aa5c765edff31dd6365d6d6d0f02fffd8322b634a0b0ca0ef879907cf469f08f58573f2c95ade9bb362140900cbfac7a2e82fbe4cf17fc20a5af20ffca39d4b056332514a1133b027c6d9e5335ddcafc9a1b80c9d60134608d34642435d39d11095a2587b6d57d9bb9a96001fc1bc9acc6cadeb23746d996e2023bcccea462362c70bf495132c817c59c0f2e2977db082e091d0340d7f9dda3a643c6fd45a7ffb18c005f8de3c1f2d0a3f2293d45e1264678374;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h39ef5e47740a762c3b9b73ca641fca17c8bc881bb727b6051b0c8d936c54313fdf9ab16fe27176df406bdd0445cab0f0478905a3e6a8c0fe2bb5392242accce2fce8505fb19f3dd49ff4bcf9ef686f93be4de05be686c11892582ac0387b6fe1f77f97e6f8933f5c46c44709aab9b4c46b23b6cdfe562a90969212559bdc7ed1f198f43bcdc3613a080f820f5681cff7b3183fba16cf89f1befd5d29ba5ade057386de84548887de7721376d93c49bae23f4ac25d0b8abb71f77b69836f7dcab833e80cc284a300f2126b49ed48e7939cbbd7cc9573de66c5c9d3b4b12d7cc2e02480807c8595e7fd665b29a3cff808e370070a1b956bb4711404d36aa9a5ca60f9ff131f8872331c87e33736cf204552c383107eeae7b6e0811588fc86db24069cb0b8136e8fd2280203e94ecdc2a13dbe67ec1ca4bd793bc57c62ba2aab3f4c2441718c7ef5a93579f5fcd8e74b69f9542bce5dbe2772584db5fceaaf1a32cc81604c401b32ec0ee9ea9b5c3ff2ac9301b1df0f23d64cb239240786d0f752aa62f95404bccd9e135007b688785f529e77c7d5fdad45546d4bc105e32f65ef47f9aa003b92364b8fba17aace8c770021b672285dd5d218f99563603ce4e90e213accb933e510580263f2a08a0a566d0bb4c8cb310ab948f89520eeee61ae1b31d942b2784d622096e264426f7a16e56c6f5d94a56bdbe88be4bd29a2dc0dd06;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h32a00108beaa628cc904d7b6652110c1e691fc64ed5bb827f611885570a336a0a7e9a52fd7438d3251433b781d0d4afcb47f85498a6adf2dd58aec4e440cf4e057bae90ea6bfa585400422796dd1baa68b52509f77ebb297aba5401a8e3b1c339fff1108a3df1d1cc3fc17da62d62ec90433986f9d3bdad533185010c004fc12342fb7e03aefee3c85a3104af081faeee42034cc6ef7108e28cbfafad6f16e9bb02b4e0fa5de550aa86298c27f18c4d383582ad9bf29eda9914cb19cac717d783be2da5ff187061b73054f8cdf6ed8925455ec64ee53da22223cd1672d42a63cb891542b28ab90e55b832781e05626a7fd0c75b3262144fd7bef543b518649d122c15cdaf810ec89187ac3747f469995a9b51cadf6753df5d0f0c7f0c7467d09ec2dd2c2032f63a25854ed27edf8b32b4d9f349e169bffc7905dd618563d7d8b153738b4dd4084736aad0de20637b1d7955786c847fe19c441c2193cd6d3a59dc9b1a841637d131abaedac5867aedc577d89c3f329e5312aaadbee0a644087495d65af4babd6b0d5f98a3277cbd03bbdcbacbeca88f53e3617b27337c826ba159a49ddf3da6c273180cea9b941412d06f721dcac875a12efebe873628b500056c286c3ddb7e3200eefb444a3d2c239976437cf6443be202d6772cc3615405f782d4901b225796b90ccc1f65404865006c907a1ecc94e4bf060616ee049d267f9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9252358ad5c7c51ed3b8e0d6248cd3eec1c8bcc95576f767a56be5361af03c8dff2126df9c5341b3b3a3744d4926ff74ae0ac7fc0ffaf895568334c6b11ca435eb69236550b13ce097184f56b9bb0bd6277b0d000e280e8887be66c5bf85fd98b36a162394fbec64140e9a761fbf76ced215a4fb0626cefc48761e3a898f57e9d0fe7a788d8ffaf0e234ce9abdf90377a5a9dfba24b5687b3675d940e31f8db6b1251d76362db530e1b05b7b676520e935c774de80bf3bb5aaff4b19fc382614f5f4eb5bd59be3c3660dfab0fed7a0a204c2e345668b938c63778de69cd8b0634a221ed604eb5779245181c5a68f91e0ef4c6d8b8b204326dd5c98525743fb9fdc41056b515bd3509d243264a24194d191252d9f119e0d3fb9477f871d64428dc5cca8bd7ebd83aa4530b9cc41237f694c9bb591aa4676ee42ad4c300ce776ec40ed7bfef3326ea0caed69d79a7c7d17cff93541d48ac3df5861fbccff68455ab128fc311737f930e39e336241214a814a975a6fc5d785eb7f221f5fb130b541fb62695310f6377bb0ff29d0b833bb5da9bc05fb7c3bcaad082a1fc78ff171c75373dfe457fe633ea522ef3e1441aefb253e1763e76d00705d5881afcd02f352b579d3fd7f87b9d9826928303d8a2b74745de79b7d8a90ad70e2e9dd09b02c4f1cf26e7ee0af0e500831c8e3f621cccbd014f9f2993e84f8d7b41de90de1a06d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he518f782f59a0185978d7fab437650fb81f20c705c076184dfead2f069e0d7d705077d2d80658dcfeb8ed9676914319b17e2b6156c0bb32930a4726dcd49fb914b7c8e6f2980aee0ea08b41fde9e3f1451254f63292120aa6d392d516bf25f2f3407511c97d454fa2beb1abc590bcb2a5c6881afa660e37a822384ecfb465a79ea0278982ef9595de24ada46483c17e57f4b17f6c75f2c0f09e7bf1f6a69b7445f83c35aeb26554ab9dc79cfd25cc3bde1fcc232eb9745cd94388d6da4f22eacaf626cd49bee149b1eb8a02c48233f97cee8ae2925ebbe7016a5e8a666d44ad7c846863e1f6d8f428f3b1cacfb0a7ed803b3741a02170ad99df0a0a06d5cdda15b4d64c4bc6f49dcf334c68c9adfa60973855e635119ee0ce4a1644b9b07fe1094bf229403f4fbb7f26640a420f4e9b5831ca190f8e09bcfe9582b4e3ab7a56352a99c294f363a1461097906890c735b65b01907c99f65065670d754f9ae7c6402a5c38c214dbdffb69eedbe14c52804db8a8137e221dec5fa5a6198aaf18432defc3a66f286b24b884cefc59b2051ab51c5bf154075b95552a1b42b838cd685d00d661ce92ad64bfd40a9cec7412520c31b5e5fe0f27ff6d47a5ef37507b64afbf24b5b471fb2d9a6c74fc451b7bcbd0575fe48eebfb7dd10b9a793b03e0f49acb1ee9a6414b844388a3a9f05328f526df5bbf1496b372db9fc413572458c65;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6bfa09207468d6865ae46b43c33a6b8554ff72860c0884f34939ca8c5ffc3d401f36d52026ea31193c15d77965ab35b4726089517c29877aabc22e2367359b815be180e943443cbb9e18c404f81ad5f99cdd1fb76626dcafc6db9ad0f005271a3d5d14d1b917b1968c22c42d857ab9d1b6f0cc5e96a60019c23d707f02be2009c7e41e0240d6fa5b2a5411f3fd2a80eab7973f002235eed0f2af40ea970b2709be554c0ee717c5090b4fe60b1bdb913764c99ea9d7ae135a0599dae6e2f9367d885e70094a61ab7f5650845dbdaf44f1d8cb20db75da1895cccff1b68f5b3de57ae207f39b98be3d509412e66b27b6a7c3cb37e3bcd23209318c3ce2fd01a7305862a266ea97c4785091c9a3dcc2cd58fecd908bd6c3861654a81681b4b748e68b3997dad7328476d1fe58fefe23db7c7aab11c40efd6daf3a3b8b5303fddf372255eb89ee472e32ca7fb4f0ead5033aff49f5d5291adda57e7fef36b53b4916dfb98ed1fcc4308b9ffae194b0e9371f50517d1c9fc64fd1fcd8a09413c12a36130ff2dcc8708312b62a5e77c9cafed4d1d9e5e972dd2d2adec66590d31c9c58dd6c85f306c7659cdf921902c22d6ba8f22435507c74a3d2e804ab825f78a8b99d9379f0252088b3dd31538551ca2eedd26a0d3908e841cb89b48064b061b973aa65f52e80f38a1460c52ca827203a8e0ff298cfe601ad50e5a9f0de742c2ad5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h39bd4e0072e4ecdd13e7b6cee4f77294b50a55d47c72029459bd34a41f6c2ee763d2bf3730113a311e4966a238e56a35c4b4725da446f082eadd4256b25cbe841f5725d23f136f07df944b7e980561e879bd29f9bb27cd6cb836b0fc5446894c1d20484eb7c88861ca799a62c74483f708b068f5b2a0a6ebade8c498a41bfca409fe86b69636904bb5e9983b3a0a12f93ca3a8150a81b392c534de8fea277f95b433023b392ac511da816d7dff007b77d80789c52d0e8d3d768cc856c976070a96734c45290188720f10f7e1054beb6d3f9738ba4a883aae73152eaf92b97c7257aec414e064a278bfb3a9d435a5b7970772af2100d4fc8a8a48e28d50cbdcd8a05408bdcabe8d3c8f4d4cf3d721c55246f2373709d1e807e63487bf0572dedc9db1946f0c7550e500d4604d95e90dc5ca7d3bff8a024b9227898a707c5c9bf03dd8db7d05c98b5c13ef0e5d18b653bbefed105c1128478f05c7d950fdb587b3063920f2e07ab93757d1acd9558cf6cb8acec1c1a12d991ca423f2830a4deccf0e71b3367a02c163a821fd10f29944daf122a525f52d01b35a4fb9ad72df62cbf4f4f0841d35c05c9f3c88ad74339e6c74b18b8512a5216207a398cb4cf9d1b970045328e1a7a1cd41e2c46089a7da728bbd4669199469178c5ad01ae675d75c75e4e3a6b42eacec02db2b16de9a06895fe21c2c9047305c07bd494b23d2569;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he85d5c31cd9e5c91d4be3d203c18a150ce3cb298e76fd40f47d22b16b2cc1f821078c6a5835e43e7b7e372e32910b8ea47bb445a3552bbfd90688cdc78754d3766b99f4967940010720c804f1349a7d3f87a4a4331753c871e42f26cfd4bd8791610e81b6bed0bca520e8478d59288735200f86a0fd792914b0cf6e96ddca0ab65db262b080256fd5122e604d4d052818e47db7aade464a510251785ca56a18ff5ab23418c129a8279c6f7de868ae2dd6d4b29de11dcdbcc3236dc90e37eead2c5413da6b339729eceef8a7abc27c68ad7cd9553593b40ad996fbc349f5c6e67fd9c06bc22def535023b598d918cdbe566922f67907af551c6118cc87c58e28e1d61f50676e27a74d4b84dfe6063ef26fc36e94dca96e91d3fbef064b71fe926c567f9fceca35597dd344b7c30b9720cd59f6f5de739fe7bf9de83c4a3d2ad884bbecee4334ce7709371741a0b9fd9ac0aa24ba332ec7433c0573c6551b186399e1ac8bf37762e97b1bf96ab6ba1a9e271438af0d93bc5a5a42649a931608110e321937197ef1cd981faedec801cccd9ac2a5669373a60ce621aeddc69db0170baa2b321568edf29c358cd8bf37f9e771d004b727e7947aefca276d2f5468666eda706005103bc87f92afbf614c804472c66baae4eff7ffb3b05eb00f14e3f2e6006b66dfb4f52e0b9b9b69ee061583e583343f60afe8ada39a37511f437e46e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h14b7ad52d48810c50d589356821398d8fa868d4d84997ae47f6d43f51fe4f4ba4eca4375363a68fee63e0676331c37acff0bd02f5d5f5d57bea19b9d0c7b2348966c5c1bd26e37c3532ea240d7bf73f2c941b6899c79159a4d7b54541be951d21997a2cea269581439b436fb696db20d16aed491cd180de7d07a170de9dbeb2c122e777a29345b95d3a0e930f047751c7fe56938b1e909f12cbf75a40738918bc6d40eb59d76284af92b096712468cc7612ca4c2350ac37ca3db43e4c14257883df1fbda27923a5eed175d72d6055380db9d1082d4209509d2c0b48bd94d4730da72725d2cf8024234a6dcde351ca345e54650fe1f04ec2db0def40b7edbb93e0e4c30533e4c7aeaa99d4093694866ec11ab2d30ac5ee76ef17d7bc46a6a71d2ed7e58f36c4dd287f281203752fac95b2ad419efbf2bdbd91ffe3696de551ff0ad09fa744d1972a19e4a1efbad26824cbcf3bdd382c5e3566dc29b970405be7dea2953c6a8eeb35cc652cec50661b4007fe57dd62f9e2f2c6e45a314a67ec5955230507369507d5dc903735eaa130e7c5f0b72d970fdb137927643d0b63cc9adf571b66b1b02765dd75fadba8533d37aa38c9c66b2a7275bf5e240efabe30dd565dced0a0d92ac97226af3408628561c752d3393efdfc50d4cef45bb298594284f2d9336bf9474d8188951cdf1cbf747f1fe8a4a7807fd88ebb4e5643d36a4ae;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6fd35acb6ba1f2802bd133f0a627e7f5ea7c430775f47edaba11d565f961effbcc3be7955c553153fb50f910c10ee114561c0739055e115662886aa486f3024c6937aa45d7dd26cab79153196d6e40855a40dd4e1bc5e9e5480419be24d51438ec0890fe50fbe5e2ae8340a32bce127d6ad2e96e73452e765ab18db43f8019747c045d20016ea078793a7f3c692f11b280f57db3d5e980029184fe584d8b5c35c27d5217ef60404577aa2e28c25961913d596580e9e3951e73cfb325ac6cb4b3a8df14fdcf2f6005e082e9986b5a0174c1dce51ce601a359f2373f750824acd26a45650dec92141c97b71a48b65744338b947ae82d9ae636bc60fe8c3f8aac6d9658f3151d290c2e3b94bb8735130028665d7ec01bf2f82a5edef6c2c9de9d2dca5fd65c89b28128952992aad3155e4ad1069fae50939eaaa1329dbcb8c9c0720ed1979c76647efe8805f651059c5d725f94eff9e8394260a5f25757538eea244ea597fd6190db622350ff772ff08043662cd04e56b54c46696674541ebf93ad99b4d8c9582eb6120648f4fc4201dbe50579cd760238c4a85d5f5dda96c45a32b942013c8394247c95fb102c7af2a8d27ffb2effe510ea8d68500c53d77739c013f14dba8ce0e32d8768ab7e39a46151c21218657f023679d4b03c7a1d1e260804b8d88f883011bda29ab7b2131a81825f71c669f98e78cf47f2813556492271;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h814e6c2666e673e6f4e872241e2d97a71cd39f19dd25c172bc90c90cabb6ae5b9a0f2c573f66d3ace2ebf5dff4270d97ba7f50b9a7d91c700c5ab1e94c3f445482dfbd407ebd539668cf45df593116106b19f3d266dd812a0c9c08674ee5aff797aedba41f2fc1cbb6398444d9ab942858b5aa6ea4603e84db9ec278ecdb84e456f3892360984fc5cdd4d5e78de473b9702518cda1450eb6c671c25a8ceebaa8bbb841c3a4415b73518b86d782b546ac3c7295252fa75b52ef43b8e65ac2af659231e67cfb35b5bda7d78159912d63f1d1ed2917a07764dd1774ed27f3e094a3529ac9225f8c65718c2a15735c1adda81f0a04f131ee1ad6ae71b09982c9f8fc42500bea29fbfd14063619574d9725042a6fe15f0c1db6287d0d3dd3147b0d0baa242f4a359d5df89d43f0b73437701e49b4704ba7ec5fb20c38925461c91a031ed49b6d464c88d46ee7152e84ee6e9da0f5e99de84dd613f758e236ad1e279bf8c29e4c643310dd48452ee875dfc33cfb23d34b07d35fdeef5d733f551cf172e2658d6996e22c6444f19aa2de774dd7e71405b5e688592a4a8e2e8a4562a1ae404a3fe6266421f5cd166e3256d4a8404616caadf84f4138f3c6d4638d792186decf715ddb5ea53815f492777d029b10c9315537be329c848e347a60ed8f623a6d531080e786642e16d9141cedb6283a1e64bcce28ac0322c8e295c94e6dd110;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd2f628ddd912b4cefa843b758cf979558c35692321c14da5c41f5bb9de54a6e2924dd7319ee04334bbae7816c3cfcbba250f55ff56a0e6a9e4fb2a48532b58e676d8991e9a38d20d8bc89a9668dc245279e751eca8be489826ffeb94bda33994facab251d2873b912d2145a00382d488340f0d65e2f7f357d445f5248394626cac6e80e1faf63ea9509ad0ac0e174bb200d82f388a419624932a147ce14dd889bb3f64dc408d402c20e95c556b7191fa4011dcfe982c5c4f972a594e5b3f27a97daadf515265501485d8b92a1a4b88159e86887e59d39a94b7c0e9b8f4fd550ecce3da85e3a36fec07b9097866eb42095f850410caa7eebfa53016329fe97a580ed6ed28c6cfceefc8196e796c13d671b68ce6e8e305d8144349c2bfc4554ea319fb6497457eaadc6fc0c400aead4e9e4dde83059087b14eb7ebb66efbf278e7a24373c31f304ecb0c13b18198911600f45d4bd3908d6392c1d1389630608dcce6dae692da5c9719ab6026c89c7b53f2b4e6d8a3c27c05a432bd8c786b454c6b9a69c0920196b5b91008f08746249a9997a681711004f7dcc9059ec086c0c4eb9211a6ec482c29d30c77748d699d7d3b0a826b353cba4821aa8553ebf82ee9e8a856b9abf3c30c06c163e35b59ae5363f339fa4693fc68e6b2f495216dd0ad5ae7726da78f9b9838c28657ef84d9e09138e3ab6038ef828dc9966103bb3e4999;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h373e6c55f7cd8b582fb7b0551f7c524e379c9fbae72f70629a8383a160babdb119e7a795e87c47f3e561f485094e3c1cafd012a72f837716619c8a998da05daf58ec986229b4efbe678efbe3625a32085fb7ff4a7425baa15adb84835733246c2181585e2ac563b9c9b7f72f6f2fb21aec3a4e8c776a02e327a455697a92db3ed694e70dffa088a5afc03ee9df5bc3464ad8d2bf50a99365ea8e0d139e78200fdcb03ab3a38b49037b77ea7593d56e5105962c62e70a7d010729f3af364e3eed22e0f78b444b9bdd2d823b11754f6e237a796f860810b8e625ce21b0f45ecea32679d34e4110450354bfa6ca0dff6bd0faf031dd975f33bd6cc16f9b4e5d18278284925191d08d7b98f438d359f66741768c4e9b107180d272b7718f32440b6cd0b8666d4c502898e815f6deedc4be2ba45b691ed394bf1b7527c1734d676af6f236ff490f008baa0b2c02a5660fcaa949cd6cf4c0584faf50ddc56543b36ce662ec9cc96bc3c858352eec67d8217a84a336e27aafe259519d1e3a13b8affb64cd7c6e7374d087e7f98a77ccf73ea39ad1b70e1e8c8655f3d73c879cd8c5f971a5ca551e566327e32ea7f0f9846d2f86bea58b061b28d41f15cf6b3db2514f515d12ec1287dc3ee03122d6cd6e7df70710626acb354a97a7c7effdc8a82d1b8f9aa9f1e43e81780d3ff9e3d6ffad508aef57c96f39add75d689e3878fe2f468d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5856e02a2bddcc04450d941574c1ffa3d02fce71a922c7e5caea5ef0d12a26541b844769c7d35a87a50e671f21637b965e3bc50ad916f4cd1775b9a12021fb98e760303f6a48972cc5975d39561c21fef1e19e1417441f47c04fb3cd5c5e1ac77060973d0dca40006f5338b69d8b58bf505463312e6e60bed9c733c37d75f92132eb7d2b228dd2b6a6ce8fedd6fdd431b728ec5a4f647270b7d32fbf209466e8e58d5d650b835cd138179005ef4ac86bbde1bb1016755a9769d218c6ccb7e58a650d8666fc5c4a8fe6416d11d3ee292b825e2a5c809842bc4bdc7eef09acc49a31982dacdbc8d599cf7429d515f89073eb7efd2f8b7de8e7401edf137f07afc72324ba5f274220c71943baa5e2195ee2b088fa547b6709cc9b4737389107a17d783ca12e607eb84eab9b891a5b15ec87504322be9cc592189544440697432534e681c131c7e255d880cd3a49819299e935c826bca69434a3ed5728b6fd8d857ae9f3b9f8ea7d76b74a17c5b7f596e649dc3251cfed0e8a6948358bf24f562c554dd685663dfa9bdec4f5b61081c1ddd316919becef621c50b393ecc475d24e42851aa944e0bc28012feef57a6441569da3b8662cb55d8218a7a30302f3d6972d386043f594fa713d50efc7c8e489ded2eb7778d5596434b4124e3889be70ea0e5c630481c71925bed8788a5633de3d91f13fca7ac40aea1f8bb2d4eb58d55466;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb915b53e187257eee57417dab14974fac10c6f177cdd2307a91120bc8a26d0c9de4feadb5eba1ae839b33eb25e6bce7d1a3eda2e5a0f1958edb3c648a3292fba3e5e45763faef813832aa30d5fa3f762f3946a1313d47e896528c79d4f76b11e5803458022ce97ab5e23cab4976e358a8e9d5c856a0ebc876b75f54aa34a3ff823f030277db14c6362ab6915846acab8531f3b9a932123fd2d19b741066455da73acc55846c92f14abd8a5ebf367919c87b1d865511e22ec3851d6cfb20da767de1a4c50bd21b1b8e7d742b74eb9c9c9bef7d6c7f19d2294cafae51055aa8c3457273080755a0d6773dd1bd3de3d496767f07b85b47ebb1e64ab98abd588ac00a6d686559d25b4367ccf4e2d7d508f4a45f3a395230fddf758cfde53d5118225e58e5a159b111e2de0763237ccedec7e04a6de26e7ef991aefd392b82cd0301c92ef76dfa8add8bfe03c7154141cfb0a9c43596ca33d26f4c7611bca1b10a3ebd32a45f392d269cab604a03380edab042b0c602dab46bc1e53e817f3d031d96cebc2572d6c869c5f053e959d8c7abba86a20248f79ab91a2ba4468a31b8dae985e61f658927cff8afcc3623c2a32abb42f9700334972ad2cc68bfd4a30bc1551be0131ae769da44dcb8538913b519690492d94a65f47beabe252988af9575b2038d1680ded051cd2d2cdaeaacbf2ebcad0f51dcc0d60e8812400f52a0e15f691;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd1e506202ca6e5290128e985fa56825a887c60c98f2743f8ef3183b7e5e0937791d51d57b1f81831530d2063886a4855a8ab6c3978df5070ef603c5fa5f5887f8a92fb3f2a880b9cad9dc0a6cfe7012f0a97bf1f7ca1c3730adecb87223bffaaeaff4a5da0cccb06a799a445cd031950cad4789469988bd04e33e41b41a597222df5bde88224c669a0426db3d798febfa440d61e6b92589dd6f59acef3ab1fb455716e7dac3ee8e40f25c751af7c0afc52fdaf0b11b55ee896b5db466cf0f9ad8058cb9691c79851e00f7f52b2b7f3c05ac38295e138ddee9620ae8a1f6a9c109bdb2a080b1c4ebc9661e448a980f89f2c3f1cee84933ddccad5961cb5bf96ecd9877f27d20da5e9bd25c3967f7fdf87633c3223ca9b6c3216d9f727f3a6bb969d4666be960e053ffda28788340e340e79e61adef79b9a05272e3703169677060d919090dc1a6782c482f4bf38771e7b9bbacfde7a98108be3f2082005c6803abe74fc96d2c099a69a0c2ed02fde87446fe28804c88d3c3c07acaf59035dcb5fc5eadbb279a0779e988804ebf3a13cd5cae0a2e799d7576795d0bf54f670b1b3c23999da60abdacf8eed4dd00f304689c63b95179a2b768a78b885c4a6cbd5c23a525b1951d3acf07afdc31300246e60c2ff7af2f4e7bda22807c0e7cb4721b88291c70c4fb6284e3f108e96b505346be43f47d0f54b8f09abc1565819d56a3f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2b5b7a441f9390a0d9218a018037965884b40f72b61dab7c35bd648a6b453376543b8c69f20710b4ac7c0c2ca71759431ec8882bee0f25cb4261f0ff8d33af4bc6c2e38e168d2cb836b2bc25ec2606e5c7a490e81b8998d8e45d8dd9448d373b484f09db956b1a4a6afcf6b5faadd9d646c6575b76d378d94970f3549f7b345d0911738949404d27501f7ed8a1ee02ee275ab5483154a8ef1820a7ef5649b7ad91ade5883bd7c58d3f0a77af954fa7b2bac0795809fb318427c4d06bd1e3bcfea69df73aad60275bfbbd6c2ab4579aaefc20e683b9a62bb3fac96ba92f4c3b842b80b7dbb5e6a69c911e99931b044ae166f8e59435b141f75c95a4e7d4c073495f95236300efdcbec21d10e7d715f184d6dc76d926b3728cf8f079f29faac37d7ead547738fda1e5afeff09bc92ed013a6a9a627c69c9bfc80c1c758b3140dd715043c1c697a0bd950b600df1f7b200726004ae328d2bceb52a6ca6e38bf61ad20c766875c1e866986e387db998e17bce97f87a5a1e362d34f67593dba2cd2937ed88d6967d351974cd4c3c30be856c89327c2173b782dd58558481be5c51b003f08f34087860def68a4047394179111c5c9775cc446ac31fa081af81775554106eed4ba8fafb50a153de5391af609157bb082d9ca654621d3e3ae113a951efb2532f5b82e16f1f4af1950d919b60544d8a3707385e5fdd63a9e097b26b37ccf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h761cf6e63cea112eb70eb6f2e1cae9077d01a6100ce3b41ae486b9943f1ae7135682a0830c0a8c1f6df6e7558c6961d80804225aa3adbb094562dfb33935bb08090c8bc686ed523175aef0f9f9e008cb5c2e7a776475e98712c6493898c38838d1c059ecadaf795f78adf793638d56543628b32a701800451ebf030bf85dd697421df30a57db107743ca7e0c703d4a34e1b622c8e7f4d29a242937e39dc12baa315c5892df62d64a8918ec4c95d98f691167bfdd390ce861779cb4c9925769af0fb237387afa8cfa6d84b2e753c5360c4e0b879bb4bfc06bf22dfeac7a826ba09a7518fe1d86f2fb6159e3c0bcd33b77721d2d2cc9261b92ac96d24f75e46a41ca36cfb190ba86110149920f31f2b0d90584a73740fa389a144cd722c9e3ea7a4756ee9dd4cb461ad406bff7710ec60185ed67a0a59d9c7dd2e3a2f81ade77e96fe7da2f46df4919f2cca75144732d930b186075571fdd465883ab0aa58f3366c80928c860563c44ab35bd4a6b80c1ee1f7827eae1e30886fd49574a2438c7154b9a1e1c889b23643bcb44d26f8f76a33700dad31a8f091b5d91f04f456ade2cf00eeb3b101be52e4c091b360c4442331613fbb804b77324d58faeeb1b8472c9f2b74b4edbe2fa9ee60dab28e4c9fd5f48d7427360755d194a98b3962d9973e2f04fa50c6432906eed4c8c74224b2fd47a3225f8b12bc4f47306d88e47f47bb2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3ecdc338d51e8e0b2a8575b258812ced8f4226c3956554e06debe44960f9ab899b112184582f1606143beaf61a7fa865ccbc5953cb5308615711e27f2e0ed3cc275a8a21abbe9164e18e85c8d32032d1c320375dfc9ba61de4cc0c064bb07cac2fe027420b8dccb2e8a05dd74171c244a9d92eb076f48649dd173ec758aea40a81c65421e3610b2fc7566a90128f66e145a08253efa60d229f2694a202a174edba36ed69f33c34845a5ff463e7c6dcdfc14e527e24619e59f748e73093a4cc6fa2829fb833be00564664b22a36eaec1bd110d0194e5191c3b95829c080aebf6f8dc35111c291bfe9acf880784dfd8f3d5e800472bd5df25bf9f84e5c0d33ec4b78e6c7dbcb0cc2f4e19c367583614c3b528d973ba8ecf0f6913ac7e9b0560495baadd8fd83ddbe2897a7bc9ec1d3a3e61f56a03154f1769d1528ea2a70ed16df3956f0f9925d62e53d919c9a91303bc795861ff42da28a9e18764c387585aec42bd9f92e078ea797827bd039b1f1b9714e599e8299a6eb02e2916d99adc01b06f82ecad7d627bc518cfe1e4eb74546995b0bc4e62619e5aee922238bff829b483c9c0b5d4fa27d8283758855f16c641db03fcc31d3586a1b106dc06bf60195eb639b90253c439951d1138e99919abda5a440755cfd14f12a2a9c3f010ca3b425d34e7bcb931302a069c2262661e0c1c5911b9a556bab78763248428dc44fa511;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb3d9918317ab57539456244568b7f730903e10f035ba24ed8d08a455f2801f17edacb665865d2a402acf049b098b7173b683c81428fe9b98822a09b54e261abd8cc397dce70bbb1a1d3653828fd56df5b669b08a4a9ac95e13e5f930d24efe5617d082858eeb0ddd38c9e633866752a06c5c5b09faac9fcf635d95de693f187e8006398bda2f2344f52d6ad68c92b584d4f94d6230f3e01c27cc61d6c50f628bd168ea41fee7602e87a4ffe56f18b37ab267efa0240a3b7c0b083a430b03398977ac0d68a92c475c3d613fe099635ef97cee065419dd6c967b7a524fc5b7144ac78de7b129a0745fb002b0c991de130c05799048a039ad684dde686bf26df9bf89c0c3e3ff6e347270419c8bbf2d3fb66cba9912b28bc336419c5a68255e04f5e4147f6af18d651182d26af42bc4b505174b1f661359ec74380ae294733e4ed8cfe0b18376d1037a3c94f5cec062ee0e0bfe924bf7a990adb1dcf049c427ba1fa28b1adbe50009f510c60c2fea8bd823463068966bb7eaae3c566b21fbf4d1f533eb2fb3d4be3bf157efc4ee9bc45ff30b60e697aaa56140aa94606e5821f74a83586ff810f8c7675ba43533f220b66476367c124502baefe58a8c1bc97e586c04d770f6ea8114ac4af1b8afa966991ec628d5d4ae904a165d258e0a26ff5fe365a2889b5972e9e5bcf36cc02c344f00b2859c9e6958ccb9741eafb9ff53592a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3aed0339b7b968071a82d8d3d72b86e133f20b32522d6a1a2049483e7e16594a2b233b851ae19412169ab1b94dcf41a430160231031174d36c98a7dce5768e943fed7f34e0328c49efcfb9a00b462f781ef53fc52c754cf99ecea54baab3eb439a07af1e5c65723cfc26e01b18d13652941b23f6afeb9b180878c47911639be368e23e95cc0aa3b3907e38a6c42761ce49d944400834fbb1fe9accda12ba50e5d04c2d8d62ccd44b2a9cc7419cf51e449427d22a92e9da81a676a62e8b893214b05b361250183f1b8fd31aa4433fb33eeaeb9f59cf5ecf17d9594c15240299b84776e00c6e0ca1165880b442875ab8f2840dd21a5d54fdf8d23fd8d5d57b389df2469b92992954511425fa225507168c9cc9034c8b31a0f46cfcb2d48e2b70fa707e76cb14fc8244753e8ef6a41498d7f2e2135cccd17135a8fc63ceaf34f04ad850160139d8842f1e05af35110c884844fb8aa3550bfb06258cca933eba706ab639afd76570d287947954ce92205d85ab33eaf2eed5ac287674f71db2aae9e48db2503e2aab22d9df30455590103835bfcdce0e10b9f647ad60b391ea072c70dc268e436e08ce45e43cbb6284c90acfad6580a72e564b414f48fc20ac578f06d00aa0cfc1b833cb6b4c0c963cf23a77c1132d0f37ae92183b14bf2e480ef05bf97fa3fa2f0430367bf0267dfcc1adf64088ae7df51c6348f34ff447c65eaa4a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2c87a7f20c3ad06cfc799fc466d152e06be9fd992e4cbe5381505ee696c61e851f7e9e14954075855a187d5e773f465c278fcef2b177d1c9f24e201bc14bbf9a73a3b9601e8b62d3656e108a94e74894434ca3eb09406d9e571d29c3a79323c28ff6212378459ae4f69e6eedc5438c7729ef19b6df3d674180f729a5356d5b30dbbf1562b25589e6b204997098d35a9d61216c90d18e22a266db55326a3253b68efc31efbc30957bc900c6fe045f48bec9c0992423d4633ae6cb251340480e298ed407ffd7e885f8587b80ff818abaf9d42a33d203bdb2657944ebb1a74666c51da9cf561f8c6bb32b1cf3bc08bfa66e5569f8ab6501a69129caf48913c1c9da28578648949db0a5d65f967b4d48ff8b894e98aeec43d56b5125c73da15bc56e256e2757764e9763e6c6fd5f789a350b6065e6dff1ac7a13b6aae00e2453a62b4c1c8fab1b101d1f4ef5a905f5c780cdfaa90a7f6819427ac7d93a580dd16ed7aac3d3ea85442703e6be13cd853efec78d2ea2fe73d76f8b85f5cbfc832e320f9da640f1f11ea07e37c3079a2bef2f88fb126026d383f5cb487b5145a2509dbc9bc99a05d4117b996f645f88064c5a22f68728c1cc2eec51fb6a44afbf9b90626fd3e49e57acbd310090a21b571b9facf8cd5e9b1d9469e88ca2f5103a6f84d79899825b6bb9f54896c0805cc7ab85bbe4ac1b0f9d7c1c632a38192f176312d0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc60836a14c0de36ad0dae11d3c6e1e41114046ddfe772d10deb6dcd8ac5f9560c0636e197f8b1b0d242d5f1d57c774fa276bbe05b5cdf865d1248cb2d35c403b8c8601203a60fcd46cb5f37c6ad8877c4cd1daa6be988d7aae62730e502da8a1d5d241c6c0b2582fa8c7ac0b721baab3e2b35056c2c509ef490f989d4ba109e8dbd465405015aba079fd3b2070e94e9b3dd0cb5ad6bfa09a44b6d98666f883316c730617fbac7867e6f0494ba061be086113bf91e346d865747efabc5e861410d047b13967a2cdd94dd289ca0ef5f51e63f892ba3f80e71ef9f35a3929a5ee04d80d0142477d24004886a2d4123e88ede909a9609b1f32cbeee59c86d8b27a08076a41eabf0a421064349593c9f84c73dbd9348e91447d9ae4ac5e8a9806b6ca76c3d4d53b646e780205100a87d58f83300dde0f61c505c2f78d086f0d2cf2b5d653c7c05cbfe2bf1710b12556fafc93dc6fd89269b6b293efdf705d4bb8f2956700f211474aa7e6abdb10eeb18ac9b5c7ee6b15cff067fa14d33daf624fc60c04e5cfab1e191aba2d6ae952c13ade8619e9da965019d224bb272d5effef3ff51fb16c6a4f1039f3d9fa7df64c563f585c39330eb76b76512c870d780e81db242c0f2510f38048cdfc6cc35eecfc68c0559af6da93d33c3a2a685778855d195c89e0b3d3d78e0e81335bc6c909296d6e5a62af96bb3abbbae6ee7cd793bdb4ab;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5b0ec9a5fe4543eded7fdf3c47b60ff8447e2da394dcd5dc282ef8272ac32080ce1a3f6115f1e53cf5642a022584332f697c73613c954dd0ba5437524e9e3bb563d63d800df2ede39319f9ee51ee855db3360062889a78dc7d2a036931142b39f8c7527026aa9534f5bfac11546c76da361b2c33a0c4fe27bab69f40803c0f0175437f18b29a95c4fc0d85e201bf07918ad44e26cf9c46bd63e7a1a5305e78ebb738af344d753e60b3e051b076058b089faa87506e42391ac7528cfaacf3a03a64fe831719593765143647cbc120f10bc1c7c2067dd072ab1e9a3050363188c240413c284e0db0e01346050931273e7370bd636f737846270e4e1f76cd49a97d5097c0b0e7f28a7e542599bf39946d221bf63172458e478f546811511b5a3048511cce5572f1645d5eb387a7e3df1153b90d793cce6cffb2631fe51766a1eb55cd969e87083519cbe7ddc4d94418eac68ce075b6890897093f48613d7a383d4a3cdfb71a12a088dbb308999d351e373654d122d03484a82534c7f58426423348d2541fc2af8d5197c987aabab55ffa9e8140c18bf5e48b534a70c40f9759935ac5b6367d05be6bfb7184daee8a1beba20782f32c47157442e4e096ae02bb4c4895811b26f3c7b282c88a58589ae0c71c93aa8512d847412590cd472e723479ec5ac38373f9c31109bccd34441567d8975e3e91e2c265ae1cc71d610d2844e1ac;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h913a66a913c59eab4cc8c0cdb0e959c864443708d58583daba1e21047ad1c1b3ea4415204771a5eb14056b6f43da80a137a3d340ef95994c63bc18a703c97ce58c1e29034ec5135667042d5100f6da27474df0e9381a6e4998cb65f2351276944fee2130b993c1210f989d4e0e67d972b23acafc3f1e2fcf1b721c8d554569c40131fd6bb0002f90e613d271f4812b23942453f2c1b511e7a9b62952a921d40c36576e1c6fc7a97e56e47a635cea20425eb3e8eb377dda028ce0af8e963784f6eabb5ae78aba14e18ab8a604d4321c2e74f7dd6ce41ee0bb93b00f6b36a066e8bedda8e4abcc0d059491f73bf3427b0a8cb376a635b0eeb53bf981f0ee3407cdedfb467ab11db502e0aa36277d1b0c5810bdbf869013bc3b4c5d999f6b734fd32d79fa7b2e01283ee3a155a3856dd7168d442b36465df97fded7259492db6c90ace8794e2f0ae2848991be4af6852b22d54a9209304fe637d6b30da0a6ad564d9ca39a1645c536e03a4a726904522a6192cd7f3c12cd9feb3a4dc8705e18feca3313f1eb94e1ac9074103de472520216900989f48fa9f6f50cb2ea06d1dd875aa0d012103c35048b2552724bdf98779716dff9e0fef52c195c18d144dafb3c36fdda70bc7ec9c887e34b762a3d011bd7168e3780c80e49edb693f2560bb003e023edc0292a60380a8f42227a89a4bda37d2de2258f4f933dead9684702119364;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5279bbf692e04356809319c17d4177e878d32b1bf86f42b805ce8cd1b9b21b312d34b2e58113306c2b7696b2a5a14540e3746e506407fd5a259c1a930ef8b34ff0a51b22069de4390865a693e1990fc2b624dac2935105a5e7241bc62b603f23c3c5590f89e861a7791a333f6eb681a333d6a376f5a0a59249c696e2db28b721e1fbbb2b51dee1545b20c3581b94506185b0c67d124bd5f5754882b0e1fbf96be8ebc85f66242f61187cb1aac679716883d98cc79cb09c3e08f36b7631bc92423bfd23907d27001a2eaeb70dbe01fcbf54066616a60eada0b9cb905f4c371c870a7d611c0d1d8ce176e1b1901fb06d0b9954127aaf1c7fad464fa9667cf330a77b0f21b8eba9a458fa33144067fc6ff4f2e211039dff1aa0afa022cfe2be823a56a1e70f84327cf6fdd495c5d6befb9fdc7cca2c00ab9b49fabe2f8a64b91639aea812272e730533337bb843b843e66aabeebc328ddc0635bf691f7372e77ebe9baa166aab368e6e2fad2c04716a6f1ba76d087d89d84514b43883d0c5340d1968b3c7ebca571e8c057ceb8b1ee47f8137d634da9dcfcbb9ade4316ea1540804ac7bec1a17933a31e7786159f0864802121be89f0c40736f94264bf497a2118fbbadf595cb7ecc805be7150c62e8529fe522cb1bbab2a0cd3ff0f417f7dcfd67d2c5b3b21f5facc558f397aaab8a052042d43ca12dba92a3b7e39bf67ecd5b84;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he2b206fadfb4de42995d3982dbb94053cbc65351fc4a58c373a4c1046076061ad95fc690a8e921811f7ac13f8cfdd35b0ff0344e48d08e466e1ff0fab2fbcc1a467158995921d3f645c0ab3a975c44d3c7f904df231df2ca220743698b7ac7ab615fd7b5806307c116f8ad2263ddef1963750cc0ca519c4ba4da5819370b92264136c545348d23e13903ae41a86210fc10b3d1151d37d395b090aef1378c8ce2e3ed840a622b02ded2acba3171aa08e655402a0f3c1b282b34ddb37b392f84e6d6772f9fd2ed31ce2db7a5f70711ebd3fe30c08e523cd561336fda33e1518fa0aff6e2e645735ad41d5982e07551fc5738317818a72582017abea70c0b9c3ab49042b3ed57371fd51b921ffa3a92532783c8ea078b05b0bac7b3cc5f3a5a8deadce496abeaf32ab06cd6be5f89100a9ed47e279187e0f25e73d6cf547209f43075c5fa8dd278593dd51ff80d9e924fffcfe207976c36c27fa789de5c9486077c65911a2993953c108b487735b5021599cdc92810800535d6aaf8d8eaafd5b0aca3faea2c822087d0ee3b93b5443c30c70cf5d51aeccc14413ffdc22867f7fa5eca6703ba61dcfb55cc70299e82ef172a599ad38e482012fb2ff79983d7ee81e389fc6bebe46c4a8bf79630e5ec06b1e33ec8fe1dd88dece36efcfea9bcf3dd116e2f76df0bbebf1d86c75160070531794a64e5667a8402a32235c945be26e32;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4f2d380b25bcd26ec4799d6f8eac029bade40f981ce24b79406d81aa8e75b06aa2c4d217adcee0db525f676e1f4cec6918e22c0c699ae9c854535238448977f8529b69ee65701bda8c3a778414cd254ac16837d9fbd05bf3528edec52437077fbdca8d09a860bf6ac705bcbbd72ebb962359ca827f763c1d30f23622efbc635c712e005b3f834beea2128768d519d97d03b16c6b35face5e43a9f4fcffa8cab85132ef65aafbdf5c96ec20c7122786aad6ca0009debb6db2d37858c31dc7a698534b96181284559e6a704281e72bde8539e9c32ad5b9ac6b529bb60e536ecda4e1e906547b954d14a6d09407d5e3bff77b393f22b0fa93c6062ca4ada246a60ab35d4fd0be4e68f64726c92e9a8caa55abf34509a438cfd87db18b5456f018778cb7aa596338262373ae8875905989f9169c3fff1c2edea853ae3daf8966614d589d10f2e8e3d1f32127c47a6dc24dcb0d990142324c69d79759d5defac0e0d1fbd397142fa16bcf96730fa6d7aae01a34b7694a543f66bdc4668f50afe53d94ea33625bf8acde81419a8ed7fe590b10e704a54e2716ad71c6486a74084000dd7e0650a591fe054ecde7da2488e023191feed4d70f83d4b63e9846e7d9f10d30e7a815f8fe5236bac056146859ae190e7735167758c1d6761785f0b1095f4b4a799147fe2fe9d69d0a39dab4e94341f08fecadc522ef16b308572a5382d21930;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h850e9ca1d639571166c7a313c1e3f1b312952864cd46725dd015d8f3bdc6cd66fc10c6fde37b483b8976a63a5008a475d786b01b0e5b8c2b2e835af9b0e896598ba342c89bf0e56630b60d4b3d21201d57bb9e1bb1b38e475a718bc25f502a616d2f2d28d15a125b3f62e52549f8f26b6dfad921722137994e035d4154f5d9aecd442d5e076665ab65627ed8b9e37062fd1a8781395e5cc63066b0c8fc3adea1ad2ab51046ba064e4fb843be9cfef84f5e051c9d60ffdb02f2b1d3ef8036368194e00cbfdf597e5d0fe7a6d82461bb767c757eeff9fb5ce633f899a737d0d09b9a69de1bb432385ff8ecd1d882b20ac77c9d206702cfa8f508a04d7adafbef6b4198378248321f9b8d9bc2eaef954448590ca55a927ac8e8583fb72987af1ac8a1650e0b0fb54cfc50d95d340256eb01c8a420d20f7ee139c25704f47fd6abd4c89a0e15ece88b47b965efdfe3f1ce371800647434919e92e4e20bac560c52e138be9ae423aae38162130d9d7fc909670fbb10494c958a48f8ef4a00a1e6da7e3de364dc8355ee6b26ca301c792dbc7ae14a2f938a76940e51c4df55fdf2a381806b5022465bb9db497fe522ce73ee13eaeb8523e58dbdcf3fb1957fa16167430e5dfd29ca77461f0eb94695ea7c9de5dedba7e477cd688d07f0ef9ba43356a1d34ddb271d73667e0758581e7a4a0a0e33f86fcaa48014a8ba49c4c4956298e1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1d788b61ce81ce143b2da3ee1b5c53360eb8e71ae74e71278856da9671d82048a421978795e1e2de44716044b48a960498de9c460d85fc738cd08f1ca34a5c1256cd549c44166edbfb52b20511156818b574e5a8d95f656ea692db8724677dd6e504d82acb79053a2e404d82e6d9d7b788bdc9b9071fca2947dbbc51040f3cf560e6d8185092c5db9cff19bbc8e50d5c9822c6b7e9fa47f99753e1cfad8c909c6f1199e43d1cacbbc3ed5ea02e3a628c8f0f49f0e6c0fb9d1af2a0e9c8f5f3fac5eb981c3a99960e88081a56733de7c768032bebcaa5b7c217188c992e202fba6259e51a0f1e36314f9b31728e3670a15d48de7b5e5bdc9d6629156b10f1ec0e9cca8093583bec751dae766024bb7da999f590c96f8bc165ee00e011fb6f5be84f3673fe9d42261675af4b193665b91d183ee62da150205280e712fda235af59fa03a91fb9d372af309a8d9f31a35f2f5e53b43663675e8def8905f0bee334e05d98a653c35ac4f0532564bfd18dc00c3644c88419efc46ab9fa0738296f7fc2c45190928ee57c64d3528c69f6ab3bc2b62375650f3c40a25647a67df0bf94eae71a7c90840690be61b67d94c79db474257daee476e5b91bd42c6c2346c177124b5f689d25508132d93639d50623dd847ed2eeed78e0f2cf371120cc789cede94b846ca9a6770c982366be52ac012b0b34a769c6bf517f87ebfdbf33f9124a03;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he53ae923e572caebcd1fd581ef7a2c538cbc5c6570ba732b2ef003fd34b893efa5fa32750d796f903ffb8caf0c1b090c4f935e4b5e67b9760d5f3b274aadaf19eaa235a9d2baa23dfe2741d46c007254675c9c542ba51921fc3089f6a96698912224daf5902693778d30a367e48e050ea31a2d2c052660b7816969e1e85d80bcf79e802dc92e453f2e737c4c677ced62727ecec68ddb076d9888e89d0d8005eb438e351ee6840a406af6200dfcdcad752e04e4043bb891b26b0bcbbdbe8ff6ce1e2474fda571c7de8f4646c8de3d174c96c87a4bb9087502aa65c2df3391395c17f8db5c60462dbcdfa3eaf1dafb82f4ee8ee432b8e79213aa2c7d3c20607812ab88056882af736ff96cea0f38e1421ddc9526c535ebbc537c8f41b0a6a29bae5d243d92c685b07912787ba1f4fefaf0fa42e9a6ba78006dcf2083538a9bca7aa44a7d01a20f709e7d877d6889ca1fbb4ac54ac9c29530f255a64160a5fcea66b4265f1c839aee014ebb2bde83d7c2d0e512029b0f4f40b860563630199d013aa6f89b231018d0cef6c162aebe1e886d8a9e077ebbba5e3076c0a87e0e169c4d6441d781e518187edcac733fb203a403d8638f1d0fd5e66c861bbda3bb5057cf3c4576fb995d990019e65ecea48da39d0eb28367a7142936a187258a70a373a689184646586970c8591966b6dee8d928f58e7e16be0c27c4b34904d87c483dc7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb5b0305e7f7f5b4347ebcd16a7db0ae2403dd33af0bf3c9004d8d6a9c96eefbd1a74ad159144f1b76b901857a06456cc652d62d17387a23a3125c9848089b3a6167a6e0dc60e15f7a13eb79d4d29c52d6b190d03221e0f7fcf48183566f03f1592a8e7559492126d0108b83e4a9c76e4e5f1433cc8961a96f088fb45be15a2ba6bcfbc5ccf2a8a8e86ea86fadec9e20b08396036bfb5c09c01a945b53c4791229c990780d213f965ba1a31a9b9e96d801ae117073484f41f541ad6be3fcf819ae269c33fdc160a30c3b920fef607b19f3d6543504febda0dd7cadbc18695af4c8bfd54b3b4ebce92090b1e305483d7aae476ec6ff831344596df840ed49b30c48817495e225513ce0164a2f5abe6d212a90b53c93df8a50991ce1891775d6a6b11f81dd02fef28a7a5b6b65302348df72cf780dba6d27abc8ae5556d9899420d07c93e893ac7ba37b39eb5bb4a5daa30431f71bd3acb990dd11bc69d6f0ad4d36a7ad7064c2e2cb0fef86ed533e594d947bc847c1451fdcad8b0255a6e93e0f99e953deb03ce1f5ead706c8156db36c3ddc73cefe9eef6fd0c2435b82c6c06f2eef14163f70586f1200d3344b87de54f4df0c73ef4c7f482518cbec4dc0289c98c565e696c452cc000c557b50956ed260ccea652251f160f103bc589c5042ca0bdeb81b20b0b418a94fa4f1582cc5b5b3fc62988b69f8fecc021949871fb954e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7fa6d76f60a13e419829f588b6475122a4c1eab2fed532d943d7a60f4423751c6b9c36e7eb254f1551dcf6d04c951f5760d4c493226ec8271e969fe0d55750ab92814e6b94bc74a9fe90c088cdde9f3b629334faf9d0070e4d4db49e2fb2cf17abf5e9fc275114fa695548009f80dc0431f496c53728c5a56e79774e17caa4dae5b0506b52885b75422969044d0c732b10c71f44ee07e6678ab271d72b15bd183cc140caf120beae69ea197a930fadf8103a18cff2e30848b7e5d7526ab3e9a3185b627f3ed0b896b062fa643571e9bda798b8625b5f69de8e1daee6149a991f2cb3696fcc61687907d01d82d5ffde788d1b2a0bba821f3c2ccf0b2f5f810cf57021feae6fd19a3ee4b07d3065703ab8f47786bf39648bf2826fb527e5b2de03d9a8ef399c68f6b2a00b4655b9af008d88d71e86dd21f98bbc16293b8418d178abb40a70b4f8b7f80f708787089b64eb54e87b9f846c7610034c1651caecd7d429660eb14dbb51a29249b6a1d479cf350d178931380ce79ece83f4275dca7658358b808fb0a0aad461c198d77d609d736f63f382aabd22355af7db4557b817d6fdb7be420695c3c5304605d12a0c54a6f3ea2f112e272737b1af3e3b43970f86646ea83466e54ca3b9ddec91ad87a80957c7e60e13b6ec570ea61bd48d4477e5980880fe069405eb362923a0ec3dc382997f04ccc09345cc29c2b000196ddb10;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hddcfd90faead4b864fb4e5a0af8d3a1e6aac54b97c86908ad6b39cade71cc0a3f820545d1b2eab3563fd5b668905c455db6e68733bc8faa8946bcdc286282f875807b51fbdabadbced1b8abf8b6f05ddc40bdf23559417c1bca51501732aef355f6fd81b5abcbbf28c934d3b2e7edccf553b037582e1f9588ee491a328b82b9bbbb9aed9b0a04985e496be15deb5e3557e0bd3473fbf9f516f40efb9ede6baa01b5d4f8a690797e16b13f342f1d91a1c207db8fe8a9d2ee5c865cc6a08d54f6f3a013968aee2129e47f44747291ade3467caec68892e755ed37520688ac5b8b620a286fd106f54e16d2544ab9bd5d4fce41d752794cccd7ed8378a2b1cdcdb9c6774e065f0d45d86f4a54d198669729bf8dd4a36b77fe8891d0d65ab4730656ec87b1d01f5a6e50ec2cc6060cf978043615e6db2b5811cf25c0a7c9d2706ade19aa3c2757160957eafb11b46956815995c35c92bdd3ef5b4448d85c7d60dd72767aa393abbebfb1276d49909e91838405df1fa42209c377ba967da07ea13f3af243363164393ea8aee1db8c8f535d93084919535dbcea81071aeec8cd9a03b0bfe925c4c3fc3b0454abfdaec0506553a46b9a13ac4b8d7b03e9526cf9599d01bb82904fec039507530a07b4816efc269783b25bc069180b147f0f02cb397b725f9469a2be801efc29475bcdefa094dda5f5d05e0778c195ec55b2c0a914b2455;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6d189e5b59bf766e8e7d2c510c9500eebcb728bb9166186d13235c64be6c48ddf2dc6d4022a72da442acf8e20874d5fd6f1235f43017424f372a34992df821d9713243636d2b9c58834d0cdc81d6e05818bbacd2cd9131d4ba4f1db9871b734a17949e19abf6586672f9571a19368f6f0af5e4a7b1a0ee55d08a0ba2508ee383038be3900112d086d74671be6afe940a0e43e2cceedf96f6491dda5c9338c1633c7e2088404ad54b900c2114554bda52e24826d5b145d6108bdbdf23774bc58e32bc411021a3f88aaa192628c1865defd9c77bc4c63913671264ea062c50f7bec8b6fcf94ba35502df810618327c9e234010e8ca8545a48bdf1476bd2b2d6e1358b2ab43b1d2cfd145bd26b7fecc0a241a9907c301814aabe5277bce5c19f9b82606f1b8918ee98a0f8d5b42705e2668fd8709560ca9ac408a45d7aec5c4d1556759c4055543733a6c821d15e22541718e8c1b785e2b9fa9c3f0a5b5978fc6b98b4e51a3c761f40f15c5e71b280ff517860d06c769441a3dc515176d15a4d7e782210dd86c1962137ca06b05360cd1a6d6255ef7c65650e740727ec9ac92df34eadb5696d1d6534407cb8afee90c5c1c0b2c67cb67e124e27aaf173393f34f5a9223f921a0c221bb202d96efec6ebddab1297259c7d481170cb3b22d4604e0d72f126fd2fc709d870346269a4905cfa3ec9dac1fec3de0745a42f77077c2c721;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he35f7f16be01a26536ebfa169db78082333c317bcf9ebf6e975d33fe9c0290616354d8f02eb478b3677a7f2ae76b3f909d6565f5541bb776729c0ab2a3efa296b519b6bb2a3ee6b61cf8dedfecd31ada7b9c7bf1c5f02b28940a04d7b1a7f0cfd1854e22ccd85c4dcebd25d6285c0edaf97d3842cf4e5e089063231ab2efd860a58de4941b2fbf76713b9f29ed1e380bbd76dd9448f57443d4b9bca6e980cc3f62c2569192b12013001cb0f5d1c82ae781f083c90e6695fc36fa8273bbe44af040040ebdc7d084ff6a14899687f4922bc91967c33077fbe8fcb1999021cb60d057cb65e8ba0568aaa61ddb644af393f442e3496c6b63266c3429228ba7e70474cc4ac276ceef1cd6719d03f685ce4bcef9175b6e5f67aebee04b33bfc2c2bfb500142ed21d2cd1b4289bd0c71acfbcdfa5a99bd8869ebd8870d305c68bac15ba324d260ebd7f38ef050420d57da1427535530a06d9aaca158603b61dfe1a0136752a6abefdac087bf7abaffba470ba60b56662caa7984afe4f66d71b1e40fefc3516ee1d7881c0e3c8e4f3a1e1886e8b2db1c0a5ce7434ca08c7639de5c3bfc5ed6295d20538f3bbf8d8b382c3280e6ab5573706dd1557ad790d80174948b3a0ec3057f375702d6a61d325c457bb2f0f9ea64751392737f18ad48aeedc78bcf9b7d5e4c71b1cebae985fc4bc99d96b850ef6735441b7ed2f48a6a71cbc41bc3a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5766830f5a20b9dbbc1422876265506fa2a1c2b64977c556967eec1df8a5488476737b343017500607f0386c1b168c78f434bf175f219d879b92f80028662fbc7d9155a6abe598b54eba0bae4cb42a0ad3b1ebc03a1954e2347eb04eb6be9494ab2dec88d59379d38878e131a97ef35add826b7e5a0bf937f55e4c8eabf91ee8f7d18475025e25c2a8a6e347adf55196a84b86473c36b1091fb6a3ebd99f9576d81435f37c5319e377dba49b91a74357d0efe0cb5fe172c208ed02b618d89d83528767e647c5065f341f7a2e252b1f6195b3b02403e816762dd5c68d7a9779efdf4dff44fe3aaa2cfe9dbe43e03bc80644e39583ef549185b1dfb788f3bdb5da9841502fd5befd0b6704d73c06b40034f676b25428623090b9615a3bf584f00b973aa5632ab2afb8ddddb6a59bc9df8314339cacc0a7bcbad9f439cbc385d9f1e51e47a51d9bcbf69f9316ca08a987348c17eb418210406fcf5e5facab90f251a8c45cd39e35bf3eb75b07503cf94fae8e59b4b38dc79c9203294c08b1f96b74a4ba4bbeb3db86a092f36881f3be61d10b0917b67ecb760793070a507a644e06b5136bd7721d10e4f9deabe43fe869454aeda67b90dc3e7dd4d1b837d51ea20132d81a238291c42067bfda7585d563053910d3d7596f8701294811821f15c638272682c7729a1cdda097781c678a6c42326932801db44dcd3e34036eb15bb3c6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h777a2b0de39845b5441a62d2b71ad59ac090151df1aa6ef801cbdf1c49e82337c16e9f20f6faaa840d82e6b9c58a0a344d3c6ab627b606233db8dd7f2d62295bad250807db109b0015a0d720cbebe63983c70ddff25ba55c29b9386de0cf4226e213d8f154c0d984ebc29a879b6818ffb9e77e3123d9ff5e46f4df9d4f5a1d2506ee665320a1578cd10a50df9e53d54e9453002e05e28ff9fffcd1b560939f999d50c3352a4b25b50a93c672218c6d1a2ee1b016ace1b65ff357270cac1591ef0dc8a9fb0afcf951bd45d32ab41aaaf8c7cfe660e5d57cadfe59d6ae6e7a34cb8269d955e270707b2d9a1cecb492f88ed01e20e40906bc0598962611ca4f48385474e0a0c8c272b7d8ccfe817137a795df83601bbb6407c7390196995df20043095d89dfb038ac4e5e92c5f21e7b25363bcf45f45fafbc9565c63e087abc168778dd79599d79b76a9d741f8d7f536e07b62fc3c352102ae070219232d53d203b4691b6bb16c16e8611166107c7a29eb15a4f8cb2c1d9ac7682d08b1a698b3f95d60bab577c532881c4461e6fa6009bb6483c4c6a4ccb1464650e3b312b62b0f4e9f8ffcbab64112e66e2ee850f43cf1f518c60465bff9f2c3265dab2400b12f4c0659cc8e2ea9efa8378a7108e94978c3af2f80e8c9469c16751a550643fd276e61904f74a651e919eae70dd32e1d9a021e422c7519f67520a9aa671dcea1723;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h90347679f24b34cb410e8e3a038b218e247c171d65c57cd592646f77fcbdb734d4a2d736537d18d0fc013ed39b32f5942ef1e9c656f2402382e6d9ce16bfd4a2b413990fd6a9ce3d45bcf844029692838f8955d7dab88bb60044c332f8bf91b2fd28aef73441b0dc6615cffb3489a13f8a8cb201caab62f80eab0633a4a4f3a033a4efb20d0f06dcb9172a5470f6549affa22878ee05492d8d09e6872b3861138b5263bc250506b0d783eefaa0d3f6eb9238c346b01f6ced00785f85a81ccb36e3874712723d4864a44e441a92be0479e9bea988fe33ce522ab90fb9fb4843636a75039c78e63f7a32ab0f51bfc32c1360343674bf4157bc0f91b9c1571cd9c219c0aa627d3bf15ae7d6aaa6c5607dcf328a25ec091f919be951f8211e9b82f7b3086afc223e865312dff5d7233a53c516299079b9763e2ead66d9e4b168625ebcbc70f6e6ec53842f46dfc624b58ba0ac0d2f8a58a180f84a196058746c9ed4e4a7f7ce3961234cf06cc5a20500c33f0114489eaa7c1899647e7ee84022f75f50cf14cd412456cb61db405a287e75eed2d3a64126638e1cdd31d5dc5b1fa670a521167897ff0cdadb798bdd0b13307cadb0c4bd3e429c83bf765ba81d891857b4c918229dff7883f0c48f94f930c7f71f1197306a2c74575d82269f8a81dcc5683bf209fcaf4c04567204a2a5ab4dfbcf76abff7268c9225c5227ee0b856be0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h62dbdf51579224d88fbdc75dd89e2be7fd22b2fa8eab412b3324b1b202bc033db03e5561a6d506cbea48bbfe35ff04990d48a60e5b5742dd2711182393fc605017acf7cd8a1600ef1128160efe4ac1eecf2d9822ca35ee1bce12171a8c5e8d4c7bbb7269548af0726c20783d0d703f403e7a7e80d2542881b2270f60814edbbe4f04b9d05a7b2e604735610bf3fe6ec16f0b9b94a66c1a09ea0f50281665f55a121178b6adff7f9a2712ea70a12d671c1d417d252581e775acd1002a905777406b4c77fb93a89f5564e444f6cfd6590dbe11a844d5454fee00d9e245a418dec1eb8fbc93aee6097157a33fe02924f15e5202227294456e84d3e05e68d20ea4816b6b7476385baae30a44cb0c5f5cf963e4d6d2c2dc273f48d81ac4650ceedc677d9b35121ec6ac09ef40fe99923d4d95a0cbadef3b1225c3d8e3748a5e3451de9cd070e43dae0c96b63d395039a33db988efd2a091b5c7c7b1786128419302a093ba26b3a8b8c8d2c02875951a55445fa6acee9d0f675ad5b3c87a1e0bfd56f36da87617ba4c331ec4804909cddfdb381df55bd358a1dbd53a1ddbc23efd75f60e36cf3010d24ff291c1502afd46651d7693d1e05dab4ae2d5848b98e324806b1d7024cc32ceba397a7de1531bed173d357be3e7bfe120a13c7fd137a3d1f8672ec9fa0b1d55a0c1bcfed664ed2faa92210acfef7f83d8de39320874f6ac257d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2d16ee2eee142471c01993fd909917f38b91385df219e326cda9fef45674bc607f902cc77dab461eef0d7758dca4dd899304863299bd3711e71a6e8cc58ef42f60d81af4468cb8f3171c5438f75a6e1218a1c7dd775f7a2ea943fa4ded61d589e4002b6cd0d9706709b4babcfeb19c64625d088566b8409ba066982a8acb44829b23aa57f62a68231b81235e00787863bbf8ddbd5fbc48724ad093376cffd35e4d1efe97302af0fb948f8119adc0405c6ef811d738b89fb07c1505b968964716b2cd063e045c40e7f8a3bd8d64a1e69bbf62827d9aab328cc01e19cb06cf1564dd0f937108b04d99dd817d6fa6067f951181df8d174c4acb827398d266f400dcd58030f4ed1769df47813c9852b4a3910f07e47621d20250410f78bfc453d5fb2ec026b92de22d2bed36e70e990746e7acf845d888550c11abeb7f46e6a116585ba13a8a5d20882150c50770f4c62b8128a2c15d822c8266dd4ecf8fe80fcf1e38da9d87f1cd28b07c18b9762a5518838b6e53d610a0d61457bcba7ba7e061ca8b20bc42571d6ba28dcf5726750ec3845fe639f0012c838e954c26ba0c028dc76e135ccd09daf76715a12bf5fe404338881ae71dcfd808ea43186ba769b5cc54e0d2827bd94bc7ad37cdf4bc6a63a0f70559edc222c3ce820312cf81313c659facd00dc6cd985cf46d847def5df4f34f94c729fffb670bcd7e5627c88614d140;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1c00f958a610f3de78efe127b96a6176a894bf597245d0280db540e1b5d52edb8b6bc1dc170e3d0352e37733be2f9e5a5bb91496bd28709b5c1d7e72311d3db4019a49bb1a1340152ab232db46e0e3914e6b3753a019d70fa7c30a872b9003e127f16cad014a88354efc4fa2da6096b688768e2dc5a67cda32e8a13a11cc22928f038ce6602e40f10d05171fd64fc3ceeca0d342040875cdb40433f1675dc0dc359dbe4f9dc4265ab54b7e894ce9bf905996fa7b5ca21a8bb6aee36ec27bd920eb51e208625b2287f7c6a6e26be3be23a8c0fed25b2f06bd000210ae1a9cbef4a38b52fd63b54f037c5527422a9aa4acf64381ea577f5170d295c747e2aa09d425278f600e943a4055d6ea197c9181b4ff445ae5277c2107ae023c136db460a61c6b9038fe4fe8fb6fbaab32f63ec89c0fddf5f6fe08cc8d9798a4a9710e29c2b0f714778bba9d37afbc44e14b37bc4e906c65f1219993be04675f224fb3ccb3d6128e632413e85fef6262470847cf73b48546a0fd737f19a82e7d559af1b2a88d939a7d250a09ed9e679e956afddfdc267b1bd39666a44a604bbeab5e345cd811c99407faadad2d4664f2f54e209f07788946799c076f2c0350f28b547b04fb6abded02de29fc23853346326584471c46608681aee90ac7189e2b9d5d6157d8400d9d95083ff219cd4f1c915b5f724e103f69a2b38fb79b1a560f0d9a0977b4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha6a668121c80c9a8fee5b4ced91de060579c587d61b3ad2185dffb3e2ea690cfb86fdd2cffdc5b81ff683f3aa76258ace5fa88d84c94418a455613dfbbf2e7c97bbd99e09c6a4dff77106241141bb28b62f50f821f400fbfde04300497f776c737e3418ae8ad06ffb228bb93e488f3f168391f1497c370bbb9edd201d10ca158d7c36c7d5ca0adef4879c5616099e5177a5bd0ced98b0a55e6ad10e54609cf01618b6bdff8227792d57c4cb46034f9c87c72d86021409a444ca29200c4e2063714bec91e6f66764cee4815e33130f64f84ecca6b351a77a283fb9ff455b2d806883a1d06f0968edd2df62ea7b8bc1558ce00fa02c023ccef0fd3aa3c024b528b602324458115770c944ee7459ad7f704964dfad1c2cbcb96837f3597ba8088913b74c6958d30ee69e88cc316fb80b3012a45245ba253bf0c3c13781ab64cf77435de966cf4e0dc9774a1c4a5c07b3e5d629ba87df3560d7b1077052983e9cd0916fb87b79a1d4dafd5c2bd865f573d2b8c4ec4a2439b099cb437bb8e3885d47ce365fca9baa4924682cef1e06fe5ff2601f872bf27f74e2f6a5fc4f65cf6504e0497c0a14c8d5289400f8256c913b2bb3d14518a115d5412f25bc52dd95790003d2d72bf43d59394d97f98577a25c3ec08ceb1f6b66bcd03f4d49183fb538c5d33a3f0555839949ebe286cfe37f05cadee4dd4e2bcd560166a953415e09339dd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h694871c8b372d3c443b3dd160392a6a486bcc83d39cd2613ded05a54e9d463bd25a5b879c6343f06929e25f2dc91e839c6fba4934c5fa37642f93274070bd9ddcb6b41a53dfeb5146fadc808df788fff339b4a15412d0eef638aaae0b9cd18f29757f02f0e11f9400d89a486c3bbb009714562ff245b085302a5f3b878faac87e5caa2b731043210a6fdd18c421146c08dd0d61ea9cf84bb49be531624133bc16f3bf2b88d71266ab30890fa49f06320af5868f4dcbb29a2d6f6dace206376fe4dcb6f1c48fc2ab0295b6d82ec909d398a6eb2eba21160cb6a76df61b31ab51ad00bff476b9cab2dd2541b6c79ae308936be515d9be9b182a69b86266008fec7f8c6a55a949edf2e316c49e48b7b9c35921e33a7b19d949dfa7708db410931cca33b8ee63f6cae46abe7a15bc75884951ed7066485da875e855dbb16a21b3635dec5f89ac0d059b04362e0364acade06218fecfc37348b353e751f8c3c4e56819bbbe9e3c8f0befe3217bc3bdab32dea7095abefa9333b86b2c455c45f73d9356972b516d87fc8843d2508d61def1b2c4f83ae8c22aacd5a957687136873729b0d7a05dda23081aab99e0039fc6f96b8ad2d25c13abe56e812adf879e33a219659c6b5bf788378cba96598e75b2be722d33d2351a93ee1160a659dbdabc06bf55a80430d327ba875ab94d17aa217a57a0806735ebae7c951e35d38e9573377b4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6c93993760035bab3794e3837af9bf70f73f0f8ece22e38546444b6e9e102c952bc0ebb790ab898dd48aac61e97f37d8f126bc5cda46009a7e13b5c128c70a8fccb3b55c51369e82a891ae80e6335f6ff84609dfe8e061f21e77b60ea5638b596ed91d2f9d2361fd5a9e643bc6d94cf2d16f1ed12a36d0097bcc7dcd16c67be2ff422dad478125164fcdd9e7b6e0a9bd03a01a8719a8656c7906ae7865577cb0326bc88b4a7a96472fa948068827d625a23cc208a1a730e2d6dfb4d9e2a2b06b7320ed6d838ffad23229d4cf029b541a84e500f25e238d12661c4b2bf41ad193f068e5aef8924200bd1557f0c0a8bee281df97b867672469a75926d337f8355488cca9217209d4ceb3112c110b59b53258e7e38a1269e2777a37656067b58cb2a15802a91725b52afa9f29a0bd68df277244dee0acbd7f3d2bc1b8d5fe10e6586486f1ae180a06ed18c1e3ced9fe5abb4643c0a9f71c5a3538f75e9e4cfae1f3d850cbcb638ffc911c45ae149f804fccfb384b68c42d39825e12cf5f8d79339bf6fc10c19387b3b7d66694a779b1380c2dbfb26bfeb432b84689e758285a7bc2cf12e1bbbb7a9f8aa57184a8e9cd0d1b121f5befbf2ebeb04a99b37476605d71e30d072b1e3b6aca4c13e785e4c08997a0abcd17c790ab025e0f6b848e2d222db278791c6cc3b8281ac0e91899109853bb6f1206866a8946214aeb3c618af68;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6db8d957b532ddbfd567fc695c4f88340cabfd5091a23c9561e930cf959bf3a7dc24e08cd44b9d264bb47180bf03d32371b9dd64849ef1399ef8360649bcb2c7986e9f37cf17d92d09ce3dfeb6d737b2dbc3054f46ca8cdca888f7674c865e5478365dc54ce92f413516b0c50199cc4417cebbe8c33f6f5bdba83d2e3078fd091ddc324893f57f29cf413b1d77c1214bcebdd78591b2f5e1bfa2272677677e1984cac8795cdfce6e7ff26ee350df34d17c3b209c901b42991d93b1321f646b3f4e8bae59f6d36653c755afc7ab357638d37d00960e4c135f9ac8c33b3fd0d70f176070cefb03caf96740e7081e23a1e205229b097ee5dab5ff5a0fff62091da3a301e3996f5f2989f51df7889381313c88ebfd047c3cc2be7a29118a16ebe038ed99bca24a759448e10d75ed91da3e5604d130b49a05bd9db0e18a772d7bde5a773d3cbb3d0d81f092adc8f09d88890403e28cad41502628e6134856c74b3d2b17fbd156bc062fdf4c2f2a72a44ca6be8c5cf128a55bc618dbc5a0b87dfd9c0e4499465314ecfe5ecd4baf5fe188566b8a8ee46a74d0b60703ef6ebe21a757ab2c1c397d3c07c27c75ebc3143a84f25e73b143c1226181025d79e8d91bb589ab03f006e09917d5d26b3ff5c79ad4e2a8336e302787b31f8b154e7b3a0494c12a6e2391481b8938c8d8d6cdc01a1ee62fc3ccc70b6ab11b38f10ccd4f2ab29d2d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1bbe06f3246cc0d74b1ac9ec7fc87e28e26bdb3a699565c017a59c26a6e810188161ab8b1bf0c1059a80686193702bd42898b46397ccc923219211845b150814f9649f27508d4818d895812d1ecf61026b4bc9876623e009e8ec84194276836e164c9e84cc4ea4db8e40928d506e9b347f8376acc716438c868249933aa264f97498290cf58da5f950d20b49d3b7969d720b9de198d28cdf6c556db83f3985c122af9a52bf0b89773a76d42974070fcac83c65a6ff134dd51289f284deda74a552398df9403ef8fc3734e5d500006a9f2b1f11dd7e83c355860beabe0f60f412e42f3e70aac8a6361f0ddaab8cccc14ca98318e985af634b377cb11a3c92e4cd2650a37ad6e4468a6bde110b97a6341d8711c9bfdc5be8a373a1ce419c714fc83e5d076ba65c22e7a93fc40748f5767d1c649f3058ef8f27db2680744d563bac3b7da1cc868897a0b6f4d1ea0f01a0f12521d77777e0d9c88906c8fc5318a08077cdb60029102269a5b6926c038a41820475ecc64addb272f96f101e74dc844e8d16b03ff49b6e6bb9fc452f78ab2d136f95b1900cad3ac708bf38fabf6fe82170c8187c8b16d616f56a516b945b724f71987fdd0bafa4063848a0c62bb69cad7919d7167ee3bb2c2d0257465eca284b72129cb765244b217d0d63363a93e8eacede1d13b5dac8151dd34de935cb46bfc5b34f10a9737f2a3a66444b266ee177;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h19dc69b60c927a354546d3c8976a2f1057ccf87d7eea151b61bf4170b1e9a0679eaeb89df615ae3cf86703f0f88f292e7e30471aad534a9f413df939482ea8aef20c0fb6b8600f61050ca68024001b7e794a22323b87fb4a3c83a58040d5ceda90ccf4d3f4aa35c76aab749fa597f023d8bbe745d731548d0f083f41e55f29a2ef776b8d8b08613c08833ed1fd3c214573a6a5f1b08bcd5811eb16c4ebb65dd408c51b3405a5c31d683a59544314779db9bba7f1b5a17299f8db08e3d865435707559486f0dada08698143f9b777ef804023c5e7a3e675e953e8452de0aa508a296633b2ca07352318963d7bba2ca2bda7f3ffdd9b08a5240e8d8ec691b60b0078c8c2b3f03b8c247aaa9e4970535678e4b8369384ef7a4fd351f0a369dfeebbf8df2184b818fc1ef2d39d233178a62b99a55f08fa81b1180cc2fb3431824cb7bedf3fecaf789a3d3884402d5d3a61f2e69b9eaaecddbc9c00d638f2808d08716f5f55b8e4370060f0acd9d108b27890ae80b1469a3032abba34f0b82e250017e6e173fee6c9d91c09d9164b69394b2dd837c395045d58c7a4749683ce4534defa05f9a32d78d8e349c0ffdfb9c0b5c5142b325ee6bf02e0160d564164809bfc444cbf36aea8ce9ba90dfa09121ca5fe80aa82e553309a2ac7103a18601a3723d0f1f2ed66984e7d5db9ca3c8d1a3ac8019e7ac7f6071e4b833f7576c075af32;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd9ce6aec877c8444c9b094852661afdaf70c0170afd7d9d0cd453e3394207f21fa320576eb1f076ed32658627f344088105b8d5986a238cf23fe4b47bfe8c090df35d2415aa33082efb52c21c94fa72293d48e7437095a6044e91a08ff555dea132804d27f350f58c3aafb9af5e05b09a0b844e645a92892b0cc1d4e8a12ffe1fbbeb97d301ed5bbc1613ed20c0e9f3d2d23a1bb8e26b51a1755323bb88434412e19009a54087f15c2c5804bf8c017781124b84e9909136d51684c8baaa8f0231b03732443baca8ebb0969e85ab9f61a55aa685155931a3fd3eb420f8da191efad539ce07403bc5c8de45c25db4773eb43b33cec3ae059dd66766708c30246bf2492034548124dd490a7ff77ed941ff0d3d7fd4d084537e99feb15cebf1ccf9adc3a0bf13a5cf9a85cac487dbc7d235dc4ebc0ded0ec0683f5224c0b0deb69487cddc745371f29281744633281735dd7e9c081185712361f3e6dd26a31e558d0f38c8e07c13c4c6724b01f3e738988740c3658b458a097ee6d682de99aaa842ce046edcab1255fa0a017b6f3097d97023b64dff5988e2bdac2461650b0e3ab451181f69749976d945a1ed0bb93709142e99e45da329ba37d916db022473d8c3ec92b5da8d80053cd9f07de503f3af0866d9b9a02c5169e04cfe5f90012c40924934802767c3db10fa6ce078e24c331fe54e0f221a7d484474604e14c22103141;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc1be71755ac5fef16e3200963f2ab51058356bec4fc6f16d246d0ca6365a88ad95dda0f75412190a83146e4c5c1a3ba7dddd41a9d6764377b72e4858c45ef4d4fb5933e171e394476d68b84c3c5464f4f3c66e37b44f5043082fbcbae470f3a568cb9c9746885a76fcd4eed80b3d6b0af9df57a0204dcaf68493b2ee0e60ea8477a2404fa5efe0508b9a337d3f2303177ac7be1497ad62f70913ca8237a5623793ea51697e41b219c141d0e05691e09504d810a4d1673d97132c4eaa2ccdb434b6d249e22bae1eb3c3d9460f3d7fb8be270b580a71a19b4043cb925828a013c35cc3b79ee86ad531bf1818e7b30d93f3edb8de462ee9e8e9677dc9af2ff9aef182fbe8328faecea73705bae9464c631cbdafb2f125babdf95736b75534b1f5ecb30920455e47ccebcf4df18863c948a00e6bd870e18d12c7a0bd7faedfa816bdbde128e6f98655fdb3cbee10f0e2bd94dd19d6ab858c23f635a78924a0a892fa4185dc0e609dab6942df0df87a8d6009e0e8e125aed7cde803e8e7884fc6f5cbecce5c9af0e480f0e83f15ae04205614c3c1c7328d28dc1f30b6c1eb28d0f535e5cbd1a6ddd18042a268dbece8f70ac3b4bc0073376015946bc72bf7aaa97bb8e433338de8bf2e792a7f9a7aca53ca60b256d4bb6e4f1f30cf67c8cfa9f41f45d0cb790cc789757bcf918ae3c2f6114dba93382aae25768666419ed9cd785939;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'haa88bf650738e59dc8259e1a483ff6a769304bd29d7f4cdac15a4a23893470cbff5714233c42a7c246d4c5e1b36a73b306dcba544f08eb333be9cda9ec25f9efd6ea0191fdff9aa04fe053d4ab448e171eb83f837a320f1147006be0f02152474ad4de1c028b5e41daf52816f6cc996d4400bc279245a9e4efae50414cb0d7aa435c3e230c732789055db24605fb49f327b09702a066acff9cd6039db8f9c742e5dc36581e515da2333d265e6cc6dffa57ad9e518a17b1a19338b17d2730cc845f3105a9bbc7e58d517e3a8296c162df1436b3958dbaddac64c8baeabcbd20bcaff8375bb9972544a1df8c775666d07369457c6bf353258b0686d036a8458b8c2826b60fdc044136a9a672f035be8b3bd7fa2981bde7d9d14d7bc2e9daede8fed420a544545721cbdb5170d2b1b557773c71aeb0aed37d859d94dc57debe6de1fcb5b613e237d0a6ee2e4f3ae84986e0dedc0f6de883d67cc1de479ceb364af6cdf784e78daaa87d09e1229f87503446cb240e61831b3bd077707bca8dc386f0e69594ab06110b9f7e94a9daf0f10a7a6c68d28f050296737502596dfc6ae6e5ad810355d6e234f47b2ddc1f26da8c00e30d1fc45a2a14eb5f5b7d3fae69c9f2d90b86eaf93decf3fef9cae1eecf2cc44eb1536355ca71709e8329d36fa80e52356c194bb29c34d0808d150c2677dd236f2d12909893333145b45c46b5f8bb00;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9e71aeacd716a4543b7c912ed588542d900527ddb91d38c9a0b863bd0b606e552e95339c7cb60329e13c38a8e4c6c26cf01615662bf4d2c7d3a8860b4f5a2e7d10f489cc6b9b1a5dcb9a9d3934d10010463f8717f3d1f0a14acbca6807c0a8c2ff55361ae42a05b2ecf5d6ce34ef131bb9f7e35f8c9edab8e54e1611c2186f778de3f00f5b61040e69a3199687b2037c1f16f7c562ab6d89d44d121997dc72b6a79eae7ea5e87ee202a16b168c7ce397a043fbdb6e399cd1f76489822a918dc2ce34583b87aae632c01334e09c2dd6a43da9640301b948b935b6558edf4931e19a176c879a4062f77ca503fd1b95d953db0f36a389eb544f0bddfb6d871511796e159165383b8ab82a83d8a88cb7922be2edf2f4ee5117ea6673a11a1d5ba166196df8f56a89330575a72bd752347ee757819ce7030ad03a7dc6a84bfd4f9237b41f5561db8618d73fbf413e4e6219c1f08ddc3ea9040ec7f1afd2525d164998340556ac311194fd812bc5d3225835e302bca51319de9310d66dc8bb3dcd2fc9ad56ce5589eed77202dc86887beaa88db3f2562af5cebb41b63aaeb88b45a5fde45a514ab2747f0c308ef8b7b8aa37f7f724c610cea8e34ca5a09c06e938d40bef8b19d0e98edb4bbf43b042c330ce6e15c8d3cdde46159b1e800c88caf718dc600e5fd147e88992f9abd50f7079960fc9c2a623e91ee83e829406c1f652755b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h705a3fd6be2c0f1bb2414b60c573bb24513a7b719669f2ff5fc8e0059255737f78b7fe8a28726656fb749adc01e46894f1c10acb63821dba8973a662a53d7524ff8ccc89331f8debf591249c9456b4fb07e8d368c11a4a36df1e5b9ad6856e8d4e73b3cdcdb6af9410bd57ac77541ffe5e7cefcaac48668978b79574da32a0961fc6087e0dbcf19e8476a59b87b20501fa2418d0fedc6af7f43829075dcea7100b3685b05bcf745f728a16cb81a78d925e322664080e5d8f24b5cfc7bc5d963659035f6eb11c63133d3aadec4852cac5924150f37ba2733a82bdbce0775cd0a01cde2b58a782a19d8f0c9bedd6dfd7197d9670674571ba8fc124e108f017023aaf45ebb90d3ff4fa0712368afef2874c97ec9935f707a1246b4ee514212ca71d7685ac82aefb093c7add882117b27d3b4dc0f3274ba95fda9b0c55510295976e9c2a86d822961d2c840d2525e14fdc39e63efd47a81b5a6821663abae65f7eda76a47bee88309106b094b45a8f53a3129ab47ea1b7b26c5ce8284d6199658c003692d4f16ddad54e61421ff6b7b804cdcf215848c0585838acfd05c39b463d2ab61ae7a0e51a8145f17f42f16414fd84c9fbd6f7afc1a79f0ef6ecc8f9ae5408302beba8ff2071fbf37b34f9b042f0e0accc05bfa8c5f8501d569c0af5556b7b03767931736283d14044f15c425aa3cb9d07ea3e96bcfd47435e51ec1e7f9c60;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7a3ee47a89cc9d67ff632461459de80c48fcd218d5bd9e8aca40435f39d63025609d51c87573b8ec9736192f193a1aa200f89567b9e5ff9386ae09c312aa98a6e3ba0b677cb624cfbc12a4efba59d6c3d2affb84dc0b8350d37d293e9a325da5ed0446480f11d974afb8d5682bd286528dd27898f2a6890b905de2d28e24787769397992b64c793be90bd5e26fd61bdc0f7e635847d0bd0f3f0c5d5cf80c3aac4cf8ce78892c4f1c06c4e20fc8aff1e089f2fc17f586e69c412932ba1a97dbbe537ff09b12a89b9e38c1e23f7197a786b0d78c4c27c4e0a5e37d23b7b2df7c64d60b4537131cafd278920c5f463c3a23c1d41c0959fbfb53cf86c7509ac9634167cdd77dc65871f9e3a27631a4c9f91cb337449e04c74d3174f7b89e38cd97862faf2e06c1090d0548cedf167bbb46b10a0c6c0965c92c550b297c7b687cbbb54ca172694b2c50fe17c9cec9cab1dcac45ac78cddd3bdceaf2202ab414e4bdd4e9e2ed8bb96ddf41329c795c131f5b2c067bd7ae5687205bf76d5fad2ac8316fd7f964a56baca1034bd7e3cf4e1065995f3fd031d76d3d7f20de48484e01bde06facebbd6e4f04fb99a1e5b4c462bc152ffffd283a84d0f3c2ee42282438f94f79a51a714d93ca6066eecfe4a1430e233413d3f2e4277de4e95eca578b7537548733b3acb22ea79c71f0aa683707a297ed4eb957d7b80247e0300c954344b683;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha0a30443dd85e6d94279a896e440aa9e40c3b5c3373da4968dd5bcf27d2f3508fa68d8a95f0c560ffa768bf4f6e9eb8a4eefe2fc2b144a497ec41c6635296653c96150020eb4541e7bfc26c92c404e6dcbf5eec0a2fe9c78c83fe5ab6e25bdcd8c779961ab4d60c653443b098772cc0ab08c22c79cd8e9ca2a584edb59565900d90c2334f2cba5b6a0b9d47454f1606a24253785cd844f14c9733ed944300a85ef0d622c43cd4ff21c752ea78c44fbc6f9e80fc9eef5953264daeb2e939a759710a6b85e4321fcccf722facedd2596d5823ec9884bf399978334a4d79f07188b728b7bdabbfe757fe459c34716382591b67da2696e1674fe3306ec216146db16c96b22b3792f5607f35695a1ebdcdae23e00a56211ac6450651278d0bcac4ad3203c6776e2e5017024bf60e1caeda331a6fed7ae118630d1ca48e89bad2e22dfe370a0a1ed32cd3637fedcc88b36ae92c15af409e7cd625c96b8ffb759d3a5537ce64969ebe87eabcb89fff887a7dec1f504a03ed444ca8b7ff00329cd1b5227d13e03ea7cb17db155e87c8226d2e6bfceec9beb78e452745d67d2ba4556e86d7ba215b7032bfa5f2d34aeb612655c74c941b10b9ee9989f665b07712b834bea732a02053415a877f219e4d21d7973ba96412df6d85192e8345af7b528bc7c11fecd7d1fe232129dd43c4b6e9c9903064510faa1f1876f28b51fafc0bf96fa51;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'heefa2046a720e18ebde0ad96a1afbb95b172e44e8f1c94e7117404db15da8779900c06c9b1af9789940b7729132a56c9a63740b42104d9f446bef5edf41e99932089fc98ae1dc41c16155997df3adf6fd6a25f3432773ca840dbda02fc351994a18c45baff8b8fec0db8c92c47e73d3e7aa2286f6615fb373df405ea3c200b22c7a7794d6d76ed3d32abc54bdac12a2fbc57e558a0e79f6d122a8e35f532847645d6fab9d836e880b70f726d72c1db959229022e92320976cbd218c909b321b0f9af424c2aad69ce4bb6b6448357bf6552eaf27d9cbbbdab7935207af8b0f041297d08c12b3446f82ae1bed537a68bc3bd43b90e935aeeecc9249a6954a54f2b0a68f4ad8fd5ee6a11b94244d9a884b610873869ee3a6006fb5e99f9124c19b4f284aa440b4eca643a426843f5ff21964b35b890ff28c95c78db3f5358914b9ddce1ca89338c444cb2eb2b2e47cc8d1cd09bd6ca3b9e3fec1454848b0c4f1c21ca3cec08a2b1e5aefa01863a476ea310f0a0aaa81e236195e7e50a154d4bc1ee582d20d81bd5c01f5b537163dad1f3f5c4484532bb2a65e9535b74f1fd5f702f2c7575432b921847948cd0282326211aa11881934baf82f5efd0056862da37537c3c3396c6882c1a585bdbf6cfd908729d44414adcb83c5ad6f90906c083b5ccd894f864e9c20c25628b4fd88fff76f821623774ef7b3c5e72f41a65af2c3f39;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h774688e92064f6ba7febc53a7b3ebd2caff8d6f00389c996c3903671520058ccd4f96fccf6e8c69219b2148f482f2f5c36dd2ce629ebf4af81d42ca758ca80c99fa0bd6a5448bbddc9b007e3718409191aa0a8f0125c6acf0609ae23d17fe30b4f878b6375e89141b73048bf4e6686eb57dae05c9a66e11e2c509ff0b04826dcf9079db9d5b0a052ed5bea0c9eced46d58f6a5b200090970f0993750434e7f765bf2a7ccd884b23f6759822f056b046c151446a7de02058804a48e580aa3e787679aa754920e3560bfc6f6af2da7b5593513086f60ca801b4025f04acbbdedab2caf22fd4734352302e31f4b1865a714dd4b06a39347006dcae7965b2c4a8633c71c95b76f3bb8e0f0c7fcda85895128ef09490b57f078e0e0f51bea750be34e7f1fec5ea5c278e2c12c6a6d23df7b2d22d059dc0f843fcbf6b99661cbd8f7fff55b518c40840ff065a31abcc7c059deeade7c7534e03bfdf8022c379d81f6829bbe3748662156e8220292312be287752f624a80bd6818d84de3b527d0e69511c714974283ef756d4f51b62ad65da0a44dd9fb4d1e18fd37b8fabae6c3d71508a1aa9a30ae777daf8de535dea12277ee3a4aeeda97ee2d14f9a2e056cc00b2783e078804fc8e1ff72fe07fe804b85ce09a06eb1237a3e3d4bf35850048b52f617db8316c7d0fae08491d38af5973b6b47b929e495db55a85f97ae6e56e4150f4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2bb8d29d4569f5fbaee728fdeb2c8c0c2dc7d7ff0aa2546457ced9d5eb49730dc86831d9326bfab473802acf2e3f932d6a8535b5a7d51a475f13f3b3f0ab60ad69c959af50edb2d33b3e9af697fba6a022aaf65cdfbbcbdd3ea794d807ceaa321402ee7448df36aa9a8defdd79ff0a6c55bc71ba662c59c702d009c9f8df9b177841f0a72bc6bf695eefbaa9d5c86d1577567388e615a34c1dafdce05ea55012aff35862749f532f0f9edfb38ade852726980ea37325ad5f3d9ef537e40f0ce17482ac78bab8c8261fef6ee5acbea6abdbd721ab6ca68162931b13f8ec8a54afa28c077d68cbf8246536d1401d047b3b7feed1c6519b1566732f27c2f77636125259fea9fc2c47cf6845843217942a5f2cd0c451ee873b5361a39739173239d372aac0a9c1913fb2ba1e05dea3f42ff31886fe6f73d65f28aa03bc46dc167be867a79a38119bdc19b2bab8202823a65030ece0a6f4b2286be682e44307101aad2acca0e3056b81e97cf319ffffb20fb2387e8b7d314525eb37db9c424bb70bb9f1862b65b2abf36f97c480e81c3ac8155c0f2adaa730b6b7fa83362e7e805056585b82b5bcbf6bb57b425f6a4c2b2585013df0c7f3aa58b9e82b85c350b480d80ebe2d3dee091e6a7adab008b7bbfc36bdea67836717d0f5c8fff1600cf8f84d1339a898fe9b4c1bfcabc6d761b2f6f700897bc0795837c32de8b46dd088d545;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc3c520de43ee6a8d52d74af79ff62e359a9ace2de569bd42e73d2355601370fd63d7da3d5848bd2e6c0004f6765d0c55e028b15c7ffb035d303113d6521d361ffc960b8b8cbf0b0c853665192e5902254a2e034792f147237c3fb160edfe0589f041d4873b1fd6948cf5e65ed62ea4e0b787475f385686b157f341a25606e325ac9338c8081622d0720b1e6296e7d87ee6b3b2e909746a8c4f2be20ffacd8ace47e5a5abf6df860892665db512d859dde6f81118f3f02141ed1d357f03ee32e4ea8ccf7626edb60bb1ba350f3591efb5cc41b46c8036e433a1b4045e8ba6355f90df3a218398c136c805b30e86d4a144153b6ed4e5e62f6732cf093c669173b329124baa0d66ee504bf6a8af561f9fd3d5b1b430fd6ad5ba9d79ae174cc495ac7d8b430612a36ccae801e265cc505f02a0c877b4f7f26033320c4635720fac79dd90798ef7bba873443bbbcd1517dfebd314de8320ae6cd1b11cf2b96c7bbc63f9e5d555d612760d1b48cdac889980a4ec4c79a74542a89cbb7ccb2b810e25ec0f302f68c4591f321b9db008a99234e009f82c9e9587a49eed43a14d95b63ebee4a65dfeb4a14c3c115fee36a133c4e854193ab8cbbedd914a90d039b0de606b530c0ac5f7344f751022de0d16dde267548f6f403dd8733a692d3170f540824d72db22909f56de8af67ad78339015e4deb5ded94e35e61a164585a3e943b1968;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h81a8c782213a9157770a988a173a5c83cd0eb7d73d4d366feaeec0151509b6b5608317a64d51f84d575d30114a15257faca0974b115653249a56f482c3f06bdb92ff53ecf357575ac79de17e6673b95b8c1d964e51c07a6f4672a82f8d934741994b2ed365053f3a41f636369660972011724ca49c077d81b494087129c0bf2e24b427c7f515bf8ff56bec4e6905d75015cee3cafa388617038c6b8ea3108c48bd83fb9cb4989b8993ab2566228634ad5c29e3b3d00fbcd5597a83230eb2ee856f86932aa226eb7e05e9026a0ef71ae10a64618da1678ca3488ea18739dd5099f5478cfb21f246903f319f88e8ce0b6e19131336391b9f4cbbf109f7fd8c97c0307aea9ca942a262bd5dbd8b1f5ce6ef0e95866386d8e1d458d1359add259ea00984e3cacbcc3d4e97e3cf7943b92103c53d9e29cb6e6295d725a3196b11e44ba2ac746d288158d40c42ea27c31ade275419586127235d3302ff41d2206ab5035a1c5cc2895b1a7e7782c67c428436ff5a37cfcd332dbb5e82d21891be6a07ef7c2c00e23eab23cc30ba6614daf73c63f59e3e75ad9895fa9daa136fdba192526f6b957200ac8ff95b0b67eb2f40f95a1f8d7f6300ed89942ddd0047432d2d6950ed717b9ddb115941c074d73d17a604376589d5c6342b2dd7091d16ea4f0a4a7dd977ad1a085f1cde3a7255c41b3ee3e42e1914aa4534d9966b8a9a4e193eb3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcf46c36c28fe0deca618f9345398f097aefd48804400867397c894e7c981122491cd1cffef03f176e6273cd80c771eddb058f316354926128615b05b7d8e5dbb8158e2355a397abee6eeec3d1120f1eab5b3d9825d22403e4a41a99e92680a9502d24d468c4c25c71ba919f22e297931618eb169419ddf3d016da5c3533902d522b7d37b680212043abd84bf3eef313efc1204326ce29fc7c71b76aa8d78a6133a6caef5f91bcab7e38226ee67ef96f5c02761eccee568364eb47ae92409a7d06ba4309fa3ca72219ebb7edb5f2d280a3bc85caf489063591f8fd79c46d920b08fb632c3a8c5aa6de5d30da09124e41241ea848f2ab18b493d4a925fe2cdb969b4928d8d235d2d21598e92dac0b3fe86df3811dcf2154ba0465506966135afc9fab96e50949fadc3076a8f38c29ce59326c53a4c8245d7c3a457dea0ab9ac4155b4887f02785050bfcc05f004080402ba0bfde0c258afb08bc6e07d5ee1eb8e93213d26427420b20d3cdfa7842d1a47481fda0ad0214ae9496296c381410d1c188c8075158c4026b8f803ec7154cf40365f9122a92cd0237391308355d04f5ab977db8af58999962298376b8d21d1cf7ef0b2a6cb6c1b2d6597e7e9dc7b8e1be5b290b03963ac0bedfa8ca2c7af6628e7b5ddf659144c37cc5d42c4793d50012df0805fa8b04951305fe0b428fa5063b2623d758ebb7602957307efae3e0f78b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1092c651013f0b408d46d773f0987eace8eb0f654a562bb59c5c7a724723d2ce17e9feca2a98a727b5f413f5e9015c7ba576ae18a11e6e840bfac3119f3747faeab69b642638eedca22d98027ce744c9f695726d1bfedbcf53ba762fcf37ab4611930bb22b7a65af599cd2395bd0831f7c2c1baeae3315d0e4acdcff6dfbdb486f3c654872cf7d2a32e8523431987dabb8be0da1eddfbb13264f9b838cedc7c92aed52b71fda63565a8763a01a9b681c20b3eea5fb3be97942d9b662c0aa053e3ff10805acbe557f0998858be51abd29d228f622b922d822e8e4a48724343f40f69489d71ecee14214db60a903e5406c8d9501a9ffb2f5a583dc49e6f3fe605856fa39175d90f1b862c7622beb96b45ec8de36cff8e4626c3cf5a71d554047a116b8420e336f2a95893f1525e188b13eb44f73da7f1b2974aa83a5e6a9818369c11eb6f666aaed4e8c38a545c421929cb56274669ad6c136a4017a784b7aae163f3573b90985e9786b1ae020893b5e8c26742b7ff8b722e9153be32c2bc51e1891dbcda8e2713d0efe73664a375429f4779ff22f03f6c92c9572191d19a6363d39dfbf447bc3e31402d04257af2a2a86ab6a99ec3cb7ec09ae599431d84a7304a4873d3df65ed90f185a278fdf5257a7d85bc737753c50c1fb28c951d04515bfb88520c54979ca8fa5b210d763d1f2c9de9f25f510f566636e18242bd8087a6f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h98e8c58008bff24f14377ccf81dc9be0c4465e858f0f28ca0191febe2f48052cb2fffb50ed985115311acbdd03cd4ea39155d4143789d2bebe361d7f086116720008a63462f13e6707033d3c072e9418fc766465a0739d4ecd369c7ea859d27c060b8798bf0764516397ab7b09fa73658ef0b5dcd22805925f85a6be5d4dff7065816cc8704e34c070743c0e52eaf114a46e4505dc65e609d5a4f3b35f40938d3205f11d1265c9d16f46aabe3ccaf1748aa5e71e8a8244ccdef184efc2392a04b323da891d9e37ddc70c5cbe519c589285911cf4d25c0882030f0b73517c5c8713666e342609b9b9b4c3eb69730295e2c299565eec3e79e99b382b35b41766ccc8a24fbae30431edba77f88267c5615963fdc2555c316caf1b23ac2fff9bf9190e548394bf5ed4f18675e56450c12a4a166964ccc205ead7faa91af370fbe7e9d92e1896ea4aea96f956d0d9276980418d81445337884d56872e9cf31a30d42f99d8ef83f8ec0f8c50d941c3504a18dea4a0c960e7ba37a4fd0cdce25086cd70ce76c31930f1bb0e1b2b536ade326eb9ed7444a3911102f3819f8816f2e1e3c8dbdfaefb4c2a593f41f274a2cae1daf1978c804e21df513c38535c7111f1f4da445625c01c4343a8a18374311e1209088b31df5c080861db76bda1934d3453bfb8cdee7450bff4e67988509bf3f321119a95b5b39e8be270e5beca016c8dcbca;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc9847ee67237843c86779354aab1138c27b30768781ff286cd2b77473ae33060847330e9ce9c07d9762218943b81fd6e086abc76eb88c3659c33b484150160c1c3c4a0441c81f828cc55442df331556bae6e9a3b534ce2837df0e38c063d0dd6a6cdc323a6ee707b6a16251fa83178e62c1bcf3e98539f63cda1e0896af9bd81c460221bfdde748152f6c9dbe76101b403c14732fbbd512fc5fbf0e936a72e414c42956f3875dd6c5f6426240d6d349c7b7ed19a9ce95bd3836eb0b14841ce9256da1088832f696b6da6438f30d7da0d9934d4b5522461dc2971ddc3de4e95251d983435e13b0918a316f38b97753ef8a6e5545769830d30329ee6b320842f1e70b50071d023de54b5ea3ec890b6b9d80d6de5b5685fc2198fd62644cacbf315de02ea0995b24dadec7264999ac20dfa6bc3990763ebe8171442afcf87e61c870827eb9181f620ee73d186387cf4aaa8b6fce2efdf14b5ad17811ef9d22116fcb2b260f9efce147f3786e2e9f312f7c46f2fa17a7c374b0b9a85557d0e6b3496f16fc077ac823c89dbaf1539300c3a47d020658a1a6787b022a6d1b52eaeca996a072db5dcf549bd4386f1e88a0cf5686ffb185e2abdc17347f6fe480309ba0b710cc4895a59feb58e57c3e72b12f37d15eda5d4b1136d4f2593593a39d99d79c4f0ec5f4cca2361cb417b15a873b01adb69d69b771fd5f2193ee5033676ce70;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he6bde9d81b5ff010195a4056f823cd1e4528c800b288ee4b82e58f5c482339bc935dd8692ba8ab50bbbd13c22b968524b7bd8858b4e70ad10abdadbdd3658684d9fe73507906804741e472216c1e9b195f2f5fe0208e9a9c67c9afa9ccb0d6595ec8e391765633325f33d36072accbac6346bb9bfd5577c8acee31895d5d9819196874e6d524cd1405b30aae78c423147ea41f56e5e235e77b3820b2a31b1e1a438afc98086003b56de13f12e52ba5bec4e5e99e52f59ef9a63fbe658b682cde6c3293ab726aacde980644b40367ee1ebe800b53b767e9fb4347f7421981cd35d16eb615d3e362c43408fae6f9c2f633224fa9a51c9b1a3e3e9c059e57251c9a918a601dd15572eebaa8e5c21e81e6795acc9f190f239dd5faec17a6f614459b05b0c8ab1e8f98e05feebc21361fa1775553de2b29f26539706f862074bea260ce28586c81f608d81cbba439be4f880f0553f1804275e0913999b2c48eca83c673296118fd8c7af9bdae0a32280fb9ce2ddbc036bc952540b16f95fd855c6ae5f27415f4d796e2b0d32316195483915eaa6ab1fef7248cbcfdc0b1cf15494ee0e649f7ffcae80cbce2ac72fe61e77dc60af707ec0bfa130cf0f4773073c364a433b0488c72ae0886ecbea74b5014643781714985f4dc6153509c6275e1fe9263938f074d373cd8972b574631104a8e0bdb8399cfd7db4b00eb70b989039aae71;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h54d1173b6df6b1432cbc9128fc2cd71223a18292b6ab9aaf71b68ead7384c760cda483385c40e661445790fdd9962620ce547acd27da987bd270bbceb610fab1dbac5cb5cd44b2fd266783df9b83e1ef95486737a4ec60f7c947c2d36d6bf56ad785df306cfcc6c279da15701a2a1ba764f503676d455cbc371a7efc53303a38d7089e3b2651ce8d520222161d5556daee78233a7111afabb50190e811880f597b9ef64e2dc52d79c7b3311798a6e980ee92cbc182498854981143d7e61b7c0c26b3afaa61858c3c4b42f25bd517097ce29f6abef5357272307131d45c00e86c5de4d313146664b8136c05fa1f4d8763ba49d71416e9cd6c047e71345314c458dc20638ab8029e4b32c76b8ce039eaf4ade6f49b5b73371692379bf9d56df3ee72ea2461fd387fc80e55954d067a2c2e2d967e1146ddf5fe679f86bbc5d5d9341496095b72a63cd9740621cfb71794eadadb6b6fa775327d72bcc2fbabd306af262e2e3b0c4195e2d0d25baf64c833bbdc1ba1d479632ac11f5f353217c99df9d4b6d1bea8fd17674ae49a8a834701e5e0e4a6b4efa367c75a9f2289261d98d94d0c126d4af1965ed0878c7a7435caa22b88e8e2a92f958e44c7ba864bf6f9c68cd4e339d17c22a05c1cacef6cace2cf32104e94ea9fafe14d84cea6745a74ae35eb68d290835eeed841ab20fefff5f22c119137ec49a8022c35adfc5ab1be91;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h412ad9e73f078ac154697117552a76bc86140cb2d02ad3e1eab8e572317ec3146d983e58e6d8f7e28816847b87aecf8e44638327a7dea723009d300b064dc0d606a667a45e4632bc12c44e18a208df2b88cd9da1db45dce103365e81298021c103a0ee301805838bac51c775b263478e549b9d430e3e234498bc6e947942064b3d089ecf3905af279911a8e53aee5f157c9b559bec16b7f783ac7498927022c560c271a5571c950cbadd842f0d20ac30cb6950cdae63d11319f08823f0e0ee74a6a2b38b641d724ae7a8e56f72eeee7934728180655bf342270da199d21c62f6c4c1d01338bd7da0e49cbcdca235fa28474a6d30a3d5a0f1ab3c8fd9485b961425f73ceb5e49f359a1e1cbb85f3dc5615e5066a0ee6a939bd5d057e8170e6ebed2d5383e69943f9688ea38a21cf869dd7d09c4a592189b771591fa2b0682d027b2bf0d9717507d315c6a0fea53aeb36e2ae11a554988080bb7494596a9beb34229b90fd265cb19b629fe3cc973fba89e22a10063da69b80979cd78b2c18c8843b688b1d7f67b9069039c788a0566ce2a40ebbe44012a0f6509c6e13eb845866e1d6adec9af4ac236dc65c67005423d2b45cc2f93aa7c7aaf33842648f623ea2f1255f8ed2841a3da8f88d7b89a0440ef396e315a729df5cb1f9329bfd42e947a8316575351bc791c89a76676dcc349509f1a461afce9a11ae8c22bee541ddc7a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4ff75c87082ceb43b97cae545daf8d0b2bcf98efdef6d796d6ca78aab96354dbf2249c063ee70205dd0ab236788f2817730441a80beb41086c96ba71a7d9c66a5c2765ab1dd9b29382ca0ece4ee9eaede74bd06dc5c94cf553ba63cab35d7e4e390dbc15d82ff4607f63976868bdfd3b0fbb9c820db332cb85e91e81c73dc4980669ae311f46afb7688e1b9d1cc8832d6658a493f58a237fd49db79ec16e6ec5eb2684f6fad1342600261f9f5e6b70b8d3a2a2c35a13956b0b8233f345dfb490db17c156447f080ef60ae559dc4c9a1528af5f5ffa003fc5d0104fc5d8d0fe0703113e31d49dabcd077cac3993a8d79b3eed0ed495bf5b9c9dd31d74c5bf9125518000fdeb466b239da803c8ca0258003492eb779343cd44938b9690723eb3eaa8071163a43be00e0b525c0f2c29ae98dcf6b47bc2f1c16057175b3c75c6329cefe9dd9e5e17ba4f2cd9dbeb9d000431f2ee954b7177b01d50a6d328bd2af0bfc1da75116612f57b42a166ec8b4ff9fe39be0a7a212fe1ff7898bbafe88f4f8d847c150b6fb736876a8f4f2d006e30c89721ab0a9dfb2c5b3ef56b5bba357ca291aff251d85c5d6e7bb976c5521e87d9a9740aadcd7a3fa070b21678bab6d9c3628ede30eb8cb3df785883eaf03c5192a4ca57901fc20d7bfeec869fe016b1b6ad6271092c2db90453f42da3ad5cedfbc40458b4ab979d482969083beac4e4bc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha4e84f4724a3a8b3c111879170e0fad853353afe50a8adce92da69615122edf1c5db4a9413969a11b2759002b56aec1e015f151a28e53b11458e315e11b79219f9f87891720fe3cd1343acf58251d25453ccddd352c9e7c1cffd47e12ec568a6828265373ef6ebf2a7fe121a191457b6b245a1343105258596a2aff547fb5a7cc497609924b9650e9193cea8633c561c88a0d12a8178bed53f7580b8769f94fef537e4525fbdc595fe2a11cc24c6d4f7f480a613159d5f2bf49ae6db534655cd12f7f55ba94c63f925d5698f1547c311a398207caf1d7699d448bb7e0d0936d857443c387927aab7a6253e8686723ec7ef21bcbbab7b7c784df74f77321ce56125733d87fdd8c41501bf104bdeb8ba015ff6efc9feefaa0eded6bba8694e8e4b383fa1516533b486873f1ee8dc7f6b6b5a8eaee1ab26e8255bca1ce9d00b6e48fcd14ef57ab02a2f42bcf5a3c00361d672ff0d2fbd8739ae8e3f3434627f9bc6e57b796a80bb8d7c0306318832aceda1449c38275ee716eabe24876e17e2c5efe07096828fbca8dc2b5407ef15d4214275bcbb1c0bd4a1ae4f2d725890d0136e49cbf495bd22c4c4fffa60c0d5e986a59f0f797c6eb722f027fa8c82639509780c80dde7109fc1fe53461d003964ecec43eee9c075a7e3e49cad8e5726aa86616d894a0d00187e91f83eab241aac856946a16b8b01f338da2e403729af54e530;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h91f92e573d2dc5a999ba88cf6f8aff0adb840502938fc0f7f20d5ef259edf31d61f7fa8ed9f38552b06a61c8dc4ddf7d7b9f88694277fcd40119dd54a7f3b5b478fa795180f9084c991c0bb5b7757815051901a29bb5cd5e134f5418303bd978239f904392774e3d2d35b64bfd26d38af38167ddbd67ddbdf64067db4b07209647e19529ec48f99dac2195e05a19b7d619d55c019e7fdaf03f674a1d41389f1f4e801530e24a6ae72adbbba37d5b74e4eb543bd54dd0edea8481a0bdd9231f54f22a55e9b481ba835303293f5535094a1090aeb2b6d36ea5e0062602ff211fe1f272bfd4c447cf82d655c010e18cfd746094b83ab604c72d4a9b5ff07c15230c688208f2611cef9f36ca3212e260813b3e1f3a3c855f50294e61b199c3e2ba8c95efd3e4d7563013caeb91b9b466eb72d5128789a49a59d6fa55d07cfdb242d9ac079caebeaa4193d2cfbf1257343e1ee08ba30bd17ec9d0da185434ab0ad275f28a9a20d43c64d79ca3507537e9c1a7757706f10445acbf3eeaaf411ccca7555baf5409c413d133f46c230a11d8a1ad996e97dbad3484b7f87c4fecdda630445cb0533939c90a909ab3050d8b876d9d5d6ff39c2e36750bc2d14467199661304dbe2b765ad9a5fbb59acf554ccaee15e96847048a4ae3475d710c9410721a84557b17e1af2b08d9910078978bde07d19f15b0b9759612d4308e5f3cf2579578;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hbb273bc375eaaf8f820502eea328f757bd6eb639c7ff23fe94aa254520d6084add4e0cf7c00d66ac3f1d98f1b5cfd66d6c76eb89ee0601c6b9e9c0d6bafa10202d32bf149c22c2fcb62f2ebd3feaeae949149bdff0dda3c5b8e67041b811e790a8d495f3934b20bec46327a42912e38fefd173ce5cb9415a4d056235b24ece693c28dec7b5f50861c021a7fe50c6ef4163fd26dfea91c2fc4ed64732be45778816ad90cfbd96208ee9f3a8ed9b33d8f2a4739ecae6cf7fbec05da295be038c893682e8b706d53f30b69a3483c6f51a3ac4eedc66e8e581ad3f33e419dbe6a8e73eae224284a1eb90f55fef63712934cff5e1e9464873b4dca541a14775ea03193302201785710be761f241d5f5a7c40534ac09c5989fd8d9a413cd2444a9d6046b4c6a2182c2a87f1ab80be9a2da8657bd6e310a929feff8923b924ef220ed23b60bdbed7b8c456472d1525889c75bc10f8c4b3de3c818bf09fa4f858948a48ee2ab3813b5e237a7ee2a33e8c312c983629054c8329f8d4324a5b7f1317b881ecfd6b34a1c9aa0b0fab8153faa2bed16f3f9eb202f3be39c46f7a88d7462e8218fd5c0c97f9e0cdfe571efea46aaa8167ad062dbb537e10fa5773eeec898a08bad1d5a62ec0f9e1337d185ae2bc1518b8ee1d66b59a6b4039ab878bc0f7f5fb08569355325f5dec0dcefac05a94eb104e1f30f27589107dd0b198628762d6f08;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3ce2678e4cf0911cd15cbc1693824829362fb915801e922aa0534cd0b2ce641966bea07351c4af945a6dafe1bc12ab87e2ea89fdd9e915123b264b2a895d9de34a02d58fe5592bcc932105fede59991054237d7eec6cfa24ae35912821b8ce6745a43010b128989d5b30c526ae35b820ce8f45b590eff199c27cb760924e2888c088c690a4fdcd5a7b8e8e8718bfb080404d370208470aea80e2c91424f0c1226f93e3dc74d26d55b226861bf8cd58c110fd72b0ff1409fd44f84fe942f9b08614d3f9deaf0da825a4585a46da3afa1f20344c34072b3a56eff20095156025c3079f7b60f8258e91f338274ea4957a6bafaef3d14d2450b6fd423cc1865c97946424b1ffde1fb00896464bd60e30b2e5570da20ad95e6da904570d3985b01bd57afb6dab3c2ef1b15b6d10ea37865e2cf8937792a3fe5251afa5cdbd193d7aefb004320d2229dd43c5c278ae38a284a5a78e3b3a74113ee2adc575ab166267e14b168c83ccf11b86e9cddb9b422f33513fc510846808a25dc337f21e2d7de149a0bbef7b4fc76f6138d0e20de7310c8d8d14bd7a30089741d80b786b3b3ac75bf2dbedf1843c46f57765d2f8421e179ce85a90820a23827323f14f08bdf7b226443ad4921fd8679e8197373123f45de4d0c662def20e1b4aa78d80cbf690f1d10b1c5247491774c8f74afd0cfb9ebf5379e9c90af8c8722f9e03fcc4607b4618;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he312e523a48dcedc75e2a0affbc0b7e36f4e15ac6822d706a9786d9101bab739765cd6828fad5f904669f2bbeabe4494d112310e6a5b2d899a4a90d90448e1651150fe2222d1b2c0c3aab2b9d04c3d6411eb14d3825a4514ed6d13c61fcbbc8e188a4ca5f34c225aa143be11e8b2813bce9eb0d2d36b14a6a887e48c5de8f74027f99b8fc2e274d1e1864adc4e50934431f7dcc00ea39c30c28b57298cc74eba2fde15462bb7ed5770c62324a65622077bf163ad38afb490d007dfc8747e8349662d3c746261441f5b99a0f0d8d8b31828a2a775a8b6e82bccdc6e4fc0bfbae7d47ae88734e82731459a3c602e6a74dc337e9bd0c4f399f9c233954b3ddf547bf042f97e900710299093b9a57f9f024a43ab9689a1ea5036728029dd7d7e5fac53db20899b4882f4d2c330da38423c537823a8663a87249a3d7d15fd6e1d3503202577ffc92ab1db93fa0130bebc512b78bca079e855c41f36b0231f153d39ffd2fb93a7a5eb588f32393ec69028bbdd6533810869487126b87371a6d7b0eecd975db3076926ef8a94b26cde35a121b20bb95d333854e2d7ca08f9e1c205617832dc273eed4a458c137bb0439ea44e9475880e5b5eb350b99e5613c274fd8e5c34ffbd5e132047affd3628d32e9c8cd189caeeddac7a5f72896040587c95c0808250c654469c927de1a9625fe7ef47045d8059c32bc3ccda9144f0c5cd82954a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h14652b579b651470e336c859fb07cf4bd3712952a427fb761b550c3026dd2d1726ac0e3e840d4f3f5ef46289d46e0c2f9efacc993d22075ae8c4076e017d41ca98126a072dfc936b2b0459d8a65d89aa19d8026bf401959276ef8a887f7d132daf60678b8324d08026bf4fc595edcdee27a02239373206201041e5f287a08671d2a44900181d4cd2930478da78d96958ef8329550d1f117cf67cb13ed03a40106fd632e5c906a99ac01b9beb806ebf4593548373cd3a8010eaa4188ae63fac55af662c56b25ac787c58bc8f3ca0b830162e9272f9430940c1215c39b611046a143d938e817498e7fb2be85f38c72daacf3540f7bc3c973a0769411fcd911fe880741c352520b936449e14cf917b3af8577fdc10158d8a971c0f0be0cba99d85388f5d0911b056dad8bef96b40589d7a0c1bf54fa39b9834f78e27ae9790ea15359eb0d0f16f655a9f23b5ddafc656e9a4787e429a5b15c0eb67ee0ec68ca89f0fa1d4575e10ef2c1b44124210b90c9b2dda7182ca27bde9e041f68af1e6ec78051b3af7a27341b2afe2e1575c223d28ac2bff4d99b19928b73cffe0dd727ecbf7eb1466d19cedaac2e9525706b80e2ef9e5b192d333fe495bfbf675d47fb2ea61411c4c4f131f0e18221ef859a490e79ee17077bf6130023ec47374a32621eeb2f40157e6c9da94adc2bc0f6f2ba5df89969c0aac62fe5ed2a21539a337e5de;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd0ae4c809f07a8e2f4fe35c5746c7ca52ea6b6a2e475a20d8780f5017cda1851f71f11e608b5ea53324ac0ddd740b688b99c9596ee46616d897b9444ed73627928e7ea5a73fbf881181d87cfb14c5a62cf2ae18c1487172100fd732eef10f343e8c20c20e4e64d7531af73f3ba37243ce27754d2bd1b09ab1efd48887eb07275eb97265175775f4bc8e1faa29aecb7f83bfb83d4f891112eaaf004f2b9c817d5e4476fed0288817af180fc9952c6eabec2d567b40884693a3ac44be2afbe2c326e9bee37fceb05c910ec6debaedf6039c47905dd038e7645089feab5de0b055ba79438c1199b9d999a147d734316a510937b018e68b10cb52ae6d9e91801e63658342fb8fb79e804aff408859bc49ad4475bf087303201247fe8775353d4539cf187ff5be5545a76d0f493ea7ee41bbeb8418ed79bc9f0ec3a9f04d4e6afbae61d97c984e5a378198e02625c11ee0035ab9c959823d8052e66d37eab412d456fd3701c15533eb0d1aa53c7d27922f5143f17547769cff460aa6e7a472620d7a9d92c59265e1aa2efcb806563ce9c7709fdb147a70eb78057761e9217428d2173558acc1adf5de18b2e083e3a863b3c38f941ae8aafdafe268b131129ae5505006ad779381ed6d5c898f79e6c7917ba72aee956b8ddb7c79fe4bb15d07de992b59d484a84b46aaf466fbbbfa354129a76ef05ec99721886453fec4972a5cf604b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hbdf002b96f57c2c660834c1dd50f8b9edda44c7dc36a9923dc8f6fce9a0689a170e32326c8ac1dd2edd15d86201fb260a6f7c6bdf7f8d013395bde7140461e312881b4aea8281b0503f4c7e76b0a8509a8c78511b18f39d9604b0468048a517ca7a53df68a5a8bc284ff5b1dca1ff3ff130d24047414b77a4eacf0e863edbd9141313f71c6f1c3c712d2fd0245e4a5338a8fedf43c989e8b30d4b1fb550c14fdf037f1e1ea467d4e28aeea70259e92655d7de8732313a285c52bffb5063fb7f3de2106705bbb8ed8329bf488f85a9d079c0372f9fe2fd3d24d034cb023b2ceade9077f69c932cd44ec6295711b8c3ed33aed9032164b16be9f154bda81f7ca74b1cff5203a37c727c8591c300fd89c18b977d020e20776d7cb3e9b40604f8fee5296619161a1b21e428e4eb8377175f87f4385ac1098075f31d1196d0222115cb7a8a67220a0f718791402da78bd8031656f01037e309ecf74ce174a31fabf798cfe6052cef421250a48f44c71d39b10c73a732753a27ee20394fc7776eaab4f747a4f7210d02da2634771f57c64d7dd669482ad2ddea5c21a18d7a6596dfd78b5822924389a977fa4aa57707115e8667600116ec3f8324726628188140de4279bfd63a47ce9f4dd24b38b73c2fd8cef398272afc215dc70197aa29c43b33e6f481c14762fd5714685edeac4de0db62f1a9cf082150ac34d464bebc87f99135;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h15312bc595d15eeec58734f829bc3a5f00984bca9b9a0129ef0dc1b58bf347afc9af55894fc35635fe1c609c07db579b1321458c40ac33a7b8cfaebde90413d6017158c37abbed354e99ec09b689bf8c8d05f534a07cd2267e0d5cc6e3ea2ea4f6031670f0f08c9686141dcc4b692e189db7e655bbcec8eb35cd67d9f7bf69b7abd42dae98fdd9667b93086fa978085f3c204e0bf07056e4d02304d286758c4aa1602d166508aafd01bfe57fdeda136c26760d132a05dce2e01b9e3cca0089ce53e8b2aba985ef637c194ccab3e3a58fd315dfd99cd600298e64c9e27fed2fdc2c99ea2840bb258a8c5992e755a1c35f502748f8044cd26a60c845ea52f93c6a495168a79531cc87e35ae64353366014c8e35a2cdcb28acb940328a65341feadd6cda1108cf1e0bbdcea71f197c585ed91d5a5767359c10dd2fc9a07421cc71ca3bdae33b55159b67881eed01dee03270be1f0d59dabeb1ee53365e07939622ebb64971c64e39fa1a9c484a183265ecd9c5670b66044985ad95d31ddaacecf3d1b42bd815c0c19a016cc7511e6ed31430932a1f5f70b241bf9fa3040114eb1fdb7d30152f27e93b97a168d572da4506d980a66d0297985fab19db22de17136417e75accd1510d527e8ecc42660fb1591ebfd8cacae712e1fbffcb9486756d2bfbffb057590a3b3ada3b2d3d86d16fd5fc4d143924c0a31f0de31118a44fcd4c2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc211caffeb642e086d3c95169351d55d47dc986307961968f58d689f3a98c5154a9db6586ea9076571b231c900d096c553036b9bf799265910f81dbcb2d4c761e4977c4788e00d1338c33a9320a4c5fc133d1b2e63d62c3076a9834f6bef65f6b3ecb1ae7dadc7c7cf8232de0d41be64c201de88c0df357a16900b6862416685261fbb8cbd3818462c0fc39651980375a3f4439c97cb20b6ea981ae3aac13cc40249ee90d97059105665176989a17ed821f5dc6400a526c5ca3c6240d866a84b8e53d3faaac605cf6bc45168ce9dd41e1436122d9f885e62b23447517e1bc5f45fbe6878fdd20be4a32ae2bac6e1586d09851a7c329342969886926accefae1b31941f70cc8d516424254eef66dce09db564c6d472f8069812f7582fc4866de80f558d2659fe108d78c57ac5bec7cb7560764ee7c6a11953150039e939919d625bea4eb7cb377525600e7d8d9c6e010b4c324e9d1d610859436f3d8c2b9441c23b4a854e974bb4003f70f2cc384b2958b7fcc119e7914c3dfa5c183e4ea8b6c29323ffd173382d639cda27239ca94972c174307444c43ef44dfac045fd6d01348b7ab91c57ff8876d45c23d8c83e6771549cabf342559fa4e5b146a7ef738b98b8923e551d60e2c3bd57b745f8568fb037b26642fea04086ab3c542ff6d928ef97d2b3e326fb85938f548dfeec2b296f3604151cf0162a8f8f14f09064876280;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6cc2b0bfca350b25692fd005bb517066e05ff85d811b4837b63b5852516ba7a2c4e9b977e1f09d3abbf6453f6220b90c8c006e557072fd23cc24ee31bb9e5db3eec1f68191d9a4efaa4ecbb8f37abcc91b2941abf0ff86fad98bd8e1a5ed265bb4a6176b751bf6cf4f5708c09f6eb72f2646d31cede4f847cb28140f7a08ac08ebd2cbf27e63bf7f70058c0f8a6b60c3d02c56e332abccf298a428657ebecf65e17f6f3a9e7ede5aa9e082a548e4ac9238f86eddc58f57b3326cf2da8b2ab4fc87193e01a5aa6600a9c7b50e3e28709337e206c0d7f48011b706493b16cc52aaa6071895f77b7f5176d1ea15cfaa6c32fc4b69c22516ed4d5844c30e94800116664f289bfcfb8b8e1538850fdfe478d353056e9e913d52a2328f22ee8fd07c5929c6d5bdbcb5e49204a3de2c4fc66786a382780a5a94f753ad8b4d76c422e6e3dea92a4fcfca31fa797d42b994e8c40382a73553c58f4be687fa3910892436a44234ec6d927d94f2c4b73628bb96ca2a2fa84b4df9fee6bbf1a06cea34353b53b7c739c78aff52ba5170ad7b74942d02dfaac3795a6644755c9286971ef5db573bc4ba519b4f048f944c4dad9d694b34c882c2b323638520d25f43fca2d6987a98165af4f27d780fd879c608fc179daa63c041454205ad070e31d3b3434ae45773d69ff15b51ac80177a0cda561ee8a0d6a694448f3a4382d68986c216bbe3db;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcdb2fd744cc5497c7421970a305b6496431d9d1f36b7307674b74ac9114aee067f71b3b96c532b2df51e6e8a34df87bfd62fbc0cf9cae076614f5ebd543afb021e6a92b748a56cc1b3a48bd0c63545a86e5feb7129e4a6c35bfbd7b7d74083800315cf4d4bc4fbce3ec1f2abf11e1e2c4fef9569b5860d7d1f64bec2c6c52c586803b6f76e42740153c6e3e76a62ea248cea6d0fe686dd575cbf6c87c920d95057c075d3d2fd5e5b576122a8d5175055a7f3ff4b2961ff937607c17f0fc69b2b6396f0013faa6ca680a02aeb3f24bd9f51a571bafb3d0317c99b8cedb0fc6ea374b559994202680e2aca8e5e2aead1f74e1872eacb68dbd2621fb10b6e4fb6e5ac54e3520caf4b05e36d83fa485ecd3b949a64cab8082372799adc0ad5fbe5460f3984d529c0ede172a111cd4f498ab1a5499bd1be600183247a89263419ea4461fea2b454534567208683d8377028d90121defe69392ab1e937dca98246114b11ac07233c8dd485ba3441a7ad3baab01a4bcf11644e12e2c3ce8793a48d9902a2b38682088a96ac8e65d74ffc1f5c6a83a214c472b24ee92107a69e1e62151db4f72f2adfc2b929e6273012bc88982429b9fc5591b69cf838d3c6d9cb171e1673a13b77658e019da82287d3afc31f176ba9962840de95539cf10a5aee0cfe5a65c6184e1acf8f9f51b9353f4bebd25334290dbd9213a3e6407c4d143b030c92;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9c95ba955d79b965ec88cecd65bb7b3deed66a18d3f17acb40c80dfabe714aac303f30f532ced68a5f7bcebe215944f8e793599f95502ba9c432a4a9f00b77aaae53c0687e570f5b0c9fcf295f25982d6718dc9d3597d28e96a8e568d8ce747eaa1978bb43c4bd958d4fd767f8e46114ac0074bc7b86e0e3d9b4da4d396aef3bf3d08f871ddc4f4826169c5a556bc046128ad5db23c9a88d18f84ff7805402440be6e0673f2482e8ab0b89bf00d5930b2ab2e8e82ecfdd04a6c8b445131c0ca057d5d87393c1564170dfbe6dc1d784f2278c85409f33864c408d338f4332710ad914e98f7f50bec196092dcfadbdf70924263e1cfeda5a003056491ee771ae7cdc6d2a84b7fb3fa81ebd8bba7cd802e15bccef0ca8797ffb42f9f48ac1d32d2e5ca28f61e4ba2e6f677fe4e4da1e0aa4bfba09d0aa08f03334953451b5440cde1116e75eb98850b7bbfdf8a801e2759063d012b4a7d3cb9e558cfbf9e9975edb70975190eac5f9056c03705ed27466de021cbb0fcb2a0cb89f6cd854414c1ea295b41ea75bd255d7f13b64991ea42002fd088af2882e84459431b28e1862d7699cc46a80ad8f3626f6fef609a6bf4bccb163fb8c8a0a08c58787038dfbd09f78b94c16d3a807608ba5ca52f1d45bce400a1eb65fc18e2239f41ba0270089ad54cc85a606e06249788d3cefd469e91c7f3ae7d32062d23b88a2c5f6c73dba95dc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3c54eddf31604326722c6d27cd36edcb81f3457aacab6c705ddcd6257b937211403a2cc86598444ee04010c45ee180bc030c2edf07d220c3e4ba8f90ac4d921409be5b94ca7ea010773e8a5dcdccde0b704f3e5281551be0fd2bea840d5a0a779212f4babc072efcaaef819176bde74021d1dce5cf3684ae5b978d2511a4e52713f8167542f44fb3d84990ca1f452fbbce1a9eae50d152ffb076c9a33eefa548971b9fc432e133377d757f3a30130b1855fa2779bd6b278ca404c0f5b53fcd6b35eb48d3b437c5b8c207b590178c2995dcd3750ef3f1c60669bf7cd6f9e217ab2abe5523e9cf3bb4603ecee89e905e29a59a6da29fa70d024c42672d510e4f6a8336e5e306b908a080c4d17f9798ce445fa7dd3b2086b4b7c96ef1ef1f345c4e54bbb4f61a57f3ac315b4e1d3504a34ce9187b9f24b54234066f516ec45f4df94a43af2d7d84da2b3afa27b2fef3c13eef69a0b9e6aee65bf05012eee0aa730179aa3012409062ab187d66d94029130a423c1b9d4f723962e58dfbf907325c40a98bb3eb945d94a493ce5d973f17e285a5ade0780aadf5f835017f98d09a89306ea7b872b12e9c718d8ebdc175fecd42a9c09310bd6f7a45ea32218a828bb2cef23bc15e6013143cf07afe50f4cc6f2e84d03404f047d84a96f12a2b0b33e766be82f436ba90b9fe54facad75967473743ac847f838e366df5c087fa541e783b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he5e35a1f0c38ecda0f6646894c5f19723cf32a04562f7e92459f83432d6e6c052419c15e1b7820028e91543f845cbb3ab52000e2c4bdce1c0ef773fb924c190a7a80e1b338bdd1a9633996cf8fac5cbcc1b4aa53a08d1986a420e69926b86a20c101ce47a9362db343eca183548d8bd573e7bcd4dd3fff8fc17e7137de7f95b5dc541e532ed15624258a89bf6d3b074e3ec76e489c7f19cebf9e1d6d55b202736799fe94da10fd98ed2f79b75f4fbf06c274e7c976379340bcec6c7cfc79a334fb2e585931ccde97161f2262496e171b3935cd529bbdef56f399733cb16ca5a2ada40e89d21e567d4895f1526f300f3c8357a9f10b5c86e8da310119fd92d2b1a73ee8e3b509b21a01ade64fa1853067d70d19fd4d1b47fde49fa7758f49b9397a00637279ef951dde5c81d0285fc833c4722b3af727f3c25315081d6b08f196e3cb35ca7a0655631d7164fd73d65fe376c259b9b8801db137f2edd7075e4b95a8157127fd28d7dd27ad9c74c5fa5ccf2619e68f332bb97eae9e5f4a02ec50cf37db79efb99e771e5f700cafbf26a13efc252b3f957b927d3f5c9f206720c5b6c19b1fec7a79575fc45a3a883664926bfa05fdd3e724fa626291191f53002960399fd9bb28e65a1b2866c5373b4bd3e313c7b566ce5af537b9fbe6a4e46c2add75658e13e918cd9e053d3b4d879ed5a450e64e07c873d9c61c3764301b84a5d1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h34258df30f9fa1bac9c265b3f2277cbea8942e34926b8bf19cabe1e456e6fe2dfe337286fb7a59aba94e781511f5ad95dd1ba37e17c126141ba1bfc038171a54509e05fe9a5274d26babd1056b31f0436ab4cd805800a31e6abb0512a2397b631964357807fd97660fe48a7ec0aa70693c555dffc557d02127de0ffd43bde79d0c375869b1363383d4cd66e27e74209bc4bf59a4dd3068bc705f26fe91c355cf345b19041b18cfaf742b440378a651ffbf36555628116a242cd267baa941daf14d30ee99c4df2ca9ff8b026b9c1217f2ecfaa1c25835d16cad246dbeb63f0f1e82f8386f3073c7a3defb68fd3176418feb7186b8d24850920549f7b7e1fc3fe966763dba6d12cacfecd3471682e27293225c257dfe4b30eb748458340ada85958c04f8f9b89a6210a2541b980feab12714dfa665830bf7af7fb99ca1bab37df474d37ab6e42d3c144c77bdde78b58269a75ea22be039d404f8357cfb920b4880597f97ef5996ae393381392f13c5ab2e1a8aa8cec616dc3d197197ed03646f5c91c7fc3de670e969b59d2bfeb988b60d0bc142b8e8c3202cc7b16b03df64b548ab7c7f52eb05ce72c4bde62b6afc3c6510a799ef15a453274d6bc6dda3aca909c04f4e97fb034480cfca4d20280e98fa0e6d0e0ddd7acc4d7efe3898e33c2abc30d58840129fca2db9f5a05de4ef949575f4d6c14c0b7317f8b804c2cd87b89a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc545f2398c07bea36e449790233fd076852156d79d11d66f47f24523f696d9d09c4ac6651a668a4726b72a801f70f54b469055ebc98e0064b557e26f05b82ee321596b532fa837d39602f195ed4e6a4b53ad3783436be706e81a506c42048efeba7b4a781081ca073259be093b5bf54a88fc56f486f426e98737d8304a6421be061f57f9aa042289c439b67e13a87da087742d2088698cde01584eb6e152e89089aebf1e6c9e63ddba4a261a739e58453a0a634812010431a2e359763238c0e9b6c7e2e2ed31c15d555ac498164024850f590b28d2100a1fd432ba2ddf456af7eecd4a46d70c30f1b59aa6f877d229f221a1f6433e67c02abf4dd069bf2caaa84ccd850e2f419e8f085805d3696216712f355dc77779de2504194f64d8400e512330b224073586366d8c2c61ae1745aa167adaa2f3cd1054ddbd8908aca1d2977f1970eb246f9c5dbee1d9654e5cd197b591fd5b36290ea9815529d31d700fc328f73dec7c755d0f5463892327e5ce56c572598656365b20c4aa471985f19387fa777ef3fb6234bc9f5a01510708ede4da56599f3bdf195c017414e00ebeea721f6c1e6bb87017997db3cd898f06936b85c208a9bb2ee0d17a7793b0dfe268fd3b7a8a224a6b7dd9037208d8f28f5ac92824f687dd073a7188db17f9c08af0c2b2e2f15662275eaf757d32c9d62fc1c7232dbd56244456e206fbeb1601b48cbc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6dc4130cc7c0ff47d5b86028f04a38d54737b54e91c43fa779a6ebc44497d06823847ae0033001eb8be70358d4584636f1e591e6c636e93a72d90fff62852f20ad67ec013742745f065073fbce2e33d87eb24671a65026cfe6da2c2b4534558127cd8584520489f6fa4780d936dd8388679d335d0d413ce746c083f1434e757af27e5f4d62bed3be2464f41ad7652c597bca6a61436c408f2678438a00c3553916a157e3dbf927bea49128b7b6c266b952bb6bc676c9f915d407a63667c6e86b0b1ffbc8d3d53416f01596ccb5ec70eb9f0d0c67d322c3085ff899600ceeff9ee81b9394dcd252ae3f47c16ecbe0c3884add72c42c9376ad5f973c0d6255bfe473437250ca39630acac267ac16cce64568fbe405e3132d225a2cbe76cda17182b79611d0c37ba9c705b7d73533c16545ac0b7acb6563990a8261e8f79cd7c33e9cc7dc2fa2953ae081f29108f4b15340075da468ff4eff75b1e13aecc82be9cab5bd4741b5afd885642598db5fc5262f4fcef6258319eb27b14ee5904b600f9f94f6bf76fba1d9975f891fdc4564f0eb9b9a6780dfce47265a31d35424496662def223b6dbb30f6600ec92c6ab5e184c32e9b096597fb9d74fd5a1e30aa53b4dfacee9b5ceb3d8788b966baef26ba92b0923b98c110819969242230a4aa8b3e3c699cecdff6dc428ae14c7fee65bb2499483144b9aee366d581e56250b5abca1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4b22896b9b35792052fce58f7abda725d9ca10e7b931d0748f36617da0a47ee2e5cb9a108f9dd38bdd359e91bba321976aab24cffbac94f014a7c456b0009e7bc666638c202a28e25fd63651952664ed5cc18c823456d4b9c03225d68b6a8c6d98cb0dd4af072e83e8b20513e241464f2d4353e34f561bf53a23610236f44b3a20292b5744cf3dc89b63e4032aee46ca8ea979a196a6bb25d274a97c1ee3985320a9607308b30243efbc9f50f0808eb087dc1b9e0cf4e0c2172743981602d89d10f378b04252a753c86ca3bd873300e299e8ffedb6709f388523447fc4a5c339f9c98be43b3eee8461eff788a62350cab2c49632cb4380c7b138122747d86ed0ec213cddb6d882de7b9feba335d2c1f777718f06945f4a5af9d3959e29ae6626a609330f46fae09f72bff2917f162e146d2ec157d2bc3290e994d3d767f148ecebfd30342cdf26de11779eff46aedd467908def94e73fb49200ccf75394a8fc5e761ead33ffec09501234a0431f142badf4bd8d8ee0a3b3b0f59b55b464e81c1e5021002f425f17217d0b662e8488396492962827ae94bebcf20a2635b4218e3a18276d8c951ee677566995bb8fa5c3b2e83c240ee29902d17fc4d2c0f3464b44c34ca6f2f57388e07c0f4e389d89d152f6d9aac4868720c8f73053a6607d3dc3b4d7c31f29ac88329aa5ed96b2877125225be96a36f71595078b796ea20565a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6dfc02131c9417493867e6ef4031aa43d748cde8bfd755a1b147d66231cc4d6a2d7f8820c4955d8f4716939342cb29cf8dc86205d6f89e5b7cb4894d7bb2f6d011ffb93a0b8860a92648c9bd07ccdadc9752dd0078efe0e3c5883b2bd7aae168978587b021d3ffa1e943325bb639492a6b64353ab01108e595d0aafb35111d1dc684568fb8e66117e2360ac4a43d98f866c74be4d5ed2281e09818bbe01bebe2aae60c4f7912dfd367dcb547893aeafa1e47a9ebad29d34bddc16ffd945aa97ccdc1a1906636dbbbfb791a55a290edb2acda7e8d859539f90b83c26b25cd63c233f9235efabbdb968d47fd494fb4ea62c4fc90a100b32eada9c43da97800640a5cff4859dd33a37d5013f545785c3f230365be65203d69211f1ddb70b17b3d45bdf0fff9e81f6d543c4ced70c25f7a40557cd7a98de8775aec6c65f5839249b28489d9a57db4a9a0b89f41976056f0f2a0ffe330d5a8959f6f629f313140e3ceba45d49f9532abaa3e9fa3d8cb3f1dbae82f34f749dda6786523bc697f7bd156d5eef3e735f77441e50e989c6f43cf4bcfaa680fb43f16cae219913b74079373208c6c42c3e51784c2c324c6cfdfd3bccf205092143e06de8b971df6804600aae8f31de4e4bf66e486e0b52eb3701298a7508d89b2ff149703ff1660553ce6dc02538a92543e9c6b1081581dad3cfe21602d76e130646ab1751201716197146;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he9485b9f80dc967ccbaf36a74c8e2070653d631dc516f045484ccea83d682e67425b3962390f004140af5e83aa08822a09638226f040a2ce7b2a1da8181925bd3f731464f91fd8fa2d62febf1ca38d0a0d904134ac9119a353888d48dd758b1b2a7e6b0ce8ff522550015d875f9e4e72a9aa18049a7ae757de79e17f4ebfd435ef4ac7c25fa126038e3dd1b12b48cf9ee3a722a4df90ef2589c4dfc32a93a249761bb22659ab6357ab3c1c6651cba3167c5019a0298513fd8321310e2cb2ad32eab0513c19d2d34d17d26580dc26c74fc87b8c2f9c3696a572dd95d587ea7d05c0ac637c426e8bfaede2532a136932964db133ae18cf097f1f36ddd398f9f878d58e74d73ea9bfaa40092410e793ea4186e067179eecdd22516095ea11ed9f7108e4278dc77e182ff7a362385031bcfb3f89006b0f596e48e471c6176032b5888f39b42193af6ba1a4dcf424330b762fb12998f2f78f09c714e7ac0bad3c558b718dcd0838abb74f75d09f1e9948ca29db0eaf0bb52970069fab843bf8ed44d7957810090f10568fc8e43aafb72916060ea03d2221d4ea034eb764c2bf29e6e928db6ee0d0d74c0d87ce7c39428d23b069ce4c7d7afecf522146fe9e7f0cc6717dbafcccbd821f48a2dd48e071e897dad261a1fb5b4a7bb8e087ad3ec5a3b370de8e147bce0d284bcbaaab6909c8bd9a8024f51d8d6143fcf9212740aa698e14;
        #1
        $finish();
    end
endmodule
