module testbench();
    reg [16:0] src0;
    reg [16:0] src1;
    reg [16:0] src2;
    reg [16:0] src3;
    reg [16:0] src4;
    reg [16:0] src5;
    reg [16:0] src6;
    reg [16:0] src7;
    reg [16:0] src8;
    reg [16:0] src9;
    reg [16:0] src10;
    reg [16:0] src11;
    reg [16:0] src12;
    reg [16:0] src13;
    reg [16:0] src14;
    reg [16:0] src15;
    reg [16:0] src16;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1655443381b307fa36365abafaf3390a9d2da3337acb0d414b1ec17702d5c106d1f3fa006;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11b6a6084c0ee78fef380f64cc740c34ae61676c47e8efcc3226355a700d7d5da099cdcbf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11b8208dd399e032b30dc1eed6b25668dd11e3f8a7bbefd36ef5a5d294a0ecf0b1e794d07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15699c7a589b0f3d74e5e72398c7dd812313e03d3b1209a7c081e8f59edbd3612fe1ba8bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h523ea8a5868406c3f1f74c1865277ddebdb42f5db317668f8e350a131f5950b0b6f7fab0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18c3f325b3c22b4d0a10273c8e595117ba3cba59647c07aeeccaab5e10ded9211cf1fd0f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11314d8a6e768f9842740c97f18ee5ec1844ebf0fd7ceebb0eecf4a6635eccb45db830b9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h56822b65a8d76e97a8a69f90a93bb7e57cc6dbdf9a212bf39c8a5adfae9d2c5b2b20856f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h919bf5524adcaa795c7e25050488c07f81116f036fa11bd95ae6beff157cc71007dc4583;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbd1c554bb44504ff7e68bcc9e68698f2665e4db80bf4d370ab86c057781d56b1b04ce346;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf4d2795f25e009094ee3dcafd8a59e39e6a5aa6a80ab00ca4e495d8231f08404db851a04;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c852a542a859e76ebab65b9c5d9316dee54ff9313f75fc1b823ad76b8f3ce09dfc1b62b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c47272fa9c2876271e85f9a2b5e8929ca78843a7b75f7f91c8a8094875b8b58e5f1b9c1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h67ed61f5b7e86e6cb644cab23e7ab953d4323ff3ee04bcd366be2304e401bf3bdf19508a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c098016613ea04e0aa640d3186bef044e141674cf895d029118918fedb918bd10fd82c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18f09792d9d38c0a339625dcc0054db7fbbf5b979149afbd945c6bebf9e6e940bb6333bfa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb87bb334a52a6d121cf68b0b1ef68ec05961cc71f96a950a89ed08dd36851f1e7543d471;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be2f8cef43a639e3aba1f4931b031af4a76bc174c5507c5bd607ab1be8b9f2edbd17ac17;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbbdf329df873599a277aee4b17101343c8a32ab9a315178956cec630763633fc49e591de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12e22e8c9ad77303a5af72d41917a611033614cec30bbd5cbd4a578a0b31c484bd3a4ff4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5fccb3eb97742b993e02be14e30b85da7d551eb7052dd3bf63dbb938936babd249e83d0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189ee97c13d4f30d755f3a381f112b2a22ffa54d5088da3c440d8ac87fdf7886fbbe4f9cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c69453861bf4f9531076477ca24966e19c4f4243df3982d2c1a5f3579ec173edfc3c3aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c72573be092c67894a77e61725d21336e0ad8af4ce8789c2140781c84e7d00351e09214;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ab101e21e22559783efe9b66828c09b77bf336615a7182eedd133b17e3fcfcca6b4f3af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h190032d9da4b1517c409fe9bfdb7c6450b398225c2dbe248b7e07927e991ee2840f74a1b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2f6560c5ca68f2d8b1ae39c02e339bc103d50cd8a6c141a602262fabf77256a37645a71e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha66fc043038f12c5c1ea0d602c2eaac88201528608b65a1a7413959f119c1f2ffb9c46ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h97f13c7b796fe96ad6bb928fc4e69365841a953b722ca8b1c59fb76a7e3f75e539605552;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf3700ea6c84fa3618e445068dc1c3d4761209943b7034d1a6405a3e08d7470b35c7aa0e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h93c83b0cdb202cc61b449195356ed8e4fc6081f98de4249168beecb81c7fe9c21e7fb4d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae22f96710306bba2de0b62fdb10c27cb6a437452e65af9edccdbf891af82a423042ba71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182269e1e2cdcfe4caf9359b9247dc3adf255beb6a0bf8bbaf4904c4beed0b6f623e7cd63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he9fed42ea7b0317170af35d363ec7f28bb68ab9c140f02c254de7cbdf1c2c9925224831f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab8713c70a0abb82e669b4a7fcf25c43df98e2e09a0439b70f948bf0b7578199ccefe37a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2841ea32b9087013d1649b188a087a73a307859feffbbe5aff3eb81f6a1d9211194f432;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf507917db4044af7e2534b27baab469b58ace542c2aac92af275a3720ebe543f017895f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4431e21397b1f0cff721de15dba8b0bd1cce49a5b9756fafb7351379f5bdf4f81efc30b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h139ddfb6c70a3d1b466e17e6dda37a5768422e610a2ef4e75ab114e625bd780a168375c1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd2a4dcdbfb53429b81259f6fabd42f831958be94980df2d6956b01bb515bb68e132bad8d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc35d0cd6ee01eafed5a612d40f06476df4be17b0c94d529ac4191178094bb8517d157dfb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd2b06c1cf3fe8cf7b60a7a62661799f857fb2fcdf5631fe8c2c752a663bdf4e0f5856009;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c238e66a152f90a14750741e85c7ecdd786e1b2fb9878223ad92c7dfc801956b05f4e131;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h35a7ed80c9d9eac726c97c093ba2badb6a6c2ac9d3764cf5520b521aaaf737a96fb751af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea4ec13457b165bdd1bdc88be1520a0be726c89a07c9111797eba68b44cb56b1bf5aac58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c9ae7f1eccf0667b303856fdb5046e562bda492f4ab7940abadefd7c62d7fe837bddd68;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2c54c801559c7f2e2158ab801127543d0b814e6edf771934c0f36f27a61a525d342475c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8998fd19bf7e47a8bc0df6cee6a03fa38b5a7e7ac3b1d4f128c57612f8721090ac8ccfc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d4aec633f4ca6c3da326b7d7b7479a9de068e46071f23ad5ce07426d4bceef6f0373809;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h130a00152e4126a500849b01920d09c5f9e29480f08b47dc779d8ad8ef4f21dd1a9c6e4ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2df3ebc2f38a0f0a08fa124fc40fdd0375fec92e73d4bd6e33516843adaec0ba7928580;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c39b8aabb4e88569e780f773c9f49ce28e8689b13342111d02872676c177f61064cfc568;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10edd42e4159409c49b56d15ae7543034390fa88469c88545cabb530c6317fd51ba184302;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f05211032db8218be2088c49d593aa43705e63b9d7b3c2591a2dbce0dddb3a1524635575;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11ffd1c5be300cf5057153af7489c4129157ead83a5aa40d1d52d17c4d7af2cc05971b826;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7233a367d9a37095d400924c0a125658b6782b179fa813cce10859a26cf4cbeb98355ce7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcf062a084ddcfbeb4b0e009f047f363e0a89a7866a7e31219c65ffb0e3c1a95f92aa576f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60666c6928d946b7a5725357517a3695d7a5d29fba9b2585849047f1b4bbc97a90eb6201;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h80cf70eebed045baba75b0a756622eeff5ec49fc4aa08e15e3b6de801288a3c2485e10db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ecbad80bb72d9848fa706e50c6a339e9cdf5b38be0e1a60619a4ea9fa9a17967159aa6d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91d936d4cc5880228123cbf508efd90b26ea61be68b23d50b3ca0724be26e03d56b098d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8f7905c2b0a3c32bfabebb12e09d6017df6b03730c6220d1e7f330f4561fcc7c998b23bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca0caadd55c66e90a6584d02d44b295dd0fd4aedae9a0dbc60ffa3756566bb30f7537706;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b9ed564a1b00ff253ae1798c40d86258c489feab086613b186b460f7c2d4d1564d656722;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h97492b1b011abf6a96b12d40feb4a9b6c0c8ef2a1f6d617f629e407589c33bb9058d2ee5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1af14c0e08bfec167e37e0df46244171edf424b4ae9a4e1285d9e4dbd715b71d697dda4ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h56aec1b493656c868ccb6b955dc1348c394c753c0e0568b790cb4a7f2fe1f2c7359d0ea9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e4add21d59bae2e075a91f33dd46c76a1b13bc2fd5973fb45c81a4d53a0ff7d61859b95;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55f97582152ef0ed8f7424d2c1fc7b52f92437cd84f64d0a72e3a8e6bb92ecaa61ae4b11;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h30906437d464c0cba292daf1d955c06ae7133ee63e0ba33d5763f3575de1559a843bcb26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'had2851c4d3133e7c74616588a2289b37383bd71e07720d326cce9bfb953b84e00c3b04f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135e098e267f848235fb5308cadce4ef7bebe23a3d6272f88dc2b96dbbb792a1748fc338c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14356094f9004b6b9a0f4db318856814fb0449fa39090f7a999fdd2fe6887e332afc54b4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7de0989328fa1de2cdb23eea214c7a7a799432c677111d99585cf3d0a8f44b370d1a35d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h266d118ed79d2137f948cb098ec7d527e576023719c28e22237ed1b3cfe33aa4c2f5c878;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8fab26609548317386685919366b4f13a931da13cc9b3a2a31d9202c21a2213ee06ecb67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc432065c96d9089924e5c98cab11999c65552c69b8059a9618812b28e149d652e6e622b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7bea9f34cd7fae71be4ba04723fa318a8c5f1ae0c0b288ada989cdcc6ae1a1106e147;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfaf465a2d17e7442504d65c6d9c5228beced9224b226c8a895210493858b22e3a7431eb0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16ac92f0650e61af98756a9e1fd9fad04b7938940fb8dd862b4ae2e8dbd339451c36f81c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h127ce51994c9660b03091aa90757e782fd34188d08620ab342384245499d17cd0eb40f07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h185d9aea330969c84114952e766e5dc1a8892ffbcc4cf53d3dd7f68ec7272459a419e987f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a6f5e35fc8d8c878248e3ef6e2a20108894f63ea15141794643508b19c445c1a5168576;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb91278c918d6e9136cd28f61d7a74562c761d7b3b33bb40d4db6647ffb5e113a9ee4452f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he56b600dbe67deee32c5cb4fb7ad4637f127c416609c1470de4977304f389ee07d5af5b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h111280e8902a0fb850223e99e6ec06a3ecdce36f0f6597255c97e274f89f27c0c734bb8ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heab925491b3eb52e0babd9d09ce5e24f546bd7e7e8a818af4bb6dad156fa2fe1d1e663f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he6396e3efb6e45d17156d501517eaa623f57880cac5a9e40946a9a3183969c13f89a2e45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd3a0103ad173d56a56c6a0db588d33eec56200c5e2a7fcd78ea40c53b51d5223e40778b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h45602a5db6a600f1fa23437debb176287a577f5e5694667f9a288a9b973deb60bd5f7549;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e954f24134ca10b38e18c392872ae33faa8d116f45a236a6829e1358ea4bf30c5cd24f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d021e692656ab705baa9881f32c96403d8a0a12adc09322c582d7a38acf02ae3b895a70;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h159bb51737ba1c22dfff8770bf87277448725cc2842f102c5e44bf14cc86f240f3bd9280f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h47112d2c37874bc54db6530331324822230f773093060aba06eb9053bf047d2dd244eecb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hadcd204ffc66857c02f9332d3b04ddc00cb850fb299aae463ad7818ba5b7c7340ef8f1f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h37b3a90a0cebd91b31e28cf23052bfa890e404b8563a1c7836161ada05df5f74399349a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h150be9aa210eecae32d054ea358fe8e9785fe940b84a56069295691df880dcea329be909e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'habf1064aa1bcf78feaeb4002fb97dd4a674afc2eabfd85d5e19a5a3feff41243719ebe57;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f19e07c919b4ea6477a1a18a610b4574221848bc3ed202aea30a51afbb367620002cd84;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc2085041aba8c219016e2fb453392e8b689fcb4e008f9e11d42abe50f85dc32b6a053110;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2ab3231fe9b0b5440d815f2982d4c99c4e8a5939393a5ae47433652da06245b6e101dce7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15dbb0f197a93751f9dfa99e9ac6bfc1917eff18cd04c1b5c577b474a6f77145b1de3ba8d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3dd3e6632a93630a1b68ebac5ad11f02b651adf8b78b32772488f2c9e46f204a8f2279c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf03cd1b8e7ac1c96d21aff62ee8ad6f9876f85e37b2fef0d7a7a4b5b9cf41cba9db043b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189bc535d99e2b71e7e7e288264814fa5cb009c39cb0782b3df34907e43acfeabd0a2c993;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a70a687b08eccf6c4fd37ad3677dd7ac3df687a4b8b9d05c3b8226cdb2c21a10572fa66e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1322ecf29ca21c7b149a870847de90d04abbea1345196c2aa3f0555123ce38e75591db5b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10e84f5a537bbad6c0422596a736bfa6949e03ae64dc1e305a9b1bc93bd57da305595b857;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8770195a9bb11fb3d637ba168bee39dd431fcf12298e6250feb8a717ced9f90dcc59113e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1581ff99feff212596fc8b7a01d815ac5715c434bb323f054f7e875994bb651f1b6ec87f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc7e50cd924aad6dbd2fa49d6ac49d5fb9d35858b6f72750c3743678c1c4d07e489204b16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'habd2940e9137919fd9305022cd221e52fccefdf0c64f8b6e7636e1f5bdbdd65496c223c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12cadd1b391e13c15ee7cd89bb17358da1dfa14be71786d4f173e9818fc49a0653c7b43b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a2fbc4d67632fdc53ec02c809573d2712dbba8b8c222a7fa5d1d1de5486caaa511b71ce3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h137d75e549ffd65ff898fa44070d7267041b3fba0d92e83e9d7f7d6b12cc6d8f5b5a6e7cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d31d0d3b90192126c587d54b225cb4150b9d9a55ea12e4f1b075829ef6b049d8393b3573;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e6282e2a8262ad096775a730d915d6bf0d666d0ade34d4eb5aea4ec6e44c2677b90286d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc04c9f96f6dc87b73a03191210d58ee918ab9d1895155fd4f555feb61cd214d5315e04d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf0714ee10f8b462fa3b35c0f1f4499ba43e9fed988dcba0db33615712595db51551570f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h473fb5e69aae48641d1192a91da23bcb2745468c7572985138929b28c9b495ffc1e61c69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e28944cba92dd8407d0a8c600c85745846767953c4b019ee11652ed22eb05e5bfe4df98;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7500e54037ac359db4f290920e99e018435ad5ca73c3b902d1cc4539d602ae838d9f50e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h281ba26fe25002339401bbd86d29a7e192259f0659bf604a8ce66a56646013142a56b9c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87ae14607ce97be7fa68ede9f8953089abfc4215af1040baf305cda44846062d7c5fe124;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f72f3421d730610821881be9f27c672b8a92df93431a4e63f7b42942ea0d1e3ff117494b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ea60797dfe59f40cbaf3852d9f9bbd951f18845cb6cdb7db3a2a41c311164c58435f0c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3812aa9e6e9f4bbbc675f1f8f20a2758525c2ff9beed682f9298ed4c5d1bb7eafc3da9cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d03d70a942eaef709cb0241027128cd0a9d769372a202626f4dbb95d3f9b141e605ca19d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h159b01be43f1f96d9d873d6601374df1d579fa189a8cf5c8d888f280ed3dbfce514f08e2e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4a1acb69251005a70bbea4ef2e1da2deb2974a4b969f535e87a84f0f4bb367eb819a96ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hacd4ca1ff09d1f8cf9682ba981ddeaf759ddfd681e6c56a0061881734a25c0bfb2b85c56;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14af48e98ca0828e2624ce473f942d06fb97cdbb9a53d17e9dfb12b77252a5495d64bc6a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha1b687b0765aab5ab286f269f7690d3a4220b920b2a8773e5eca5c8d618e9671e85485a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1df5c9bfc7c7feed26d347f2933c574bd464287216362db181af8d137d3661c19b6d9ddb6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d4eb75bd97a558b2b83c96469c54ab5a1f10a0c6c5d0a7c6910565439950483e8c75f8d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5996d286f445a960609ac28784343f1ba56a1fe73961445072d72808a93a4a750d21284a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c1abb3d45a7abe784593f3b443fc7d995404221696bb94fa9d8f4b2f3bf17663fd20a1d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4bb03fbefd17fc57345ceee3e039779248c01297f560eb87308431e06cf852ae8e35e46c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b14d736c754b996394e0c4e307e6f2550dd09999bdce8efac771c645dde618a7fcaed5a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50f49fb160c17b55aa583fa14fd0acd62626e155be8ea58a91cedffb70d7a6c3763c28e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e7cb94c8c8a772d58e9997c45f391ebe7b32ed31e3f78840c33b863c610f97a75aaf0d85;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4ea91f3b3edf9c2a98f83c53aff16d184c3c9753ea207e9d7efe0ca2d8f4e4acc0cf26f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a00cb1f8a2afe56bc22fb0cfd264dff4bb0bc4575c6f9335a4fd81b03a93a8e6ef21dba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17b2c9ff70ee4dbdfc2e145f6cd6e28051bc76761c00f9f95f1d552dc1db2474da2360dbc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7837e531bee6ddcaf9c025f4ab5000b4f60841e291077ceda727b33f1c7b0abbdd40fc3c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha22f065d5b66f4d0e15839f2d5956491fd0430dd78cda171e929743edc4accf7d3733e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc3c05dcc762a3c97227124314067540732b28b3c3bf26cc713c2fff187f323a92c12ce67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he136e970bfc85d76ed44530e44bb5894a9862cc58d2b132e01e2e74eb6524eb28abf98f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b0dfd570f00b4143fc8d00903a6d562690f5ffcd2c44a4362e0018d9ce691d9376855230;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a83629893d7e3a1e2e3e66e224dbb58e20d4c48fdac75daaa5756e20691e99b171c0b78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h140390476d0c26d904c48f286728549dd68c95ad7641481e0d2c6e651778424db360bbe68;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13f4b0765c6d8966da14e02fadf26d9a854b21aa2e1582e1e789e4b20a048d9e7a453d7f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13fcc68fb5119e55d3283afa1ba5e69cc46d57b728ecf9cd2068320ab33cb225f734c6c9d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1669ea08dbefa539c914bd01285ba9da1b52f5bb089e0103c90c39a47c3fab14fdc387bb0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc5738ec351ff41780ef652210d8d1b635491e8d578c6e6ea6404ea1d7a1588693c3f9aa5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c303d81ff0b2fdf82524125de4693746107a5d4eaaea200ea5e12591ce6d8293f0741d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e91d3496b435a76d8e1d4c907179611e19ad48a3687bdaca6ddab4058dc87e4d486aa0db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e11786dc856c67cc22bc005079ef6f73e5f1c0549fbea76c21a5672fec403ac15f43d1f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1607ec6942c493b43c3ac9e220f5fdfb94143c2849bfdf920f3fab56cfb072b16a12e7ade;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18a89e26fba669366067df5aaf8ebc10fea58e5a7f6c795b44e30c8e11f8cd3c9fe040c2b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1319f59995d952148d27ca7fffebb8ddd49a7a268610e3977e4d262215b16abe5f47be819;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec689294ddf73b960ee112bce4657efe6d6c9650bc88f62b402def6602104fb712d8cfe1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfdd0cad5217888c9478ab529b04c9488c2c1d17b7be1b0de5fbb51e0b32282963f4ac7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h90918902db395b59422b88a4eb53c0a2eafb1d7eda658403644323436505b1444acd1784;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h184a69e913d42604915e3d2d86751b65505ffc7d405821e0f13f5c68a120de161ce9c043f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f380e966741337184d0a6146f8430500ca38d02385699e3a913fd6c307f31acab5c0aac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h756e5920cfa9230c32da686ece8474ac6ee1d5f6d01c1d58abe02fc0371d22a6324a70e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h130d435208af7a1f27ff7c256861298c27a83b86a8b235fe033ac003985cda4bdd8b57022;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc67aaa5cd8f125e8badb8e15f7e549942bacc71c5a30d68a7b9ad1782422c05bb7032dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14e5bdd32da80a5db25cca06904b78a8923f5480469d27423da92bcf105682ea78a7fd397;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d74ff420e902857b0af35b549363d1bea0538ab075bd20bc44cba3ae9edd2a85814d3467;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d55da60c08511d90f890cb2e5925f80e8a923241a774b8172be75be4859fe1fa88ce6deb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a9528c2edfda47234fd6e7f4d1ad767739165f10178b0b07f3b0788d432995e0715604cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2181d1bb20081f16e30e0386cc1531af8db2e6015e6384c9049b19a2e2149504b4964a3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc155b8717b538477635934d000d2462122beaacdd842fb93080065bc27534cf860a6f81b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h90f7588f313e531555c6dcf6ce75af4d540e08e2cab41be4610985dd8c2c6592bda36d05;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1551b3994ffdacb3c11278958262da4f71873edcec6261c4efe68907a6750de2e9c71fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12de9f4235ee898aa044c2065defc9a12487930fee5dabbc589bf5548a2f9d46c16928868;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h111821199e7b4f1ea513a07b7b9a0c95ebd539b5d10ad0b1826046636e0b9c48bdb6d9756;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h25cb99df59f53cbf5144604954f925903101daf3cf79bafa95a828b0de1ecf60e45843d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc888db8565200f6e111ab22d24b73787c6eec65e2a6605fb73b8d05fb628aeee8ffe774;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h619cc6a007519906264f4026051407337085dbf7f4572b2bbb2b9e78bc33b7f4b5c09406;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4515ea6ee9ba4a15c25c8b67c7072d3e0147ad8094e00fb22d6b78cda8c4d668b09babf5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1600291e1ead6d4e5fe6dc93dc0240c297591029f343dc73a069e38c6abaa6009e2ff9526;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12db55955c3d9e93ed9a281dc7b94e653feb25f35663fda1130f4db086ca8ca9337d3aaaf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h110f378ef9185a4000260c5669afe0bbad2ae6f8b7af7c886c4344dfadc61f36cb61cdf7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1d4d91b00fdbda11e1ac9d631c2164694f2a96423b750db45f08aa15db48209c8495fb8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h992d956f665638d377ca1deeae06c0483f8851f34f189c56b54048f205699ca1d64de6e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h747b9fa3554647f060a1b94dd34378c7c32c1bd5e47ce7fc6b6a9d486ea5811e4f54629a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8fd23b8630f0cd1ec5af5675216dd5437017acf238be20724e24dd0486c92300494ca782;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b06743568de44665ae3ebe51aa3451175234dec4b23393e01f904820762b711a45d18b6c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dc4645ef20bd27cbb813cc500114fb2f00654474253becc28b00677c1560ad0bf06f864d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b0d10fe34beff9c9b651cccc5895da3b1924683847a135f47f41483acf1abfd6ef8260b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e539c5a813e99700fda52038223a53ab6ac278f1eb4e36c977ab7c5536a84db8446b5348;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h119f3935176b1d467a1ddc6224c675c7407a990aed215d781f8dfd2f1cadedf76341d8a84;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfae3b7b25c47eadbe930e2be3eeff983715279ee5ee786a7f6937dc84f12d5d78110a188;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h491d43428f66d102fe107c52d14305c5962cc72dfdff5baa4d707e24887b86d2d274a0bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h43220eab473a3022536506add1254bace2f99e21f910a978a2324a5d1ae46660c2f3021e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be5bec8871b55832564064c18ee51160f5f33093de15ec4b36bd5b94ddceb0ee59f678f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc3098d49c513c233c88ec12a32debf4212bec3819166acd5b82e0d039e6601a2776f5e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1538f97165cd4846472bff78e6d247351546b9e8652b71e7ef4a30c37ecb92c078a7b2454;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h498f8b591e62abfdf33fd386d38a47e22e7c2537f4d7b22d73f11c1e04de37f0cf0cc1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15bce3c50c06599d5355ae91858f3b943c72100b27ffb53e40c1ca58b4e40e383c7bdfbcd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55fdd759cffd6448867f2375d65b5f995cb9184426242f6a4bd14879c4b8841d72dfc40;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cd9c960b216cae342bc572d3b8571ba887a90923c77ea7b3e37218bf873949f1031225f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1307d760c48690e0134611eecda8552933b0c57c82f6d5a6875e1b45ffd4a52d86531ebec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6fef8f96899b55e89ca8e129f00ec8a2fa3f6a830aaa933d4c847a1298170d70b9412b7b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h188a38941836a523bc28554aaff011998d99fe9f65018883b5acebf2c3b1f35d800b592bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1810d0726fe12098e58f715dca532ed78e055f91439ccea510521b3649ca8125776b47fb4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ebfe8acbe0fbdb9f6efd5abeb588416c507985084ef5d8e2e94af92ad5a3066d03518057;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10454571a0b474a65723b1f5e7cde576769a266489f2788ca69ae92b3ae134e3cc746392f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h760d1eca2f8b1b1ef401245b0dd59d268b91fbd026401bc582436028be467abcb3782180;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91f47119e18a1dec8cfc61d39b7074723bcdbe657cb3fd70bc5b0aeccce30af385275b7b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fb15165041536ec1ca874d046c84f17d1e66dce372c1fac8617f8cdc031880674802e868;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe36ebfdf0423caef83e2014ddedf4533ee9fc75a47958a227023bef3ecb7e954298ad9a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd6b6ac624e7fe67850f0c946b4da2d146250346af2b6a3976b3215b3c12cede1b42f9eff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h188db28a188191e7f249d67f83bc7f1b882a60af3732e715221991d6ceea2e0bb4230b90f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h522ac90cf4469a1d0d01c9383ed708a18540a6ba46dcc9716104cb165e65d0bebc085beb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12dffacf9e038c54830d536fae3e27e77e92d4a8d25a953d7faa61227bd184a348e63f99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf26c518a75eebdf70e033ef9436bad182297bd780d1c707946e070fa6eaa8334d7d93d96;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d619d131e30f4898dc5c55976fda434e4223ee919bfaa7808e2c152930957a19badb1103;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11ae6ffae38ebeee606b02d9781351de540623f9c2dd41c942aae5a70ae967f50d088ad5f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h64c565f91afea7b616301513125c0f93d0fc29298e37367b4133d1274b2a7459dfab3d86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13353b48e2736106d40c0769a2c6bfa222990eab844c7e0433d6a421d0f1086a80c339fb5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c5160eb80fac76132046fe178e3d12d9878fc06c896cb03b00bc808b88608fa377269b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10a64716d083e13e5c40387b4f7603ea365eb570213c89e12af8ffad88b4688cf2d136fa7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1463a1dee434048ea816d5067a6b72940bdf4f58104fdcbe382cffaf7d3e4d40171036b6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14370f5a1fc7b4b6fae4c24bf3db52de74eb8f59830403c068c9759ca470ba5ab58d61a9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbaedff853c1b4b17467d6ef500a7274f4f61ff7e92fe60043e86302f538fffee121e2ec0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5285aca309ab7197224563adf2fa580effbc0a630a0f2c5466be79c525d214598a77b99d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hce0e4d7c0213b2ab4c186e2374c21a9df6427e7a720943ab9f05bb67a6195b6c6c83941b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9546e68b135e12d2657536dd92620fe8d47db5ff66694e6135aab2ae5be85a9087120a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb30236c8b92991838b9fbe4d4f02abd62cda9ef61e1f0058739e3e4ef22bc61ed8cc4162;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4acda5cee432bc3000978d2366d006a8aebe953f34bf62a30968d7641fccbd479c55478a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ebb979dac52e4582d9e5997f9d40f1ef40709993ccbaf59da34fdd281ba1b1164584e48;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e8b4de98808b72ad69c0dcce377632f23ed2f8c4ec616e06c5c16451678b9435028bbf8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d2504cef79dd3a85be756819f278595e30cd970e3ff6dbf1c0db3cee642813554dfbb81;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b63c82a507e66d2451a1b0fcf2f208a061c6461f9e2f155bf44e1091ceb3d7a7686a391;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166266b31ecf83f2c24e2b39962da4286140150f22a9ee4bf2e217a9fa885cf6a085bca1e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he950c1367b70f5a2f472515773a795abccaf50734d0619476882b8f34c0c5b08c89ef51e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12fc749a63c5960ce9434daa7ff7e09bdeb386203a5a97cc40bff9b449489c5199e317082;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124c449d6a8b4153b1a18b7a2df8a060be013b281190958bd43a73e8435d006d6fbd36ed9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10f8dcbc681eaa43c284f477c92258d84bffba44c4ddd41c9efbeb6d0eb9ca2e9a3b23f65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15621ef3321a9fb765004408f7d2690b268f1ad0c1c96f33688a2f95359dea8f20114c891;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he52db154a96b96ffb6e7310155a1eb9ff3838963a350c63342d56d40db205b3fed55f5ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3bcf9ae7103d104357e661aaa787bfb5c28bccbd6a64d51c36d121ca2cb1942b758446ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dd6b0cf236eba72f0b71be74731c45c760a95133624df1450bd5aae2813fba7200580fad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a172d5f7981fc1ecc321ab9153bbaf3dd6882927baeb63555ae5542b7398bf0d68053f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e621f9888092f2b824ee304676e50b2fdede6cbec4fae6d8e4d344f34cf1d0f6bfec8ab9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h160f4c07139ed95e764e39510599db003b736209754df45617b1445d1c74a609d3312244a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h28d9edae7d465fd715f29981446b78e23441e50acef20277ef8a866ad71c7d1821a4af6d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hce4513e15bd8b16b2b1e95e83472076f77f9990f55b79c0ace26e9a62813a78c539badb1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h99e377a3b2dd2bef0037055dd3a28c55ee4736ca062f7a62313c5fd4c016bec0598edfe9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7cbb301db6962392c5fdc2288f3b5e66f26523fcaa961cebebeb89f1427fd7b8a246d4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd5d3679638694a3760bc6384ba10f127d27422980b89eff430a4fa36300fc1979606518;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10efd4c9fe1ea235c3ad52d434d742c690d5bf267518ed0ce31d75a7b054cc39035eb07a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h401561c9e57be3be101878f240645a16294395a0c24f6aa949ce308f4fc275d15efa5013;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h69e2ba763fa7fbe048a886b6efd7bd8eb4139bbffc734da900adf0a277055b521a14657b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59cc06f99136518f20cd37eb8f9d8848ffe59c6a4075ee22d13b9006956d570d5abdf52d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he14b3e634ee6cd42e94e3d7c8d0615dfb2eef4cf7e640ca6c889835f76588628579bee0d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18ef700ef4d03ce1ccc5e8abce32a930df7b4482cad39f69dd2dbd22dd28303c6c99add7e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a66e360fec0f6aac2a4a9aa9935161de2edce024986004e9c758254e7ce725dc092a168;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6fbd8c6413d1f4a98471f965398d1c1a893b5daa32bf103b624c5727f465c9bee5a9e30c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h35afd792db934445705bd591b0f99d392086feec76ff7279e9e5c9511f99ee307ebf41e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h40576b1379a93c5f8213a77fad2dffbb83ab3cc10c17e6d7c6403363ce5f4d2cabbf233d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a090484b3856ca0fce04b3cbe0a47fec712ccaf0fa1cfd28900e92751ae3e8ed4096f82;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h44bac61d63968b592981d5b4df58874107e6753cf798a2cf0dd494ed2be8bbd1a45e42e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb062200593dd3c41c90113bcdb4bb548581569f63ed0138674180a1cccd77488d04634c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h81ccbd86cb47879e018de89a3d25826ffe7dcb218cef3da387a7b2152a70f3fdd1392e4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bb667149c941f5a2f74e5e521933f9b57cf9325e7314f8c6b55ecae94cdcf939a780ce5b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2213134bd16a457820289fbc5b7896ca9511769fa234a9f3a3dc337d2b151ab2d6c1e068;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e4484cdb77c3e8ae1e547807b42c26f7c803478cef7ba4eb4b0d8c9faf69766746d18442;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h57f6b38ddfdfe065a9a9ab0de6f080419b449ceeac0c01b6685f017e2c007e16b659371b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha163249177950dadc633ee61ab54c3cd763e8699fb2de819d3827c9720bab54971baafae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf400d59f96f58b9bed3c1bd1c930e06e629dec3f6c0519ed3c9d715fe7b10ada33ab4233;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb81e00ece90d60976571495f630dc098cea31509413304f9b3e64a04fcf9aeea4cdee48;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13f2638c5a4756a5069cd3d41a7061c8fc01d3ba343abb887704ecad6776b26455674fcb1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4c86a3ca390931414ccb8d1171676570f269a429defa1f87611c921dcaccfc2e1a24fe50;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha864ce88a4c23161557edb3b76518eb0d300be9ea3b26c9598d10926a75903d05e856932;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb8f0a8e56757e826932945f0c954c3e985fddf4c299a71d4d6c19f35dccbee8da04058a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcfdc69c148d496799d28a5036482bb7a96c2035f735a337887e10279b00fb9096ca65312;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1243ad1c6f95a602e16cceba15682dc592fddc576b437031760efc70e8c05f807ecf98a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h481778598be0fb1c5e3bebdb8a77d6ce23202973d46b42e1b80e1fb6253dbda47dbcf09f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h45111c86829705f0ed7f7e3b74397c5a552f365f8eb552ae6038ea81c3b860a87262851c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha2a8f14034b3bffe362aa58fb7bad4b02a1242abfd8f20f8c606fa3a1f0fd4c274bf8347;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h246deb64337d339a5fe3aea8a8507003ac0a0f72f6d7cf1f9ae7476c87997d0e748e80f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ffb6d5dbfd900aec9b8044c028bbb3de814e6379fc1a4b9c4bb2279395e06b56b5a80ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h152c6c2bd70c91eeefc307c5c3b8ceabddcb5233d5d678aaaebd283de989b19992fe07b08;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c81a38f4ca54f4dace7be12890a109b465a6f6c086fe648be47c6899a09c630bfae237b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd544c801de169b7f89912fc835740a34f06b8fabba4aae34f27c1c2b3d59a4656a2261d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15c814133f3ac558fcf034630a48d5d8d875a9719fb2fb14e670a20fa0e92179097adb348;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1288de032d3d4bb68ca676a1259e2661615623c56e9460617a58cefc73ccac189d678ee76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb9a3e34f2529dea8bededbfa7c06c412c3f5ea89db07d1cc3cf82ce061e60404a5160e71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d44d3bbb7cb6fc37499bf9ccf43a178fa9385b146aa0e89da9546372433d398f11a18b7f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h129b952afc41d12c00cffb4885336280e8e00c3fc960376ef61c8c32280c9b677c0bb1363;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha49d12955a47d75bbc4088844aa718f9d8f2656196cc18eb0649e1e9c0df2705c04d0dd7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb5429e64d3816c7a82eb4789d9ba3e3c79bb137969d455032d0c0e56914d1ca81cfb640c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcbedbcba0c3494827737a6d2ab31765e57347b6db5d7c035756d9ce62d8cc849b142fea5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e3fea4ca1727c2bf1a895580d58fde7b0869aefa241e7a1c3a1a0f0b0b109d93095dbb9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hceb7c5c1b0ac0f582081b589eeccf6db36d9986b182c83fa7847025efa77cb0b0e82fb69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha7b2af140ad18706b275f20b8497148524c71656a0b0d5e9165c1d2c9db5b0a99b3b1778;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b0a703175085aea2fe7448cc21799ce38e699168456917e391c84da211893390043f2291;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h193a57b5c9ad767127404cdc9b41575ecc20477ecf7be2c61dfdfbe1493ad0e495696bf62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f013d011ba280afa083d266ada468035dcf6b4951bff73b91fb0c169fabad175b24441dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h149daee1f9404ad764af0004d2449415ff21a45832d4c95d7013f5a6ab3193c8380e4810f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h68e9595daaed47b1c24c04ee3526a03a67984512e79ffbc576488077f7836271768034a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d64b5e27497c4d5222bab3bc48df4628a1cae06e9173b136e95521521a89359dc16e057;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hacfff7dc4f06cea558e47ef8827d9d846daad21c8ce1a7f53b6c8cb61086bc442da0369f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8f2601e57030390210650aff4e5d08a8ada2a97212625f21fb2ff35600fe1361914531c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h119a56231b029f7ad0e8c87bd95f87f0e5aaeb341d6b4a63e1ac22aa3a8060163589bebe6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2a6909d62dd0d0dfe6a6fb34ac03b57fa8a4ead5c11eb4a21ea7a7c57b15f6cda1f69998;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13791243d552c83b729737d72a2a45477a77b1be47ad89327cacf22548a795437f958af3c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h188955cc7d6cd5b6428ed0445531c00b810802fb60279dee6adf0b694a6a75a95157c9c68;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h74b3175df55684935559f5b06ee83c88a75251d054393d4de5a19dd4bf10f5b70c71e274;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ff6dc34e65102d18e1035b0895a2119e471daa7909c9815483cadf1070c740ac3b67708;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19873a40f66093eb38fb8a76b65b1c734fc6a84ac3df373ceb094be782d8860e406995d0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1590e5f8e536a6c2e90df2f46dafe5cfa802fa4b9a547542063a29ae3b7cbbdf9b4a5d4a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h120bba337630e81c3da6beeef21091610b52028f4d4260298e835ca6da2c821b769218b6b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8502c187b230bb0f05e50e4019da335ba0d9fa56e466f328d2d04c462a06ee9684544b29;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87396d5519d266845649e00240b100f1378f5ead135d8467450bd9392a39e2d8da15db7a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h285b68730ed838be4ac30b1009e031960e91e0ccaddd57d53205c3cc21c2104e420496c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107510928bbce779b6f458c793e3e5e74134906510bd3a0fa433d3fbda452db517a19bbd7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h173e844f7f7625450ae53a6cc2faae6bef357511c30de819245227ee656133b5fce370135;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h85921a5588d7545f7acc69181cdf68d19840d5e5729a448d847e7830715d9b347767e31a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7d7efe1023294b36af4a6a7d6766014a877eeb2d72ffe9752818ccfcca2727a4283c924e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fb0b01f81ce8d2219a7bbf703dd4cec263f01eb761277951b5f646711e871b9a7a0e57dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8759d948b35772a59e6dd1b712f6d89479e090127f0e7b18f5ec94fd37c9c48187c42a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ece70f13effeeb55645e6009a6a9a2742de13c389f9e01955586b41d6aa04b47f837414;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd9926c9d19aa4a8c4f88497e299f4228fb6df6195da4f3299d10c04a11bdbc575d8f90a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e238652492ac2560e5dbb41a2af52ceb54e9eea48b3f8b4e2789f480ade90df7654461c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5bb4d275e43db07d6be577c9bed756c8500971e2b755a38ca71342718f34fa7af7c4673;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d944be329fd075e9eea10913766b2bf63a1d2209aef609866d2f76dc5df26745c9833c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcea56daefe747a8de441f9261423c1fd3ea9f05f4654224dc77fe1930dc0aeff3a9f8ddf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf03490fb4082b00ebc3f31a8a10aecc267fea4b3eaa503011ebe1dfdf10635daba5fd44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a9de78f381a72b61e895a266b7e04265b064b42910bfd81765090eb479b9c9241551ad41;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h835ac57628f218440022a0ab9c11b29ca7ac16a4e056e1dad431248b5b1754e3e23a5dbc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15f95f484c7d41cadcc947d18e9a8bbf2c20d5737bd726ba013095560f6a09e32f3b057c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1093babcdfdf9295166476f4ece281f2ca377b47ca53bf48db7f3a69535afa891eb037226;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a0d083e88a28ce4676443c778e747f68a4450f00cbd201248517c9e9697b3b80d0d830f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1876a91fc1ae3a8b4dabaff46752f455c48ac75437529bf962d01afe671c112e9efb5f63d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c1dff8801081b82610c2b8ff07892572622443301ba0a2ea692f9e5f91fab6a684284f22;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h156579c953e9f775c9b64458706e69d7b76a964d81b827b9151b7555d7b8d45ee6b1bd6bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h80f5ac4088469096cfccd0d6146096d7038d6d48846daf7cb6b7025825a36786187c9305;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h130e6cbc760afb6bb1c44f2fa200e398f889507981a527111c89f7024046976271ed30d4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15ac23fe06f780f32e78c1531c945c766a0f8bdc8b5e1cff0bf57d94bfa75c131b295b156;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11dbd01079f3d091a9ab4cd1b7ede906dbd4ecabd4a16e71bcd07869eeb80e4110f37efc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h139b9bfe271f8f3645f1f36b5135edaf8ad3c51a0526bc0ac79205f6e0a6e43ed3473f1b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd00119378351603821361a3faf8795d62294fd3e4a36a7a3234a7517870a7ed800d1e7df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113a15a9ec5c31e8461312718791f0958c694f2ad02ce843b78e307b7a6a16e3974af29bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8acd862ff59ab10a39d7e932fb9a8d990079849e24f6f8c9a523b567054e39849469df5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h998ac08bc2916e0a5664bbe61f714fe65ba6f34aef55e8947bff34cbc15807fbe22cf140;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h39dfe895f389f768d99331e258bb650f74d4c51b448e4eb3a0dc43c8b58855245930ac58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e211de61f17b06be32cbd2533a25a0df4e6bf5f47d15a50c2ff1e1ab5c00f81ace47ccc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b70366396ed00967bae86401694471323da4373091dfb0a956a258157e1847911c903c1e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1750b149dcd7a05a6b162a4c54a90f28309cd1dfa532f54138676e13572d47892713125c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h104ec6d360efd3b12c99224f9fc78a9ace847213a371a0cbc17eecf2b3dc4ef63d0c3266b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13ffeaf0e53c302db9bb7d5beb46bd02ccbe5c2b2dc864e604ceeb2b7623bc6f1a9787795;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee9de678dabf736f3911a7dc93529be6db444cf9cb71e056bbab218d59b066c1bbb3af90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f3898321180f017287bb07ede769606b4bc4f0c0a5f66a609d5e04f6554c3fe1bec35df0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162a63d566955d5e01a5fc383b71ff7b4a43257737f222fc22da64f94ed40fe0cafdea132;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1794ad52aa9a462b2961baaa50f4ab2e7a7a651e0275794f64397d94bc37565d95c3f48cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135bcdfd947e8413ab89372d70e2ed76e0ce6cde6089d9782075aa5554369a5d5cf9e093b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17327592b5bc0a5f52fe50ab32ad144027c22e4adb2784048131743b44c79a44b9a741c7f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1900b02aacc3a51c03fd124dad03ab5526cabc12ceb3d8fb0e3be8dcfcb6f9ccecb0d2e74;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91c39b7083f8335b6c9ee6d67102bfd2920d6e888651c637991763cc976f70593cde04b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ec80c7cf5a7bc6fbea0dc46c3505c36b3977367a2a745b58479702be9d9f7468a03071aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe31ddba65729b09c729a42afe87ac1e0aef8b07238e0971386f155b8ba3f32f58fd5be0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124b047337cddf72fd2886c39314870628b0ee0e90aa0d29a6a7911c3e8c88c7b1991e4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef232ea96bfaaeaea3e3fa513541b83208233cfc837314b75924722150e7ce8acce588d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3045fa7762e8253724c71d68ba814c350947e04fdf28d621a89d57ef0a04a1f8c853d3de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8f6da4f3e494516a2dfe32196faf48c4bab91b96cbd0eadb8c8742eecdab0eebc355861;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19285aefc8b8b339d856b24ae125eddb97048bb3ed7d9060736a80f9b7cb853d5e3ffd6f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa6667f0a70a6e5e4d31bd2e9bcca609d9d1b808b235fc1b10c6dd3aa3d16122cab134ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc66ffb3f24344100861dc228006fd3e53bf11bf50349bb28ae2e8a8bab23b35a648308e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h139f7edc085f13a99b277db6e4dff47297dafbc1f85eb9a07bbf1a0a576f5f84acbbcb7f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1154186657fd49ce093134055634e7b6f10dfd27a6d7dd58d69bcefec9e9d14393511c6cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f4348e7bee5b671c26360db5b7c4bf647b74a7ef3aea62db102ff7cbe73a2f7c43a8d119;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a61fd400aa1f663d39dc922fef2a69db1b573e1508b68b2595c9ab20b1851b6a8a040b36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13fe5d2d782b14870feee6c767fabaf2ee88b9504e72499fedf92024aab209ee74d12bc4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hce5394cd05c834f80c16eef9b41d640d83fefc75367658cf8b3295e7ab5d67835ad192f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf79cb457c32efffff70f91e412782390cb5f63bf1942377fa03878e9f39da6e7ce5252e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a283b694b81c098a85dde13290151ae38ef0c696021ea2d2246e12028c4801b73bbd09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h836940154f957a77ce3145b2649589a6e37fff956663cc2b9b4e1f840b903c9b5292dd39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb7ef63b0f3aef6d9db0ac510731668b6487f53d95c8470da46a71cffd3f86871349aa63c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd2d9f273097f2d8a098656a125ec5f880d281735b4d991b7ef42d823b820fddcdf08bb82;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6198aa2d7c63ce18699919f8be79d184e75e89a96a92fc36e845b3372b2fd09adb5f961c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4de51f24f3f6dfd018742b7d44cd30bfd60963ce8b5f784fbde7501ce31bee99c007c44e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha287b298860d6ce95877dfc686056ceb524bc8d3db3137aa890806e7b1d84ca74d1f96c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc1fbd49f0dfcf3543a81133b0678f0cfc9abb1a191bc5e99dd5442d89d90072782d3ef00;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17a7ff463e5de02a993253541c374792413ea3c58a88cb21be69637925b85801025f7b1ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5d69eaad8a690194647b58181359d093b6259773a14c7164369febc39a4562f0950579f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a8b6f94e29e07f19d4a67082157681fe374e980692b3394abc76e7ba900d944a9a91d11;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cc20031ecf279d6520f7f841885fba41c74e01c79fc7e8430e4930c648fb180d6603cfa1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14e0228102e97e9cdad20c5ccb36224519fe98e46c1647e71bfb0a8e335e85cf85eb79bcd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee9a7b7250c523d6e1769a55a329aa3c4b1a6e1b95a21aee2c05d65c28269176dd63837;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hebac3632de4c7b1c5d8342932f99bc8a45d607190889a4750f6476efde09f0140402a961;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e6384f6e4d901475501b0b8816f0bb68cefc42b6fb09535d9175f800d9a99e90c2c73d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b02ed799724457a3dffc84e95ed9d3b41808caf2ab9c41b999655117da9946a0d0f31a0b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7942e07ed3c3c44e0ae77912da240e9ab17f97f11722559b608e56ddc215e4f8e8ce8267;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107dcd7e45233ec285a606ff83ab60b4b80dceccd9a36908fc32f02b2448a7f125c3861cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8526cec857a08a6486371a5b6b95a2df768626d5325bd67f95405691e50918713fac0603;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13409934e4ce32fddeb3b21555182890dd3471c1621e15a021aeb05944cd51ecf1f3b9b0e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha0d13328994392801e79e1a76a74ba3f7270bb52d546caf480de7b0c632537e6885282ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8290e6f588ea8882417ca33e72222a5011e061f199ce03cc89bc4343794a2a53eb5bb1b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18963cd3902c15349c5dea6289c8ecbf384db2522f9af011f331b4bb92cbd7e70ded5f653;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he97ec6ec9dcaacee5cd43ed179726ff890aa04d8d70dd7b139e3fa83a2894345ece3d108;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hed0731db5fe1b9c60219314c7581ddf8c20768c270d713ae0891ff34c1bc613ff3df6f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0daa7aebfad5b01d5c82d662b472215fd5b8517900964d28b750ed73bb895c394510425;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a559f024c3094b6c35e5ccb2ba1e7cadcd5366ff0acb295112fa8186773b5b5d70c63b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c5ec7cbb70aabd21f5d310dc68ac7f1365d0fe493f1a99cb9d67ce5871a9d02b3be9f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a44cd35ed0f00be536c8ff1586c794e8d5c42edaea64921d0b319deaf4686d655432633c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ab5dc1207081a55ab20ceb6c30aa8ecf1642f3be307e71eb2d0525f7f1d43eeec45b922;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11230c9537d045d0967b5c4c867b823fcd1df6664a145b344c99186b508b26c9c1a1afbcc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d034f22318840f39e9daba82a2e7ef96b81ac6a09f9ab97a0718a34cb39bc57d13b6be8a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe2d8587d17a246bb6b4ae65867ff4751c15a61b4d01be8f56e9bfac87385719d8ff7665;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b43b4c147ec56f7d04d82b584789c7454ece4f606541b8cad9682f6dfe34f414a246307;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h141c1495fc3e4582eb1829eeb676f5875b6ce8be24bafda27e1577975b930e58576e2b68e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h144bc986560d3775968028ed4e6e9cf53473e09b90a7de4429a98d70de465a6319adbb5b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h320b0ccc2bcd802a1903ffa254c206919b5909e4ef2c5da4eb2df39b9f9d766f48cdcd7f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h76575b921e1e929dd3cbab8880538ba1ca40c259062cb5bce95541ab24fdaf11a102a21f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1048dd3ea50c7a57e1e871abd5fbeb85fd9440b0fe9790c9c32bbb94f87fe5b1e96f75fbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h614343fb13f00a7ae8ca0cb0a4bc5b04163caf11d27bae04cfae171b5a78f4932e93b184;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h85766304dfb38a5494977d885eda48163751fc0dd688e43ef22fec636c33f82a1e45938f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15caad991587013f0adb26f0393ec88494cbd77481be98f98246fe7eb45f1aea7927fa524;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb159e2b61fd42a40820c6b894b230ead4400e66d33775757d7accd2e91f524c8b376329;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea7825d9e791c1943545d6da46d6070a7079545ab18daa2acaffb9a1645e37c9e04d3b81;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fb412d2d4c380cfed4f6dd7dbb1cbd72216b65004ac2cf4e8a9403b8172434bee41da0fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55d3836f765f8b7599bb0a561ac61eaf840f31be0666f98d5777a66c8b63f533dd795370;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13483664ff308a0112ec0a88ce251c78156c0874ce5a8b4c675fa20f5134e74b592470155;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5af054321a4d4cd2b52c1591d35366fc6b890f2d66c5a2ed6e2d8cd9c2f325c2d2055f79;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hedad4738eda284fb5a43aad8cc944ddf5e0b9c2521faa783cac5cd1c66589b0bcc50cb9f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13126e7e62279e08c7ad70c248adaf9d17706852f83dd304c6282a552633ee072547cb472;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fadd6939062c23802cf7f3cd41ffaea3767c1f740603edfdcffe12b6dd9213527c509900;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h115e57835fac1a4d2cac4ad0afa9da09083c7ced95ee179a6815d7f822bd448c1f3486c02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162fab9f0323acad3a447af9c5eeddde91c865b74bdc412d741b620494478999640b25675;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9e2b6ba67c13af9e29d7024b467731990b39911c173a0853e2e3a220aed580d59243d5f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h24a03701a074c04e32fc84d618981efbf5c122b2dff93de8c409e889db3800dfd0c757cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4cc512194292eb44b9fb1a78e9011b58c8e43c08a99985118e2b1bd5e3b506136f582ccc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h84d035efd8152dd54049e4942732618a44dbe12e0134f2a551fb21c01e99caf3bcd4cebc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h158b885493be5f375f91d51eb492312d649b8a05aab87fa0122914750efcdc8999c0fc34d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124e10fd12559165dbd31cf8329ab6a3e53d51c6a700257e15f2bb11d6f0cbceab0fc23d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb68e780bd2c6492ff7bffbd69c5a0b849bca85c613fc6a0b8e93bb1c2dfa867b2f646389;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc93f5adb4d3500dbcc0cc86d1ac8e1137e2047f7b2e1c07d7cfbd0064478713347ad40fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12f944cd6797430a5e179b6b8ac2dd6be1be58c6e1fdd98006425785c335e9b47453b351b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b02ea2b6644aa3a446c4de67437fa8d3cf86199f7b280d7f5084bedca71cefff45d84a20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d8b69551c90912580691bfb0f5e9f40b82708b962d986201c147e16a79382f9c6bcbbc6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c35b343adf2e0b85ebbab4d4dadcab57475fd5cc9680b4a932946bb3c8eedf43a456925;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h193e38edf1dbaeb6deabfebf43a00e752056a834440b2ad49b1073fe88bdfe1633610744f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h143f413caf36751dd37b960a33197187bb212d8baa7856d0808e0420d5a20891e35797305;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h244a95b294c151ace1580599ad567299a5ad92965e33baa219a8594337e2f082fab2dc62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe0fff1c8c4867c7fd7118f79e18b2cdcb7cebac7e5cce2be72b75dbcc1b4c8ede522723;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h104aa2853705fc7c791d4720ea1e28a4b410de3da46c2e0673c87f96207b404e97b860389;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h524580d32fcd9def3ab184b83c27483ab167cc205a4678592f66dbd3c0c2eaaffae69ac6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1530716dd840810e6de2a7570595bc14ec783694eb65e56ae35ed86eef924aa25691f9789;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166368cf7cade348c9f8720296cede315909fd52df47bcd45342664734a27628100df3d74;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf089ed6448dacc1b51c796f7e62b747ee6a4331d8438269add5550086a8c1b39102dc8b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c42c9ed58cfac9ea03975d147ab54aaeab7ac1a7ec3d6ab3e258c63417dcc8d0b01a0db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h705710e5f0ea2e1af61b4f50d5ba6c6cfbc29b253015dbb7c7f038af93dabb0dce9a1e8d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a923425adcbf2c420d0d3dedcd8b8d7a67bd9740f9a979ef5757edc7722077bdf77a3a88;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16ee9c18e83efd37f3733b852d00394eb135013ea970629b3316c0c48c9fbae5a30ad6c2e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha02ac3526ce7f9934d33bb53ac909cf3c0c47f6384557c95bc5e5bbdf7f4d98ae34f90fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbafd7436dd1cdf134febd6e29263d3f840dc7b55420bd2baaa4030014b601d54399fc486;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h168a7e918b5626791454e1ed175d9df0b01be138e83c083536bc39a4e3212a4e8aaeecce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea8b0aa9be2f4b42f7971a465cf15dfa8a0f8ff6b500f51e46551813c451f031c26d5cad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h123a2a9a1e62639e15b5f8f10a27d7729686b5cb93555e30234f6d2f7a7f63cf9a20976de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12a3be8895e2e9a71a34e49334c01ede808f9d3080249f0696da9066f83d84142a2608e03;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hde66b2b796c2e9fdfeabd8b8df685c0e70247b78266bbdc9424288834a54a3652e1c8037;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc4c011a85587c59b9f9cf52ca101968a2ba0fd0b64fb37db7bff06a6fa3db1bf7e9dee2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1448c8147617b2541dd1048053518d2a986762a3d217b97a4afe776d9c35e49c69ac93a18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5315eb20dff31040668a38a5889e579b69fde25eea95840c910af8305ed3c83e2957f463;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc74b4cb1228135324bafdacd3f5ec4069e4c7df1cab8fe1503ef984e6f29dd6413d328b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de441966f75cc8d76e3b04cab418e2d0edb89a0c1b97ad4b34c0ebee4ec889899f8d7b5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10cdb0a331e53539d1db49cfa28e1cbc53e12b616ff7a8b34fcdf1f1d47d0758258f90ffb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h491b3f22a9a3cc36bf2b683ad1adfb2b47ceee320ce8100ef9ca80289a9d0a9b29b7fb09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4eb3b396318d0013caf5c2108508cade3e0dbbc2eca19d586b9fb9798321503224b86cd1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1791d38e2cfb29609c6843030333e221437e4363022d155900d8b27942a5d4216c3766d72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h948154377416cecf156596c4edeb8c5de728e5a8ec13b1029af7a97f8d7719b51b1b509e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c338c61c33787a94aede60742185e7ec8c1246d5a6dc00d3fafdc8df5f61b424ed14eba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h142a42e8d64a9e67dbad5819051bbe6cae01d9a35bfd93c355de1345360c1584c6f39d237;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd3b94a6048d19b8d30d91efdea7ccaf454c359344857e70eb0b3ab36e1ef949f9752102;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he846239e5eed7875a282dd61c7c013598219ad4e469a04404a6172b914364402ce3f0b5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13cbe3b4fa8c322ae727cc6cc72c8d49f980dabd237740fe8a2b2deb1b379b829e41e036f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3d4242863b172af4e4301b33798a8d8bf7cd1d5730e0c527cb260f0b06c79823b808536c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7d28eb48b14e1c57fc51d79d45e4652e329ab884af644a4a76a8ec8bc80a865ce1389461;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c3593382e097a4fa18d792416973f5bb4db2601ec0bd1a77fd98bf58bc89c8872fea0b6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f99e5a78b53ea54ca739f246366fe2f80336710729deac5f1966a1d32856b999ce725999;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h69ba2156f439d2b6103204388a62676c61c4fc53fd9cac5873eb7a5168f95abae45c9ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16f2940ebd921c2928f32e7b6f3cd564314acc148fd2ced1573c47e52136197421dc0e3c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h126a4cbdd5f9c321d31f4b34cf57d31a34989a6e0fb893d3dfdeaff971b511e15d2f0eada;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h129bc61f5e72658918f1889716d3a8d9bfea66107ae3eae24b0c5ed69038caf6561522500;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h84ff0434ec99f12c4f76fca05d522aa39add97c60293b4de07c795eebc3c5c56714bb589;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2682b230c297aafec07726822da7ab4b106c1ff2a84e245a769db61ab6d0961d93fd99c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h178f15e11bc39fc819d8fb065c7e497d6fb09c81109d8b4803421e25ad01b7fb64214f6ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4decb92367c346af50992a91fb23b71ca0e78387dd42f58cb12a3c1ca34ec0f667b6bec6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcaa42399e04c5db893a4611a538c68983eea98d7e8f24fcd0228ede9af7d4a084e97c67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf573d48d077a4989014a654d71c5541cd5091667dac501806e85ce508b916f05feebe62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5d7538d02691a635e7e6fcb124f4d6141c6f68c38d55637dc2bfa76eb5327a9f35866090;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f40daa58a4625a50471192613570e899f8b08b27215a088c28e00d6538e93742c0ef88e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fa066f0ccee74b56cd9dda5b1b234d976e686e7d34dbfda40a0e7fcf8f7aff1029f81835;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c3cca34e743e5ae07ec7a81b3fe796da1d53978d93dc26e28d9a34f22279db3fe36c685;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he08edae46e2871635118344df62c5a6db959acdda95320fe9c1a414c9aa606b6d7a79e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17a0ce455786be9a29e607d9c91db0825233b885ae801045d7a389bb6aed0bab17bb0a2f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h154da69ebc96bff3fe198bf4f05ae8443c36ec48231711466767e16942e49ca22bb231a63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h483628ce8a5384ebdee074038837f29e18cea5d57cc641437a2d3769f3fd055f0de9f041;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a62561b0f4f8d16c2f2f00d300d4212ceccd017d063290ed8ae382fb5daf909b98c187b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he41a2a057acf91f4e1d1299537e4557d6908b97203d4519aa07aef618203b2a1d11ed936;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dfe058fc9f8df705b454aadb69dac3817e5a4d529223ed712004a28c2ffc0289e92188bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h114d872f0062c8ced54a1784c81cd7f645cac8b4c3578280e5d405e739b68d62bf9fe665d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h92c7b6d2d6b019e6448708a814eb25a76cb2b6309bc8d3fa56b01de9f4e17a67a4327383;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb44aa34d5a21a7b9f3cff36269baa2f2457716b57ac0986f5b882a4cb60ff48b5629608;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c5cf655213c45fabe67a10455246c83978c039e574c5c5f3f8f001004e0fb4c33bef6335;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bdc4340903e5e9541b89e9c7017a85d6ca8997b0c685db7d1ef69d212bc4405e754387d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a72180872437a36a6ea8e7ab35442b0969da8b24bfef969d996b966af112043aea3bdf69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7178430c8370289ff35fb176bb7767c5cbe8a933f5b03d9e949901497c88d03c92e0979;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15efd11e965cc8ab25f570d0e155217673c2b52f058ff5f8a965b906867c6652e82764e93;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4e24e79af22b6b7bc638b4422ddecebc0abcd73039e1d9a97c15a64171a4c2c4529ffbf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117c543d68f326884aca46caf47ce89fa90a131ebcccade7bb2a457092514c46f307f4de3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h164c84b81135e35046b7fae64651bb5451f235608b246063d1e90bd8b97708381d3a5d584;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107b94d03b41dcdb63d1eb350acbdd9aa5e01f14b16894366efa81c5b0e8842147b19fb46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc80924a8f8d43eedc0027c9d2855e7dfc56a3b4a3146128a13baaffa9cce4f3b9a71d501;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1ce13f9101700c168b02e562a76d5b453d81cbf59a5db92ea11a2270b10643d9174f3b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ecb5e59a916be53372c713aaa77d8950d334e5b06a55de604831e66929c12c986bf72774;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189d2c64deb5977300b1e7380ad592a935cc83980437433b5d74bd46699c07ef296b84846;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcf29f9fa1371b6e29ad4c7f1faf604c223c1e0cbde9f4fb3016652bd368dbbc886cdc8c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6bf7cc6b851eca4247d3d473874930f4d8da7606ff2f8ef751e7e8a043b00d0a020adb9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f27a637cd123f2d727ad6c71dd41ce9800993051474df62942619cf2fa8f25383d2262f1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3ab535a72f10be346d502a159f56ca519c355aadd062097c950b2fc68a684cf7a0642591;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a07c68c299c84b14b44ec5b469ae4379faee3a886c4e4db58f9245d817c6876432385072;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e693fea7bed3253a58760ad83da6f67480b027ed91717de13e63e0f52e9b2b34e25cadeb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h20887f220d46eca768591a5d9ae5777001641007fa1dba0fdad5c7a9c704c5fbcdd39acc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b90929e1e3da3fc50f86c23ec6304a6f923b3152a561da4e814831ce8a9aeedc0433bdc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1581f333f134cfe2655c512215f5b931ff658327207329f9e685ffcdb45b05c9657dabb45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h118739c3f453d6ce1e82771659163832894192c69cdd8e61e3a838a7e269c1e8175b5ae2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h70788562c0733c26e8c5638c2821bbda16e40fde70fcb2b7bba00d6e84e184539f8679ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e544bcc6f63c66afc71b5bcef90091cd0a1df1d424649dbf04d3eec842aa96ccafca3420;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a3b604a3359dec28c7c7bd43bd34111b3ebfa477ad30619a4000953c1e90741774ac2092;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e20f777ef6645bff4d56e13e3a5869e087b4e63f8bb86ee038107196e756d2f1a874f533;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4d4a8011c8a8bc951fbd7a9526242a3a385ef52ee37a85d7a27bb8e540a6f155216e76d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13cb0a3d514678976b4884283004823743cfbad4dd0d1941204244a0711ffe5d02b905d80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf1e43472b3c45b295ac0cb4378725270bfbd24ca499e151cb56136c33e3f3978511cc4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1513daf5cba73e9a90ab16f1ab4d02e97fac71e68b1ad2cad879531b8ddcec7a6bbb2429;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcb82fda4d52793b3b47d6fbcc133e43e0b6392ec4909b9a56c8c1d925eabf1ff4bb3f345;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ed86ba662500eb01c869651cb1d66cd2e8cb6395174516cc1f416d517689f9b04a243fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h46def8de00af523148a5e3af4d9a836c6dd929a715846ff733b5e84b08c7d3eca85d9f30;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a48f7414e351a4019f6f085e4e24a789efa18d4bf99a71fda029ea32490ea128d2896eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5531aa802bb8c52509bc268f8e2c05c03a9ea9e31d13f2142d4576331c1e96472b0af519;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17792edaa7a45f2121df837ce6d7b80ec520534f09cb45039685e788bc288471f6bfd059c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h76d61e5979425ff4947659ada8eff11fcddbea454083ee812e41f2ff3f46a4266f15a85d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1ab4a9dda6daa475f1f31d2ba19168fdf63df0a33fa82bd9e787521da276195d5ed0e8b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1529b23a941ebcd185bd622cbf6e60ea1f082eb4f3cbf617915d10bfdd2460ee321b65b21;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d6e4f874dc3b08ea084f6a1e290972095dbbc8eaacb056aec522317c879ba8c4afa7f90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a304f727e974d15c8dcec21c3bbb0dab9c0402687b06e68b17c35b1f63ec167bbdc64431;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h82a59a32f3a6f9fa8f41ad930668613232663d1b5bb36d674566541d8e738cc07ec515e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd7d08a901a0824f942cda06aba5f2aa22fba29dd631ddf184791f03407745e50823d2149;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f55c282bc838e5b958a67ebcb6b16739fa11276623ea6bc6c958cd19b9c313850900d670;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8e9067b2f812cb6f33f328c34d9a433f3fbe3b89c8def9a88f86b555146039bf9bb6c8f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1caede497858054f03272e3f54d1896b59ac80ae1bd109e3e6e47bbfa2a6f691b28904ebb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h115cbb9df4d6a246764ef8895ee384e1ff4209ba39ec852acc74f5d8525263ed81dcc67ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha55b7bdf61a9a850518e2732f2a8eea80a9c629866b927258245e06996caf97615e02f1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14f85994b70c602d8105b0761d53c0767b4fb9bc0bdd3445d15740b40b6d802432bbd707a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc3a2a2c8394af2be9a2ca968e74f594c6ac3a5ec49a4bb44003a0aa9f9de0a8909a4a4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h44f43f017a53ccde7c864d6cade88d9cc842d9c134f58e4b8b03d5752fdfe211b8ec6aef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h174bcc9c142b4fb3b9d2ee13b7544cd8b1d8f30bf25087b52928caf299de4619fef5819ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2a0644e2b985b2cd44d2f4d282eea16777fc188686a049d87bb1718e2a1c53d145c079c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbd9d4e58193e5ec88fe3abdff1e601c119617b660f5bfc4ec64704bcbba26e544d5488e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb95914edc6be29a7a13ad55fb3da6b246788da0ce6aee2e05530b773cc1273c40d75168e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ec3af39325b551c57a5552c210000c18f74472d540f22e2baec04cc070bed2e10ae01be0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h873119fd09ac9a9d1c22f9fefbe0def1d176c03031f7e52814b5a63a858c8cdd759ff7e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h163f021dab1f45df86dc82b5cd47a03b533eb9f339c551881e5600b821c2e70dbebe47a34;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h171e745a5f1d95dfbca1e0241ee4762bac41670298cf2159d24381b546449f10c04424136;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e0954e1d0fc4aa64a10085ed42877377895addc519fe3f9946c4fbfc1101c11c828d83f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a9f66dba44ca52181664af723e869c53a7613f4a55278db73d9d47306655f062062c9993;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he26cc4b2f4c26fd62723199c9f663a37b70b495e377f97681b76f67aaf472ca1159748d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b534837c645149ea088b4145a2215619ea57fa1f84d4d69a3f1120e0a89333c941541a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he3769a0957785bbfbd8a2cbf67db0d1a9e5d5d7067e7e5a3d8b1c611639ba6cc6afa783d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdbacb513a303330d2b868915ca289e256f985b993154312e020457df777f68e2f79e1b7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haa70cfdb844a4b63ed3e34eeee2c52934e906a1a1cc95f99c622934e703c57f636907910;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11829e2f2f278e2539e8c03434e766536e70235d1e4c724579316ecae7c0c52bc37d387c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a11761925f23da57a321e4c86596b9d75e897d83bc87126d8581b6b10cf6be57bea5f6b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14d4b09c5d0c4bbb148276bba2a8baaf66a244e8487b06e3d3ed40d3d90659e08b1bf1c15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1935e3d920a368941cdb3dfd2c7d691238f11e75f36eb1724b7455aa6d112439a16ab5e4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17718ea959f7dfc2c615a84125ad3181482bacf495bc6734946811248096c1888e431c46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9ca151777720cdb2f9da2f499a72dc0e6e1a18a3af2283ffb278de1dfc7b7c27d0437f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4fff6afd92052cec51598a713bbeceaf529c2dbd77781eadff880ef66a71fdce1e0d7e1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12decd080a7656228cbbc0c0dc48dcad975f2ac71a2e19901741d1b19542406fa6658c223;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162179d7838af45e7a9f764b69f2a45dea292c12272f4d873eac85f167cd6b73d3df6385a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e87fe4c102719401a49a670ab5b0c93d3f9a11cfd25e651090035534a7270d8cc1fd9798;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f31fcfe49677c593039f810e2b65714567e691ed0c3376c343f04f798d0f51389cd296f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h100ac494d10898f443e66c10ac16c638699f91435ac6533d23c2b4c93ebfcd2fc6ebd3aec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c700461e776e76a7c77a0f5a23de932e3ebfcc44ebaf6097668ec772b23f147658368c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he2e2d769b02d633827b76bde7bc31ef703b04433024ef28506c43756815501c87da6bb3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h139bf13ebd758f6b3244d550935ab92210719ed08ff973fbb4daaf6b3ea4674897dfbed86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha4a472babedacaba31114ea788acb4a0633d8569029837c6b155d545843e2bb6c244f69e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h192302751e6ee39385668d437946962f29f6189a90042713732d167369d762550cafd4cc3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7ead3eecb233a96239a0b60ac04faf6da83898c18b852fbeeebcb01a4c3658767ff53353;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1455cb57a49cd8a13f07b67ea10de65b262d5ad372590d92d94596e1dce5662a5c430d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c16dcc4aa7b82dba064ed856a7d2c7a0668bc715a34fc66b5e55482ec200a0be03e4bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bb9144f53ffcb0fa5adf7f807bc58774bfc411971b1dfab5fe36e22cea29861f2ba862ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd9cd489d2b511c475b18c63e1662d4fd110e0b721816fa941e7300c7c5fa3cdda6299;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6e22dcb12616cd1c3da9aad92d922d68824dfa194cdb8d23f22931daf79512db6100725a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h74a6df12dd5755df7bc91f432b3d291bae23716e3e8132a5d32fc93a8ecd4f87dd085d3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199576de4a097c58e1a1edac77f018a5611876c56e465654dc377416b42a13795b2d350c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha8a1aec604f0189640e2d6f9dc6c113e87fce6e6a539df475040f464b47e4e4b7390451f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf5d345938d1122d29fc31950a58fc34d555c75587d383131e777b9a4ae5671c263a97f09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha8e7d41cd9f4c361cf39c947174abc8c83e8e96e4e6885d97e764517533e3d003a83db88;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h143a56d226b555ad5b62cba5588c4b749ef3b2575c30a8fdd6a566b1cfdc368cf9f52753;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1191a555a700c538f25e41fee2745c63aa26fc6c868bfb761c4067c80e9533b8c0f160eab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h25d6be96497c0f29592fc9c54414e9be768f8a6c43cea12ae2b45d4f2795bebc884c1ba5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a291708f646bda359ea95039dba8c784a9c44d2774c6e47c01fd73e6248e2e7089ca8cde;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h179632e6c3e9dc26d7a383653da537ceac945811491db15499cb16ba8ed0807c2895bcba6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e87056e192a53a9d7cb9b35ba2159e522482017531b6ef8593e5d7feda8d7740b05d4e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf80068fea29c4585d2a80c838b945f08b4cd027f78a76e1e8a5657571c6b026454f6eb25;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1529eacc1a35e4758811424e108af5ed87bf9cf3a86eabae92a841caadd891b5de7c97028;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dab62ffd628f21f9a5e42c96aacbf1cc1aabd195a4139c055d61c610591c2fa24d5dc035;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6c9f450d51f7d15805691bb5694d5bb6a3c33bc30b5b0ad6834461a67362f970307e9ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b53c11f75831c4e9ac79d06c1cc280ecb293268d99cf4b8c63dc946ded9ed71fefbf30c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50144f9d1bf9c3b4a2482f60109df34857002a19802470a27f078b534bbad70fbde571b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e43319ff59af3abbda6f1c3bb4739f7124db5e7a7de0f59e0b61f0876abbdc8692ce5d90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcf83149b4912af84ea9f852f2f6efe5dd94373515ca642ff393e98e547bf51804f6d363f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h154162ff6666e9102b96c88301e603e17db3180ea938f49368a71bbee89e68d14518810f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h121facf07f4db89c40ba762d5f0aa7246cec39e26ef8f9c00e9ba0ee67583e2127f1c7dce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12386aecf8c82b44a7b1b277a1f9d368b58025e4f1b1cf9d33d1bc3e679aa75a401d70cda;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b4de25319a936f1fb135d81e79dfe096b5a8a854c838fd44cc1f9be580c30ccba227cd50;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he978ee4ee56a19e3a282320992c134a05bc72b2ea16bd580e0c4f361698784f3dd752679;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17b6e89ebbed8c2d40e7de62395048d295ced204ced98f89c9f4e7f7de9223127033b7aae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1412204c1458497d4c498e4954ed0f904e72be0aa5fc361438b4312df2e47c864b7276963;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c0c95c13216bd2bf5d44de2b44732c01d0ca152e9a2666b543bd31db67847ba15dc8adec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199aca5af168c2424b917a332f67d278bea8ccb4a47082fcc409decdb707c359e7397ba43;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a66f8620f8fd414909bc916b7bb48105e856c1151d48b589e35db4a715eca73904358f09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a24be41ffa24ff93237d8a18c26c7dd4c85f1b8a5b823f0e1d35b53c4ebbfcf295039e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h177ddb7a3d756526ca95618d045af0f0da3f6cd8dfea748b9c5fba08dc26f1fc108a53778;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1426385bd0d578092281ec6fa5ac4d09f62e5ecbcc05978376d076c75be82b82efe598be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51053ca155c17c64ce3e0be1ce48be01784e74dc2f3bfc725fb46ca11bf5f7ace6d432e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha01223640d9b92c32cd6d2610f4cb5657315836912b65480a13764a3376619afd16a109b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12aa3bfb1f2469af3bd5c6c004cc997d4224ea2cc453b0ab087aa7d0cf7a70df8c05e1a26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb63c948954eec4af5dd0f4817809e0e8d6aa709c09dacc5bd856a8a7a59d449a3aa9fbf4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13df1c681716a6a360e68a056964bf1c0a0564313746d711583ce828b622b2cc088be9425;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c1d7302a977892bfef97d5106fa1aa2f0469f039f7b394637790134d0a1759f6e7f34acb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h129a24e026fea9a166963ed6a40272c98068e2ee95b8aaab9ce2255d85c18e74c37260bf0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ac131ac442163593ac9bf71f9ff50d8430c151beb86f6d70011a92ccedae4249c4f32212;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bae6e14fe0d7645d7c27e3864d4082c7d33caced344c89456db4263a739d92f0fa9572fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11ac8ee54b23bdbe3dd14a8fc3002119b8eac5a8d48eb69aaa953d574809e5a2d4b912b1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h96e289cb5ea9b3f9506a81b9950ce416fbfb3cdeb352d676bebe06ac16b729e4c7073e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ae3aee5caf574791a20a52deb1e5109178e18a6d9b8acfca47624eb46ff165858675f3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h77f5162ca3df1cc5405b59bd8b9afd2dca10149e3dc29054a72fed65810f45c334d266d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha882274716415edb66d71a4098efa6691c558dbfa6ccc4f44ec9c3789902b962bfce0ffa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c94d885e05a43fa2443007b56cc3466aee7b2e931edd6bdfdb25c5edc0569ddd4a8dfa68;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b56bd49354378ea20ca9f8216c653bdad358687879e2edfe6d8223bebb39313ba00cc65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee15b60e7bcac4433829e9142a76736b16a348de6466db5648c66bb52f6ae849dd204bda;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7451448bde2c40d2144276cd7fedc48e0c2516c7c8c27a9d9af09444705fd59871bb702b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'habe065e1454bdd9e4570059b3107ba82d2f9cf616d181e410c6833c89f8b1baab4d64593;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dcedaf25897b4d520c7a69a5b8b7b56ad991391a94d0b55ab18d99b94ee5986446f510be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1125818492298493bc69729136d1c3bbc537f3ec7633e204d9cf93e1bd546798346fdd5e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6881af4ca53130f56095731e20f5d3515b56686ffa3330b67b23fb2405708e52b016a6aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef169e3175c9729888717f4ab32e7bddc3f0c7064eb0976837f7b207d0edb1c0e384a537;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a6fc157e78debef482c418a680b799d8aee086b57b04a9bfe2fe2d0f51886ab1c8052951;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ae918015adfcbd63d00d8e88552ece04bd956720acc312e25c672f53c607acda3e4c59e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91fb638dde217c74212189da829a6d72134af6deaa4d20feee2ad5f437f3be1076973fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd338ee910b1a4e27a3206d70d674e31a921b07ea5153c0f103ac0d4cdfda773a53923d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc6821055695ed8060df9dfb1ac0c527053b87ea5d8bd0f0cfd82d5f63345a688ad658c78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dbb47a8629532cc76d4833f5d1f0971b6538995945ade0ed97a94b20a06d607af7b163d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c66cf3e082df8f9d40106b29b4e28bad1ba3b8f1ea928cccce59b3c43b6e14bedbb4e7b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be2ff6f7835184f5d95021f85213c4dea428561f94df09da28aef2d6b250e3c0b95814ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha01838f4ddd44c77d2f5c690c96bf19ef5831de32deb37c91f7942a3749580198da3778;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1fc4bd8421d575bedfeb93ae8513c5ea1176df5669a6bd6cce7f6c53325c80381bdd7de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h143129dc3dfca99fa237375cee5db72277a42a3b408a4a275659e47726e0dc42e107b6a12;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd3dca90d001918a79052f467774766556cebab9342a29881143502631c6f6ccb16cc0581;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bf1bd85856dec683d3cf5cfa921e070cbd7adb3f4651164891bd7fd0e5c721f6df0407d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1526f553963141eec0b3a8a96f63a031a695bb16dd7a554b85668b32c304e34b8de7f9c94;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h173bb4f17bcb14aaf9432eca34c1f57c32babe67f7031d36909d3ea502c28d9baae69bce6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h70eaf669911a49307c70406c14ef2ceba4640372728d5f7de684a1b464c34b4cf8ef26bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36dc2ecd8139173ecfd9d90a891fca678dbdf17b90ed4355390d6850938f234818877732;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc18b0fffc34ff3ca6e0023eeb62a38c085b9ec703b0b6269c8ecda08d6739d0b8edce27;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h184b63d47bbde70654a7078dbbe38aa7034783901e3b6d6ebb0884f32e88035e4e8aba38a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5b949cb9dd7af6206c11cbd87a70109ff817483a5bf21f9b2fa2e75b0a3f69a9a4485906;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187b07ce39cf0ab6d317c2d1d224425cc2b9bf44b83935c9376539a4e51eb53644e86782b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10a3542440017fe6cbe6407db9aedabb573c1db2235b5b63c0e2779e1c86ebc20cf3d962e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ff163b937ea577db90cb0da5c99b8fa3f375ceafdd1c39535a372a6af9647693a10ed08;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h373601188c49156d04153178baa209c8c5b07b622265e335c0c7f7b8b3acacbb077d1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf8f531947caf939c916d642fa0187c4949cb83bb0d583fd87dce220ef8e213db3964e650;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135634bda6678a090964ea4abdd3a7f26bb286f06ed256dbeaa220842aaeb6c1af5163627;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc98525ae3e13392a468a019dbdd719f0f345fc557f645114af72c9c4d77c8a061842a86d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h445a78acd1e905c1ccbf25bb002efd5afd3f7a7997ef21478b4a6656e3bd8ead508ec39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h122cd1cb6ba129c78de03546f32940336f4e9512775ce3f15cdb062d83003dc990b3b6f93;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1025d8774273a07d4c48273df0f79221ee09cd0ce9f3c215c604d46b8204471d976eebb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e09109d9788fd51eccb149c380d138c3025a18deb9760f2b57b9cf463f9859de210b6d13;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e49c6add5a782f079b7b5f57911a117e73c04566eb87fd759ac10330e6e66395356ed1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h114161f956bbf0bcc3bf7c229860dffca4558a858351b3c843ea29a8e874786d5b73b5e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da181f06f2e0dd64e4b9466901293d96c0b7628fa6f7780fe98c77c8ffd7080570424c58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eca2c880065cac893b872ee5bb13fa27eba9fd939d4e6e51c3a120e9490f65eaf81a8bce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha22cc8bb998984fe2a3e95c785020a7be05dff32f8e924139f6a2cba3efa72a51db26ece;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4ebb58296dc39ab628d2f5352246b6155283a11037158d780e18b210cb480fb345acb006;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11345f359be713e380843d01d07ce6f10d97baeeef4026ff0a0e1e6f45bf0b031653a5d54;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcef7bc6205709a5d515c99cabc71bd9aaa02b18417eddbadbf151d80e87bbfd66f65cad3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a1299cc4de58fd90fd627871edec408ed92b9fcf4f13376c35407bd2fee140d43957743;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h45d7fed8f5dc3887a77019f1fb718b7490c475482faea4d7396f3724bf5994ff83a3797b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb78d3a1dc6b8915d95532d2ea4d90fa8ec651f8bbde904d857b66c00d5fd6e14b6b3f935;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc5bfefdf43bfe3b8528f9a1e70a1d8d4d9339661418bb61a9e466fa7b5391e8ad8a552c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9fc35ce48fed5d0584c691601a55c3258638342ac00e96dc22aaab0ae8a739dbcacffccc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19992528d8eed4636dae45c33a67a09ad7caf9632173c52b348d5a32dcb45b6b6eb4fd03;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he03223deb997e63527a24361c1dc397bd5de724ab97cd59240e3b44178248cca1904619f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h168fb6936bc988d7cc7ef88d43e582c5cd86aa4196217d1c4b57bb7dfeadfe0ffe6d2b4f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc00c2c64cf47aad6192d46d1e43a3790a867dee280f0c6a98f787c7defdbdbcc6c090504;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19532f0a5b4814b88a55195817cdb20d5036241ea116cc4e2b7e754ab23c7ad1ddb11293a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16067b75f265848d14a6708656ae08b0869c58f164a67344864b2f8f928058e8c72ea075a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19b9cf22a37709ea6d9639e87407bd2c08e71bfbbd4030f8f22cb240c675c665359b315c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac366245dbf7e1c46df8331fb33249db47d62883470a9a46ed5a4d4ae81d31bab02054c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155f238c21e8acabbd7bad8b1ccd0664a3f976403da4337ea973f4012ab699ae8b824bbd9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbaf664b0391cad72a83f2891a23a4d23d7548d5f76390495c55dc5e1bb65c2452df16ec2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h152ac7e2005854b003120317f98de7a14fe1d4c3c0f8abf8c9f35b155a6200d8692d264ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f0b5cd282a3f8fe5c9de7c4dbf5f5b8f0bc711fccbaad9347c82c8153ad5d10fbfee667e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17a5aefec969ea84e9a36f4f9b21a031271c567347b4b8c40b15825a0d76f8071c4ad30c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9b925eed8f8cbe8bb72f1398a54a1fb0dd8815ecade7039338f89607bf8d52df1d987c6c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hafea436928298dc7906baa267f506f37f6f391ec2b35108600e7fa376f9e7c7e4efed9a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdfabc4b4b07f331388f9268a1a89b7c886df7316eae88fc8308bb539dbf9c1b3319dcfe1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50e12cf38d57d9c0694888f59090d57ce0b715a601791a33851810bba35727b48ee1ba3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he2108a00e4e3d7f83e720966df1a99ff816eb2284987c1460c0b2cb3aa509689669ca7ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h152dcb6a3cda095eb3fb3dc5ddd1c88b8464b811c6f798d121aa9f6dba9703655d94f237;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ede716ba5150afcf89e15762f90b6c9c71f10d2a2a8061bcc391376096e6b79aaa7cbd7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h84ccfae7c33b76faaf5782d6b276513abb523ee46f190a5579d84ed43d70b959446a25aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8b1340b6cfbe37f38b4ded55630594b2dca149552d3c269649fc63abe3fb377b71368b31;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2c9859ab4e2c5d90e9def78c2882b272e1abef417584d0dc85ab640cb1b23b37f13bdb0c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183917df5ccc1cb4e57e2d8c57e5a98269d72a500d3ccbb64b903e970760f6437e23a8e62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2cbb95e1513c6e5c1c5551561eb5d384fd53937ae0003b225f3e04e8d7e675190070fe4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec6ef2cd53a7a1f20afe3318d5a5ddc935d481838b72c8095337978c55e16ab8a21b7826;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2de383377d0fe0d5b8d45f027c6d486d8d81063e1d887e31c25431b0e6db4c5e22c3992f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c0e88577b2d119a8237afde85d5fcf0dda238971edc8aa2385373ab22fb4fd672c4af3c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h462e8506fa11683cc44098443efaa08a4fe3bd6c0702064d13079f9c704e822e31d372ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18f1b60f07e15a460b536868fb50918eaa469368f7b2724ec594c892010dfd4207d45bea7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1faf690bc9fbccc3bbe67d8c7efb8cfaa35c80846f80f10b6c2fedc7abea5cd095dd1a02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9e5e427f819562e5193ce60695309139562f8c73fe2438a99231b0349036964bf99cbc31;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d3d25951be3ad42cf50d24f2cd950f7e3f36ca5d32a708c61fa7dfe1657b485648e18ee6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18aec53fab9bdc64b7a6b2aa4d9b65ef13a3d20528661c610086cb3e1e84537d26b5f9e29;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb43e8669932096a9e2388e49e0a57e1beed496c5f2c540fe93eac38b745b018e19250952;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12bdc16bbf4fa21dcb40a9d32c33c41d6b5d8ca7ba19e8184364ae64934b1e9c80f683afa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb78d8115f85259534767c36c680ef6605211182e44e34ebc17862cee1ebfa7d7d8dbd2c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7cba60f6ebc9a1605489f41e3f9180bae606c44a15761442b2ac0b17bed410d73cd04ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb8f9a93913d80afc501fd61179c6e852625b85a47d371cc3711e8ac3c276dabfd7436b9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36b8e9b15cc94c031f0d0cf6cb31acf46b33ec45a5d6cafb52dbb7deaab87fff0f5c08f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7d5b3fd822d2aa070c6651cab26e957a68de1552d8ef6043e84354576719bb4e91ca4a02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h857166e2514b542c48c79caa707e4b725325a6aa3b33c7975d238b584346fc3aa9f0febe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1081472fa5bdd4a5de701b1e928edd79e4948da34582ca348e79ea5141824af78d131a1ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c0f7aa7fbcfa161f5887c0c917f5262ed0e45cb4628db65c0603cde85b327d7f19eccf6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf4cd12c51f7af14cb22758cf50e6774d89b277c971be8f12faadd88b51245d7c289bf643;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdeb6e39fb6d1da4a84e5846b37f88869dff871b3d27e718609f85f846cda8ccb57053681;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0f293c05e479feb5297730d44962ccd3cad56a722edaa43b287bad0239e7c7dddb4faae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd5abaf7c0e050ff3edc3247ec20a264e6e15bbc36f67cd3d68aeaf1c2ab8c5fd0aeb52e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10edbba4c2afcda431c77f0030af89db1e9d2158891b0372b0ab2f404247fe6405b9c5e59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h35488a880e460b8adbf8b11f530064f9ecfae2862cfbd52668ef1b8298826c0498002368;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17b9b18ec382f4d52ef4b56aa948fd06908f052292ad16c25267ca68d2d910157e6f96f4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcae524a30ddbdbe8abc75f427c95ff5a9b3d157565d53f1865dcf2dcf7261767d696325c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h634b4253e48c5fa9861dc9146583dd2b05e985f1f3e02656f28e6b1de49d4ac66dfdb14d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he94e4d916ae912e8395ed66b22c41ee8851948953952ac9a1792f46d6378fb23b2c22525;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1b3332c5f73ea3d4c4a414eccc80dc5f8b4e94b5cdafdbc6b3bf912b12e997f0b67029a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbaa8a3fa7e49f085edeed1af1e8d4c248f69a931c71e8dcdfdf9ffb17c2b6a12556aed82;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hff13eaa2ccbbba5fbdf601736f8b3a37919517395168e23e21c3f6d89e72ca8eaf887a72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h180511dc9d739b289b26319150a46c9c4390a9c91bbad1c5a907a1312fb4bd2f5610c9a5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e6d7b685b6e4c9dbaad3d7864cea6d822626b2aab613f74b88c59406059e0f7be4349ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h63e3e57decce2f2a75f245c0638e023f2e000e3db39b13b0ae8abe5625a53949467d8ab2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h64a0960ba3b5abd538377fa6dbaf880f6f20ef86eb14ecb19181d4925db56c9e7423715e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ddd6097f12ba1b3ce310d46b882d459d01951016d30e0da3359ac7239d16ded4abd1fe75;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4edc883fe3a68cca82342e09e109767699102c7d1d8fd25fd9965351f0558ebc9d669116;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9d57ad3332801a0fd3c584b1e6155ff2764f6ed3eb531cdc5844a38aaee824f2c0df4d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf9e2b57e8648f988760a79bf178ff9f51d0a39b85a6dee107abc19b11f99f5df05ffebaf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124179c6fc35acb7d74d055f62f0839e7153dfd0d1da7d1a9bc55816039b8734b1be937a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3f27bd3edca778a270a44e2e8647602af4efbf43f3a5799dad0c9f56d5a11852be13ee1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h40a0a98d33b0850771a8d6ac059650bbbda06b15421357c7f936389ac720bc6f54c9a115;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1003fefcb11d82bf3cf1c73fb1863e2fbacc512190a743cb4824fbb3dda46f6fe1b0cb57e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b52122033de94c719e8c469296ab480a00b13bb3a863ed8f8bd1a4cd793b8cbb66fb344f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e1334b8954b07bb7043d96c67990e339b0a95a68e4c8a68357b44cd584a20b2a6144feff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15ab736d6a102d0f6a5d7d221dfd8fc641657cb0877b6bb495dfaca80c1e2f07eafcc4a5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h160198baf16ff887e07eb91f55d1dac56a6141ff696c4ad771f01ee11f38b1e211b284ebb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h48902097cdc57d3ae74c12d89dcd5643c51c4b81fe29ff7e568f2a2bd510c1c3708a774;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6c5b9dc11769d91f85c87bccb9bfc984dd6b6abf7950cacba26f4832e78985bca925fd5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h76f55948c2c0efbc6803f22a230371f84df7a13bded787e37ffd0efe23915952db98d5cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h75aba15a238dec28d6be9691af98a96e479fcb290acac11cc933e96b6ad0d6d7fcb6ef09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef1ebcd83e66c34b8247d4cc4f4795b294cc77419b89f85a0d1914dbe2c5f79eb7c50eb5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8e00541a24ec647fccc4cb7e85fd2047478d8dbdf2721046b14648754eea1247eda97ebb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1df2ab1d7c0599cd62df1ca47970588ec0b340520e4265a6820404a16382a024f3b2aac30;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59271edfd9b85168a83729a6c84d930a29ab68cf6d6fd435f935f2a4a5bc788c0b83c20a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb94dec871e2f860588cd131e35e1d0afa5bacb7b670b52e7c58e8c0e8903d9c3dbc4267e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee91981be905ca050cf1aa6f1b05cdeb5451c41d89b0ff75a964240b61092b839057bc8c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h160973fc2628f5c97831c09f353cf652bf077608f4f4a1d9aca93976f2056cebd2f3935b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13bd59a05e74f09fbde5ab992151890551fe2ab2cc816aa51fb854b7d707cb5b3d9eca62d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19dde640ccfde2f86facd22e6278a6f3c0aa40b7556cedd87d1684b327503c96e16f90854;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb04ac8f94d84794fea4fd0b19e63344779e4c30554a073ee307d80ed24808611a8b28346;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd49ac7169d3217ca196a5bb61e0e8e5f451616d78719c609aa4d550ee749fa92ddd6a1c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135a6eae649403c26d6881d311f05916ec855cab79116a6fa9c9f82ad6be114456e696562;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1abc625b6ce2bf0c04cbb2d43d8419d8b041901060a108c9f40a1ae5448fd47b9db7fcdfe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7cb8319e0715e87318728bf031d82ec5ce15cff00835392abdaaf5cff0bc48f272ced0bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdde5b04329d942dcc876d712a8144c4aff227d5ac17ef4695b4d43cc11409e786fd37302;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h161f3cac09ac485d9e35ad7493782e850c17ac00f2017b57778be3a809447ae8246f947db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4ca569793239c5a784ffc47be3dd154c064d33c0fb0acb0f7f39e0e7fea7364fb70e80a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c1f7c900a911595950a178fd3b183c76677e419e1b2c7ece9ea3788b471505bad03605b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13b0a39cd49c709576fd06f13fa1833f99e2e069e8dd19fb72b421aa4ff3cb922886aaf80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h25363e03492155255c65e4ad8b32f8dbf6034477d84cabaac0e1ab3dd103da6113e4470a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16511018209c5d4756cc2f207561acdd5febe7da5bef6c945dbf2c12539c1ef4ccb13a135;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he1ba6466abbbed333f420edbdcabb5718903c832ee4f46446cb2fa8fd3b45c827920b450;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15c3d6c6ed20d876928ab17a470a14b6b5dce828f4a4fd931ea8d10c22968c35d4fc312b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h52b5d31d9c04da4b4d0de07fff99fd1ad97197f5cc3c52bef94ad815ad0065abbeb4b3c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1184942f6ea841211bc39cf14744b83012619fbea04ff9cc43f581f6e503c8e91672ce2b1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12bcea93f61ce89d252340b8f6c3ad78b09c05d40670260bd4a30979ccdcd6c80ac80ca34;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ec83515ef41f12b2242f145b1868d78dcc44be0bcf4842f14febb61b85c32022cb0dbc15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c536518841c04eb7d52996eccaa78dddc57f88102b411d702171fa11228d35b380e5625;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f072638f1e45b3fa7636ce460add67b3f7452318e1e6b514d5eeeabec6d13003e49d5d43;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13cc3b861fd3417a8b466243bf2cb36f6b80e1730eed5c1996ccbb1aa49ed18d9c78bbdfe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e99a6bd4c5cb9e214a6ec129861f943cb3be81405cd7946cba592e2bbfcef67b96019e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38a55d3611f57519aeab8e7744cae0ec9b4feb873878e471d3f9b46aad339305f17a4fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13936beb8e045b4fb156f79c110b8d266655b944cb8bed2f363bb04b2735a598ded683f07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h119d977cc6b1ebe39af59746494995b85f1e72cade9022f89660da8563026e58438457034;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18565534f6795da7a35a76596bf89d4f51a8fa239979bd554801d0daf1df0670ada2a2cff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de8363e6f9bf8bef4dd678a80e1a0f09a6451c99f7a3903ff7963b3612f139165ce54b2f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f08d196b9c9786e9764bc75a3c533d6e4f8ad9caf9d375fcda1246b24ae3c5e45f7c0587;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h26c264d64368e4cb3044c3bf0539c61d7e4ac5dc140ced72c58a76393ba98e2f143fdfa2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e6e2c70624d7596885c4b8df2277714af4b3db39e98aef3ebb7b032449e74b098c19262b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8dd4b6c627a19f89c219cf04b727d3d363f0ffe1fc9d22f565ce1bbd59e306e40848582d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a5a022563dce57210747b9861e4fc8256c8158c2d9131d745616056b7ebe156b756a87;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bbee9cc20fd5bdee263c5ee3d1e0180d213660d2e456ac80d407cdc568b004bdd9a980c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a6907af11454646d2ed48a178c2724bd112b2a5d586e09b16c3d424848310058dac4428;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h81c254c54280a6fdfe957644ed9394db02142b7ac81b3f0cf4b118a9652c2d6365b89cfb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hebe511e3faba41131b01bb09b73efa361192029088e2089743f1b771d7a2cdea164115c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h927fdc7fd0165586c2fa240b3df2e1f3502bddfa8ff67d6c8de86ec807e5232a98ed3949;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h123ca49441f522ef7b4188dcb213df3faba54bbf8ef11613347784dfbf5d172b12f3cd5e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c8d55725f7085840af0de56426353a9e8a844e9b0540751bb752cb419c0e37ce8f9e4df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199671a3e039a936ea5e381ecb41478e7f008dcb3029c83324fdb61e098254f0ba536d3e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a21ef9b372d207ee35e6a4da4fce25a47583ffe559598da4a997c9445344524020c50796;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc5756636d7dd3fdad31fea16bd615db9665957739e6b09fc851a012bf90ae48a8967a9bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h76a99215a4ee0d46d7f70922625ec850bcd01e87ae430288086dbe305a4b9688ee1d8a6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1659cef4b928309b29d5c6dcf24f6413b19eb1ebf3d7ffbb41fa9decb153a1660e20fcbe4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8eb0484f1055fea95905b18b048492539f33bd1aec801a676f35748947831be0b7b6306a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18999680c62d63df098844c43275f53791977b5527e02c5c0fd4acfd1953ee76b23d724e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h103f14b61bdb87a065f14e63669ebd12274bfc5a350065d68eaa38003df4bd52b17758f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h119361b0379b5c281863d5dda1a2818c55de83f394dc14156d1beb725826059c029399bc0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h66dff1315caf3a3eda6a5ab90ec14a22aff5971daf8d1f05941a770634a10e1d8e6b070d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e079d3fd06f65999c525a4bb46703e202492a50451a04c2613eda13beff1941142cf4811;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ae1862eb15963c26f3aa980910ef621847eef2ec51592b3b1d6accc989317ecfd5f11031;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b37dac72fe1552d92908f5b2c19b25375cd744ff02511f55d207cc6651c39b9fdc277b2f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c28d164611e10cd0c7f44efb840fe93a1b744af0affcc8afca0965a0c1f58a2077ebf4d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13199d3d6af8160ccddc390885ca6acb3e9d714147c947a23389cf4583736bae06f513744;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h32815e1d7fcacb8c1cc0cac1528053983916f441653c58faa994562e6c09319908a96b57;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e81e06bb5a2b10e06472cb67d3071f6a9168a15fa2ef306373e479fa28c34e31f78903c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h512deaa1b38da694b7ec87abf4253f4cbacc825902560e7638fdd9d1b16248c540f3ecb8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18a296edfe39851cdd748c6a0c540718b6b75e85b32d71c7e7a7b26d16a9253444c5fc33;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h175b5249b482e9d56ad249b8b931dc4fd168e89d13ad76e5315892ee068647ec415f84c7b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d573d319a7b71b37c471f8739cffca1c9a7cb03127139c4778b42ad048859105b9e2594;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd6534a35562afbee8628606bf4183a168446835b0bd4fe6106a3cb6f163b99c4649fd5be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8738e80b1a656faf981fe8b4ea78b1027eef49d4b57be81b12834e9f7a5140d2018acdc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bcd5ba8c4f0d52bab62c28e7938f080e6aacaf6161ea3dcb320c909184d1007c8e710f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a324fe2b950d4f75f2715abd490717b46e8f8f1e773243e9c8a6668f931a3fdcebfbd77;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8c83590c18cccb67ce893864a2075e5a68643ec888d24c1cdc235bdfd4fb29a4f7bd99c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b8e0e59ac1fac16d4e103ab855808bf12185b70d4e59d8befec484a4414f6bcbb978316;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h495a03137bfedefa1361664b2245d99da0ea87c8f0ab0fbab99168d720757c87bfa0c501;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7352a7fd32f2ab08e47868ae17f2b48a8e6c016a6f7b5f8def12319ad42bc55306e437e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d9d25fb843d95768b46b7e615f9c3abc96c3af02d46bd804aff82ad274ee6c2c53064c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e88feab551eb73b6de6b50b2719b8bdec381eee5b99f5229c13ad06fe76a5b85463ecff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de7388c9656a3264ae7f02b568fe6e2729d8e1a9d483bde390e68e0a03371277e1b4931;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha360451c4bc7eebba6d3cee6908ffa7439feaa373dce1db3db3df2dedd837eb2feb0ca4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10ae5312ec9b98d85a88e5aa83085346dd8f20cb8c5f0a4ad9834f8d689b90971fd56124e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f545dd3d709a85267630cc33342a37a4dc39d7eaa5398175ecc9f2daa3d1ce5b99dc5617;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13ecfb994c9dd27c3f67a4cfcd0229e62daaaa26d378c12556e5116d5c4200d0558173af3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b56fd734a1b70088362c2a17c4a47ce786ab4bbe63f1693cab58261b4111a0ed417fe55;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8f54564ba953bf4a16c2d397e17758b3b176b295f8d093a0ca9cc0a6047e6135b1d8d945;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f39acc5adc7fcb66cdd1c1c038fd7a2ffd758f8fa9f52fb30e7bc6d8155c2d2622c20aa5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13689a6660981a9243be0eb65c0ca125aeaa56f259ca811180405173b7544a7294bc9e66e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e481e9a83d2f26827b1678d8f535838702c61320415e2f708a7ca61abed89ef43175af38;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h899c343f9cb11a67141b3689c7003a5c80e7add37e01c875f561c800d0a3b6ed1c9f6680;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a8922d544c86759f292b3cfa1ebe07a686bc3ae36074015a90c7a82ad56a3849879e0c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18334120710cc9cd4b624a3d13ced8a2a616cdd1e82d5a4b78ead3fd70e2ae8a62a203608;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbea9c95dbd0b25195c20b6d62c320d668e47f9959e5809815f2f2b5e6da6c63cebc7629f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6c07d5cd16238aa2c6716458b30b525824b233ca9bca67d1af8289bced19841c9c400610;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5cc1d9146cf02f24c08b9262b6f562939d38cc211292107602a11d3db7f05d8ac389b4d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h159d8ae7196e0fe9a552c578c83c45399000c58772a8f1d29c39edb7aeba6d7a2a2e1643f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h827aa35a9138b819f84b955cdf38069aa516bbd6aa8d0c4ff3725606f0a37e8ea9610997;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb8da7d0617bc175699d098ee1f90de0f15c262e239967679af3937a446db3f26973df7e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1938cb8548aee5878f48c7ea61ae8045d968bb54b900256f2b455a2242ab2f92f0675d748;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da77d305497461342e1c4989c85a99ef04de61f9e44e5f0480a0492b3dd370c771788324;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12290c10f365832f402d5e182c78fe0b5e117cfd0409fd5d6b864bca7c5550db58349e7ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a80d68e11cca4967a9fbb13984662169ad475147a048eb6cd3774b14995e82fc1a3c470;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3ecce77904bbdc28c7bbee7f923103ced21d22871f896093eba23c528135f79ffa7b585e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd1856e50b2704e1140424fc432157b144e5f6408916fae6f674bf0c01c0ffd826623cc81;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h134f5a0f6aac83a9c5b14894f17091f15e1741575acd6f033851db73c7a5ae9251cb5a679;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17b7f8dd1de892c09933d4d2797d4a7a44a6a9f60e8ad8817ab8110e00fecf7abac2acae9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h281d39d92e7e3b4e390ef79e9d9a998f2722d1337cb0b98499e9f326d10f41db8df87b0b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h194ca5ea9ac30a932b96797164c0a82858ffe6b3f0b50d720a2be587cb03d56a6e7ab5ce1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4a0edd552733b5010366cd8c8e57b23fc70d62c8365161034b4acd3c2df2f27f4002f5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16841da19f36bd4775f3f355bc7e4c15b1c382eb2146e9c0f3e74d9c496bc64b62366a6b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1999e0e3132d8daa948042e611699ddaa6f5ca857b9573eb7ed1b9331a0bb87b36b9d3cbc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2f915df6e134b0ab2a99aa5ee94ebce33c6f512f9f341c4444108bf7a8084f0333acf48;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3992e93bcfc8753765b1e5fb96acd80adea1803733d3deaaebe07f12283e74294c9947e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f87798354b6803cda0e727556fb3c8b7e4682049f84b47185c531ec2ccd2214112f3f609;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f84b83dc5e07927aaff492a58cf255305fe10d577ac90f776cbac3b5fcf6b98b6c75641;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1662482b8da3200ffe7810d99c0cc964274360b66f31a66bfd7c74dd87915e4525ac9cfde;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h149480a90fb48cfc02fecca226fdbd796694aa5436b4771d06dee1c83220386387045f8aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14280c2e5649ce7ad9af117829233d31ed84859f049efbd6d176539aca79c73741b2396b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h497b5226b5cd93e935301b3c54e1437aa6f01c79b0bca649a13a3689448aa95320a3e375;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd90af54c39abd6cddd129a7dafd81bc5900fe6859d016c78daf41a6ba48387adaef52ab2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c622c64552ba2c96d8330408b7e2777c5ec3971cd5177a599ae9a76d941c9cd672d2b81e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98f58558ed0bb3d8968eea2c5c44a44f213d13c62b084f456ec67285eb1f8e88685c17d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c374e833570e52e2719d0d175d56e20b4d1996cf97873499d4af89543706e1c54cdd592f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91032d8097633b6f75105803f635949101bc5d40dd817e403aaf31b1f3d477c6b1feab92;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd01a5cbebc42df08ad2415d498a31e993f1eb892e353a5a3b12a0aa725a2ffe0113292e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc9969710c56f89c3d5a0bad95b551fe58f034efeebee801d05d253e078e201c4fabde1f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h831e49a2543c2cb508043a2a38a50cb7d8b0776ef34caaa5c11962522358079d5c7d673b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60024c69944b6d80b8c4feb67f9299e0058b0cf15a23348b1ce51f3ffb5ec7e71c6285af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1abf225f1dd8a6663d4aeb3611ef26bb9ba269f9a512c40ef6d51121ed5df6598a6fb8f64;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aea1a190ad47be50be964e491986eface1ac47a170b3899351c0acd1640f18f76b81b0b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha9b7a8ed1f64200ac3fa1d10f5567cdc6936bf9bc7dd5c817768b1e92f52f8f74f8d4706;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c3725429b6ea1ee6c62bc21eec3e7f001e01381205bdb1d62be5cbec56dc078a4fe98903;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a44329db0d14f4975c0700794edf425ae0cf022b4db6d1a1dbd61b0967981c4638710792;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13ff5df5338ba0a712fc147eee61ac9b4829a2053458d72eefa503384a922b56085535933;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4a2c0da58a5e34402a06ab71df4eb998931be0c432bd61001d294c6f6cd07ceb3f923b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eca99aa849d17bf68268dd4b08dac70a2bd341ae477cb338e6d5e00f7c00ab93bc85a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h703774ad384d91099085f4db5170a9cec20e3fd673c1bed39e04f6f9308bc1f5ff0de0d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a7697be06ff295ed9f7f26729b9c0749373f9bcd56d661b7830d77d48b177ddcb2528a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d22cc09f10c5d472bb1161011fa8d7963ce7107fe743d81bfb9f3003432bd21df62d86d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d5c01307e1e63a2d8ea29fed48eb328e2fb43fb0a3d20dd64b875d13c36165103316f15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f7503890ec75ce903dcd38fdf9c4a3666a15413887969c41b5ecd5f20cbd9cd547366e10;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h355d8c158743b6288575effacb95870e982fb4455cfd9873c516423ac69ece7ccac0aeea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h521e0f8967cd85a130d7a2273292452abe0791f4daa6663b62a1372ff3371b5199e75402;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13eac2c2d70396d1c2346add2b06abbafa48183b8a0ff4af7580b7773d75f27295e3486cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1959a9b9064e926bdd8b56e99e7e196205048df62de2a93ac749ef6094eb05b886dd995f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hab5e8c3ac3b0d8265fa2d1c6bbbcd1f29378ae6a3bf8b9655665e3afbc12ab0ad28fab65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6bb908c66ffd27a0f83221992f9b53c1f56f880c32526db92313d163fdb0d199184e5044;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b660f8b0a682cbff0108381b95efa783c89b54506d0bcedaab1f94a75d30b596b25083a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18bbca1c6280833648c92ffdce9906561dc061f478266c316028f6dc6119535927e9907a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hce4366db827c38bfffe1f93e0be81981698680b426316cc6aceef486bbdb53482ec701cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3da508626747f90afd638ad443cc7b4b3518f4ea757ddb4b4896bdf450e6a30fdd823df3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e3ca8b0f4c37cce3af2fe4336056f8a0bba99ffd074e18e019ed4e38a55e4fabfcf0235;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1870970ea7a7c117eb7cfcb1565ad87694c108f51f3a60d54463410eed3b852ce5cee9b9c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1286d4c87dc155015f3d7543ec2a84f57f1f77ef6b82192e42dc81ff28d634d18782bdac6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1027b0cd464872ef10121984321db97f7d2e785daa9791ae5def6d383b4412beb1d97a0ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bd94a7c2e79ae7ee6691de3b62a0441b13b0a5b18fe41d2c57bb2da4b33c99da8552757c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162849bb150b7b6aa6bfb429cd9e64fd99407df9467682d3b3941890aa4c380842f572c28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h718596a2d05751bc6b3c62cf718fee9fdedf46d70aef73dd1505dbdf5ea59c1735767819;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he9f0c980b4e1dc3a0a93b1d75e9397736e6ba69d823a1a4ca820be6ccd58ded718631335;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e837caaaddf48b785c73db8a759ec557bae56a70f53c32bb088991bc40205f33944d662;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3c8d9c6674e8788c513a386339a79c5f4092de5129c5b2e762ee35f942664cbdf057a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124d85e29b97f216c22e2407047e983448978562d18b6afe9c45e50fc647b1040396f8602;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183ee05df0bf675d9be0f5d3d0a574f559b7a482afb9f9c385b6b515a0ac5947b9cbf271c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h39d10a9f4128d6c6be8a2fd338c531b16d43b33823502efccccfb1226dbdef4e3e47419c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd1ed8a041061d84a18f7abfc32d0881708a849e975fd9eb638dd702eac96bc4676af584;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17bb8e1b6eb291ae15b4e5445c3c0fc3b9133003128b0cc07143bcab1a4dacf522b58b367;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc1009f01a6a4a789ab4d09f9291401db8e0de7d20a2669510b4ad83a67af3b78cf3a9c73;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h28beef7fd985680846ab14918f9bc670276b18879d9887ffd55c7f0b5d912830eb10d857;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d28876727edfdfa0c5aaabe7e5766224df7a3e8bd44f049d4cd26126a35959473f3ff4f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfccb2eb700537e3945499a2b64b9fce78451f6a437c376b80911e1a47af13f1eb9f12953;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b6212f0955fb72b90b04c5ce8932d92c3c384264600dfb0731e9dc5a936ffaac79f2ef4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf9ce917e46bfd9199b0134e9acc6c035708d0399a65b2f10b90d3a0498da07616d7aaa91;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h419bd49f009b44a64651ecff9f748b1ec5ddd3328d04c3abc61ec4e98e586067ce89844b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a060a35969fe44da330b96ae03fb1f320dce7101cfe2d13fbb08036410894a7cccc824e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf767ee54c10bd20bc055d51f167c51ca40c63c85ecd5f600ddceb3ad52292591b4833318;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b923d167211a3c53ffd4655909f8e2b53d6282692cfff6115939a8f2323d6110f7c06c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd4c33d20fc203b744f26e38c443d1fb6cfdac668502981575eb8445ab9168a200ac23a58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18c8a6d04e6bcc452480465ff2a5ac2c7ebde7a458ce633d51573ca8414e044822ed2f876;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h175542c34d2621d03fbea87f62160d4d234c16e9c0ed2ff41b4399a8f13495a42fa6415de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e3a99faa02780048464bd2ef642dac9549ecda9034f524a578d81858cad3cd13f6fc8880;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d8ddb804d4167a0a1a35113b209cb8c58751298191b0f88fafe73673cd14a7114181078;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8352e51aadbc746d176faeef3ea15f355b55982d207f2cab386c29c14f914e38d703071e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3932612c6da6ccaca3394fb2d5c84a1ea5c44fba31f02812fed1a44fc9c2ccc61b03b0f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4508108bb6494de0beccd1846e383411060c228fbaec91298dd7f9e025e326ed49ccbc62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16cbc42783a646b105b4b6d0b41096770eebf9997cf0048a738431955b23efed582f0ca4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eabaa0551f99df18be2832771dc95cf0bf387c6a3964f24d3d8e1cab22e7dc78197a61d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd5bd606f6ed1c3f31c4fb73bf1306ecdc077d4fd337e3719645efbeb6a7d05c90c21f853;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he3124dd5f967eb9f328bfb5e8cd215c091b442a7ae3bbc079ea84abad5f8489c1cd5243e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1daf9c53c136855b1e5ce790fee36cfa32031d86b657e734047febdb0f945e4bddadc80bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12187c65b32595f25f88a484349d2b0b2d1fb7af63f256499df90399273531a53a0c2bf2b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dbf89fbe2e16d065858e71f1590a0188ea882ddcb5a2adcbee474fad7429cb1d3586272c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e41d47390af79ac1fb68c340680f6906170340c87273be672e3324f446d7eac317324374;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heed62924d49298e2775f842f317f8eab9f551df327f1c0c792f3464e866225f5f11f1a54;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7c4e340eeb5ae6eb96f536c0e7bfc047234a0f36678ac8e77745b2b819cdbba93049557c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ada57a28b569c2f12256f0a5429095cc62d152d596afa91dd1e2647426316bb9fb6777ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c48183cd248ccac6530fdc54864940c2e76bd5fd908a533c2e5c0fcfaa95f2ac5ba3689a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d6d67f8a779115c791a5b72c6f2163b15630c8981b618b5c501373fda50467981d0289b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h830fdc4453c292f55e290d910becfaa44d77221da4db90e8182fc23e111616dd3146badd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1993f7124f8d6d10af2696d53226eb8d379b0c132bc78cc39c566363f253a7930528cb73a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbd04dbafc3b2b7c705ba7ca100511ffc1ec1f20441c18423a34f1c32f8a3171e77311d4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h196ed3563de70fa5b7fd3a1580450ea92b96c2c5c5b4e6a1369d8a507e04e574ee78c740f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdf697def29613b85acc2efbe8b36ea8358511feac3d7fbb9a993cca4da8122ed59a0ddde;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e656da045bc5a496b5fa1b136e6015cf93e566cb5475856d1a53d0cfab44c33e4a5ed345;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he9cd84f8e59b99ec090f14493b417d6f3d5bcbb406438e3b54892499ab48e9575397f47f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9accc0ed130d41be8717be024fb2bfd45bfe807c25f454cf7b55a06dabc132541f36709;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h154f28183c3a55c2b3fed44fe214cbb99d43320386d738844a0346074a4c9dba521f3b96c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e392e0e995ef66fad1b045a2253ba2e373ce56005ffb78272cf2254b82e9a4973cb227b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a3a8ebf10dc257bbc018bf3f3b00ed5067893b9a1cb88c1e67e444cd9030ada3c67d2ea9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h181ec44419154ae9de1b4bddc693886b704c15976ab3abbe4d0d23f7d0a433c5abcbf636f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h567958bd2898f8345461f91c4fb190f0cc30950a37418bc3c2565ab498ef2ac1c384c693;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a95f653b2dee7f2f25e24a1bc5b5d60b6ee6ae1321a77021fd4d53e5b1abf28773f58a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h62a21b5ec8437d7ff829dc9dc4fecc075b252af35086f61499632b2ebfcae362a500d1d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1952528bb2705515ec9d825887f5728999fae366ddb4a25b339906716ed7a5ab3a880524e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcb97b8ae8b3317893826640db54acb41748dd9325d6a79b317af97f03eca433dad6986a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hebe10bf0fbac6c48ac7028b840ea6567e21f0197fefeb34dadd2f9577a6e18f99dad0c0c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h789d8f4b3babc98574c74e251845506ce164b9c35a72a1515c04ff544483932f2c5368ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38c199bdd27f15a172fc405a93831dced7fa46962a4e4ba660b0a1c62aaf4de90b02b880;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f62593349215be87f9cec30d4fb6ea808938d1d1c436a4e1ce34ec109aac56d28050af5b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14d34987523dbf1194251e308e86bcc7f5f8bd32f09e4a6a923c942905579faffd66af643;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he1d4369cef72746c80e203552c4dc29964081bb0ef54b2c8597a68effa173022cfe0f03a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b8d6edd5b0a99fe585fbffddcbb0f85b94b7ec088f5f8bc4cf14b42813f165a508232109;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8198a09d1939139919d9a4425e37a30579af0f05c028a1511e204243a1a42efb111a8e9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15c0bfe053bbfe261539f6f2129c8cc44be3809dee15091b64e29df39f654c259a6b53f98;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3d6d876b05dd82d63cb65d74f71a61f5359f716795181532ca8c5b5c22a8183d02f71605;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e9e1ff3c335563bb7109c530ba2ee72054d36cd24d496f751bb8aab56204ecb7dc65612;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9eb27ba473007744997a1b39bbbcddd4a945f6bc6f9f6c95a6075e7b5ac6a9ff0db584f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f4e349aedbb19971967d5709e294b1c2a83b39f4892660307856c5a53a27f9460bd787b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1092c793eaf7692f69e9628a65c8bd864beda7feb1c4087a4fdfaa5fb9414cb84b2a4c674;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14603d1e04d7e76092ed3e504dccb4045d259846a9d3939c1cd406010a2ac49e1c6790359;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h123824bddff9ec7bdbdea8bd31069c996291a89b2847a74832bb6ed7fe9e4d4ac869fc74c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haff7d602278f370b58c0dcf124238e6327c2797848c8715d4ff65708d895239827aa2f9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b42ac000fca31bd6fffebe1b90a9195e0d814330407a65bf36bc312774ea32b60fe7d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h495c70f61c8dfe70e048d369a27d271e5e7927f6c893859cc020fa220722086d74f5167b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14d9283c5019a653a4d94516242286e0b2eea1fbca65b2439edace650d5cbdfcca9aee403;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc89146a0ea632ba49041e03dc3cf3878aa3e94527ce3d102e6241826225cc3275abec58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f2c22335d6e6e061d0220023e21ed09c0e0a00b003715fe529ffc07dd52bfacdb5389e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a388ca5c129704df1d45adc2daff1fb9a3d3ebe66ac47d1b171f993b726632727496bde;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe912087c126062b3e05294be3d623ad89e9aea250436b46263496ffbe6661a20a2ff318;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h945d5636ee5f72cdf10c7f4e52341b6ead0e4bb47cc57e101554a7f24aaa997024d1fc35;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2315ab4a0cee132bac0b62ad6bc3d0d284d53955add2b461555bb42c36b80044c48aadb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18eda2de73a6b3576bbcb93271aa4149837daceaf35e41dc4d3d47e404e3358c91678f8a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de45f1b82dc13067258299e6adf5c667a0c59fdcaa7e4eeebc1c8a2ab8e140f749c6c558;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f281198671b83bde49ca1ba393a16862c4630aa301b3842601d4fabb51313e0f6401822;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17135a86be3fae1ae1c5106001843c36b6e1102ebad326bb460e6b2ae9126aeb8e0a22781;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ccc402f17eb6f40656aa3410c79d2c66c518970cc96effd778981de7a5dfa27e0e6c250;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1123ba1de08b0c185dd0b4b63a22c5b70e9f275e626a8d45b15028577e6a5464d094230a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc2c55faed25f3abdddbf5ee8f5b7eca69cbd77fd6a5894ee1f4d69365e850e6a5cfd3b01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e25d22c984dc31b5c83b6997ff38be8e6b08dacc9f9fb0c47b812c8e0cb9c2d3d604bd63;
        #1
        $finish();
    end
endmodule
