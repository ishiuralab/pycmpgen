module testbench();
    reg [8:0] src0;
    reg [8:0] src1;
    reg [8:0] src2;
    reg [8:0] src3;
    reg [8:0] src4;
    reg [8:0] src5;
    reg [8:0] src6;
    reg [8:0] src7;
    reg [8:0] src8;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [12:0] srcsum;
    wire [12:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffffffffffffffffffff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb90660605dcdb40d962a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19860f2faad5e891f36a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he6c02d782911e5c1736e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f795690c959b64673aeb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h172e6e03fce8f3f2a1a67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf90f6489534188e0c04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9bd4d0816542df9e31e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c4f379a60664645141d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ee2112ab2bf4f0a1021;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h78bfb779f96f61869ceb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1856e4702067ad47f4be3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ad2e6c6e0b54914be121;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e053060f2d82e65e5f51;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdee3aa3580557bdf06d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5cc328af87af443dee13;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1458febce5ab954dcad72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c83f31b3c8d19aee77d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dfd5a50e647e2b0afcdd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123b14a71e5ce88ce40c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1664f1790816081bfd6fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15405fa6e4f650267694b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb4154ad232ce8d10a656;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a6f7bf6c1df9a6ac039;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cd70d779386a4b74e87f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16dbc61a47093abdbc0af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbb5037ad1fbbb600cff2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he496752e7e58f8e5aae4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2bff97c286b6b22dc3af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc24b5c204bb71fc50912;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h627feec5a9647af10208;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f698c088799850207aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d5f0991f30858848b12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he313d1b22cb9fa18319;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h49293dd93a76dfe19be2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f9cdd6bd22be131d5c9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9ba153345ac6da0dd3e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc0c09298d32ab3c6396a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h138ce0eb8bb67838bd0a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1deb19bca12e9e891f1e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc7a89e1f4d8062f0e2ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11492b959d1fc70028e04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h159bccdac69163332f34c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h169b96ee6c285e508472d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d3b8866c73098224e37;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e891c417051c158e4288;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14a3e18c07b3d876d66a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ebc0fd3acc35b45a7987;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e344ad56317183920225;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h939f3c08fe417f57e5be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5c39623384936ae8b7f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc6725d172111264cd344;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123eb325e1e90d951d721;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114163672995170fa14e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114dac7e56de6af35fb8e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7110f58a0f1e16a0217;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb993f9c963fcab9af60f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bdc41a54922d429d442b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h117d75ed6315d96f94243;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1055fe93a9085d84f5167;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed5c59c84c3923406db7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1509d595faa4f221fd4da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8caa437b50701bcd62cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a8469911f2b908621afe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h176f21afaee227335da0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16bb86aa28fcb1b322df4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4b2a4f2d338a744a8dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12bcfeaf2ecbcdce69de7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10ced2ec86697fdf2361a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h82b3162fe18e7b94199e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12943fe92bdd2a0d784c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h127fcb213913d812ffb68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1508774c6a1f8c80d6911;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a127bf42fc4e431afb90;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5c41395a7f95bdfdfe81;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10afcf0ecd29e0d651aae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1743dfb8821987e8ac52e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16bb05fdc2b03616ee285;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1817546fe9b068b2e990b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h190022859d4c8fe6e7b80;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fde5a3742ede56b85c30;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h586c1fe4357659d5ee45;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfeca122af653895fb95;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fad7900d2f789f4d32cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57411a292cc4cf45bf76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h127cb50053f173e4377e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7dd9f9bd9d1ceb3a1993;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h181d4b83343c506ff8fc3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ded0b4a78628d4b95dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h112ca05f483da8e5b1c73;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h88a251b41346029998a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7969a313276ebc188768;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd3653cfb9ec4c9f0220;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h155e2491539be19d236d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83e02aacc27b3b9fbd40;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1516296ad6556885f924d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a491f3e8843df783b04e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h175821df791a14bc47c2c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h307082ce75911bbaa9a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5027e508b01ab773ae3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd94075f8cf0d53573f17;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d43aa8ff8ba819e9b4d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h146513e8af14fb8af4a26;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6ea9bf6c286085dc47e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b60419597651b45f28a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa31b0d5c1a73d3fa19c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h87f2daffa499841bee56;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18e6d4f6597bb50d7b25e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa135ac5a9443509c300;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8840d5ce6bf696442a89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ad0b083f1b7fd1459bc1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9cbff203275ba6487587;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12754afe7a9cb1311f75c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6e457bc17abe7b645ee0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4e9bbe814f92e1314fc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h179c75b86c1df60cb773f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h573e879e59f24c0c1a1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf46fbfb43cb31a11f953;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h177402e5e4dc8d679b151;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1adf71a37b3130c7f281d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c925ee49857c05f5a0a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1edd8fbc05d7c72e163a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17e59af2bd79b290b08ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57dee923a0541b3ae744;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2a771ba8f1ea3e476c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he6db3824adac11bc4862;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c6425f89db0140cc9be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he2f114e3f9535c57b51;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4bd755459091238b61be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13c70a5801241150a9b28;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19ad65d5eed7b4a8aa133;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h33958bc9059c07629059;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h169414cb274cb10be123e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c739f72da18bc8fe661;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef80808451d7322bd2b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2b61710df28f03e1560e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea56ce5c9e57ac978ea9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha95522c8d9c1ee84acdd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f1aab4c7a3f66d52c03;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16e7131393fd9c90262b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7463eb37d8f30e27b7f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a0c9c4b85a0a87daad79;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h65942ec8943c96fcb2f7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124f930e4148981be5c68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h55b10329a6c87806cdf9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h459af1c1603d25400ade;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104196c3ef2081fb0aa7c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5f7f2fe0fdfdadffafc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d950963c18cd655d7f72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15a0d213697958dc812df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd1b52278717de1ac3cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ebe96501f46efe13005c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3539b80cd8c1f3b87dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d939767b21969b405e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b2acad7051e375c16f0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fc0a97904bd8a642a14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13864ae97a734da9d6ea3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a98f28a990e30b7217e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha34c6f6dd0dfc665b9f0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1441d0b9606caf510c06c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1beea67da01bc03026683;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13f7da9020c08399869ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1595930e74cf62df1383e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f581a70b9064c8454e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h90934b0903116a5eab41;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e777aa386f8ffa99765d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfa8af2eee1a818404b85;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16085edf415efd273a161;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h303bdcd54d8cb33b84d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1efbd43ed8b76d172e822;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9453d30b919a0fec3495;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h120defcd85a207cb2601e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e236b25a4dd3bb8b9a3a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc78a5012396f865a80b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e66c4008bd9ca595fe5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf55fcbd05df2177148a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h116adf2577734006fa2e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h37c1dbeccc711fa40861;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2b370b7e1b3ee948766f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h595e7e4ea3732188862a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7632f54f820e179bf3e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11d09546b806252881084;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f81efb2fb3d303cb73f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f3b9f7db52430d7f4b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3f5a204684949619085a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cc57608396ce13559c89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b7d07b2ffd5ffd5fe6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196a14bfa1daeb804e21b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5535b1389d0b358ea55;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6cb7a3ea6ae006fa1d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1951613be786fa0ae76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h107134bb2357a9b268abb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eba4140806788a72d3c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd415c3785a19f50a4bcd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1217d1604d7d1c65731;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf1f6c2dd389708931b3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heb8c2cfedbc9784399de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc314f480a472355dc1f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2c4dd04d734bf93132a9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4e731d671a079ac2db0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc7af04078c1af1c46863;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfff69b100eae2816a717;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd86df5c5d41a17e14f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60dbcd5593dcd8e3c31c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h55902e1f6e9b1e3bdffa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1194a0a186090739b25af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6fb66d255ee88e1df711;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e7290fcb09ac270e1cfa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ab35d225de0ce594b60c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h23e19e8a27f72276bd0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h109190e3c466b75508f9d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f7135b1a957fae27efef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec1cc1315f1fa450004;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9b90cc4f42a450d3727;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h364d9ef1c466669c4023;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd16b8f1512b7c2fafd0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18a81303318f5472a1b50;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb831c65339d8e91832f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf0bed06e242cccba3b85;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f1dd7f407f07d58966d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h199cf636df3c1ce8d36b3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16aed1191486b6226c5aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123b5fd3f7da72f113e8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h222221e9e616c08d3b93;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h129f4591a773531e54258;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h170e878dd960fe870b7f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf596061d198ad090af4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10b05ba6cafa6188ceb22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13ba2e69ab770540ace78;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11a6013f49ce68991d22b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57ebe6ba65862bff8de6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11adf5c14e6f0a72b25c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7f6590ef81defa9c4fbc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbcfbfad0ab996a948fb9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbca812bd436202cc6ef1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h329df991ac4b3cd24da0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16672a8870c13dd04efe5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d6188b5c158a60c69fc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d377d501111e6a8a529;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ab1a138ab62571822caf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bdfe1425476058ad363e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1961e114c5dd2722d5f72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h50aa296b6304e496d68b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f0dec26ece9b80a3201e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h146f38967917719b71b44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c7b33cddc4620f79102;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11633b9dfe01d08a6ebcb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c6878fe8d7df345db9e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h332ba2b17620466c4716;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2209b090f653954a5667;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18398fa01be5200441b39;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14617e135d75dd7ceaeb9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9564561b71843158033e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18fc9085429fe50eca795;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d63104d92b7fa746888;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h127abc37d2a8afb52975a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd8cf1bf2e96f479caf0d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he816786b22a983e7d58d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e00b2ef030cb8d67d1d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h113354933ca9d693afe31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd86bdd330359d0e5cadc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h173973bb07400a8b08c0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3175363156e5e2fd8b9c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d55f8301fe0628d52f0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf86cb3824fc80e4b03f6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd1dbbf1d9cf6e29bdba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h127029c17b3c158181577;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h181ced97c380017fa9163;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3953632327892ffa0079;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha6bc3336771100cd43e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c5f9e80724f7b9eb5e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h127b379530a6cba253722;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fdc2505709f8ef0f6fcc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h72d7ca843b9ee29d95;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h126c66afcef6b24249e7a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h197b7e61b85381384e6c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1badbfed0da435cc7918;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b6f51fe5ff5aee033db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4e88b45f63d355042335;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15a4f2651b8ccdd502166;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb64d150274d5f92c0ce6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17504d8aef83b75464f5e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1617622d285d2b08d1213;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f630b078c4ab9c1e1b17;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb71f0e7393208b6cb716;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfa9152a07454fae2926e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16fe9c2fdf4bfb4222556;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44867d04bc161a04605e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d244e0c2ada1539d275;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c34eb846b128e55a5148;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bcaa4f1acfc65207ebbe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e6b40a96d0116e89fb5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ea40251d124bb9021a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11801517921794ba8aa1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b86e9038b4d205228dd8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h141e07e970bc87530e7ca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h72a6697f5b093582b23f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19639fb0dfb7bcb2f91ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha0f0ff233d8d0c1d0dbb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18f165a02e1abcba7c97e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2b7fb33c1c74f3ea5e7b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f645c133a49c50ed7a0a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150ea1c7917316ae1b71d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115a74d9786975348ecc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6714fb70092651bd0a16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9496793958203184921b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103a0c5a7f42c0c7a139e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc59cf59b5ea5b3a438c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h484650fdf0d41e434ce5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ddf44e05218ccb57ec52;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb34ffaf3986e497831ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d04aa3d0d82602d69db9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b7496f41acf026ba2ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h144db42b454e80c1ce9b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb7a582bf0012535f2f9c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1347a389331438c5da1db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d7c5a8cffa8090e2b25;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6bc2f362da22a39e4d7d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e0d0a40c200fff562091;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38e3b63bdc2259ab578b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38087a460b880b2d8e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha5f0a4d1a6511f1656be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha77403db7558fddf2002;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b2711a1b74eaf748577;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h938957db5bce2a02eb23;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6cd1582184ccfb17df1e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2755f1b44e211e3e38;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68ac298c625b69495b12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5114373f58acc78c1d59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17761e1fd42c9a271d880;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h555e7642e0cb8bcf14ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aec671c3155d5e499acf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12bfc8fa530a540a08419;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be4b34a84ad95dba51ac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h199af511572dd4f3f67b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a8740c5a63fe8181c4d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h72195937c29d55eca743;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d91107b3e4bc1903c36;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbb55df19a5c863e4fafe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cae25a48ccdc372119e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc516cb10e08bda56825d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h257806c2e92c37ae04cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc58de5888785b1c1df5d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c48f97b7cf38df98f36;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7e55a030cbec3e3bc44e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h127927363422b560d77a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be5dac0141605776cc0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8319a40c335f6115adc9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16a7b45d44e27b0d05822;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bc38d4d027574b626137;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14fddf2e8bf82ebe88bdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hacb9b1585974b78ae55f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc24a3c7eada97b054d99;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dbb2ced0dc8d1322fc7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h64cc5df91a5dce1d577b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc3ee3a3e7abe00240fc4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11db0e99f97e25e7eb3f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1deb7cc328ff9067a627e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfb65ccf0936247228a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e4c18d249c9a8522593b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb55a24c51c45f8ff5877;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb71462c434953af243cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e55a5042ef1fae195233;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af0886c752ae02301773;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94be88306ca365ecff75;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1711d7ae38b380133d7ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcbdf747c763696279e1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h61d6a99baaeaebc23760;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e8e0b695d8915a8352e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dfa2034c71f401cbed6e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1638fd0946b6c1403354a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7731dfa9744664ae036;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb88b2d69df0ad6385b23;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cd22cabe4d861ada2789;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c6beb3f64e71947d521;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c610b4cc595b99f3abf5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf0d942624614b952a5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h865183ea2b526c0cb63e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60391fe97613e96d0234;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1973820f4b712721cfb83;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc6537ad9448981b0cd4b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c45ef328f530869e51;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16bce036374946b82bec7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af33f7184ef2d7802abf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fe29044b52503f62b6e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14434435b1ae30d781e86;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ba79cb7ae9b82384758;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15073d1feda92d57e56cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c106747720a72104635b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196d408fd25eca167d0dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1937ca474bfddbe5222c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h666c4cd2aa532734471e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfafa73c4ba243209b481;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ab5f0a1ce8b0ee0dd59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a04d4a68cbeb282f26e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b02d86993e2e4e72aefb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114ca2fc3c6d98cf3d88a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc0d5b7a6bdb29b0c923;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea50310b8eac4631501d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hca08da1f2c2589907c8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22d8d7bcdeb0ee8c8e3e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h194851f4fd4ec495baf05;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140bd8cf92e30609f8974;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1538cba36bce0cf6bc53f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18442171bf9603b4852bf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hee6265acca9686be4415;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d3f5a20f590d78437478;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13dd9e3cb5c8828666e98;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114df230743e2b5ddf69a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h152f5880c5039cb2d145c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf03667db84d488c80d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de67283440f0b2756709;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10980f496fb57fd041fb8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hee5682309b5c9259ce8b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h826e3f66c2c6a46eb7c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8470b5847a703cb7b266;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ec4bb7ebc76ff061df0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1363c9583ea1806125a27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he84b0cc5b07f834b9c9e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e84296be7c47c8aad85c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f532806e5a67fbdf801;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8990da41d3fa32b30b22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a421e000f0419284c23f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4fb7f6accbffd7383871;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1df81121507e455c38296;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd2a9d70cb2e94924957;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf28ce1f9d4e98798d2c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h129fe638877578cd9f537;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16624c39589abd4c69898;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h69b3822d504c71c95748;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h108b45f59413024c9938a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d4e774ad73d7bfbec319;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13ff0bab6524569da3cf5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a79ccbe973cbab556eed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h764565eb797ffb06ce07;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b30ad6f542477deef2a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5423913990096277f2b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14a27295909608bda0ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h126e1868b8c74294e8f66;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf45cafe3f1a4395519e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6aec28a9ef7606474e0d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1246f6d31f86dc34bbdf4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19756b2ffb7513c1c3a96;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec8651c91304e06fef8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15704be403202655df12b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb106250e55e4e16fed1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h76751335e82f4b2aac69;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8b0539bb0f8eb8a0b3ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13db4b89d4b8d2e3e094f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2715d0f77bc7304d3a63;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f5fe3d436c4c3d8f75cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11a14121cecd846fe08e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h69bacad784ca044f1ad5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he8e0edec86d63bc4d2ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ec85f4156e402a3c8cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a205f3dc10036d755af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18aae039f1534fc3a441c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1084e8b38c361156fef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3699a6f2c697b1187583;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8956f663a21cf303ef12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbaa09ab06dd6a5a65fde;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1323eb11fcf07b3282816;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b003c9695dd9d0f8d381;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6401c50417210d2c7354;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c689b8141664396e99e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9b5257854db80796df5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h139ff213bc9d115a65b3b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5cf3e23e67bb732424b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f714505e57a67643da07;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5614a38b33085eaeed02;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfc4be4beb4be1696a4bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8f022ab3411e42499c80;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54f50ea624c6ba0ae447;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c59c3498bb8bc757558;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hff4e89537443e0eb4d73;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8397f5269f4b54cb9178;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17e8ed62815c4cf0c9ab6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd3101975916b572bf86;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f15ad1f225eebec67fe6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d5f966122e95eb524b76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6ac9b164064df0e769d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h953a0c3d133904d5dec7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h43947800d574c3435b0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6bdc7ebd0293a631f9da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h43b0fae7fde2ec438dca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he000c7ea7434c26d81e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b78727e1bca1d3b8aeb6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1514f87b36daf2c25c1f7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fda1a9d8ba315e1b19d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d38331a30aa08c0c8e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h680d3f6aceacf10cebb2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114c4ffdae38b7232e88e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h100b814e2934d1c0340dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h982c84a6ebf16fabfd8a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57e4ee62ff46ada5c1e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h120dfca7895994c9df379;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda7ad48bcb91477d87b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hceeb23de2cee2b89a978;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a104376d0dc94896fb4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1adc59d317692492395dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92d4ebeb25156ef587dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb632fe4de79319538b7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c82b503efff927380139;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14fde271679bb7a3e93f0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h79e2c77039bfc5f51c9e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12654e8a8e20077543afb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf8a95fd1b9f21dd59b0b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h904104004d853443b5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h230521b797907d8cf2d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc37bf29984fd83b258af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h129da2ba55b2556e6d7e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af53379361e06d4d48dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc45a3aacaf5fe03d889a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f18554fe1c4867e39872;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h23604887af2957f4d534;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b4a429dfa708329c9abd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14912405cd8f13afa09c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h855d752b278a3efaf9d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he10e798bcefcbaefa3f9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1cee1ba4ad5049953cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4fac4da45b7ad2871af4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ef5c5d1c1672333d5d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b5c53614c26a1b0d74e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2b0e1ccea87837a0d05;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h47421529f28b581514b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc49effc51f30605e89f0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he739ea6efe38747dfee0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h26515f1d60ce21a4554;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hff3c3ee8aa8cb1e27565;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d68c4d2d88c1d5f95dfe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b7e94cb2e3f4f45b2ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a8f44d1d0ec660c492c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f476c02ac33e033e912;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92a51cc944735e8ff349;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e0edcf80cceecbd6a96;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1926aa50299c0284f42ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f4148b3a3efbe03041f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc15f7eede69fafee00c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ce3646156483fa91905;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c26ff7b35c3503f4cdb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3a83c5480a78297ab662;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bd98104ccadff5184d6a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16cfaed8145a708548025;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda66b3fe6eb1b2fcd24e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c81b5505924a259026;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hddf62153867c0288cabd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h93cae0328234c6067c1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h73f0659d5ed139a888f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h964ac15eacdc8d308bfc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb804eb0c970d8e94b88;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6254dc1b08faa73d38e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h95a50ed598ecc2352db4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf87026cbbfebf48c6a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha3753eef41b042dfb59a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b6ec7327a76df4f36bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h111b85b5be380326decb4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15215518d7de93d753153;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1f98d2cf066c6f1dca2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d6a0a7353b26011a85d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140716d199e6cc3e4de48;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda311e0b04b1cf7ada46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h122b2e17c9feee150828e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he08ea1b9e20c8dae1517;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1979aaef04cb26f4b30ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4017a3919c9d3e08f8e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83008a66ff912fccac4e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb83eab7ef6624946276e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha1be123b371adf3319c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hff85f9b210785e453c6b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14459d12693b53e15fe38;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8120eeaf7e789bcc87c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1687dde8893e8db8f8c86;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h705f566d79e00618f26;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c5d1443ce75b76a51c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h40c1f21afec91e017cde;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ca1aed48fb047db4a57;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h933dbc652f5fbe69ace9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a19028f96b120fe69b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha116988f991b0f3002f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be720a790fa37149ccdf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e063665770cb47f147a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3513b96e87797376870;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d84f6a7e998555ceacb8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db59ba349f9ec9af234f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6daa6a145fd92def15d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf604b5d1811c4529e2c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fb1018120eb5d686919b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef5af97312d728c31770;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d3283db38349d710f5cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8c0e1aeed551661e4f6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8df3db90b5a9cf8d7009;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19932c80e996e180acb37;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6ccc28c4bf20e24fe32b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h47e11bb9eed3db512da7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ab75d301f3d307b8112;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa3647743284c1869d10;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he3a3f8e7943820e7e7e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150fe67647156bbf14d7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115eb4c1d8e45fcd31764;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1579bc745c266e0c961fd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b389073862d071e3b085;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb4e24dcfeab4cf7edeb3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e7858d790578227dedf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h137bcac877f8480141426;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15a16c0a327417bbbb18;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d6f93d2e8609f79c5f9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf83e6c4c1438b1cfa66a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c0769f3d9bb3d326d630;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb46c8e185aef596839d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1df0e902f1a7727252439;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6595595624cd94b195b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h164bee66b15f145efe6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10033dfadb83617db22d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5bf5746f8a1d51dccb18;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h75edffc7f5f5cc795a3e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11aa816dbd3c1e279a561;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he875d53075f74cb25f0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h120aa1aa06b63f9ac4caf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h108a756bfa6945221678b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13c28658297136b4e8ca5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a80efb474b7678b54c16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2f5751d1e231d99a510;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1359328198565056ff67f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a0d743850214466de1fd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103e5c002acf431031ff8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1866fa4845e964f1abd15;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f6eda2c3f78a4c238dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b3e1264ed0ef554be803;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e21fa960e267ef82f43c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda14810d061977ae2adf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h283e14628d4ee4c7865;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'had63e01cc65ea5d89592;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15265be1f34b67c8ae053;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11d2297e51e27099a3196;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b3547a647d21368d8197;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c7a02f12c2b0f4e28d31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4927ebd3229ec31bf05d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h167d748e6800c6a575634;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1402fa4bf2a37b0594c72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e0506e4fbb00cd85c6f0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f1361d5989fbe1ad77c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf8ccc1a51cc2d0b091ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h59917c92d8a466b6c437;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea9ee1f6523dc2c51ea7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1673eae3bc3e58de365b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb7dc36a3aa3bbd287319;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1799dd0fbe845735771;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc6278764c7265eae6b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf8c687b43aab16fec8d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d32c0c727614adfd2b94;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ff4e42a07032a3bd069c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f67ce2bbd396385f842;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b06037bdc59720371d73;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2818ffdb82f6fca7cbe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c74d1998329da18eb3a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17bce847faa6d87f25a13;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8889964e35a3700884d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h141635e4b69e2d6956728;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1186ccb8d874fd6ffdcb3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d1a4e18e887ca909343;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda814e5ef53ce4c1f89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h191a285d693b881db9bb7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7b08e476902aff64a9de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h72a9980f464340f542da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8ccd466d7ec32a2c7c97;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1faf1ba8f37765bf9e888;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b145b075c069e0c4d6e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f3aa11c6e1179b7eb937;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42b2f0fe03864ff5ce85;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he7e47843e5b68c3a2cd7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c451fa0761f868d244d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h335588787f82cb3c8a0d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h73298ac7883785a7e625;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12d6df0b0d91ee33b98ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eddc5a88f6e6fbc68367;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e8025d357e98a0be4d5d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9478e27df162c6b5d0da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1544728d3d229a88f6c6e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae36d4964fd1dd5b70a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf3d2db3573d1e968a54;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcc4e350560691e3c51e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'habc46f83ecb6c62ff9f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd0ce7b8e47a34b438bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d20c2dcc57619f1f5c16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13052b5dda458af5abd15;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h378097f3f7d354025000;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be7a8895ea791ababcaa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d8db698e1b4ebd0b4c3d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hedb707ea56198b50f726;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7f8938dfd988ad341888;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1edc0cde3957e484ff36;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11a5004f44ac5ad2d2dec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19a347480aa392ed0e4ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfa00c75f5f66375a8a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h169aff478364a7c39ba58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde2c54c35d1f0b37ef81;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c45ffd1fc878adae9a11;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1824aed5c09cb30f56a67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19a8b199ea5323e80161;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'habaedb0b085774266c6b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ad715d69b206082125f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h84dcd588f5c31824502b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc2cfa9b1f3ead9f9d2ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ccc249dfd5666a6e83eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h125ffd185a20fefceffec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11354d4a44331f641dce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heeeba1ae3239ed963b6e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ce4adde0fcab3e593934;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8ec6e183bb545067ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1df9992cce1db7d9ef168;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3143bee4959484f8b840;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h122bcd5ee45a112d976c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e4e9a854c073922ddbac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18e1416f2fe321ab40d8b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1726c9fdbc12edabf60c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2b916cb64b2e47975f9d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h86fdf76a54870bc66351;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd6dc5488dc98ac3cdc96;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22542fb21bb224b4d97;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f9a207044e1e6bab4cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h819bb303c07e4e44e81;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10010b9d9053c61f9f778;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8fdfdb56853b65699cad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h58070dd3af22de3433c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ab2100330d11b6e5aab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f144d7b7ee0d9108d10;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f6b136336636f63f72ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he5063ce66fe4c9c2a4e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4fc7eaa561593a41fb9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b66ec3c33ca4bab2f5ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d39e939ff679b18dba31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h168cb81cc80ad7924db16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h93f0029f79cd0787c760;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1721ad687d4ffd6c6348;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd6c9b917c01ce5d926c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b84f53af1c371535dcc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb06c980213825d180aeb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hafce578a5dc04f9783b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10fedfb9dd181ca4d0444;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f3ddf3250fcf2bb5ab8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6afd91f22a717dabfbca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h126628a7220b825ba5acd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c4f3807e0362b8ae2cf0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h48b7ac5490fa814214b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be75ef6144b47e75b477;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4fb5d39a83a0b83bd1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1799cb7fdc900d6da7685;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d35e70a513ed3ca11aa0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbed9f41aae746a925f9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7696e9a020d622ade8e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcc389403895ebedf9969;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5ba1ca989429921198ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d83600a0128810419e0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h64616f514217a1047553;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed87c19b682b7d1eb2b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha78da7942f1ec9e42190;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d935f56c7d66ed7a6c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h613bcb4c979665eeed92;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h191a7920635a981acf66a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h156c3e81b7428fc3d1f2c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf1d0f52c05c49503311;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb27827559c48a97c3189;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3b9bcf6684405399ce2b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdde1d9485ed0d2363c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcfed34d7907915b78b97;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h24189c39b01e2cfd0834;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h151ffe783b8ce0dadeca8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h313bc6966cac83471db9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c15f4f7ad1dee13685f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7419d29cffe6cee27eb6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7cd49fce9457da2bf7be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6759c024b7e10e4f8e04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7231e44143f247d0c906;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11565b9bacc9c56bd1ffb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hddc6c877c543ac15f98;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94c8f6b407e17befc58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d892d66c222763fd69a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2adca50af551b6443a0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148780f3955f2a30b0945;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h45f4ecc70856a07e2c11;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f162c8c9daa7126ce495;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103dafa459acde3c4dda6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e21329d6a09497b3e5e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h742e4a5d9f09cbe6d24c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17311d81777584d157975;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15bc06dd1c872884a1ccb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf69320b67e13cacfd4a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1452e53d802ddfa72be12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b4c6dac6dcfe1fa4097;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h49724ddd6dec9721851b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b4800789a83849e117db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb91cff6c545f5a17ef4f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31ecd6cd7ce5a066ed2e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60f7a878d0334077f085;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d32ab7f468239148352;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39266c43d2fc5e358c18;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8c8186ce4a778bfbfb4c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h177136ad3c2864a91fafd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h518ca7f96c43b2981cd6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bd3094871da2b4fa150d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cfff44c7ea3d8d5fca69;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc493210adbc2f67f1235;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12937dd547bd945139efc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1adec92a1a28bca11408a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h26f17a43f7636a641874;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16423012a23041ead1763;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15aa8f6b7d6286de4d36f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18e5a9ec511d9a212d81f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf51bc46b7a5d509c9ac5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15590f677411f572eb353;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9fcb01560cb09d7da7f9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf26a0fbddcce2823bb9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a5ec95494bf04179deb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb2e113bbfe95d5b05d08;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124f21aef4b026d0c4fdc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hca36359a70f2902bf26d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17e69869459148bf098b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h588a24f1430414c36ec0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15b3023c63c48486450ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15fcd0ce6fb9dabc715c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7c3f0ce9a477615a8f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha6b046db7e87170469d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ee3fc90064bc8686fe1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83cc4ab8db875557eef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf0f327a08c0ffafaf4e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1293bbd08299e0f1960bf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h46ab9ae38f0563e5fb37;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf2404a624dcbfd5f87c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfded5af46afc207ac34f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13e91c976b36a98cbf1bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f7b21ca6ed75a127d94f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17dc725edc09f6bb213ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfe5f5b19c8527aa6a50;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h95649678c42194d5086a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h189c77e246696129e5b69;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16121e9af3b3ddb37071b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hca303f4c64928ecf2862;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h95852c99d31ae4f2b268;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16f0a10878b67fc6024c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1add4f845378caaa63476;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca0bf16e5cd28922cf8c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c4ec0217a3c407250fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54154818f12621140576;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h74d72e0445c52be16b63;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103460459d6b1b3575d64;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f179272e43f6f616b7e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4fc0cb8eb13d81bb7ea0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h773c97bb2e0f61caf4ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c7827c30798896be2cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2000b059b6c41893266c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4580c3b813fe663e42f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he6ba051ad4182678718;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf2db36685fff940bfe5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6d4e0e7e854769f78f7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14367977b531ac93a5542;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10545bfb4146e60f3a71f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb4cdc3d6d51cc1392a61;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8063b130c54bdeb529fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc944cc161174a5629592;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e7acf3abbc3a9dd9750b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2a471aced29d572a28e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h657d0cda5425c868cc37;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14361cf25c7d8457dc7ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13c4b01efdb396b612ef8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda78ceaefaf2041e8255;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1298d3c77d4fa29e99846;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he74db1cba5473f7539f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ab72245ada542231ef9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac5fdd1e01bf7d397448;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcc40b4c291884aecc9dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h911e55b79b942188d2c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h193a11bf32f1db09bc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha0bf0edc8b51741a4366;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h176cffdb2e3011526e9e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e878ce210db8a7cbcdd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b4b9c9100ab0563500c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h99de34ec0c5aab62289b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haf73c4ed91a244c5d73f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7e977d789df4229f1110;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22c8f16666c06dfa898b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19918135f3d82807c94a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf18f0db5d875ed3086c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e9dfc274b0bb5b65fbd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h25209f74fbfa0fd02e34;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d60ed9696fec593d2b31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd44255135bc837315005;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h63f251d27cbad3f32157;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a84247e034c64c2e88e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17399cff61438471b7aa5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f16b3c639b2ba1663719;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1533fb015a75108a10373;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h162a5522a91cbf1b3eec8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15cb026d41c5d2c93147c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13a8bd2aef80ad82c2354;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hafed4028cf9b0079557;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ba7d917e25751bba8bb8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1adcebf1c0a40c9d1efca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18fa6aa639fda2e1427b7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h108e0193e757c5462459a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h163ed1e470ce68d0048dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h149cc9209efcb71d472c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h102bacbb624afc726d318;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he37e49270ece46233157;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ebc74f42e1bf9ae6baf3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc59fb1ccd690048b00a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h133df9ef9cc8399391535;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h95b83cc10cac3d75cf2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89088382d0c5b22dba8b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h647096900504e23d5a10;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1da2a3bcd42133b87485c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha14ab46a6b5b84e682c9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aeb9cf6b6689c15b06f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8803ac447490662918c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc8f7cbb562dfa919ec4a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2f3782ef5c701976101;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10dd74862fdbec9e4c913;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38154a398680f04c439e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h732b515555b7919a271e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d25597cc820f9c3afd3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b965c3d48059042a5045;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h71014e746dfc70491fd4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5fa34b94fb1fe8ade3d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc6d74723afb56e90d2ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18fab05b8cffd377ec78e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e5a029a4efa214af4d3f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d84e15632f7d8bf3777;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd338d688c591249d5433;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15cb57d2423bd702be36c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13291b60d2e018f1b3da4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h90affe73405732aa0dea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44c6a3b6aa0eb05091f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ac598db5ee811b7fda7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1458416982afa44d29e08;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5240de2b533741c71104;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h116c45fa17fe0c04a299a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h33872737861f101b9861;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e84caf5118f10b5f7533;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h669c48d9710de40f2800;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a474c7347ee27b2c7c13;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haba78746be31bdc5d1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfe7bf2ab2d1c097c7c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f6740d514b913ab0b28d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1abab2bdf1afaa8ee7dc4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fdbd16ff319375c020c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf18711d8708124d1cfb6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dfcbc6062681ffe2d811;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e7235db77ebaf4de5da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38fdade463a0c3cba429;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfffdd7e340ad9d313aea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hce29dea461e0649bbfee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e57607bf712d51894f44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h155ed898f5467b8b56a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ff0b83291c4dff4df60;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1329920d42148d4f111c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54251be50d2af404b4f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d488034ca77d5b2023c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7afd6aa5171978478530;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea4f52b72fa9249e508c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60d1079e4264217155b3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105711ff4a15fbfd6f92e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf32328394b396c33059;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h76b92a6fec1e5e85206d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h74551b25cf92bcc37d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b36192ee1fac097b3cf8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd97db6f0461cd728097;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a654a105b66393492b71;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2fcaf02bc128197367b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44b8dd5819fe0ab3a943;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h157c388cd270c2d9f8d27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e562ef7708cdd0bf3385;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb98aa0ae9ecbc1bc3895;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e71169fbc9fcfa80341;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb78869f7b2776074c12a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8f27fe296fb0bffc1fc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c6008ccd307319b7c912;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e6891ca5fe53d285c6f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ed1777090aeaa670b4ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h87f3fe7a3ced597c6f60;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb529b451add8fe4fbf8c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h93cb2c36fa2cf85fb52b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h71f16ed638ce5219748;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h132881abf0de9ae86d7db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4dfe3b9e588c9f511762;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd0314022c64d535438cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6ce7fd7f8041038724e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15fb8366c3ac58ad5effc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16162bef2d3948db57e3f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d23d26b372481c3bf87e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heb93420129d01802235b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h29538278994d3be59725;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h146c12fcbe9f47f14f2b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eef4ed409a398b5db55d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb18206da67f222bf1bf2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d93e01356562e647554c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ca92fec1342116bd79e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h111693aeae5ba531be8ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16fae3cae362190cbfcd6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8358d0666425131ef92;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf5f13d1785406d64767;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18f0619201da8f39dee3e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13927167e2dd33501467d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e192e7d823526ce8c651;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a276a2398701f70549c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f35114d4933024ff894a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16892687c70cd660b5879;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb01496e8ccebff0323ca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5ca2c741e95346480520;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42c887bab2631dc837fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fcf727138aeb98bf469f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h800358edc590bd1eeac0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2fda44d2a7e142c7d22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h915f9501b2f56ddf73fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h369e5cae707514bb9bf9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d742afa13d3d028e25e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16eed3d03735ca7204b67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17b0668992e410d11118b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cc50078558954cf4b4d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h245c38b597757a762caa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7796a6a89425a270dd8b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h112af44690c1055d749d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h53b26f3ac66b3410f7f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19bc7f49415e65cdae6eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcad0bb85fc018ee59ee3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d7895c8e1c04acc7a2d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fbcdd4c3c431f72dcb89;
        #1
        $finish();
    end
endmodule
