module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [30:0] src30;
    reg [29:0] src31;
    reg [28:0] src32;
    reg [27:0] src33;
    reg [26:0] src34;
    reg [25:0] src35;
    reg [24:0] src36;
    reg [23:0] src37;
    reg [22:0] src38;
    reg [21:0] src39;
    reg [20:0] src40;
    reg [19:0] src41;
    reg [18:0] src42;
    reg [17:0] src43;
    reg [16:0] src44;
    reg [15:0] src45;
    reg [14:0] src46;
    reg [13:0] src47;
    reg [12:0] src48;
    reg [11:0] src49;
    reg [10:0] src50;
    reg [9:0] src51;
    reg [8:0] src52;
    reg [7:0] src53;
    reg [6:0] src54;
    reg [5:0] src55;
    reg [4:0] src56;
    reg [3:0] src57;
    reg [2:0] src58;
    reg [1:0] src59;
    reg [0:0] src60;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [61:0] srcsum;
    wire [61:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3])<<57) + ((src58[0] + src58[1] + src58[2])<<58) + ((src59[0] + src59[1])<<59) + ((src60[0])<<60);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h311a245f78c7b71c28dd8294d7318a603f3f6bd6a8278bf0b06523c12e960eddc70db024222e729db25c52cad648ceb1eb426a54c5966fe49613b0a6609461e2e9ef6e42d997e8604df433ada5dfe074d4ebb28d25bc2b4635da6b03418d7eec195826e0df6039b16eb0119bedbb560e01a86c18e7be8769;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h110482d33f6acfb4f0cba5ef2d0f811255f6d4f9466306cd2e93132eb07ca8a9fda27fd3726715c016a4cd0cfc0a152681468e77869bb1bdb3af6fcbef3b738dfcdf2eae6dab69545406966faaf4b4f3244a31ab17b7dd500b3885a3524770280e9a1fc47ff6525e09689683afd6bca0c7c84c89f76da4b97;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1312123cf4c2e7417dce56b3575c0c81e1d76a46b448b7c7b59036c1c01e4857d5ed8a4f3a357ce72d5df43537c971d4d43ad66c4e7c36c0227e2edd8bac4d225bd6ae924dd327da83d199bfabae6e1297dcae720d39839ecc9dcb44171a2bbedf79f6418047db28f577de9e891d82cd5fa91b939fbcb5c16;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ba47e4937b54d09d0a04bb0c51a91e4370ac56ab4d39aaa33e5fedb85380aa312481ab326b72dea710dcd95c83e352e0849c2191bd61563e36feea12503335f00873b547427e0c6dac1d865ce0b16a78a999d03f89e153eda5e13c3324db59e1ce002fff25c0c6729d27616ebab56a900506664b7394276;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b7dff5d6696bcbcd05eea8a0fa218744101ccb0b995c331fb5cf7205d35a601ff1c9e90866a50149433ca1be3839f3e803387cd3b40c90b32ca8c707898b7736b1b4eac4f7e6d8a3bde2040c3a079def89191f2b1768ccddf85d5343326e78fb00f8f726759740fd87af21e7b08c2a70ca157ea5469a8d91;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb8fa6295004e8ca65035ff18fb346fa0ca31344cc4887aa03e06440feecc7c373dc45b31a390ee3ce6083c4d092546859ecee44604d990620af9c8dc5291a1d01edbf7b61801c43de62df7617e101f1a209957ead6a6bef2601246fc4ad8a3cfbd9a4c0ed73918cf6697bdee00b8b695084b05422fb36fc6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ca75c5a4feed19f8b90c68f35b81fb5f65e59ff0fc1527f092d908213aa3cb8bbad5ae0bb1d7084cf2c1b62658810a4e59927a9ab42daa757b3718540e3cf48178ef53a3c7cfe9fa8fb5cf2d6ee1ab6bc0259a9131edf70c61983fcc796864cb5611dd54edbeb0fd3c57a08c9b53a5aba10f114102be99a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7d09b9f07ce8c48892e50f829ea2ab0c8df9e5d07afe9ab918b377657818beb66045068fac7c834dcd7d115d3537aea7321b40c754f271278af1ad85f55ae1f6bf6737ed4731dd426e099c3c706f63de579a6279ee9fe896173bbab99b873dda543fecf648f07b2c96b842a158340f9fea4670219fa14d01;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116495bc48e2f9cc93ebd0427b5f925bd9f97bb7387abbe6ea8590d5446fd4124c76c3f828fae7059d907b1c5af4de32dd42bf69afcaf7fca49e3cf0820e5bd8638a379be4e56bf497a1ace7f2a3dfdbbacc6479c80e647b9a96299c3483a2864eb30900c1ac7df773a8f1b0e54cedd3ab1c7a161f9804c48;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b341bd2c6dec76128a6304daa321640e7a9409790d19ab3c82c735ce4c5753545d68bc261a5245a511e8f313ef5fc3ce5ad7852150c1456b7c7a5f3e87f091173735b34dd444bf6d3f21b3315968a75bd69ae3ea6b005352a587de62d524d257cf89bef986b4eceecbb441bf31efd482bcdaff3d77e634;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c63a08c0a35b60a930f6eea0155daa5717b5d9b11e3f964b63147aa9b78b3995d9d6b5515a871c24b919d23d34243cfff21d1e74b3a0eee51986b92b6858a75400b4b557ddf2a08851fa6d397f465e5a98dcb329269dd3ab8330e1c4584d82f4ee72508d61ec2ec7072968969d2a592fe4e27a8a5409c1aa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113c84df244706f014cb7fa3afb1b82501c6146dfbe1135164b0307d050cce8847080c478e2ac2ec0f4023b98ca3ec378973b6ee6f4687dbd180cfb72c71c7b0b2d1fa47dd8c325dbbf6627025246818a0168de69166867de64680b96d27add21714c0be2bbc0e091fd62b8d4c4dd0d6049c7baf73097761b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11036394877e321f0203126cfe5b5bb81d54072643f23eae8edc9394d40e1c620af15a24becb208dba18a3e8c57cdad2be78e2e783d9a701a7ffc96013752b7c60f361385d65cbe00a2653dd05e6b2edf17f6e6b253f2b026e1e2bdef359c9b15261fa2efd2ed6dae9da0a5ab82846ea20fddb00361a27a7f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e9a410b4da0619b5282baeffe33db24a641c866729738d435eb55c2bd4c67802b23b397d8467ed8023a6fd989747a40eb9e4385283e18b45412b057402202dc4dbb2b3aab050ff604b3ae83c869e8c8bb8374cbc16a4dd0e75034842085475c237b24eb276761be56016cabc8c3f7f4eeb546bd73e1005d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h37e614e43382d37f1a7c8d426d583e2d75bae98d1085666eec714af6e6c27f6567fa93a4bc00f8a34d44362b6336a8ace224a67b1ea8ed1096c593e5071a140885b0b8876cfde402ff987eca883c7b9f236653450eb5e7f03ccff5e0a73003447b2437d2f9633554b5322b0be5618755b42c9620595cff36;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2522799d125cbdce1176205ae904223c1dc513bf0bc0c0633185999ca0da4bf38f2e8a30a69500464310036d00fb3bbbdc7fab0afad20a0f9010cf084ddc5e667a671365eeb5133f0d2e1be2ab2e7e5e821ed7819d1e960f5319e62b8eee52bba448dfe8aa212f780c8b4efe8968dc223e016eec209de823;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h190023eb72bec45694d6c2763ff29f317e898164422db59f275851357ffec4160691c71c1aaaaedad0bcb8a64a9b55d956f9238bfb2b3202c293dee215b3832988c321152fcfdd5e15d8cedd1dd54ec098a848a7a88b09903cff92b8e3102043247a215e5abeb97bf4a912c58f8aa25fd9b85f3b3719fe367;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c17d93bf0162dce7d41493827290d1d2ac5a36f77f9c16e25ae6155c3b5720726c47e51bd228aac0be147f722d7d6a12515484632f49875c826cf01a256dfe8afcccf4f12b5a52e33b6d52c9da93c2b2b5989e8c314b09207e6e9c89e9b023a1ee6076d181948a8720ca150fe66e3e544e4970dd16b86423;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he3bc9fd632daa00c55bb1888fb5d731d5d33f1428a64f0da485a88200a20454d31ed1755369d8032079d7cbd6626b2e6d49b4b87fc54b2d89f2078a0ccc32e0b3e9e4a2ac3ae68b7aa1272f2cd27ad7b9e7dc9d48047faae4dd3f3b16de6553773bffaf89947c5056f81d0ad9b89eb3a4dce45144fccc5e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10e90c4d341075f6b194dface48dab68e6beba8c9c4b81b24bbb3b465a3b8b2262895e60530f9759107f62718e4fde621fb28b3f90b8e1d132e0c7030723d2e47d10e9c3262fac537f6ab67aaa610688d969a44c7322292be57276c05807020c32637c3222e0d6ab835404b09af653514182639b35b03f7b0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eea3db37246fd97aef2302ee4a5e56b39cf1a9cf3916f68529b893e402fa6b2df9fe5dd784bbd367a95ac0de5fb7bcbb57f315ed2e03c5d6a218fc5aee3282249b1c2e57e5c720a370e390977332668f1dc80e2aaee3bb7604c3383511b07dbf51491107e585351d7c0cadc8fca36209da804075477aaba3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h354f333bad546c6e0dd66a689173d7d993cf677e2052681d7900e75b0d47be1576e0d69aafef545bbd3f47f02f2098fddd3926f10b38b8746ce3220738e35d0d30e8c09ee79011ac9fd92052aaec96ed136079b42f460edcd9911f8e6c9ff08b19833490e309efc048c83e20b08800974db9be5203837973;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f5fff18be6ed4db56188c306e263645d18400d68f636e62c80bbc76bfcf358f5d01a38de8fdc2e8532a40567acc6abef7ea3e93619e5128e3a5d43ae818af27447c13369f25ae8c247f1a6182777f2244a9748aefa7e2d4edab58c02ae06a0a1cba34c18a51864f0caae0b386e9be27746a3bf97b5ace1be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ddf0ccb693f95f2de53a6b77334c046231549c972a3b17e97ea310393e0f6855f636cb00e12e0adea4abe111caf53886afe3fe65ba7fd040ae2eb5e7567859de33138c220b00c6dc962352123ce98f52a5ebc6308f45102a33c7d6d4f75e7d6309b59eb9b7def7d5edd5e0fd4b892a9d835c236ffa89c433;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149f03b8487987383bd60d95a3f42453528dc412d8753ba732097947012289b68cd81b5675f9ae7975269706684404c06951cb5a81bb55a51207fe8a268003065f4a577d0a666b281fae68a0f17a5b63158dc84d45309dde85d3de34f86f9f80d27bdd7c7a8e8e3f572bf49fef0791ec671e5c9b932c5cea9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a59b1f94b2d1540dc0e9c39b12095abb35f1ab6f4b6d6e07ff9c957411ea7ef1015f40bc5ead8525488020d3aa9c6978ef4a87c4c7f0b0d660c1bb8c6a1d5bfacb2bfa37d18d1ad6cba309947d245ffca70fe2538ce342a7169b0767a9d480961170e81fade072df463d57d18a5b5e15cad951214c31da95;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146aa486b6fbb333cf0129d7b69f73779f4a8b1fef225b2c82b5fdf0b73387512f60fe6a5a8f3a8691b7ab86621e2ecbae1ee8610c684f4baf4a7bf108cab25755eea14a2cc7625abe7969c7d6d1682e09a46370369cbbd10f7d4c62541c1fab8cedc14aff4e85a7ff261355a479dfedf5201c3943e7f9371;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a05a2dc4f7d3dd4371042a7a62c9a7657f6bfa03c31cac6ab6b1567eefa51098fbed7bc388dddd4104af6730e7af0f954d5a7708c710699c2abf2d3b364e7e42305a54079b273fcb3a7898d1400edd8f17b36ad20a805f09cb1cf1050ea0eaf27e269e4ac8eb0de4b2e75561f8a66c1fe52fbf1e666a912;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h85f93d08fd9be155999493d1c170f774f019b9f30443b23477110c5729c623b8699041076dade315e0e6eb558e3c3a7dc805c224be8c6c3a8ed08a3a338e968eca1427aeec29976f4d96c4917f36ad334dd1689f212b4933fa164cf4894bbb2e85ad4b92b5ed7045b30591fca6a5a34ee82f716a44cb3374;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd55b7f7038c224fb544c917cc5483dd2b532d69c7ae351543b9ebb02a91db8b8fb9f257f9f1b2f362abd40e4e43da109961c1c36ab09305e5f912a245cb7468e963682353d1328953ada00e1070cb47c653fb5e14ac768795014a7e20048425b74a7b53292a2bc0407a5e6cb62fa39c5ed15ad0135b64ae5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h46d0634f5fa0626d7e3b2e7eac7fa2044c3ac505f164e3011a08e41b821e157d670ddafacca0e56962a8e17828ddc87bd5cdc789650cb97be5c02a70c613cff17f1296b77ee637dd21979232541e8f7371b13fea36079cc68c785ad2b9a3356cdd11e56189b5d63d126fc03882c37e4f0e52db777b47f3f6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h424a17e64f26cd8036c155034f44228da553455a7bdb5b28467bde9ab4259143a17a51984cea63507b17ac79fa421aa0f3acb17ec18a2401089ce0bea670b41529881bc6af2967d7198f60b2864e1684b70244ea287a093b7e9e7af7d63ef7ac0c68cd067c504f96906747b08481360fe7dfd4747d50a45a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f66d4adddc65662f2cb3be488e477610eadb9074604f1eaa12e216a689a7e9e032dababa7c5e1c80739908ac708f3c4da3872dfb08499e713180931ed8f6c594ec6a3f1d2a2196ab37e77ca63142b980d2d9cebaea5ea3996a2f5fcc073ca716387afefe689f4ea29b9c233fd3cad23c4948985b4d254cc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b3ee33d4f29481dfb0cbf705785334c674564d37c830bb333f30a05d37b178d5b73c20cb72e7511b138350900545ebfe5b689668278d389e6bdfbb109ff0e230768d1fa14b96d4a4787cf68fa0131b0d720977e2d490d33601a09e9be306433ef495d9382e10c40f40d108dc83fd9870f5577fcb439f739;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he0c1949cf5d267d2d765ee5fc8282d6a7304ec5e30380c7bc2fbe8e28d9583e59959c314254ec7113062b838c7452ce672bb595b4fd72d0482c0d14713c138357ffaf602d28da7005ad553175cf44af4a0e425afe32dc8f543d5279214e615e14e18f448d50f4dc25b17eb232c94810f4cc279f0239c23a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf1c60e768cf377e395b1a44d01f5c8cd7dcac2214adf20a15fcdf2479451a4001f54126a33e275b8f7af83ecbaf6bcaea0550d30e3eb932c2cf38ad2ffb359a564b674d62d4ccf2fb0d67047da7328d9ae68dcd5d8e5dcdd5e143f0463e7ff446244bb1c5c6c5e3ea727802f57cb241b2235a0225ebee3b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc56f41506dcb951a92fe8dd073dcb9e05e42c67c28b73fbbcfaf8504ef993f0016836675e6b1ae29f1c94019f0112a89913f1f0e4e2caf2c6ddf0ec35edf14d3aaa114618e92166e99ba96a4f41c5b3b042f9854736ac55dc80c9de14aa9286cf02288f1e9d82f4e33eefc1e47f8ca8eeda2a2499d2e7b0d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c019a71f6b43b45d00537f9b44fa00eb3e8f9c706ef616b2e608d08034453ac38f45fe385be74975aaee67bb975bb3d738d3a030295cc09c7df508d7cd59969e2ef8c71216500c919213bdd25706cb5e15bcdde132d211fbe35a78fb84e26c6aabe51776a0884390da40df9392c10e51ed482b149151385;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ba4390f1bec6633e7734d4973c588aad85d40332fc96afb7e38b3fcc2046fb03c4203127386597938d274dad4995c2c84247363329a4e47b031971ac028a70efe81ad4563ad6e2e06cb25692450ae73676ec13b39cd1bc69a7eb8bff626cab4de179c3052c532c1b3e7a5a6d732b24c2154e54f2735cf34;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h840a10863c625c5b6abca184daf4fc2fdaec45c652eb6dcdffa0e403582d768fd58644e46f980c2c086930c5bca86345809763c7cbea829d339ded6a068ab8653dff8aeb96e4dd67d97a1378f273d85cf5fa11a136f1f6cf7981f816088e396a6c71dacd5b9b5a5d68f39b90512311a2d0dff4b8ce9823e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17aaf70cf0aca87bac882f0f66dfb0ffbda949250413923b4a30de5f29a4283e65613611a0fc324824782214e385913d8c34e2063d104539ab79cbced2e6fc7532f78ecf5a18ef5f4f494b567cbceab0407ce826a4463d3d2513125c5a91b10764754b51840611769ce33971723c93dae8fe23157347fdb79;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5bb9ebcbb48615c3e66dae497784510f0ccd32cb39d61cbeb5ecb9c3781b68d90223e20c60cd3d2f6fbe4ef14fb1ab934b77aae36c0197d0eecf6c77d2c531740b53fdccc70a611000d958a87cc875d8a312b24b9281a63e9cf729d509b8bc63f59dcccf99bddb92e70e5c33b5b39e55619128796c04edde;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147f8942a341706e9a20935ce82859901c8b3e06243e8ce33a00812e1f7773d243de117821fd2a7e09df18ee8ad5a924bce9b79deaa311a20474e673972347addd193bf8743122b6014b9ec000195990af65aacd881514544bc254f49f486ab966c4a0cba40b1b571c1604fd422ff28388f0287e0d5b8e794;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h492b8640fbad708507b1fcd93153dd3938cdb14fb1130cfb7e1e4a4137395a553dbcce520b92df391ba96a84b5b9496a541a5a71e2658176712e31f40aa2ea8044714ef52cd9a36d498a2569bd241b107c134eda9b33b92be11154451777263fc7376eecf0a2c5319c8cdf47f3d9ad324dcfb0fabd1d051b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3eb39dc5504ebfd839de1ac282f367a9015a3ef709ece48dcad326e2aec47c5064ec00a0529e64481149a2057ca4b5988607cbcef8cced2a70d5938be3e9f63550bf97a22ab5792c48d34963ae31d72cd4e501757622cc7902f7ad27e58294ab91822d9c7f6be9a737626ff888d32ab94b574d601690426;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11c41d1993e0bf468c9135c49d611383a8c27ba8dda5fd8351cac661468300fe2af20d9fca08031d8e3845a99004bc5568a70850747bf4c6dd9712f1008b7eef23495a90186d76c9fc44301f074d2c85455dc64fd3e03995b27292513f53e5d44943214a4f72ede79e50de084f9121f29e44c16fc35d64f3a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'habab949c1959d51af1d00d2154125085ff10c5a1d61f6621d131a9acd3d381633ad8a9318f14a351b013f0210039b0bdca3f01bc7b6114f9e13f369429af2087fce2be77fba01af2e789818aeded00dbee7a0bb12e1575c04b575502a3184853b811f72e476fb277f6adefbba5ec051b73309738941b00d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156a47fa81fb99877025a1e15484e014cc5e6510da86a98c74775340a89cddc7bf4f367258ae3ee4b5613e3a10ac5cd3ee581ac34bb850432e710910c66e4869c7fc31f488045c28d8bb05b9375bb0063d2f666239704e4f62d08b2ffd696f630f91210a204bbd48b7f4294f311fb49d2abb20b887fe88494;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5b65509b4a98cb186974484ac01fbf563c6ff61cf9a865390163af4a9fa4dbf012ef1582901363ee3fee25c440fed9c676227fc0255e7a90c470a2307d5f369673f0feaeedd3f53d55901406b3bc9989bf579f2ea9f6b62cf0fe536a2f978f88781e570880b95a0c0b96f1e04c3624ef7d54071ac213baf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he11c92e5b8e09955dcec80602e4566f88e987983cdb044ef6c0e19f96beca7c0b884d1b07b8c5b7a2833f575d1b9735f918f60d356bf9fdf500ab8298c478e7ea9b24781a8c19c947104a516f1fc08672a3899ff6ab085c9e5d6544b19ff4b3a9df40c14c8f37d737972d5572b737ba8824fadb8816f0d5b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3785052997658d0d196d43cb7d60aa7bb41cc6176d0f82e75e3b84b372582fb42531517f6bf93646c70b5a6cdcecbb4e2935b972b5d73ed209fd86bb38a588685b13b7948651ed016ce6288ee07de461b9f98d0682b0d309dfa8bed7e94b6f217584ae6904c4c9598d998ffc2fbf38093aed19d4a52d60f1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h510828ce3322c272957ecee7ca9e985df5afe458a9d0ee2d56139b0e3e9052e1651445ef7078fcf3335073cb3cd9e54c8882141e660851ecbe2834749a3e052057a0a446cf5196049496248d8796a1def80e9af83b941af63bfdf803227440d627368d78a8c3d0d52cc01b001645a8245344fb162d8459e2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2721e466801c0e15960a9cee7f38c74dac72a9667a2ada16a95e84c4e5e237519c1d480192d84d2b5e86b1c6c40c053edba78c8d35c0730810bc2ef3c5d7c37fabacd675f28bdb85cc10aa7438a9b91cbdd4e6759f532819a89fa9ca3165a373c6f8ae84187c246d64de6249fcd333370c9c1092e2bcc1ee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h191636ff1aa199510a869118eaf467159d982d33e665ed14cc669dc34b3b1fecba3817d3032b854c3dc8ec04d9fffbb6f8fd069e2346b082701c65fca844b0603d4cb4b4e1728b8d092648a73ce65beb94b1db59a72822a476b11bcd13d4d094552a0cf5705722cba3c4c87d2df2f81a1a083d87ed318953e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h127d1d4937414994310bbb7ae9dd849b3440971c35312c6ae2e4d083a0fe8c25869813c5d6c1a4826487b7574ac6e9bb50cec41f8e8d85d287c62ad78bda01a171a41efc5adec33253ab54d6c90b218ca59dbb9ebf0d84b4bb33eb83b3e6c3e6bb3ee0ab54ff381bc133c147cf14fee9f4e0fb4bfd947af0d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h85f16c44b08cb5dc90dd94cb3b4cf8bde34ab4308872a40cc5dabd141755cfcedc1bc89dac425e627ae119f90de0d1139584906a200e7c3b624169bfbee5adbbcc90afa3ae557fd3ce51ff8c1b99a8c2bfe231a194af8eab9289e77b1fc961eecdf3ac6a565e448d81c4565d2a756601a1cc28ee95585108;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd142a43eac0b9d3cd26762883bb18fba8c13b6fdfc3c35715717d554e06bae46f65e3d0c7adf4361b9e61a00370f64eb946785ead4c922c9993d27b9049189dd6bf7225adc0b4e21884c3051d6ac2544319b5443f5c4a1830f3295087a604afcbdccf9c0e8fd80bfbe0cd8bee5e9374d824d10f7e1dad205;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146eb87d50a0a03e3688ea5e382c6531b5ea446045322166064b073a2d1a65f5aaec8586411a2c2c3e81071be333c57ec8c47c51473fc68bf06ec3753bd271f2aed9654567cea9af6cde3791d0053bb6187545b35847f2708f73f3aaa61dec37e0cdae72ac988b03644e50f10b1528b5740e9d75d24c40224;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h242aa83c12ebe954e573ff826844184fa85d8e0ff43a9493bcf350437ce9e0794052705dc7cf69d836dd7cf404f0610f241b34ce443189c98086fcb8bd2a714e2fe7d7f076bc6eb98bd322f15539d0b974bccea74d50fa0d35e765aa478c0992808d84d80e4362d2ecb8e46b2b76c788e59d28cee9fef6cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc686943a9f2033d80029d932c800ada2d95ab8fbb0181fbed2dec139d2ee4d55d0f520e57ae23dc4884cb8f94bb2df2e511f28583fda4e463260df0f87619dfdb745f5ab986f916910ffaa471978847f0f87e061d136d437a83ee93073416d35015908124759ea50d21716b3d8c718c390316e2252fe4e14;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfce6fed50db7b52f16dbf5ea3327d714b17ca7b67733f18c635710c7edd75d87aa2dacf4837424e4dd10af1cb8f1c3988d66a3dc669f4605aa2289731fd4f8f28685c23139314665d4a155333e88ae99652cb041c1a8b980e553f35e4cf5b7e16500ad2c2f346c438dc4e1524ffb2f3f8cbfc8a2db1f14aa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10312c193fa0b8cba3b55b6b2dfe521a562f362fd8020659114b140dbf557937525980188eb08faca58550f12843b25f0023d8b0a9ef05562f4f63bd6d226f84219a919178eed8eb15766e6bceb44ef1e73d59b0449a89543dc9f47036a3ce6dbe4b6dba18d9285309c8bfdb27a0f8ace1bd45407274ca10f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106388410e07c6896a8486f6577db15a169b34ddb773b596a53600433ee0c30929d833e13e59be71db91244a319b9afefc10521d58e3d4f6a99223bd1dff4a3da35ff6d7d1ed9f94462dca33608c0262b39488d97b1e5e2ac0fd9e15500599192577554a98e6453b9417ef08aefabfbd01c14cc47d8411ef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h29b555c8fdbc8de7312a38429aaf452c32a228fb4eb886c90adb01045ec25b4b60ab653470d9a578116a3e1aae63d763a5655ed6fdcc1fd57ab2db16c0b40f5e25109e12230f3a247f4a7509083596ec709c0cc249c64805ad1f96fef07fc523266f5411d2ee332211b1e6c75c6620867dd8a15ca0aa9231;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17d1db1be86db8ef0aa373349e1ff1410c6a523c66862b897d7c399fdcb8d6c095cf6b5adf161069b7b46af3c51c9420ce8125ee8e5a85ff4c252bcf2e88c7e7ba2fbf97503ff7a97af11ccf6c3142db5b87531ef0703553a0de73cf9a01b0a275f2ea44dcbb3c66381be545e0f508193e8512a6a89541055;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10fca3a7a485bd9111b0d4619af4f6f76ce23c71161f2c80800f022b002639fe92cd5f90c3f02dec6ece10fe893647ae584bd3d09e1523246d5b76821b810c820974b61c1fc4df85862b96af9afc70a6088ba795ecf4721b439ef5ea90c9e4daacd50311be6d5c81274841b7a9ac2e5f6a988d919bd763f9c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd9d5dbc065cdce10e548f03ec777e7d9eade6f2bdab3c74ac950089f4a65c6e4b6a4bc058a879857de2ff1c94c9b75130e0df97c8dbb5efe896b84916c54b0ad9a079830a5d00814975d9457aac1b793491eacb761243657a2e6b99b6373f69633249b0d5e86bca9ad9906afe4a0c2d0177739e5cd23206e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdda76a9eed3d154bda4027cba5939265373a3e30ffeed5be7d6ffbb8dbe078071c241c69d76bf6b38985fc27f12b7c9fc8f544d7b58a7ea2e0687a89df5e7d26b9cab5af946023ffc0eabf083f076bfb6b2544910add8e9d82b4c88cf481ece5748eee392d1c8bdda1aa8566fcc67570e8b3775ceefa1425;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d1f1dbb378ca93d91136715942cb7fd720c3f9b80b03e652323bbd7e6e3b0ae8d1c7b1283f63ed13034c58529eba04e672303f07dfc69f1b2a480dcb5b19b2f266fc3bfb5559bd0fdec0f050099783f6e7dd7d4fcb456e08eb4fa046425ed00518d75bda7bdfaebc82643f056a1d838df14edb0d6a223d6c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae1cbd3bfdef271377bdd996b40e50daa65135cc4ccae906d0987c1af61ce753230af9912044aeae913c7765d0f1998469f307e770c7cead9c6ac6ec906a1ba999323b2ddb84f02f503e68cc1131ef5af6b8f3d1f612f7031dc4fcf3d1e49cea0ca51e1e127e59127035acfff429a3e8169bbdb37c7bdc56;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae8a7b5f66788efc6008298469cb0304ceeeaa4faba84791f99fcbd33b9d56c7dc70440e5e8c93709b7db08693c5dd4639b0856863d7e139b7aac7ae2a3ad736f2fd216943b709c67963616638cfceca64cc6574e864a7a72d897712c4bca4a33caddf6000019e2a06e83a5d61feb20d52025c67176aa942;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a27271abe6d87a3ed0091b4dc23fba14b2b8fe1b9de4eaeb82e54af6607c5231fb550619126ab1401d179b64af9a34be22f993661e4f099f87caafe9695eaa747e23f0c779a11c62f106f34f4b25e78dcdf84d75d8e024bf28ca0dae94919cef92f176f1a82774ab117739a1fb2fbd6889dba763f5910705;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb70301e8d304e3b26329311ff7331db73023e2dfdd52b14f629a0e7092039ac83cbaedfa1edb9acb6d478ddecf7f18cf3bc7894fb19b5793b757ff279d5aba8e614a1b08abc5d2338a442e82ed19a5890f96255551bc7eaff8a6f5e898fd9a63cde27232b24dc8e2e72d697e4516c6e614b0323b0880a052;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1170f6b2a0a3a665f34a91f7a6d6aeb7924135f8aa2947289811139dcff3ab41de8b955c36228ca4f560eb573acc3ece8b385af81f0aa23f341800a84da70e6a247e8eca66437563fa430e10af3560bdd59dcca30066a36a8558ababae2ee694e7a8eb4c4183a7c3046b5bab62e81deffe77d0233c481c241;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef512bebdd1d8b05d24159b30778d19a59b0e74888091afa49fda04e2cf8415c5093fa61019e7b67a09c5914d5fdc894c174f7eeff75b988c6978f66fd07f422d21eedf1c962d3a6a163bb1bf04a46837bcd77400c5865aeda9d3a5dd5d0eadc44eab7aa210cd003437fb2df7b32deb83a12262252e8b32c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4bdf319782dee57f99f0fc18486054bc3a06baa310077acd9d806888007efa48f5b24059ce1ae32c746f1952489376ec5789672a490c96354f97e9c51be755e8f24df42cfd6d2d558c5ea944953d4406bf3854a247a0ab22ce755cf0f7aa8abda8238a7cd23a5b802a8474082255a54c1bd04ecbdddce055;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e2d94006e61f4ff515be2a0b318943d28936db0537f333445d3142aa79df98efd80a61e4831a0a9519685e05f5ce43e3a07105368c677c610aaa2b623bebb506cf47b062256f07ceee4f8702d585addc3dc85122a967068c4d38b63ba7ead6ff4494dc6937dd87543cdeaa541302f9d345be1530034f07d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h499e48b42050a74b3b26833e0e0b2ee5be8693b504478359f4ce61a1330b9c445cb30c1aca497064cad61a5f6da79919a72a007802d0c47579128f6c3e67a61a5e8f136af9c4cd6094faa7e6c93d42c808d67a572bdacacdfe5a95d84821f9dced268a1cbaf463d53f1515e42dabeb156d24146b0af10f68;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16346154fb061aad3a2c9398019dad12e56a0bd42108167e64b4ae18d69510c57aae8f9dec8d53ddbbbd4cb677fad683b5a399148647575b1a47f2857e6bfd4e846f33e6b0a79979e483b7e1613aa2df0541b694ebe7e8b8282b79188b3f4f82a5b616d8235d0ecfe8bd94eec4b3ce51c3f933802dda4519d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186d92841e01632339509691076c0799fd8be1095dbcd2529c8208fc656efbedf51fcb7d3604890c95abd23fb53a4e54a024490adfa268fe5348c2724698b24e30916c083bce5775312924d9bcf41b34e50d9192914416ee89070e83b526a348594c358f98d114beb3239136558f6038ffdd6a43e04d68f21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h264513ae2dde3f0635f300071732b01759d9762ea972ce81534f1fdad4fe80c77ca578a336c5b6c29c360f9a8f2b621da9bda52930c2a334a4b11ba038ff190f0155b02a3e810738cdb55a731abb9ea2034d5045a6f522b66a6177d7888113b127372f1b5195bd9bb8053ed6d9f18b2953e318fa6ac2fc63;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e997eee5d25564187b2209d10123659cf91345a6f3c02ff8fa9d12d15761213117f0c5bbae91ac76e1db3208111d0184920b6d1e2f8d8df10f3f5f059f95efaa03dc1edf5c9c1e50b524f92b3861d066cf67c7e9afa47d35a3c75926aedbac44d608e26bcb2b679bc7618622a0fabf51d2d6c1f46bd5280;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17bbf8f87fa6ce21285f3fea2c8cf30b7b11b9ef0e62bb53583c68341f78c8055fba06e8a4326a4da22efd48f511190a49caf5d1a28777d4ef9ba0f1f85e6c0f6e3811e8d68ff9691d8b71e737e2cefcc970c7dfdd665f154494fbb2b33e6a2f600ece6b86b8ee0cfa8cccfb1b5de2a8d721a123d4587a925;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b6f03f9a0c144474a2f9731461d9ce74bc6959aa5904cfcf2b504249afdcc64bec8a0ee110b336d718da2163a6d2ec0cc47b8bbd2ab6f21ee1d8632f69b1e8ced9553eeed67c48fe2ec43404b72297186f40fe1ae688e6d147009b3d08031a4c04204727baf153afaecdf04e26e47d9eed8f816401c4614;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8620b17fe55db8af4b35dabe1e2e7dbe2f40a939917dce049d095cd74f282be376df1ac143cc072d5bfe21d1397ccdf5f93e5948ace1e004635041fea02637a0362f5465f0abae6de59bd0a33fd36552af6301d8794fb395672725a13cee95728f0d81633bc863beb95f23a1734bc05e40616a7dcba6dddf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52e26d3f1dcf68d2b9ca0023e8a03941ca948c254c5ab26bf4086b2bea361ee1107008e8ffebcfaa984f11800ea41c6c4915b9da4a7eea0670b75c320a91c7ecfb60d10b22c68736581658a8485eb09bb5c8d247bb2adaf5fcda54cae0ba8e543b498c2d8cc86f552392ae072302501a36cad864b59ff2dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16965f8ba6ff233105fbdcde49db6f50fefba0c971838a8f213ff150cac9e72d2200533408e1619ec328f603d7dfae56c9dd3bfb077ecd857597ad5de610d0f703853eb70ef8a43e942c41840a092860bcb3e968b4994afa6e91288c491039639c38377f8e256b8ebe79e209e56a3d983ce5b35ad260071fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hafd7070cf140156e3eac95c1baaacaf1f884ebb920c92f4d0e4d0ad07af043512111d1909643df6132d12702e952a351f4df4b16cf332c2fdc2d211e86460582ddaadf53d5e7dff3c0f856ee3a6a7b360e11b9cc1c0eda7d876c5b27b57a34c113e5daca1993f1cb5e6aa01a3891ee36aed4482d080b9ccc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1edeebfc68227b569d383578755df09d5aa85715291028bfa6d223f0b3d64548a54684df27edb79e6e35fe013a1878ed499d80e31807d8473892a53dc6476271d07475eadd5c56dacaaa2f42bb26421d6228e7b5d483ab966385711f3b55e598d0dd046e0fdaa739e37b2ee4b8af1cda7272be8d8f88ce487;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12041d07e633552b72f0c3af9ce22c146fe4d1fbfc0131ba75f31a3d85a2d6037347bf4f0661fbc13d76c9d25d41c1ba72115af794c3895724793847f874712f70a02e54ef8abfa26b990379ee112c1800938d59dc752bbd7ef79f608856aebd12728cf07b5774cc26b7dc301a3f31c20e9ae3256286bc135;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19827b0ad0ff1492602e93312d495a835295a47d4828ae43bbf63970295f49c946094eba1af01a7e2e3c55b9c2e3b67be373a7fed5e178fdcb4f564490f4e60fee8de65ee8423d5035c45ae454cca1738413b0734e77f08668338232d30983864eb528649a2ba31b3b0d9ffa6005c2ba7f3d155c629369bfd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h704817cdf0eeca6ccf8a618c2bfacf1effdaa47b6d8227a9ca2587f7d64571f16218ca80f6798ca86b50098ecfbabafe6659b596e1ee48b403d8a203205ecbd122fed2944dd1c35fddd183ac5b8db39e668694f39794b4a4f267bd0a9ed260147aeeb27a1381b518051a1d5ab2b32f6abf2ab2eca6cd81be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a500caeb7b35293f524a15cee477523ec9a30419145765a6d338bacc211572874d6f1d4870bc0ca07161ca391e7ece4d38cbb852e35d0d2d7011969ad7c3eae62019d982cbcaac3368921ce98793b512ae7e40210c71b76ef0e00306342d95503a5b87dc32dc2483c92d320308faa8eef0da8b1c5513ede1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6ca9cacf36e527aecfbda17f7f05c1ac61eb3e5282b8e6f16bd5fe2b53f82bc77e5450848e3fab08f22188ff89a7bf85af85487aef4f29fd8784c1c7fc01af647d267fb42cff3919d36bf5c9d1789d3acbb2957668ac1eaf09922afe6a1c4ae87932acd43c5a1c2eb3ecd2b0f01199a0afaaf6d07bb6fa7d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h808158a61b4081f7029d3636e80aa3b60abb4063c5f63fcc15b7f191840d9ac4a2add91124b5953a1779b9492ae41060b8e2d590fd1034a106e37eb228a1123aa75a56db2ab711606a9fddda2f8d59fb941ef6b7ce66b9a8e1a3b009958aad498eb1b88aa9f82132fa3e019b1b579eb7cad4ce07859734e9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c340b1bb91687aaa4ff2e77451cd279c0106987c0895e3308e6ea31af622df7c6c693aff7406bee7b9ed61befd67d110ea6c77a881a56f8a9742019a737553ca528c63a80507cda0db4656ac39a8a4b9289dbc27905aa139c19f716a3791bcc03a438d6de1495bd8d7430f49ce9e702e1bc0e17c4429fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c5f33e03aea5c1d4c326bbd780a1ed555a7c93a97c6f869520905903692c9e0101d1e59a6d3f8b291b18030d15a4f702cf90d975e173838f927d3ddc37eaac5394b1880a5651e726429b9f6f21296c90610c60d8335d261f3a551894fd08593842de2386e897ce13a99efce96aa500fb4f3b181c19963599;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117f61d37b6f7cf11be1561e0f8d4fa06f416d61503917eb3fef86622b5a3150e908d6edbb422c12ab513f2d2bca57b2b35ea974424f27a7a0892b6bf2975e23a9952a859394d6c6451454bfdc9eb4b5d48f7fed20976e800ca8dcfebd1437ebdfd104c8aac0b02182b5ee9397b8df22d7848316b15ddb798;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d96cc28c6937512b7324d91f922a61b991cd2db2d2ba08070467a02d1fd8239ef716a8d91470473f4a68370b59ebe840130170d82a235648751677b37cb8854ff3beee0c3a6db5638091893529929bcd14ae77fc6d0187bc511dcdd07dc49caa3fe78936bcf8da06bcd7c6fc024f1f8c17272660c09b383;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dd08d441e0ef5d0a77af729a1a403aaeb7f803a6e472a9726968ad1eff3fbbd9890be653cfa65594ee0f2ba5102c2b1b9a5985892fbef48989afa0d1952118dcce8362c0a8e623c69c795d150ee49c4237376d35687f63008f025c59c747d74e21abc339f63c6cdbf24e638e1eb8f226437afff9f4ecf7f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f048b19a899c4128ff25948e880b026ed603f42d47407c7a3a863d427e90aaed2a4d4fc872431df55a062847be7ad88ccbf7483e191037f5ce4f1bc6d4821409e14c6aacb070e6bd8fb67c42c480bdc9a1ec528f4513882f184262e0475c3dacad6e1c66aa5cf755a36ada0e69c9a2fcf73610fcdc4cc796;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e080b0e34b8b52ed1c1766d18f7231846293aca640f3886d95985d75b7887585138aba5f2d267d9601ef8d573f3468b47ee8745ffc7ecd52a841bcbf6fd3a50c8fb9ae7a60b4098ca952b58fd22961dfa9e9b46a4269104132508365dc7f5c88ac7b21e6746cf90b9ea4f857e81b05867646878db509e31;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ad5442c34d98eb1e367fd29bdff3ea89d28a4cf82faf153cdd36f1097dd72232a6886b4925131d7d606c898835e28931bb73ebea3efd6b85d6ff92a2b025e58b18bd78bfeca31d5d690be6d19db134eb03192fe231861275460381b400078b3c0733d29151091a88c2b9f5cb3be7fe86a1f61d7be7a53f1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bcc8269410371695f14018ced499d6c95e986e50f39567bac3eea07c6c5102b67070e491296cf9f6a4ea84a5583b2ee2077cf1a2acda5ec44cd1fa11d846471e60c8ce6991506233eb21cf0d61835a192e31bee882f4eb992e3d70b01fabf8483644aa95cf5d69046bb660181d227d92402311f2255f55b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6c21c88a67d909af7749509c086f4960046d6983726815b6bde170ea47240857d441408333603593a37a42d76859e5cdf5695761e4eaaddd9c34bee0fb1ba46fa0579449f9d4e9256c18349cbc49aa93c01868c6af7cfed08fbed24cb99dac5024ae3e4dc4b860ef9de72c5534ceb864a1d5dfaa67dab213;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16671bca49ab60bed2a84086c038ea54830b976dea72b8394dc3ab4428294b8212b93c1f7d6c11d187493eef94ae8a2f994a08c05d8f0501d1c02e5e48b0cbdecc80d9373eca66e63d73d68d3d67e6e5a6fcb78b97f9de3c8f08677cfed692805b8559886dc272a0a67759fa2218aa1c6ef52fc9e9613d3ef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h126b781a1be4fc83278628030b87b0a21ecbd1c517099fe3b21138753c0ea97cd5e2b98f9cefa28b7944e7477993c25de4f0e5226f2ba04747cbe2cbba9341c2193ff3945abfaff2d244e902047f2f92b40a6f4387fd6c54454a076bf5519bef779910a746383a12ebc80f4ea3c565b4e303cafb9999b0561;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf50345d878bd511cefd85cf8cd225a5be9f679fdc3faa937f9d6f05cb629351dc33098f6bf71ea39eb976d49cfd593f6e99efb1699c772fa4e07cdb3ab8d56093e2d406d2846b511707e396e40f06cf9859fa88dd31da95de249a785883a4f0dd97e832416a9178ed99b839da73e581d6c7c5bfb18a0cb9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda77e0fd101e46e5463ce3e171a2d711f26d31f84598a8fc3dfd5ddeea3dcca70870a3f968211c0d6c9a2f5cf1a8c0cde3be6e49a48eeff7544cc0db3a4277dd8a61214355e6535eaad37fb309b515abd0779c34e1f835201ee317c5ee4ef0b592b6d639f1764a69705a57e14871100539756bd6321e502f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f23ca02d8a1269db7f467470159812a2221bf7ed0a964524be0237a64eab9a7248f829a5702255718a794c781a29b48200cb5cc770af0c742fcc7ed466bfdaa45b1eac87fac3b41575a19718a0781f931521fa5fc24438a81d8779ed6013f36a817c8c1ad47efd6b57423ce8b52e3db2d2ec5a9a97051a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa93eb74a858f963133a6925c9fa0d84f6fc879e95277ba2cd1cf3749b7cbf04d7b9b7b02967e5d9cc6e5a55a6be49a2d9818a6c83caa2130feece5e8b861fd3b603b13d5956919eb4f78deda1d8cdcbb6d9f7500b286f829fa0807fb1b97add51b6f49dd65bce297f06db5bfa3b8d9c2db3ae223a8732d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h59a8484c1ff2de0ef5f995e969480906d19815af797a81eb8069355feec7b0850b088c3476ff9aa16c4a734e9b001523a392b155da59e616823afe0078bd74934d957293bb36092ce3629b9ac4025049fc8d537e86eb3011edc6c03a4fc714ecfbd5fc619517011249851dcb906834d18ffca5920ac2f61f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e03fdb9d5149ec74456725c12d6b95ef1d9474332ac740d757269087e43f73b4cbf15e4874c45433415fc23036355e3768a12188628a824f3e174cfc7866cd7a8922a01de2ccefff0e0e7e25abd1a0f58204f69f2615ead57e664e9a51bf62455e7720c5bcc913ea29299c0b45459a600d7235dbbaf70ff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfaeb45745e8ba0da41dd07df33a68b6e0b06677a4e467916bfae6ae8534834bcb4545314bfe1a86c5b6a7351176dd9b7b685342d4eef6519c27964a40b8c0ec4061b4cf3455a3b2ab4b74248253808c0eeec91a254d2da3e9068daee1c33b349280fb6ad42ef4121f0df7af3a052ecf7ce2dcf1e887f15ca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd9e96e2f458938bf25cc5cad9ccc0770427c5fe3f1a5d3cda2772a571cf335c5e370182e1ede0fb0165618f73b2ab9c206c31100afa91403cffeb0dab9cb3dce8e4c47b82bda30b687af3a6d3e4d26726b84ed8b90a20be6834ba37b91e52cf938b8e36bd8b65726361ced75fbcc48881e1d8ed35caa955a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h107ccced80bbfe348b1ecaf65de4a6912de19c29dca4dd006bfe3cc8a85e624e352eb40d7e7f85410109e774cf5fd309431873ab24a60678724f47fa1b88d4bf89ca3e0fb238a1bc6c8ceb99af0d58d2828693a0f5a8bb9f68a7c75abb1251741fa508d64c745a15545de47205dead7e6e4d79218fdedcfbd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3815035b636dc58b6fafd1941df81eee72b0def058401bb01edce7185c16521e0ae69b43d1ddb2654272b60ca086ab965401204f310f48945950160b23f3883a7deb59e21f1519ebb7a9ddfbc3ce86673549934dcafc31de131fd74da7123b08450b68c16042743578a698911eaf9e568de9768163dcd25b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h976a447c6ee12174bce3fe70036e7b135c1173d5eea87afdbeb723e11461f2375345e04ea5196dc4bf36b9cf7d4c139ed1743ab039a4788a5fb633c694ca5e4ba25e75bbb384f8928e61d2a7c9c4157fbad6c402da85b8e82962f1ac9f48d3426e992d6f7cce2d1c8dfb81d5d13f05c1ef2c776f69df348b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18e4f00f4b1250427ab028eb4c411ed1205478cab4ce204c6393b4c8d682c1742328c68790d0305626163f2d4a6feecf262f975c93b279454168b312fbd35bb22212e57c954a87f1f72c6483c1e24866c1da92a868f84e7ac313808e494d7ec84a1dcb7ed8a9d2fa0b053b70ca720dfa29bd358aace237a28;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h781aef8bca52b85b2980e101ef196462a92b19ce5d8c00c4982dc37fb37348eea757de7dd169c2c26148b3d4ff5bd83990cf3e85c85ba0293d47b059fd33b31e0b48a0e7ad7c3455e18f15fb9459363872d901d48d12ea80e5464fd26e6686e83045c1c368cdb50c9dc3894b14b1c80fac544d73cfaed399;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h176e89682abbc54bcfb8c15d51f65cf88caa197217c1f0d71bc98040c4ba5ff14cb15b905975a90e5c96c6f2bb6feec235fb4f3e5ff593bf27c8f4b153cac91cab54745da857cc793976d5a7d6d5cafbd2bd63aa4919d48433c35cfc58dfc6bc8ba4af41f23270b674b317f7cd421ed4460163a4d603676c8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18330fd27a949f737b3316f0e456535072fa5a290cbe682b4b2855a991a2eb5d96604e2f9f478f5a1db36f1ed61833806ecdd7af39184252418d0101d3f3026b2ff1e17259b04e10ae7126b64ba19ac33467488bf305360ecb30bdb6582d66b05d15b31a94acf855875e1f3bdc3003b056e8ceeefe18f478d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h207daa64bb2c98b453b1cda7b0a7cef597ec9131e663f122964a679bfabd712465228d1c81fe7bf45d872d4f7f1131e9ddb3c9de1f0c5aa03ce57f3fa0db2aa295f433d9afba5d75912cb1dd75e7072d060d63c47c7f6b92170409c72037dacce32e4244424c2bb3082723e00086460203928893ea65b253;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1d8f9029ae1d89ad1eaebf9d15bd845cab5aed35a445c1ba4bb4945b8d3d1b37eb6332b6867a2ba29a2f187eaf9328f022e345c6dcb5617784d9107f70939b598ed2ef93d38b9e58778afdfca20b5fbd0ddcf296fd2734819a83cba6a506271b8e8ec971a13b6270258b44b884791ba9a4a27af23eafc14;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf854dc1bb15717db8c69af0284228c10628c2c5de585bcaeb5d1ee156ea7973e3dc31c5f5b218b50202a61b9763a9a67a744122bda5330385beb83887fdd2f3e48ff7a6f7cbf8c86515387b1bdc28426f081fa410fcb2d663c2a0952bd34409c26aa90616d2785509fd54a7f351f46dcf7fecba350dfeb66;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1204f68e97c891586e34ac112885b17f52710cd4978f87d2006ba7829e874e9d521797d2817fd47791d29104dc9de6ce599297abcc71d6ecacd1515d55a54840eb60412fb5ec79e6205f037c30605417883e1cb6fbe0e815e7dc74b00faa5df6246f2dd16941ddaf9060c1e7d812214e710955ef91d6ff97a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3797ccf00af72748bbe07aefd13fcf693d23e5f44787ab3ae59407cf387f78c7056f95a637aae4027133a839b2731cf61c8046d56a91ad0f34e5fc35f06667d6088542b4d2126bb11bb16ffa597fc07076ea68eb7592b6d911a1ed03ffd548d1057f848aed6db6c00dec9eff7aff474954e4f2cc11ebfd5f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3094d72b20d87ab950ffbe3a7008e0824b07cda042cd383dbfced7bbcad1d22e374d98568ff500d60bbceb0cf9947e0b24f0d732213e6a7fb887e1acad3f77affd5c473a89fdb2e166e87ee0f958966573a5a682a4b17113c7a0e6f13daaf6b5008fe899f022a6e3028f480ca7afdf04f16c8b1bc80dd66e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16432aab6dccdfbde61e002c11fc9792e3becfdc45929b5f535f7ff1378a719bc82c76d61b0e508c678f48713059c31bdc010d071d9b1ee94d5e6ec20acc2b8bd5b8ac6a6fb36c81c018ba1dd0a6b4e1897bbf1a55aecfa37fa5229f43cc8ce5aae2b82d77dfaea9ff1f3bf157198d192e5bf8acb56c22dd1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193a3ab4221e2f0c268afc6ff2b5a17b4ea4c8e54153cbd129c774fefc2bcf2fd30752d84219c56a81a4bceb4a59268256dbbdbaac811b459facb71a8f84854b3e430a1bc449e5d1370edb183c0c61ba3c802e7a35dc36e118205bdbe0d86ba821fd580ca598016a4c4589cb46636867a9543c6fe348e3ffe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bcdba581639147ba910c13c9bcfc2935abe1ad1017db8d9d0cccc83704bf5f152667736935d3c5690469690c23763866f9d5f1a0cba80a8fb024b1867c206cdc7dff9b494010a60475907cbe22900e1dc61afa7d2d6095a69f9cca004fcd63bf8abb74f82e2e65a9784bb1dcf09bd0a61b208c53eaa536f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h48c0ba8efeb007c268cbd20ae025658324e29f2bd3f93a3a68bf5157fe83007d3c2a61b77a204b04abd4b46960ffbb7a1c614e31e29e0f36accc8347591778c86e65fdff317d9fc51f32bdf219885c6790e3078f0f6d598ba6b0a8007628dd83f0218aaec52a08607e7a6fbaaf98497ef0e2d9607e2f48cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h130bfe0eda5ccfb99573a5f7ba9a7c00582d591cf34afe42b4e055db54555f3738d1241d0cab2e89b2297ec950f23fc6cbd6b7a3afef372e65430bfd0bb68b72bb67107c6a3d8f2711f26dad22080e9607d57d693d05fb1e9fa192c7d0ac0cb46faac8f3298e8405286d18499ee6657caa454f74b2af8b175;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfcb22533ecfbd9cc2c707e2d31eec5dd7746d7978039ca41df6c0b55e73e300157451a2832218116e0ce68fb270e14078447d07faddf4d1314c7ac2df71d54e74b8365127937707ac4328fa4d5e9d5127ced48f317ac1d8884fcd26b07398e95ce3e9004ec6e545caef88462d12234caaba89df414284f73;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1902bbeca577efc629ef98e1c8b4713909038663d86ebbfee485be339deb5500942ed34b04d89e912d74644d9c0b36a19034d019a66f38cae3e0fbb99903ef0d28f51426cf16ea7bd2753b54f07da81383879b674a14a4c7ec8e2c1626b8342f95895e72d34436d0428e733f3cd7f3c6b35886c222ad4199c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6d5cabeb9147f8efde351798b20737fc29d338a4e114243ce9e622643bd981cb936c81cb2162723fc8fa662bc1360721ccb953635caa37490edb6bab3f5bb71f2bb829aa51dac213ef3f0a1d11b8c6cff9d7d9c8ca4da5e4c3bd79e035e6177f89af97144c885df125a701e29307af1e42fda378411bd900;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17008851e3455a8a61eb69e089b9c4cca4f7605aa7eb746e3969c1750ffe05d1c03cfc7dc0b725772f11a154a4764c903adf6c063cebb920f35fde84c2f3b80ed8989b8762881d0b7a13b010125cd775db290a5e196056dce90a655a5af44818f5f51d6de52a6aa168aa5b771f71bf7edeb6fd57ace56ba57;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0b70fd850871933f7e8fbbdce33e7268f339fd2d4504cb2afffab69e6ac4e7cddb3f1c32acb5fc657cf7663fbd1f87afb487144aa29435472732c9162573b06ebdf9ff1b6914fce1091bd797961b2bf27a53d3d99c847a0cd9de045e4d4f201a1c341bea33705b927af598ea7a62d5231580a3178288726;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d296c5ab3bd4b18ec1ff1afe5173c5f0779e6a3932fbc125651663a2697d9ee141f5751ac1a91496d90e1593aa038d460e7cb2ef510fdc6d4e46d81aeeb3c99605ffaa512ed5b2b1410a5512973af2cb6daa7e693676a61d3a03236e94f711bc98f577abbdc90eec33c308ed553a15f8c4414369cac19d3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14fa57687e8093a81bd8ca0c4edcea215315aaeceeff898a3ac48af5a45af115934535f550816d866f0098bad7c9e49467224cd6719cfbf374b22e7805eaeb7c89dee5d00fc0543d06c9fbe7f7709b054a14f64b68553b7f7c863254253aadb47d39eea27c307131cf542b12d85b9c08ae2e4bdf548e54a0d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h309b3091ce42e1416c99c8af0eb45f8df98dc8e427052df30957fda57f88789ffabc7e5677db2922057be5f6e002947742e21e5555a8a77c1dc40197dc3f87640fef0016cf0438d639b28a04031e1f12aec4bcc187a2191a86af73e1ddf7172c8c5752c2b8af5dc7bad386c3a6e319a9aa4eb139744d37f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd58298e6b8f3f611be126bcc45cffc38f721cd69f0480bcca24c4382af445af0483fe583e19b1db16fdec297071acb11276e7fe86d144a4e26179fe80d304ffdf54f1d368b9cb4d2dafade9bcea8c6366366eb967d6973708253117bc36866bacba47e7d211a31f639db95fc60622f8d1f6a3beaace132a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7cf3e1a7de2171ea40557e5a87df533b14ae793ed89af86e4d9b7275354ce4f69b60ae38ce0c9dfb032de1ebe3733edba961f1c4fb4980f1f0fde22dde89908e88a9e8a07ff6251d8fa2e41ecdffed9f7ea9c5df410075b331d384ce8ff6b26d8740eb8f47c1af660c1ac9a181a8c48380b658de2cb29;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc06cbd3998db4cc2d6e1b38de5f43c4f8abe23b04caadef2a15650c6c34ce1150162f8f4a88f5e9d188dc18b5eda1fb97fb953142d60d23ea3bebda6a0afce5f4bdc3011675f048e3f426227e2d546aae8b31927ccf74adfdbfac80045d52504e2ac766d6a07c2b65ec6b9c901a93d31170fa967f1d7beca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11962d3a50b10a6e7595f05f0a5a9f6a9d62be94d4ddf35bd8f71fe1f59b6d790ecd920fd35a0da0e72e0293af5107b2305b74148b8ac009590fa2b8f01f110f66b2d63b094eb91013024db3cf4a83e6ca7fe76045c6d989e80db75c15f0ce0ce04729deb51a58c05e6b849a3c0dbbc59b0f78cb2d6ae6047;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h144c3c104eb333c055265d879bb4a127f379df6850daf0f88c8b33239711cd4d6d7e39ac8d489dc3fddc8d5166e57db313faaf154b5445f6a2ab4eddec6784047653d788439d9490e2b87e22ce4611ab62c9811c3fde456bdb5980a3d58b5e0d3aba6b1c5fea6eff554338ae7bdefa2c0b2db33a766a85740;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f6db5b6ebb74d5ede049dbfc0fb17a2bde59045af2d4e46e7233fd40610fddd996fdf67574b20c9e9b4a71c9cce23a92879932159a3a7350c18041ccf4e8ac87bf8109a7b1f07f976d0554f29069981c2faebbc0773160265bdb6f36e2a4c641614c0632397d3ba5a0dca76f6b71b8f3f6685e61c86c7796;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17568df8072a5de2851c11a567de8db900ede826013688e6eaffa45ae7713db72781119298f1b5424ea9715e4fc23385fec521753f32873552375e2260835f87bc612eb792ea1163d9456db7ad77b4a3624004d964f5ffd8046365784a171ba2e6ed2d3ad4a806371c693403345cb9bbaa739c54959bb54d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d31bbef582f03310b78c21a48e56048c02c0b05af0122ccec88433114f7f844fcc8ab5c6ab231a68949c3ba29b7239a4586624ee95768655b929fe7f1fdbb46ffb72fddd741dbd0cb418d05e5749e740615f896aaaa873323444262761c41b75f137b1f7316c4c91c4c38aab04de47288c3509c78abdb9e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15e23151001f4f3e39d11dabedd39b3fbcf3fde28680c976711216f5f7b68d746b6e6b0f3657c6d080ed0e0d414e35a2840df535deb3118584038ff48ef5d12fd2ef8f78ea1de06a3af1c9413192f35a89f7dd9f8eabb19f7b777a4192728acbf4c428f08ca310786776e49b458ada40a0a298cc912c903e3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5db2798c29f4dd8f63eab5fd5ca87d9a68e60a149475811b3581baa41cf32d6756a0620dd32d49537995c8afccbb67730114998d33051c6051ae5e2d1603e02e0b773aee4738eeb0f634803162748cc0151f22d471737e328a3ee06c0b6bf95b66c1c3714dc51cf7e480dde65d0b084d0e37bfdc5c330fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd07c25594c457fd414f78b7211759efa61b0f7c8d40624c8c43a531ae08657f5fc31e04f396160d4f9941a11a3d79643ea3f6ec37825b60727a2ab6ac8fd4759841a61753040ee450094a0db11c9208c73b95617513c2d6c4875a2cd9a0bf4319ce9b3ae98b30f6a03cf132383477b04de8cc033ef6f395c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a9bdafba806f8f6516b525b65d238cc9e1cef125f97e0dd9dd4fb6c462cce625f731301a26f361d39e9483abad509d61b3aee9e701532ba3879983f91f3a2c3fc271c48163c07ae3e03303fe49101eb8504cbe57c5d9072487c5d301fdb3109b69b559d362f564c757e985c698fbae4bcae705a9cac7d769;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7735908d6f29252d93cd1511510e4cd3370ec14de4e58d27a21133e736f907782c0a86ff2965ec8a4b0220fecae2de56ff45dcfa8497a72842da2f51005c8b54ac2a19dffdb803571cf62b0844ebb1f17894b39996cbe1c495c191bbc82971adf5617047ca286c8a80bdb44bc6bf7af375f2ad2646076f4c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cedd07ae3a3e58daad43cc2701d0678b61d10c5391979a5441ab25432d052b1ddd366769b150907081a4550ef987b7f3fab831062f5988f5d58277b8d4ae059a008372b1d6b2d178fff8dcd305c3a2f5751de8a94c4a053bff21f084d721a41732b10feb436a128f028be85031580fd48b6fbd40557f47ed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ce5e670a4967dd311391607b453c39b021c4dd15fea14e6e1922658bd8e5c556ac57843ffefc25f372574eae77dab14d6c6bd2e82452d9b923292e515120d3e57a1153b7c3722252113efc161a52629bd5c4be0185b7bd8666a7a536e6cef829b5e0df122bfd0f2bb8397ab3898d3d16ed35b66e4956628e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17d7b047157b2749300db90f832cba24a14a5ab3b7545796ec425a8cbc49e5e89367e95d0b0050254cbd2b695374171efb4b29398a4bd24cc560e7501e135724dd6dec68e53c87663c3459fc220aaf136fae207a48d0e023578aca82074ba57ff472f7fc5149e9b84fb524c6bffacb5f56f392e7fbcec2fe2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbbc210360607abfbf5c35dbe31e1eaac711301277f753af8d42702793eedb49c76f943b59ad87d2c07945043dcc729739b46a90354a4cc043bbf31934fc8eb2aca79a4e54e4c4d23b7f11aa87873cd1b90be6229589351ff169c39db2bbf7506e00dc21794ca037ca6d04a67ee42084e69b4d37be1813dc3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcbe8170df3e2f0b6750d391d211c9472e702b09315636dce89a70a432380c125e6099267cb138739994069edb391a01cfc51cb4ebfdfefad7b01c9263d58f5674dd99a02899f98cc5e4fd27cab33020cf3ccd2eef5c0d93139588aef44877f8586653179708c26fac050d03bec7a97094d8542247b11559c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c26a23bbb96e2b9999f9837b4cad52fd2379fefc5d2ff60029e7a38d66ae5346fe1eacbbe06e6473bc1cda9884784a5758005f73c468faf7c9136341851e440c942d0c03f18e4d4956d1ebd452bfeaf6a46ab0fffb1dc7d3f42b2142227a959d40f96fd34ff0f343bc1d6886795b0ac0938fcb1cecb52817;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0511c194cb0ea831d0fd71d62a01a469dd1e0c62a1c7e5dd51965c99657d5befc96966565c9da28f7abee0608897998650de4ea9dfccdc36379ac5645e93adefa17ba080943cb367de55756b5af82842c1c805cf51467e1a61c411c53df67227cb95044dee19a8fa2c9aab245f071c68ae46eb2bb09e6b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de90b19fd375d59b4778b3c4bea82f08fcb56043b747235b9f0f9e83a265f6a3b713826f75fd22e6a357f1780dfbbfb353ed70ce3a270bd099eb1aad7fd649073ed34dc32b23c92cee53e9af60ca0bec0838a1e7f3abed6695029f509f90bac2c8f52c438bcef51175b46d82c34d3edf9664f700667184e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f749ca84cb9793d2617d70cb05344281ee12bf0d287c2d0d0c3d71326c269288be3d134274f983392b8d45d1786af3d320b6f99149ce58e48e1d352d3ba7488e6a2f91babd44d429bf3f74cd46b28a944c4de276bc71bd6f590f0a15b840e461c7464b27fa85355914fd5506cbe63a93b78bd1ca6f6d307;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113e97f80cb2a8c99d3f161617be6b2809b68530771282c1abd719d50ef32c9bb314fbebccdbc5cb28aac39a51717d52d2a8f8dd0561a20d0857bc61d3cc224db59babef23873ca22167d0eeca79b4a128ecdeaa718efef428d375ba1dd20a34c01b0ddbb3d3b7f932294d2022967a70717e314b2f0b5a0f1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1572d6317ede0a090af76d3e1c06fe7d84225f75d07bcde56622cc40bd637137d2b746fc9424a0b31f20aead9ff4292ac28128595a6c4c43a6040f52f8842cf93df1581cd6a61028ce29df00cb68f117659c1cf5ca36d336d601cca1971d00caef07a0dd6b08ec2d2cba4ab96f995f384edcd181ba365baf7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb582f355aad9cb9219c8b3b7ce4295c14e75a8d8779e7b87cc2e77f966ff1ee5c2284887a1ba9b56a5f2e8004202cff4eeab5c2ca204897232b3b5d86cc68fb8617e20a178540a8c1de93dc45f59f076b08b2ca88cdcbb9961e39f724c83122cf464b85902f47bb2896d58f8a8904a8cc7d1c554604279c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193981e9415f941a1070f287935c78cfa05557d17a34a04aa2c769f09618fc066146678205b00ad180101c1ac3b874c831d8eba029e8a694d272bcb8f87df11505eb2467ff961070c9960ddf43e93223abd57dd85f57055dbb49c38396018ab0d42238071aa2b4c56857b57d9dd20726c8f66a64a93e72a6c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15e846d9fa6c9c354a2745bfc5ef0affb55e90956373b1466b87625f59891e95a014af90a95d414cd4b898774a2cd3a633c8a6d8caeceaa79e16d8a7b67916dc1d9d024131f2bd0534b79e649ab6b53ddda58462fe3a6c3a01aff74bec0f2accfb0381699ddc1298ada73fa52f27739278345800717943676;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f2de1ad17c9dcf51e44376f4b90b2b1a2a88ecfe077c697525a10e77a870e2a7a9be393131ec4e74ea0dd6f780351c40ed90ca46f59ed227caaacdd442bee1d93c390eccdbc87792a6fab20933df2c7c45d488097f5b9819fc81b23713cbe8ca8b18ca09c382897c78b0348a7c48b004cb000fd509cbf13;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc696947349c5ab6ac9a4e0e9c6811d8f6347689e1f3d4dc5f27124c5e1c506698cd355ea72724e939b9671cd50d961cbc6a3a315c79aad58f3ebce7e813cbf0efdac6c65706e6a378b6fc9c6c54a5a82911db61899e3ed721add648138b802646ab31057f83c4779082116bdec327b8d1dc3636d7e417685;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd1b7183fc12bfd71f47b5bdb317feb3764e00ba8a3a1c9a6ffbd0e58d3a24803f14a16a31d984925d2314b4b8dd4b1b685c41df40d9273696d793694a9051403d0f819c7e6504ddd75c79cb0b700c69135f69515cd13c70dc641bea6641bb88ab1d696f9b0da44ff8fb269fff42ef110315a6adcf1673635;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h62229cf3df3f35ccd34f0e8630ae5483e7d5c89f0ab400b7913cb6e826c8e4ea1273e4ebd8f40d92a139622e7676ebe70fca37cb546effb099134f027614beb48ccfc8ae403484aff241b57a9b284e18ac07d397595aa0897b730f12de9255eb0f21dac7a5fb154e567e93c96ae1deb948be796c64fa8459;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1df232cec638a0d64cd2da49208a886f17719079dfc43618225c18e5d13ea6845c8d23f4343b66719cc1f5464361f2c598c7511b254f655d677b81b06d4d9d59bcf74e878f67089e001fa6e4b7258f267944e7725fccb4baca90def8b29e1777de707c2d75ea62a57bf82852fcc0a379da562ac9269f19a99;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc82e3e8d29de8ea9243f85fe32ded60ffaad3246bb8b52373d7de46cb52cde15656aa0440b9ac85c9656db4cc3f3ade73b801fe4c906bc6dedcc3e0505cc5600935d089c263faa21f4d9efa8f967fd1056afb5960229c4c2453298b8a05c056d6233e21d43a06ff54a9bb4d6d0f802ffd3582a632c6250f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h23fa23be72ab949af4286ecac6060082ca2a2a723731d82878d80449110142b9c89fae8bc08f78ef0ca96f6b5a0732a166900838e62b71c0a6e13dcac8552be9b29ce70be1aa7b5845feca1d06866145218f8ea70f6cb02a3416f58dbb7541a5e64190654cb6404c24b02856b8b782f7dbb787c29b94bf3f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h160bb59a12cc6d0c72442489e819f8531a66bf9d64f76dd693130e5855c835bc69cdd58d67526355d52913e8841e47b99e06d8cb92c9d28bf8b0e26543ba786b0f0d3af95798255569b34823b7efaf4953ebf01a5b53a4757821f8faa38c185bf93faff792973f65a2bf9f38a651ba59547da131d29697be4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef26f934bb06ae8544b6125dba61955f1ba4f2e8c5170b557760f99275eb260ac34b552af87546ea44d9e23b39a6d536000eac9e82c2b3b25edcdb7631a01bfc00e6c6d5e198e7db248a44d52183e54d657666b45a16f0076caaf5ae3b4d5fbd1fc1d8ae88d5df268597a9882b864b5423149acc2581f72a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a9851019aaf8910185c04e30a9ff87bf649904ca907af082bf429b849c02a0868f09804df3e2c4c583961921f8ac7370230fe4d6dea23ccf02cd44eae37d369a73d328098582b7840958f6fbbe123ee494dd4bf25346579bdb89d9f2f52526c54eb23f905275ac02e210e0f5d939028451cd4ec63bc64848;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cffba9f12e16df5e3103b26e9f2c3a2ba0a5a43b7f4d0450ececc08a2916e2994e9661b108d02a169916ee35bbaa40c81fed329dd61ab44eba41aa9cac1f9e55365f1fe7b9426b889307f51425a372fed924760a0251d4e529a1ecf3cd1871d2fe96d42e8fa2034af89ad82246f595aee85e9d73574a1e23;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5e3e04484e838832262e14febe6be9d07c4a8cb1f999a5a09488e0f6476c4b03cf413b94af5ee200407bf079cc4e00cb10edd1b93ccaf68bcb8c86beccb6494ac8421e3f45db17f48d82812247d348a521c80ebdd517a4cfad7e7f01cdf80497b005dd9ee8b5dfdb0e73539b95075ee4bdf5edd62c583553;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1122dbfd330f580641966eab4536c5b41e984ae145993fc9d4bdf571177b66825d77008a3ebb369c63ba9e73a6fe8f8bc57fa562565defb7165b40e4c56ea9dab8bfc83f0ac96f61e63e4216308dc6271fd153825fa10c9c972b2ab08009e2fe768cc005cdbc488867f2b08329373cdd411702da85d51bdf6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6ef01b6f93e34ab66feeadb881a7488bca4af4f7d754d5bac0b528af62cd16da0aa9a288a5893fa89c2821b137eeac0a345aa85feb65b5b22bb8d201873f0c7176606f6bbb97b9bdc7c28811012cbf84024eb289e48eb15f56cb86ebef2837209ee3f401fdf79b13d8dcc7a63971a7a67e9472b2a66bd2ec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d00e441f8e296d58456672b0c5d63489479c45c9a392763e3a2644ec43e49b036dba148fdfe44651695d2717ee4f2d48b515e3981fafe9229e7bcfcf476e4448b1a0053fec2545420b1048ea0300034387961234309f690cabc3dccb79c23b69b57692771a34ade2aac8e8efc498b3812a4f92c37e166f8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc08d29817a63f98be68421cef2c4f0475787f1b3f6393f8606873581a50887941ed3e4f1f000b163d5fceb2981e79f262077124103a7c380249d02a581b8b7f568ea3f11aaf1febeb182ade8792fb1ed05f180af270ad298cbe9635ab3db245cc2c9fcc3b9140cd451a51b599276ce173cbf1cd4a50dfbef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d766ab6dd0f010e78640fe220464db938d6dab032d5c3e6c657bdbc3dfd8579465add7646b71c80a923bd6c2cc564684582c9f7ecc64086ca0d1914fdd7bb4114eb4fe9d7799a2f47de3303cadf2e57f39f6d48b5cf6670eadc8bdad98dfc93fadc2d17f526b187c0fad3cfa115101b0dc37207e5035c17;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa5ada52302f2aef63f20ebec8ac6cd6087c62274d8043a922b826b5d535985f29ef03fe70c756848f4473fc7c2b7c67d39f6fde4b7b657c90d7b2b05f331e27257dcc986cb2f0a3f9f5d4df7fa8218710ab43fac0f68b4fe87ca7cabe28481e715a69f8e35fd36e2e0e671f4369bb80eb487e16be2d43c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha65ba30e9f83091860c8f13a2b32324be4c32067153ee60ddc25e44174da12a8e2f69933223b3106cb505c8695fadb22c0b918f475d24be874af3945bed225a872be72e83a78c0d060c8f3ad5bb5bbd97bd74843a0f45effd20218dbc855838610bca76c7385281b3c1a3b0f42cc0ef0ba98efa9ae7ec6eb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e6783e47693073f14e1369b706158972da84ae58cb36a72c2d3963609ba0468a1a976a5e918c134fcf32c724a6b62a4db8e5aab734740f7ff98d72f9481d5c91925d2dce0142a0de94863bbd9843ba0fe72ebb2bbb1e068b79e9a2681c0c64b86dc36f972937adbe094221fe4649c87ddc345279e8bd6a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137df965610b597cb9c9e8d4927c8b6238e49e50e247e52fafde7c2abac63fa1a606f187c34eaa4e57ef4edb45f5273a23e758c556520589b399a8177bf3e51edc4f864b5dbc285b8dad8bdbc61202bdd1175082af4fb33b7fe383b9c4c1796f8da977467e180ba588ca83f5ed0d5de20e899ad7ec10cadab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2c2eb6a509ea40ded779239057e573711615f9dde4af786f87a94e8bcb47d5d35a9358103baded980162b0a48916105797c849a5ec0632176feef43e417d0c8b0eff2e415fdc4636a1044676b0d2af20e8c6ec977616b20ac0f070c876eee5d9ed9d8f5fb745323b23fd58b7234a071357c3fdd6f0ba492;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f6c7e147905f12304db9b0afe5bf0a59154e9de23f9e3c3a2cf095d7d8b8fc559e594ef917ec559a195352f07c73cc2d60c9398214e0d006304c66fc1078812697fb8996f67fcb8cbfd0985360f10e3970bf0c12f95e67aa98e057a28c3db19a8460801d718fbaad51932cf550bf0a5b3ee6555c0af1b08;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a2b9f48339070418e784d29e8289be4b8c6d5e60b27f53179b02f733feced5700ae4c5e1e0d74503690469116b03125fd0c00f188831b915720eec1a20be0f7383f4b39900f8dca42a47b16384e5198a021bffd82573c836716650960b5006eb23f7ae4f5136c70b0189d6720a9923dadc076f450810bbd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146759f7d9a4a20db0d4940212efa78fce7892fc8433ac7b561c6bfa3492598f608d68669fe96a8a22e65e5cc52846d12850dc0e91e46dc1dac8c4ddb7c5edc3810be307ebe909ccf408cc508220fc8a2a9678529de9fa2af173b7743f56b0b99c32075a9dad7b8c6487ae804f9b73f66a718163eafea3100;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h831e775976aa9ed21f9fe7dc2f48359ceb9120c9c13f032529bf477f9f574226840e0cdcef869a439f9782fdc863dac5fc570a5fff485f52e4f490953742efc6805344a4ca35367db15475f3c3f83a2bc9d29416b1592d8df81a688247e0f730aedf9c8577b8312d4f604d28008085d64deeff6f7d9ae978;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c1c8bcf61a3cd3981aa8a002a5fbffabc16167d46580707316c589f930f0e4ffaa0f344c6addfe8a1733328e31e359585611a4c32a998b4752835cf1fe7353c626e2e121953f7d0eeba4cc036d7a562fca266a399b925f0ee6b136bd277a88642b8341a62c7424c43eafd3e9df98cedcf8b20b8795e62eb6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b9b3b6f7e721217c0714c409f7f715b06e987fdd9a6e8e5aafdbebd745bfaf6a16f3b04166cd2affd4173de69dde03121c6b95a3bce4f6f0f12a702fd041ced7660560727de8a8af7fcbe64841a501333febe73204e444c761368da8749525f7cfc3d3f4d0e17cf01912266646fb4779a6692dfcd44e24b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf7d856f5a4a3801d4d374cc0bea3d5aaea2ff485eac4c4efee15a273f67526d60bfbb7b70daa7079136f606882a0019c3c084ac2e7352184e01785facbe02e987dd238daef2c0f87139775e02c2f027222531bf435d21e75bdd531fa77447b7ba28ca1a44821de418ae96bc9c5d4f52da487fdd916091cc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c5a0bc6799743687c506aaee16a7be1cdb0441ea70ea37923762c30a832074d696fca4b0104044d535655abf0d7b2e79ebc1402f6230c231ee02e2627c738a6b426ff201247709325e24256e6dd1abb3eb1ab6ce8e4125d6405660d2fae9bc4a53b0e70b847c943b5c2415998b465d28a632c9ef8b9a6a03;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e611dd208e9f94f8c4b149866275b97038ac81f5fb379233eab909a37cede2213a271af53195d36b2b7fd64b456f0f9562387252b42d4a91356e22e054a5076009e4016b470e06b3d168b0241fbace673bd2d6d269c69d32c0d0170cd6322023b54a5ca5ccceafe85344e8c9e9f388036c008f343a2f6ead;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha70d02eef3ffefbbbca7d1f4e85552039c03495233f5923f2431cd0d9e6100c1e596c57b31a10d4c8e1007594828a3d667b377b9c0076e498c038790954efda1a0f80f1ac210094db951fc020854c1f6973bf0a23e974fcd982351035305ca573c2baa82c316daeb64bd8dee81a1097e7866ae5293ae652e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e183e95f86688818031e01c3efec07a853cd699a4c5a2eb032d8a6f4b4e7113f097bf02dddcf262047e5a2083068318e0fbe7c11a4da52237fdf2476ee91f68538a2b37b571b5780902696de0c32bf045527b40387cc03810c3d60bd76fd592e34cf2eb4840a0b93e8fe56ae3a0cdb81c29fb31822b2c876;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcfdf589f1a0ea463fc0bf4ea789802d01ad41b9ae574f16f84403fc8be095310ffac2bad7619952528704e8a4e4c3d6f67a1e454aab99054a0ce07e0586ab2a16cde8985184cdc1450a917ada4bf827bd3d0277fcc836bfaae099849deb831e639ab8d143c1bf36356e34028b8134061f26bc7136b8ac76e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6739f33f322a7787e88565ecca7b06a97cfd1b5e868511bc04d5554480d3aa5ab6fc6e3321ac9d45964eee4e5261043501369b25d311f314924569657f9382b3b0662eb08219d416898378a0aae5c398ae1c998e7a170d93e42740756919214959a77c4933159d5e774263e01deac08fa22a63f1144bf335;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc524dfa8cb2ab6cbeb2d6d425a9aaaeaaa6ec3170bd9b2eb80f98dbdbb8177837d65e4fc5dfa1a258a138332672544476687d3ecc9b60f51288f539e793aaf876eafbfe40f73111460ab1fc2618fc962acd76fce6165387f81f7276264fc51b8672cf1b1b608fc323fcd2592c9828eb5a1c741d82ccd193;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10a94f8ec1d5c3fcf2b665c031f9ad360b7e6ba76e2352ae1c7dcf4200298f5fb9d50c417d63b61c67757b328ee24298ed3fb4e8846ef1a55818f839d68c69300fc489540751e131f2bbebc8f3b13b3c52fe764e76f28b8e9839ca996a56a81fca6e9ff85566b5bb312e3d668afed31486852f61e4464a070;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1469a902c2a1876c72e68ec1b508c2e68ae221c113ebc3ab67c26ac180b38b18c43dd0aa69aed5a28564fc53ea645691246dd9a1c77fa420e9b997db215cac1b03d878b4cd7fc24e574c62a6add5dfa8443a00b38abe4880c2e40381af5f73d0fd54199fbb591462f8d751300413038bcd6f35a1b19848a70;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d67a43f093cf56fe5c87f23369d426d83243b4b3f95dca8a6132ef4f62332e43ddd642a89aee0b9863df6925594ca03227066f57557df529f3820f1865491da6614d9ff3087eb52ce4b6e9612b663521ad2b0fd530d798e0be00cb01c693d0a95f6eee49dfaba3976b9eba5b31706c334725b78698b0c330;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14abf0b894d4abb2526331bfdcb81af769f0558884591d893caff9bfac7ae0f1dfd30dd736cb566d1d6f4180260b2b5bc91aa1670c16644a25776c8e39d00f409172c9e82ce4c852db49c0d26ff7fba41718e65aa2fbcf9e9e3c589047f9849de6943c626673519442c3da397430d37fe7ae409b86a8c27a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a23d5fd96e18a5a7492909e907d5dd2fb94a2354b5db187e55687cfc92858566c7bf90a35103d17707c64fb2e06c81df3648031fa467a6e30a1deeaaf6946535c727e7c9595c007681480e172929562ad0b134c6da20b2cf6f3ea732305fea016a4a9c3d2f07bd6c4eb696d23ace54b488ddb0f38c6b1b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c65c75c010d99709edda7f8f03c2e866ff89558492fc687a0c6cc7461ceb7d1d302ddb7ea8986941fa4ee28ded5ae9303030e2f30e0b7c9986685b05a6d055c725a67398650924d7b5bac7e226bff74a0a45f297b8158589375dd5e97236c5d6f753943caa028c7f1bc0edf56df0282c4e89b2d3f221d83;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h21c3d1157506f9ed8f1877c79bc7110f2b6d823d71e37fee17ef8e2f1b5bb54585a72adb02c4f76cfd1d95e583061a4e7536acaad5fb2c1136bb5b1a851cce3325a3e5afe18ac6276179d6e5735b37cb8f0b1a081058571ffc55be3cc0894e993b83151c294fdfa4c93224e486bfbe549f4752d3b857d336;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h107157039c041e17e7609b8b83e4c5555819a912a59a810b8d46fab793975c2e74b1591ef7f00236569c8722fa7e7bfe5d850f17758fd2430b1a3b5ba249f2eed7ac1fc20133a23f1c90cc7207a75b0260cd3d5f247a1429ba29ea57912da4ff58c15b07a178b2b6eb9ea576c9cb797dcb3c18fb4ee70a8c5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4001f721c2da2d8193777752f3eac41ca622c4b9a5b7bd1d2794f64953f3ec557205d85daf9d89990396e1e4b031cb9f004866b91c68eb3b94e5df1cfd3af5bb2db777d9eea0cfb56c71c727558c07b9f6b15a426c8ffa6d64e49cd8fa33c2a00eb42c1e2b9d3aa2d04a56bda52124d830690b46bc7aa06;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2029f0cf48c8408699755f0a380c04ad52f9a7399cccacea87afad8ae64763c1a64c544a9390625d1da8395a17edb1ada6c398a2187d5c5f6e680d896badcb945a8faa85863ef246e38aa0d9a422f45fe0e60d3363c598d5c3b7c9e3c9b5a1237e88cd5e9b2e1af91c5ce1a9c347a993387c6c512918936c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd992e130325db0a39bba80045bc08bd7dd181c198cbf31273d4c4c9b94b6892890877a4c749b7ac3eaa663e462b7a5488e00060a9d7fc827f8d07996add02aee577757a7078890a8210bee68046409964a55d72d40e22b2e0fadcb1d4cc4355b064def283245d2287c9417a9633368284847963fe2ad7bb0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd69249764071a26f61dc3ebae3381b095263a925f9f029d67ac36d127bee81e5235aafebe0c7979dfb858d1eaeff1c7ff7e8135dcb87a69cc6fb717f9cbc7c08ffb668ec73c635e93c569a897383c58660b8a5e876925a2bf355f615174dac10f33b3a983c0d2c6c2d2f38813e5fc0aec9d6c0fa0f6e356b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175a73b1d2e85a429ebefce9117260b1022479b79d5af2ae609109cb9d4a75b1170f7f5074a604191f4e9589977264beaccea619c91ebd4fac5d47d8c111c98e7cf7da595e31e9052930c9ff8a65e4b75b0b92a80cd8c04b7263abf5e10d9c208824f4d68b74fc357a14d8da31387308c303efb46b0286102;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a0acce8f6ea260742fb06c27f7f6041ad67469e0740519b4749ffeb15062fbd156c6ba7334c1f57effb5739303abdefeccd1ed98f7bd331564c02193f12d4c2306d5108984d650bae5372f9b74da59ba7b6dabfaf46d1dcc83d7f63a5bddc264e1de2c96293a0bd81173f98a45b6c27dba142e3e63b5e7c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1491729fb1357aec77e2c4f1c23e4b976213f2a92e1f9c9415fe93246cb20fa3ccad88fbb9d0f9199d2d32a31ab7f688168aa7a8929d707f35f91d945cbee93248d8fb6477077e6272bc697a50c7fa3abeaf69e0499ffebaf0a0d26ecab03969b255bed9fa07adcd2f2be24179bd50baa8785e8b051ff13e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3baf4756424a1586dd91b1e53e1e7eb6b77ec0d6fe200a934170c1a96256ea2ecdabcf601e61944096ae4c6883959dbc12aff8f7b52e9b5a98d04bda360f31d1394a238b27cc47533de3b69cb85949725fb4132a66ad5ac6795070a10979eacad49f904af594328d06d075431720c1e77d3f719d7fff0c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a06ded6d93f3a4648cedfd858ffea3bb0b4a07697e66486d82079f0772c6625178e5a89ad77dbada2879d0502f9ebb3eabf40eb5904d2fa1bad30e7f76a8ebe9af75bf89f0f202592c69fd335017163c17f0eb9d418d0dad3291dd2c1943af697ffbab138fb362eccf0a564d877a2d10f977d6a03318d88;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1188577204bc9416b73cdf9b18c3142d979c620c1023203fb0c6538837007ee21e03eaadec5f2bfd4aca818381c758ce0cfb7a4e35910cc0136e0dea1d25a6a8f7c4129e72c4a728470c10a1a33b405fd2f4fe29bc5c1c93718422db53454b80b8d91f488a8b639eb558fefbf2fc4c5579215f4d5f9a93050;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heb5549e41bcb1e91163ff1d41c910c3038f0d72ab8424ed71d2e5a2363cde55a8606dc4bc12327cbfaaef5d4029b9d88a45746e346983a318ffca49f1608398a2b22906e6ec3fa758ca5917ee69637b6ea9c5bd25f564529d9ff0748143ef4c81ee1a52930112d915ded615c1354ce16e2633d967dfb426b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbf24f9abb720ed7d05b7df4315d69b0ae583a38d99865f967acd3272c6426cca9c675d89e250a09d6d4632dc36c23cbd1a6e5b11fe50bdf8fc6c45c7825b45e133fa0d16b8e33d879b1e796b27299231c861bd0b6b2862801c40a420a34c5ead88e9f9ec8e6708a6613695b4d138b173daa0ce61d27243b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14cf517c1f9163dc3ed03f79a25b4ba65ce7ceb479d9ad2e9ba04d0831e145b5d5eebb7739a55a0f37c32568e8dc474b1f912c54f5be9b30874aaeebb7a32a9a2964a198848c20eca4e0b19e36ac926d95b4a15f7479043e11db6104082f908ab0055c1ca10afa91dd4e9afb8b621214c4281a0dfe7a3a902;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ea339f513ff8130a78c0cb0dfa052d55aa04e1d6718bf7b91478f7a3fa681ca21a86a6e589a7b103bc5cad4d4fb84b1df2be76515cf4c7cc78d041674ca3077e3c93ac96c68190b812bdcf36e42e9f1b1b0b18a12ea0a64630fa9c2a0bfb72d1cd99c11b3b359885dff67e8d32029f5af82a52156fb975b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e94a36de593e109995920a90b94bb578c3c00b259e33aa4ffa43eb9924d8264ded05270002ef058a78d580e80e50c40d69b3064c10a21aef23d2106f0bbebe0bde3dff9eec7e40e57c3479e26cf1899aeb77202bdda3742b6c23b5a4c44b35a65e8a3f301e422360999f8d3ce7163524ce65ede375ee1bf6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f6e40e9f7e581fc1e8ffd83bc90ca2c9a6bcd417d9aa4208f087bf78cc045cdfb844f7f76cbf603108f86bbd65805dae03d2a25c5647c4f53a69dc83bb8634a0474e6a1a1ee31f7bfb57c0db5cbe603821f52e838ab92097087b7ca20a6a6a1ba60140dd178b3626a519cdcb34cf19680352461692bdc21c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha9ed4650654b20c5a067977fd83112fc1f6f0b656313060a2ab226bc839766010c32bc61bcb5759e005c397420298ee962efa5f6848d75449337ec36331b3a74215d187eb98c96d81057d4e70469eb3811e5a95538a3f64e67ae87b2f7c93ae3059819dda08da8729c157059e037a8ac74c99bb93b60791b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hff8b02c487b6874dd3d6f23db7a6922e9c67e742ac18436cd1b53fdb7d48a5c0dafc1f16d77d2cd8a6447af831035d8ecec35f97d3cc42f83ffd3356a59524a1d87749102428ea7042d3a6421ca61e74ca2f2a8f21081702c0e1fd24903334c427d3645e16054d47caa10835d860cac6e8e50f7868d1efb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f99d498ce5409a83bae1e2d1d5cba58a0665d793579a1a86b7c49b47438bf0f3ec28cf03ec20a404502ecaa72ec74e715a0a75611bbd713ebac504148e616f4c5932831a09912f25c11649480f55fe5f9f8febc55c8b93efe20c1eb5c8ef22b87a690794a1541af60a359291895b53c7de2f33f0a330d55e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b0d81ddf35fd2459ff4cf37df308af66d2eb544ef7f895e884421012ac66934a50d1df270aa91be4bcb8d461de28ac291ba418f0001606763ed448263f205ae2c0a83901bc292a23b63c4dc20c4fbe7e826ab79e31d8e06f8c5ce963f9b3b410e2f88249630842417550e041313b7ce63ccc69b0499dc50;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16373d6e9f55578e4937132062d035c04b19e8453d78463a15ac3d47405e34c3d1fa780215efcfba4bf6b845bdd3fe8516f9baa217a2f0efe630260cb7da76a7bf45c9dee5d1e751c180bb92c5a2e38e9179ed0ecace66a97594d3d932210e885087563a0d21db63fa405021f2ffa769dba76d43e45ad6c92;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e8baaa9f4d8793ce690a5804a904e042669088ef25b620db5afb05e24ae3107a766d585be2ea871f1f89eecac1f74de9418f4bb20f4b6931d145680717736f57e1338afec7183efcde6998a849463dce83557377fecc36caeddba083aacdb28a9d7caf037db51dfce8246bc6b825b4668ee63fd6e7c18d0c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12370a8f91fbdbc7577c3cde47f7166ba88289b2da42d173c773e959b9c0c10eb9c71c193a58c35c66bc705fa96d45429e0ab9632377bd5f601ba8d3276ac95b9e2b3c61401c231b4bb3709112bdc7e78de68a8480ca921deb12a2b2d8ed0072161de1bb56add833083fc2967671f0815226b12906fa1bae8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f22f014147cef1d4412c6a4ab85d3657ad1ee96dfb0d6fae2142b9d2358e0fb7b8f0cf9f8f1251d2a54769db2baa59d1441bf6d93827fe2810d11f91aac08158cbed87928d5e2a03ac101df01aeb27d230b7796e578e441dc2a7d91f012fe00a5c0eeb4b901ec9883395237b30b60846f426159967fe27c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c1e2f761d526e175cb79b0619bd992f78391a3f5be9e019ef7fe18a1a6ef26f079c895955902dc58c73c907f65aab8318e94ee36e2cbfa30e33a313fbce76aad1c604293d1dba8d92350630b10c0b444e7d22ad97569c322de184fe916b679271093695c6fee9d75790f09e310cabe46dcc441c1bcd47f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1696d835186c09497adceb8d10ca8e332018aa81f77745cb15d52b10ebe4e029cd52eeacd485c2962397b21da7c9c56880a9a37c1bfd1f027ee5f96f765f0fc84a13ebf2467b36d62cf8da4f23fc1b86ec08740572b0598f6c2eaf539427ad11b4fe523bbae6cd82c2b2c5d476dfc8ba5029d1a0538a47cf6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ab6da76453c28ccd33e7cd4506c8307e0c5f95b458b3c646e867e4efc4c3080c93f909f5598626148049f2f146cd0c946ceb9fdc1c9413349fc48b0df5aa05ae88071010a7d67cc6c364acf1142bdb9456e78bbf102486590618f7ee789f15e79fadc40492970e451c9607fabbc47d03f79d63eb276d8cc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c0753735edcbcb321b6b7efe0bc9be06acd36cc42898f2c25ecfd8a2ab63343a05f5d4535629d5ed622e0fbbb6ed0c110c0f308883ca6a9bfc07c4ee2751a7996002f2f20917e32994061c92d638ef3020d3e668e0ab4a38e88cf9216f3316121abfe7eae23b7c8ebd7bb8ac0184756669b79e6bd8a15ce1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9037b8d579b8055846ec7bb3f0c8d28db5a056a28452a7f9b9c9af52068b423dc82ffaf337254666b2c35463d1ca5cbd4e385275cec3e1bd68ff909eb6d80920ae6676bd591d79d508a9c35038fc00a1eabeda049451b1581ba8d7910b8a3595fb3c8e0e56550c7d0bf25de1d7b970fb371507b3f0791d27;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f1dc00854ba6714eb1a94cd7f54bc48d2d62e7d07a5a5851d3c35317499ee21f5de7e819e848f3b918efaef4a2aef73d9a7c7d3a79643f868dcb18a304a1e0d09e2701438d5a5d81df8df68bae5e15092b7abec3bd11e6db1cb153c405227e651d0626eca1703f8c5deb1e00ae342aaf52ef124008696906;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h89abb2ed4787330922a308a92eb3fd58337a39ec5bdda83e5ea0a8db1be74dc730837a3d94ab1d3c9ae0281d9594de127b1099e13cc3125fb0fe72e84776b1aad421d37075c2adfea3a88f16d10a40a3101bc7781ffc74c99738de42275edb11ff932117d18250e9df5c04345c7dc8910aee200d05758307;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc161835cee2c0d06c8c37a1b65c220a60ce780a3ec35d975eb004b72a63337f3fb5b2cc214fc330e0e0de209fc3a96e85a28c494cdca85876645012a4a9dd52cb64f5266d6a90db9512e02e660c2bc3f83510dddd25d93c4cb5fafd16c6ad3d1d0e91098d37e055daa022429e9bc538d4300fbac7888358d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd8310b803b35c960be05cb3ca7e23ab91a0a1daa7137788a6c7b3d7dca32870ad1fa902ddb2ae32f1821b809d80886d66fcaa746d3f4adbdde76aa1d08af255dfbe5bc64a0401ba49507fc21d51948a7622d25edd87cf399732fea60a368937a92a953108b742e2341f6f0e2af1b2991842ff63de76c4e58;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a121bb2fda13e82b6abda881adcd7b9053eec2337c7d32e567d4cf146bf29476d90bb9e7f78a7c3490975f13999974440d19d215ed6914fe75eef282c82e7dbc906e4b7380f0c051a4a2d598510962dccd32a11face8336646984245dbb040838fefa1d80ee8894fb9d70f8eb4e5420f96fb95bd2b706082;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he47416f07a935c1680cdc7cc86b744758da283de366c39abfcff96ae129080f0d1f00fa915b81a6e75fe59ce1ce7cb82a4b18e9d020979316131a451940db9fff6288e2804f9dceeb3ddceefcfa3802622c37493e3dbacf718d2c70c266a9086a542700ade758496885dcac461be03a50b64804034cf0eaf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5466be7ab8a5fcdedb1bd220ce4588477eff407e1a0ca8d77b32a060e4e905ad3cbe77c830881801fc6748044e89617e41a948492e9a1a08c0a86ba486498c0e2342a173c9515ae6ec60d547b5b475c82bfd77583257856134b970e48b31e906c38bf8ad26e612391053f10d02a7065f201db780de436a21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h198fd5d66b56dbd5c5489a077e58f0fff3779b94cc7c92856f2e757ff7e7937229309751c0de6dd07ccd6721e623e7f43b74a6488138b6fe1c4edb9cfbf40a2d03af25cb38dd677a9a1b191486cff412d689faeced7652a8b7903c5f82cc4e7cd58739ea316a7b7770a602d507c7950d26aa2fadaaafa997;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19ffbdc7ef7d5a8d79ecc903b44f310ca8e27e27e879f81696857f76da1c373c44095f7d07c506fa628aebd13019854cce66ab08f8e7854625f478fd55727f75737f11eadf5012f06e500056730e5a80fa2a0265527962e4310f5f4d2a5414061adbfcd532c49cce6ab68af197536c1f7c6cb298e7308b151;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h337ad8773b08ba346c4d08d3c766ac8d92a7fb3c3580eef0cc91d273b517c19d9d360ce46cf89ba7441d859ea1a1e4627d1bf186e9511dbf05d71499e942a41db64a1f38be943f734bf63258417490476eac838d638be69a3bb1bed0c828c1734cb07df9623948b16edbb127abb407722f6198d4dbc8aaf9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h130bfdd12528749d0e63776f220b7a1e7ac3d93bcf5b5ae0d43d919c37369b030ed830eb9b9ca9f41f2c9639a483db2522a53429ae7b8218d00d52615e694f63cd6e9c4c00dcfe8c160ea4a7b9348e0d3c34fbee1244cfbe64029bd154b282e113e1ffc4027fb1ccbb6277353628dbbe2903bbbd71e3048bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h108fda8e496262603ccd2cd15f672c3f37fd8111621a9863df535c2c93d02d6ae396a305ff6c6110155b78864130afbae7e2dbf6d756b57dba4be582a55b96fb21d0b6cfca75ad15fd2eb6dfffd29cd2a4aa0ee9125529029194f6045e64c2c425da29bd2aee41a7eefddb675eab586f693532b22ab622af6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e19d0599fc8747bdecfece1a1f2e98ca0374b455650942c70db42f07c38d954888355887f6ef897db8ca18fe747004fff084897af89af18dde90cf08daaf0fe2a2b0c0959a00e9295f07c81abca05826b2117d1b8be57ea3100ec34a50e90eed33166b4e7c3dd2b4fdeea378ef6602adf1dfae40cb79a916;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b8a02a5b389d0bea9e531b674b962b0786426f5f4ea6b4fbca107254fe835a9eb349b480489af05afc5e53fb9f375a6e5826577dac4f9a26889e08b4482880cd6cd97522ff0e623c4e825264f12437cac088bc9937e4aa77b4fd2641571ccc193daf5d37f83398a0f306902890470beceeae1a0e6e0be27;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13521a8cfa3a6f67190cc16f54a24b8261b16e4caef1acf85e0d4813dbdb9fe0c40a361752ddad393d55ea849ca2320954c6e2328dd886e68a34f3e1e91c87c1dd35df343a9218ed01c627a6345bb4c7cfdedf5e6c96a0e60160f6aeb533f9cc7f59578ad706be213cfcdd93bf4f6cb3c2c6033aa66fcc406;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5a967c131f7332f513d4fa118585382524937a264446881f915a16fb271ad4aa5aa8af8f348a515a16306c92a109c273e15bcbc752af747806314195317902f49da519291ecece926a5df2e2b663ec35b733bf85581f64860cde5a2a2628425af4b326aa70d1e9d048069cddd957eb69e64b32c379340ff8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4d8c5a5810614271c56c937b8e0803f6d73b18b9178e627ba8e20de9cacd7764446b09e596e8ddcfa7047f261655c7d312c29fc611d110bf68ff86b11e1c7c329d86e25f553a6bf29d948b181ebf123261ae61495ef254b69e557c25ca42d5c5c45735616c5ded36764eb36b6d24c7ec1176703a3fe3c8e1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3a20d8190eb954b4c2165026e6b44b959f5b9fb5378653df7f94f0e49dc268f40aa256c12f4ec2be0fc4cf0b3428bc4431724f26f3ae50130f324165378f920d771d4f1cd5a49ba548a6d55983b4413369c01927d9ac340cf3c5d70daf690254b733b3cca4ad2cc56a658fe0d627f05392c7725cae03d3a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70cf5b904320a131460415ffa0b86b7e557ed417e16f4bfa0dc1b3d79d193b578b5b78da1606099993fa5c72569e461a6ec15ab0bb687c42f467687ec29035e4c1a5ad78db56a3ba2e645a918e58ba32c9e282b0ae3c700440bdbea50a092b337dc79791df7fe8b94718cb2d849309122db6d5067c3b4a30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h966b67b85861ac342430a7ec72eb91d4a8711c6bfee23b25eceee9c89f550083e619914dd9239b09bb0794606c178117f11fc8ce8652f6e9f10b8229f454aea10fee381d2e1197012615735277c340ee44a31eb7a7c218526830077f7a322bf06ccea7e1bbf2e72fe6451ef1511872b49d758532bad5ae9c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1727bc077e2596efb7d33cffc170c6bc8771e731cc1f5fb9121bca127802852f170d87d195faa2bc9756c99628fc93620ae7673d23a9656607b79da2e678adfe408949a8e77dafe59541a7a1e7058fa675a3779f4acf130f31d5e44f744c941ab9327e925dd9e18a0d8af14250a123a4d0b2125ac24699421;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f6eec95da56749294fb4b2e38c99888828a96342d0b07510ee3b786f1aa61077a2d0deca9892b941fc50b7040a83096c08eec694c37bcaf21eae9b0bf2faa03e8d7f35d6ac0fb984c778d094fae966064d97c27334309991868b4af348e92e85d797f5cab97623add5b56060ba9c3daa89827a2c524848fc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e1e5673ed2b769a1b2db415fa5402e87b1101eb85e47e17f5e1c7a8fae1f79c7f98f6cf9c45cd1868ef19951394d4b38cbf61cd15d5cf76d1bbc49cecaa3da951cd81e39dbb66e43456d4a31c5d46c13559ad4d5754594a390f38739b6a79caf1944c33abecccdd3b102eea31bb720da0817bef944d23ec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17fc92c8d43ea0f66e8ed511acd12f8bdd1a73a331b1f8dd402984e72f351ab5e7c061cd1c8205bcfa4a29ffb445b6fdb5000c9cde2998b101dd598a22d9a558109d91a56fef9b942e50e89b1fadf84635e66cba529ffa6e17747cd088f19d0d5f1ca34cad399bfa01ebbb39a184caef0ee6b42ae58f718e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2732851e6350f407fbbe6ba78305bd5be8d01c3b25e5faadb0d053eabc0268e95fb8a1ae40f69e8d7694d675c27a7a543b0f37ff328e0653427d04ea500827f68e907d75e4ac2dcfea9ea4c3bb1e2f7bea36c573dbc9989350082ddcdba4ea67bdff018f1c5515c331554d5283add538f9848a343244ef16;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18e70f11b6a08bc91ce2c025beb639dd27cd34171cbd62221403e17a55eb19a6e4bd3abb395eee61cc8948a4649a32a231ab2767f220e20d405317bc22c9e22909cd89622eb8cfc05262bd1737e94fc7efe81c5e84142d40bf7ff8c955a4328fd347b1e4f17ec4da2dc8c842092323afe3e4f349a562234d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13924f54ce1899025fa80bd298272bc6332888198726b50442f381963dc0be9a206a764c03686956f9fc6596516015f4c663b86580e4a1488e95a34bf210e39717206b19bb8394987b17eafdc8f80e0554c613f83d08b8a25f313f91db680dd3a8c6418ec531072c938a73c1bd49dbf69338cd547e5018b9b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18ceae0417ecb84922198f17296a792c5d447008eacacd9ca7bc3d195d5307bbf2af4ded19338abd3d4fee44fba05516c3e0f8dfa4bf54b26e09003eb982c1080841b65a9bb2dee4ca690e8dce7fbc0e36ab19bb724f07df1ac67d0fa4864003b0f4d737c302844d04a24aaf8895250c39df49be6866f860f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h32bf629e3ac230d28068090f5c4bfdc810d98b00d5d069c9fcdde52cdc73bb6ac1e8e8c831541620c7688fa1199b54be9b9b5c0648d436b9e5bfb36fd12d0f6c050e55a58fd8a264370bffd271fa1786740e39bc5f29d1a1dfc8d4a3b4719dfe73a7763d8a72ea3aa10a9152f634347a0051a9c6aa9a2dca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10fdc9c16baa53388db08a27fd484472f7ae1480cde942d0d0af4d8331ac8eb28f628f7d88676c55dc91149ac2a9d633be0a4fc4f0d455e58eb457506fc9c266ab7b186b870316e7d8210486eb0f0f7f28f77d0971026eeff050adc7622c2f119b8b71b7b4144a5c32a767a30e26d6b3b410347105c3fad0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6e89b42eee0a6f853a047c51bba9474c3999198af903307a37c601532844f4c020590d25f84ad07ca5d3f480c777cd4ea324e8ea5b26ba47ff036994bcae53fc599f91301c48b827cfebb41c4adaf517d958717e6e53a77147da4ad5ef128ecde9f0c80a4b92e161aad66721bccecef89a4cf8a05816cbe6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h94a7f0c9fba7e836d0de98b5ea80dde39e2232ce4af67e7efe1d98acf47a27625daccb87080eec9d32a8ccb6db3ad92ed5febd5e25e3a46b62a1fdac7d11c05eced34976fbe2288e488947225aa345450331fe6f10f925493afa5058958e3def31ad733b286b18b6acf8f4772443240599ec2f78c714361a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1adca7d75372c6437e38bd4280be630930638744020b4812ab7b3f62303e4e9598cefe8ccb7e8dd259b34c67351a8b24433bd1a5e9abfac66c5896006b7b2f034c58d1bfa5c5861b0aa211ebb7d81a3c929220e49446c44310997cd55c7387a452612b360cae56b5acd8f7f1490e6b15163227727312d6900;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11465d389777e02c9075d419d61704b96a808a0f981da9b385c657e4eb821fca9be03285386c30bfd1bed72f12a0a479e0ff881b2d13a9a08356e59851be0a376673fd79dac29b041bd9156ed75108f3caa4130095e741068a70452e9e6a228a50e430dcca99e12960a368a2871558a819c5e4bbe0267e05c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1330acfff6e7183ee2aa41f23316b10824257f6d0b7d088cb2a56438d848389a3e4a7993973fff66c9bc56136e31feb4ea194a2fb2cf7f652bcbe8c865062d0eb3b1b8d9bc116a755eb30a28d6cc7c3211d15bf3c388e91b1973365105d939bb639f417be2842adb8e033fd9818f8f2dc0d1e80e804d121f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4432bdc1675786d24343220a46fb38085b3cc20d3a37c8c1d0e6c2681e263e7eb9882394fb256e55d252bc305995a8a5c24c21b0839b13a2b569c1c4881e852030ce0a28246d28423a1ca154608e94f7abdca26b266a0746505967dc314050c1b3d8cde537b3fbc77bae3143c35051269be8fac8e9f667c5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d8e25093b91c4e5ace3bce2e293c0795843116bcbddaff9c242ae2a97dc556bae30c7a8c5f2b74f696e91a2f2a82f6264fc934795053a014bd4eb8e2934e9146e7f0219f79461895e9283e73b091b51e787f0776d28efdaea5b5d13202ce7680135948bb974ad67e7815c9f46f8287189a5219870c8d0d06;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h190c29731d4154c7fecf86b299e0aad5dac0ebd37bcfeed5a0115573bf58384c5ef0a9397354b0b90635486907c635506f0d4a71ceb42b61fd53e7c2f8f0dae68aa524a793cb808cb8694b089a738fa293bcfa56774ba8874f5b12cbc074938c9f53adbe3a1e738ed6d32ba22508733d964de678916f16116;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dbb9658ddc146e97dd4b9ed2ab60cb334f606bcadf4f66b0033166a20c4322b496c6f5d566a044c87146976e7664924211feb0f02a6a40f29e4c1a192d7351fc8ce74a18f81ad57bc17dbd4c8f1106e8471cc01eaf197d3c5b13914846e99c31dc92e89c31e1f3a3b916cfbd13d11fd651b0dbb0f2ccbef0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c27ee2a6035d5542de93ce56e1ac0fefb1139f357821147287c0014b43ba98a49602c5c8b7a8c695fb67a3942b4ee57b1c27eddc6b09e10371999fd95b9cfa451496733a4801e4fc6c568ee21bf9cf99447e5c18158a0d4140eb70d83887bf000c50db607efb97e40900f780ce3e5fc475a220d6c0cbca2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hce7cf7c09371f9b84857235726b4de7290e6967cbe82a9fecb5c1aa0bb61351e583abea52aced563d084983e56495d1acf44a8874e8df1e440b646b4ca30823708a5e5429cece2972cc180f3aeaf1ddf90fd82ef02f766aa08260fa04aace25897b2ed3122e4eb91caa150f034c6b46e6b9c0d95be21f604;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fe7600f2b000492baf2d7a22b58b75bc2d28839dbcf3092ff0ff4a5f331515f7ff286db1b61ce2071d5599a155b046ef714e2ad3f180b6c07f03820da2e942748227dc55f89f9152baba67a87d3677abd7d58537286bd6851f1d46f69f010c50551fb421297a5b30eaa666929103ed2ed68ec0682eb4145e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbfa7c98ad7ea67d55d5b736850dbf66540aec396f7464585051842f7a9791cd4f23d9145f8dc6a71551682cddf3171d342b26d41e0a45bdcaaf983fcfd281e9319d55888844e175ebb3e137f45e67d5716ea5071681f0e8c32e5f3ce8590764ce128a2c17058b807d4a2d012c059f69d86062e555c43bb6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb2f966b64952dff9c56f2298ba15cd4b7e6c4bcf9a49f4673419493c47df3614df07245035c4e28f7f9faf48b0b60100a84a71cf1a7e694a655aaae38ca111d6f6fb62d87b952082ac7f6988e4565837372ca7fc4ce6b3140e792acbb45f87aeecf02b1e791b177daacbbbc0e165d06f262d55f42d3c5d4b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h51d8917b8c04fd1f8c382763e4dffadf26d5531710ed819c07754cef4133b16c4c5c686f07e0ea897101a12b447a22dddc06dcc24e77d6216e24649a8cdb5792e1473a0e161bc652f6e8ce3d7727ef57bfcefe9cba7a44b1d1d0bfcad1b0e9fb10c9d66e18809d8296b6cdbdef68bee36e284d75a37532b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f589d08967e1324878df231bed5445eb4e10e87bff68d0367fb4dffdff04c44ece8d7423366ac980df239cd8ce75b073318efe7e7c63eee0f1692113c6c1076399a28bba6714ee4be1588d50f5058621edd799ab366f89e9a41690455ddeaaf5e79086898054cf24a8e51e6ebfb8c1cbe8e41c5e3fd91d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h241e1f195eb0c3f9093b16387437eb6fe7a5761bd5e263227b4a6770d27abd9ce28d543a51c6f45f9ef18c2b6660538505babbf1512b7196fb300171b7c709271721cdf63417d1487f07e4e31ee02e20e38acde45662f92c78ccd1ef10b9945bcaee5b4d6902d4deaecac11ddd393850388d5ec58a989ba9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18b65e38349330acb91ba85982018600cda9d26e316a81507f226a40688cb2c350b517eec5ea50b30ba8c07b387cb9c5b95b57035bcfdcad89418fee6227653c372545a654e22ce86a99f9effcb8a980d555299af05b94e9e1ce732c9aa949d6f7891c2d265f8bbcd2e840b3dd2aaa3b83857ea2d8368c94e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c45e56134e0e8321266483cdb06e1ccee19313bca04d93148d1f88776d4c1554379d5e73c2f50a2722c2aa440323c187c7eb110056fdac499c121d62283ee576e06b9d7e17b9036c4678b47222661cc3924ce2250ffc4ec786169a07c79745c321ffd82c03386f74ec1b4d2083a303251bd03eb53005a20;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ef7cbeaa0b562577d1fe2f933e01e4fd531deed40a5db2ec548103b01bf42df4db1a5c12ac57cda73cd26d91aad393d759ecbe5627ab0cc9329c16fd6b17ae462b410fa4f2a877ac97686da8133b9db409f302b495113c920a4947e57ed3bbdfe83747e5115055c141a5031224193fbffb3ed718ea67d98;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47311fc9e115e4b538883bdcbf05a0c5f74c6bcddb0a42af27af6ca34b1ac02608cd5f9aec390fea14a06a4073711cc5d8fe5632d001b40af2fc0e6ca5f94ae008ead89fb465517d6049310da1e99a379a451dbafe0362acb0aad1c2830d1581e477d1c62ba7af4fdfe7f152cc0dd34b7a77793e78d1e23a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h229c6f4652f5682757c0cc41b341e993fb6a5bfc3aa5995e4d312f8c3f3506451af5ea07742873d0aed02257da4a84966be0a51f4d137405575ac959cf784665ce95fa0ea12e86b62b795ace5a158475d51ec0feaf2cb516de01eb0b3f061cf7c1a5695806bb816fa1d519ec2a1cf6e3ebff72aa0fe17b05;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79903161e3a86f0e0db1a2473a42d63e7be031a2211a9ca99b92d0eb31524d6c21056100c58dde02a47effe807d2d31a5acda0015dbc916661cfd6f49b938f261c2dfde1be063ca39779d956824f8940a71565921c0aae32435ef06df92e5fbdb70efa608c68582ddc9032c5dbe8d477a0c0d52181de0c71;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5f04e7d0e8ec5d497d0aa88cc3f460de55920883ca42456bb3453ad447568e277afd86348bc03c400aca2eab0483d1213d302fa2cdf96468f8674177d66d86069ad105119db4c916977748fdbb44cae02d880f3d700c92174100f3bb46205dfd12c71c6cb2d9468081ecb6b0463571e9d00dff84a444dfd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0a7bead8e0f172a90011935d34e5144babb5ea6e9d471e7932162a7a50f69b2db9d219c371c453cf012f2a06d13979f6f55b6b861d1c98518fdc9d03ddda226118d83f9c0cdde780b75ee210d47868f4c4b357099dd7f141efa2915dd1abb96f6b58bc7c6a9eeaf6270eae761c70f30edba428a9143ceff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdefb3d0c73a8f3ae5bd71854626e852d8d8eb2585150f57aa679c759414686d765ca6b57cf5e39d572e8ce3c5bfac9376d6bf71fa8b4f6f5a49dce415dcba712c900b32c1acdceef0aed63294941ba45c73f34bf0331fdfc9daf4840926d7c64336030b32b58d7c8f79397d84ed5c0b1c344c60f3b6569b5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h171c8f0a500c7c9da250237e788dbce3366e9ddc059d41eae3c0c9db9bd33cfba53998df659f3df003863a7ba1a6c5eb43d149f5e9b6f3921b6b84500b8301477437e1207b2c8abda74bc95ceef0c631baf64ce8dec2ca1cd02070e3aea06b773de6b588b4e1978d1b20eddc62bc9db62f076435b7581821d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc057a172fbfcb4c1a57cc6fe0c02b9a6ed0fce785634bc5c7ef85e9a87c6c2dc691c7b724d951e00851cb5e3670ce645b5f819469d31198a25a7f7e391a285437938319b624b7f295de745d5d9b72dfb5942c3b47fbc2ee90e0d59077678dabd7e0aaf8c53188d48d482faf4d11c5896bbd7f38dd6621408;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2eaa1d1eeefe8a8856a40a24abc0154bb16ee00b4c16213057249aec38e18b5e4de9d90b5dbea1217e918502706061b11d0b186b00cadd5c097199026bb389e6fc0200fea1ba83c6e81cbfa699a9be36ea5b392dd3d8ac4d00062e745f5d4c700c0f9726574f1e66bd61d51f4633606921d5bb34b2d76151;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106b4f93a3a5b076288fe5095b51c5bf48a91d27189365382f7159e155a868b19e9797c451cf78009f2cb162bf7407aaf0b05587c6e81080741eb0e7419ddce52b9c853d630a75d9df2d3bfa92084a3e731657c1c89a038de384978745fb7564f670a6b13970b1170c4e347ed07af4794259e94edce6019b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14426951758e0fc34b5270896f70d7c79e550c6e4bb460f45bdc728f4df0c934e1a0e5245d4bf5b9e62ea2a3996dde7ff83bcb04f1fa747964787f16299e438b1b529cbcedbfb0cfe3f481b6a0c759bb1b8e246604e5a85449d6d4dff62afa7e1f3070517e6245230e01eb66294585dc5a0a61f27d7af9d68;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bbaa6469ecd0b1e336d539a5e22bc2a01eda1df183f961d915c28abb92008dec1429a848e87368034728037e291a45b586e20caeb9486cb39af087f7b1c2fc18e6763b4446f0c2e10364478a5654e1edb4d91f4adf4f234f5875af5e037c6abedd7a9ca6786a38fd77c1072ebe389e4c0336fc551e3a33c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h73f46ed4f44cffdb6da5234505277d6fd44e84058ce9bf74e1fe787ae2ab73d2200796d238658ca3b785200b4e6a38bda4a702405896b90f429f615e2cdb068d3e85b62b7c1e4453c08b09315d34a9cad1adce501b414b629423b7841fa0d0866e00423c6d80b272ace34914280ae4302c630700a008e848;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h60a15303f8b09cfd3cf422dde407fe5efc5842a593320b3bfa0223882b938ac14cee87d4c2e488a1682267e31125df1c1f99b3d9c69eb22fde154bbf24cc5812311286722971eb31b6ebd922157ef3135b4bec266bf1baa077121392ce95537a8543d94bc191cb953b7e1974632587d6f37224f623467470;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h167d478bdd1b90de0032f4654bee88d61d21d503d2ab0f2f06b9b8a599d2ea7b691ec948f2e8b8248d1829cbd4ed75d8736fcb3543149d70aa926b4ad94c06a8f61d37e779ebf7f6015a300b9ad7885294e6a9454e35920eceace5d5d8b426ea6852ab7ddb2cdf23ebb2da083245c013d810392ef619b13b3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h141ba0f24496220fdbe718f761e3615c3930fc61395bf1bfd741d5ec7f86d7f1f1f25caf731d66d0137d3bc7a9282926e11d0c0b49ab0a156905029dc4eb9d0819ffd2263e9f8bffeb235fc23c226bc01b437073c16fa417845352b61737630c7caafc16aa6bf923cee81bb0a6e55ac0e798f1caca482af9e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h33ed8b113769faa9a494f565118934134f588ed30704076d6f24c1ca7a2fbec620586147b7c98c708b0dbf86fd401c3e2d050acb03923cefd05570bd1d5baa07c4ee2b717c70f161237fa38c248484166be0af3c7d5b0ef98c923a7daa8efa703b500d38d4c0d47a40d0facc2203724cf370016641650931;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cbe035670142ce37ea3169e707138ca064e5c3fc5eb9214ead265f49982f3fd00eba85f0998de2aed5de7938f833e1160762cce1a04961f4d986a4ea91a0b58ecaadae883d9e2b66887cf07be31ca12b6106485e1b9b8e786ecf37a08ea84bb7af741762ed2e030ac548e232bdde1e965963c7bdaed334e9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ce565134cc4563106941a1747c1367489d466a04eff1a2a09f4d2111e4df3bc5f6b2949f18a87fdb88f172024ae809a7e6f3cec1de719a86cac5bfcd5f44ce45793c83970ea4783a89d2d1c5a8505886495a52c38caec8cb522266050491133c53fff6c1fb33c8c5b1c84351f0ebf04487c52ae26592c62;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1428aa3275015893f765cc9fa2e753cf3309b195c7ac4805fdfb38bcea08cc4bb06d70185624f2d9faee927bf01cd59621b7b1d0f5e750eeb107c39237e742d7716299d4c644d5c6b97ca5bde8af8fad4cac4d44f1bf06135c7fac81b511e8e735908385148fd18a67e475533b2aab37796d0046ec8d1a2ee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c95eabf0981d926c2ac44130e73a60e8c147acaedff38e3a3c2f53ab0422a7372787e7139270fcafce960bb90f38bb926142fc3374090f84b3f749bb1b83bce54b38b8c108b2f6844aa5fb5716f417ff9216fab0b6d8193d7bcfc5bcb8a40e909817b4549d7377485fb3dfbd5043ebcc7586288aed277be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f7d154565f37de7580d5c536fee758bf2715e97200cf65752da92b80121cafd3e7856daa2af4ed567b465f788fc4e06c37823edcd11b4fe045edfa7d167abf7bf0d9952c0bd018a9fd3479ec2b362a2b6d00f23fed115036ca4b6dea66a0192a09eeef503f0f47c27822316b3227a5c2f847b6194e782b9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ca3e5c50ae90baf74164d42f6d0b0376e5202881cc2e0f010a47778a40fdab32f7bbead87f312a5237f2215e5e0394f5f3790f26f5061b30e307bb31c366c209b009ed6ac7127fc454892be82fc6a624282f5e666e51e732c259714728a435cc675aa07cf9049c5e77c31be321f14baf71dac55ff166bd99;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4f48536b7335a7e785295796eee14f3d02e283d24b9c2dc529ce6f7d66a37c33ae9679fe4ef7bc5e1fa68b40249b7096b3eb4cadee13816a420b438404a8c6d83fb9c276b712547d1f2e5d7e3226c11fe63a5903120eb5d5db2f3caf963599e5c0967eca31a6b204b8a86d0cffdd3175b0c15882a62cfdce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102abf5e5595cef70af7a29079be7c7cfeb1675a2e1e100615174031fcbfd9dd3ae2a10ef220bf6daa071345cc5007416cd8855c88217d9c7e181d90c2365542c5e0b2dda8290970b2a5c53bcc261ab13992079eb8a738001b1f62f88f9d7ba4bea1bbfa0c71b5c1d596dddbd8ba882f1baaae5dfa07dd32;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11109415a345a5d98b8a36b7b876e883ccdb0cdacf6f2cf42c62f08e1223e95ba8c8d310340a80e3f8c81c588f46e3687add32d258b979a6a8372092b14dc2e2083e04de87c2e20544c6a568c74e1062023e1c4435c64deb3f01114ac3d3a174c6be951e82e5e5c41eb4207d936c9a60b0c85a4286938181;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137ac01a4fe9230b2974141c7a16b179b22e5af835d67c0423f8d5189329b6e0434ed84620e16d2f970275cd80d578a91b4b37947b2ebbf8a28f06cf24a3cace80e569ae3fc30a290f1fdaec229d14995d81b11a7d4f9049a11ff154deb7a8beefe97e9feae3c3cf3c80be7fa1c843cc15dbce446481acd63;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b0b688c5fb546e20087394c678e7a5d24f4d685b6fd7c119decccceef9c195fa8275edcf2ad6fe2361bb61c2e23168f07aadaeb0fd9211a865ab1874d244005637bded118bc98120ccaee2a2b775ba26137a805c66f9fc0cf2eb46761c3cbd6a16c8f6d47916b9cc48ce9425bf659579e2988d4651759b54;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h65479104c0bf6964f093df238c1046731fb5ffac6ce00aab331d98222885be170356dd701a3ffe9940ad6a358e5509dabd08268d9beee1762fd94f53d7384c3650ab9fa8a5cc8ea596c0abb1d7d053380b70c4ca9e144fe48e63b6bcda11c47108cebc708dff3a7bba51bed5c1ffe1560dfd8a07c8c9cff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb71a9f402a6ef24204fc8070d5a257530ae3244881fea258281225b4befb2111f3dceb1e325a7bc1b284de92eed8133c689b0aee3343f0e482ba8ddfa8abb19f36ad11117538d874abec23ef403ef7cc205708a442be8ac66b6f2beed074538c69e20dc0ac0537a1f07a7e6f9589cad0c6ce46676087bd71;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3249dabe1b0e6bef7f11c2e6f008aae391e915f30a246b023d1aa50eff39b31c10582196333d8e130684084b673d6f669ccf55f37d68f4aa49ae9b3d9ad7d12df23e4b14c28c182bacdb857769f2dd2ae642b059e4c6ff8ed912f1c7333bdda474970ef9e4967cc85bc72050fac4d2d3e874f295f19c31b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc325f0fb0e7c64a864b5a26304455b3265909e70a6b4ea2d6697108ca5dfa3ca2d20d8dd381ae60ce31a3d97364d39c814be92e78662a1dfceb06548e278c7b7bab14fe539a0be126b0ab115c3380126acdfa5a9141521e54f36f5635894dd906687259b0caaf8283f95d0bfb0ba5df732ea1055715ebfb5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c94a32fcb4b4aadf8e4509d7dc06654ba6860c09b87b7da7c3248babb9562063efe0ef688cda6c9c15a7bfb26dea06dc0b734c8040e5e27c0b5de4ba0138afe5d16f338fa7b383678a7de8c980812f819515c59b7b593fb6a92c5230d6dc16aa883d7ab780871f70a15b0845b6ffa23e185ca7b14e559a56;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h265351aaf4d0818d7b0a2ada4f59a313e116ca538caa51859a67a932d9e62e339126a7ba16a1e60e3dcbbcb4dbee1bd4690d3a9adf18f1f3959047405143e25b95be7252920127a546f91a85196b6c6a38ea24888dc0d783ef89f3b591e9c85a2320635480d01005b0801d241db519d52d61b2ff91b3a352;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146eadd71f8c1843072c244eb6831c5334243fe68a131a1e7db8a4f3726c7bb8c86b1a487ec8ecab7e61541c840d81d328eb7c89d58a2f00be5a94835ca610091cf8b7ddc2c26959e7a568bb16b4df368660c90b81c3569fc2e0e0a743aba446991c27c710abcc5b88c8301e322d243267ade6399cb8909f3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c6b762db2306fbdbb7c08c2ca11237caca3e7dad2c08ff7d58c97a6f2d069fd6527974585f0dae326ddef845cca10bdd94079329abbf0e2331e8c36c5bb274a1fdaf02c235a66c2705e36f6824daac958c30a7244e8bd1be7e02212b87a6ce873b4032de65324ee5547ddc296da177d72b0079614ef6dda;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h129a9dacff0bd8e520bbdc5381e51e2bcdecfdb6fcb0db2d1f0387a3e01a3c95e3b072652adab382b7ad6381086c6fe9abcd52e05a2300804b246e0d3aaa72ffca3b6a3720cd20173d5df6eb129ab8e2a550a21b91edce16a35846a3be0f42fa7ad5cdc9bd5594076c10c098deafb8d5a3d9af9f88f866991;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9fb53a022c8ccee5974cb22ff64b7096f23ac1f96888310f1e5f2360c8bb9d2941050f37ca2d7f3769f236323629b5de567894662d3ce89d2d54ce6352a73087e4a356942413ece689d21cd01d347c75b472ea3007a183043da7f930462dbdecaca6336cfcb3d5cb6b585f1acc31db731fcc87a454f84cc3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1243f3e9d43701132262209f4b9c9f6a8bea9f787ca09fafbff11a844fe1eeb46ee14c576347eb7c970bbb103080c81d4225cb6310e5654ba70d777f44326979bc54178adbbf4bc5701693f787242c0dc6949ca2f86420994037f1c2ebf1803ae77351e68ad66cb0e32bf937d87dfca7ab7106541830a2eab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ff3cdca3e3a1fb04c002d15c94198678bdccdd21378a3df7833aa8c454e870aa4f58638b4f4c69f8a84cc5364080aa176d021e12655e3920e6632647a772290fa764ec684b10ffa482966150678665facea496d88a843c66c12be6552ba909842f4d35e2c728897810918e294f0a7d08d6e2e884ad37311;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e646a9c303a67b9c928b96189261b85e169ac82efacbb9259e20888dabf2e3110f421a53348e0280abc33b32a093de3756b10ef9f599fdacbcb9c46b5343d405170119a62646fdf8df6ace0115f45bf4aee047412885613e129c4426b3c4811fabacc9f30b1fdc270c0f9b59d1d578552db9cf0180aa9e3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h187430676eb6cfd5eb1792d44340eba40bbcad74f779a72ba70ba437a11a26669bfcd8ea1e5b22b4f5edc68ecebf311b1b4b0fc168d6ff768ff10abfc933d8fdb8830177267ce91953ec058e2f0ad2e1da9b31cf244c61798490fce26a3b245699342240151566978717887a5f7eedc70485c0fcb072e1ac6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13fb06ec1710e2856312b1112f8207e9aabf8e1c52b58c9db94f8a466b087debcff9464d1330db9fbda256d30a3cdcfa9bdeac521a35b9b57cea65b7c6692468e816f44c70e8646f5cb167aa4f53dd9d2c89681b34b834284c3ed5ca3bfe27528621131aff2ebee0da653c33c49d2eeb1cac612696eb32316;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hea27f5ce7f9fd6bd9654e0eadb929cc15c0e7c1a73d833b440d158609cbbd6217b3afd9fc58a2992fc0ea7728ea31e7ccc461462ea93b1ff5ac6e758d4ffbb845d41fe5de353249988bf84e52fceca6ae6ed3ea2c23a3ecff283eafcfb692d365b539c3cdda516a9fe9e520eed01b714794f98210d0c82c7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd9b15c536de82236004ad5906b424293a74b1421fdf3785ac2131177b39dcf6580cc19e819b693ccc5ddcf8c8fbbcfb5bd959eea3f62aea3af71e255d2d3436703e07c0a507439927207f33a53101e015a09f95bfdc7aee798641a59da4bdc939b0b795ff12f5fec3ba8d4e629a6184ea7be78edf77e0a4b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h126f1fed2cd45aa53a8e1479d6c2e9d0f41cf0cbd120573c9e852500478bc2a589566bbd2a8b5a6f8f22bb6ce3456d3355399f519eac43911dc02bbca37c20ccc1e5c0ae89414600ff86e57c6a9ab43176ae0da53d3d4d5f1d851c8429c8dc32cd2aa304056518eb1eaa4fecde6bc8f6658726fbb8b0e09f9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h152882dbf4e894bd4b2e291b6ea86c8e210bebe9b51dffca57f11991298c9077a6db5beaaa5b382b915be2b4dc8323e92e4642ea2a7d519cab8f3901dfd07bd5cbc0a79408bf5f44d8d98c47e5e0eca6c44ed3cddb832c246871e4637bfc4c03c2714e20e951b602a1d13696b4acc2606b82f2d9dd505839;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1417a045f90592a20b3d010af96a3e23b49af9fde79a82bb7c0106d83020ef876e07b851fb737ee1a2500df10d8144b580f9034f8124c335f4cdb83058d8d4f2e623b4e7de48a8b4835a82d8be87c663a97f55f7a570667df94876d4192920b348acf6de7e4d19bbbbf81426bf76f79bee0a3f91823002299;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6050449b2eb02fd65f9b4273c195e53cdbfb4e32485db4559483d411d2be8c9c0e8f36beb49bdc618d113e380dbaa1180658496a443f53965a9359723ec65d7bbc1f960cc33bc85da7e201bafca5c995b1e80b34664e562c02826a40f380fe22a2e70360c734b68d855ba0c71ec6041098f6e5ed14a3e28c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f9ff8c4b51fe834501fd378c215a8e70861c128c6eb84dbaf6144c28cee6ef49f8fd390b443a9917e1fe05ebf8f1ad25da6c7127673da5963c3ea2f8720fc1eae3e57aa3aff7b1fbec57f06a7c5c1dc3d3de31812f7d3a38e18fa99bbb3f9edf94daca96a08025173cdac4ec3b0b45b4219c243dc65d4bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8649ed40160b0cf0aa0cc60a062fad000ab71819ec72a47df3c30f8c6563062ce43b000cf559177951ea2a8fd3ce059d999cbeb4581778ccfb65c06e492000d52f09c733f0ad282e7533dc4f78d0daaf937542e701a71c888e7efafe02858a6e7af045ab8c03db47da71e18fa5bed56802f46694eb574c88;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hddea379bdf04b8d52fec6fd20da2a3534f9646af4827f3051ae8491d68a70de5369895b5e6dd1242d0722fee48a41a9107e5a1041ae9903e47f789b495120f2501b81834b8015b7d869dc00513f814c1c6a758f163902da0f7d950a0b006c08a37e270c8b001625e303577c37a44d35ad28723180535a261;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2a2ea390038c973d56b2537507f6d689ea541affe1245d43d899898da19e9d716aecaa44dffe288eb1241bccac6abf36949f4cf7a41b74a14116ae225af5a225f1c4e4a8047afd34f678da5e2c9ecdde4778919f0d1979c7a47d141df47b5eb63e6005b2cb4c15378723ba93c1535799616509a68e7dee65;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fb873eb203ba63d57673a0ab6678e791591806b5815f843c4113d3f6946ebe8e65ad36952813c5d8d2c1d07247d894f4926935533cf38b48a779489fb458e1d87a0215faceac3914193ea1fc446712902aaaa0ff25cff10a9d3ffd35ac6ea31053caab1727fed6631cef1e3dce789b6800cc5d1f82dda7c6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156e44aebfc4df69114f30e0fd65ed3550a84e42d2dd92fafed58c55f399c299a56a169112117c820735f52755d112dae48a3dc09d91bc9133650d71ebb20c0499e0e50414da822bf57c11faa99f7e149df8dc01689f8774d28a768dd3a65eb3f9bf81bfe8663103730ca7bce1cddb575c7101b7c87fab9b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h90d4226fcd5968b43002dd915b791650535e5a47e80a6266bba3c8a4913df1ca1badaf962faaf83b05eb5162a64232ccea9781b222a67836b272a0dbfb68890be64d9ca96ed6091a36c3981475b03b47f9f0dac3572bd1914b3e455248e1b1950dbc210466620196d92960f89f1374f6d55f1cce3cda4d64;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5091de5645a9c5c67168bc61972672a81321608f62588724301a82c088ba6386099091a2377c8944011525d43ce3ce1fcaddedbd6c1460c04f3c19558f0071ee42b69c6d994502986fdfbd7c61d51975b30fa54b191b36c1013438ed5d30f3d8b555eefc2d683582c1dd1fcbbacf2c1e09d6b39018e54dbe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c2b1f8948528b2191641cce8fdb29de1547db282c54cba44a6117bf1ed6c4ebdb04f825edc6a24f5ffb99406f30a406cd611a0c06770d5bfada4c9e5e762ff9fa7ef7999c5978fbbbdff225b08c02e038375853c17e883d2f981a14efcebfbc102a95a03da9c63eb1bd784807fb4f4f5f2e9a7e93b157cd5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h269b3a4640e0b2ad0221a93da2a45531c20ae0390548ccb1080f59f67a77316f82b50488a6197c6814678d34b3cf8208a3424571e90f37913cef3a8a029ceb148605bda5e4b8279662f4703b2f91941fe3cc79306a22251c12dc9f9f810b243acde538ec3b1776379555fff41ea486a4999e2b91d90b7cd8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b8a844b8d8e29ec6c845b9eed570fc49aa96fe7b16b27171721374917ad9dc8e2c56bf890cb6ac50e9f6be79bd68736406a43c8f4b02730ca39ba6e85a784e211e0c2e5e2f0fbc147b121a04c43ac3bf06b9ead365b369e988a2241deb8ced2e56611115adf89ade89d238d2f1cd04461cff3afde89e697a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3cf8e78cfe2db1949882f4e07f210714fba67d2dc7bd19b23935f4e7abaf71fae3efb7baca834ccc751a625550d67c92da53e9af0e037bf487f73ed6b06f202202bd10f6b35bd4d18a0a3e58eab2f087d96b361158dea6d958c9ae2bbe905fa5f50890a41b46954ebd0f87ce4d1849ffe89078634d27e12d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8ca601a31f17a58c70084f1369da00d69a043785950febf58852d6797abbd7f003220f48b5ca866db613d133c783d183d94bbad62bbf6fb93229f894a1a70456d6947c78adf93ca367258c32f01a69e294069e6242d59265baaf6edd56a69bb1162bb2fe00c1668e9329265afc4aa4eddc05eaee99991839;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157644544c16265f3f957395ada00bf95a3c68de218abc59d1530b1a55b025f0dae7b0d6901b5b505af29685cb5247e04e772824ec92d630a541ae9d171b3325760e48aaf802b4c835fcc470e6277350d17a47902f464348d8b9aa2150aff9a066fee25afe78a8b97df03f34c53ced8b49c915b3ce5d61e4e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5350680bc732f9312b4737537af0773f0ac1cf21d52f303a1ed57e721e01fdbdebb3b24846a556620a4d70b5fb337cb9e9748e4a5c9d485732d8df5b2ba0cc7feca42060b2611cf54e7e12a1de250454d82968845a00e110c900575d811124f21b4c9005a1ece7f1279cf354ac98cab20389dee5661c71bf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18cc123adb27f253ddc33facfc8402361bfd2b2e3ec389d102481523688f5c691c1832b559c4ac504f700ec8119549456ed899b029cd3adc56580f4099a87c74927470fe56c36d42a9e849de524ee6b44bf166c2801dc2f68db80fe5b1f67eda502552ddabe4c3ee113e0857a7c96a2ce22710cbb3418d545;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82e8f29f45e1a4aff58506037891ef9af38acabe9fa2366c225a087b8daba837e12c76a36ac9fc65fb0185e6eac23977c93e3769872542c6c5127c90581731dd004e79749d2b1fc8d1494a8f7f0d226abb0fe470e6febd958ac362c3bf9872410b047ffc174edcac024286cfb1fa86a36f18706a77de1bb4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef42821200025148c17f984ebce6b5ae5b17dddc28e1b7be62638854f2a6bd0433af10098efd5c987e9f269567a9d6e735e7beed04c919301e793b647356388dcc4b5ce3ac73a173916f35f5c75db805ef529ed7c9bc8a1a299154dbe71808f72bbfa5fc260ed22fb5fc797e6b31124251de0da9a088040b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha6144c4c475590a89554f6738c86ba0601d9978d166e6aeec2beee2a038f189d3475de58df93bb61459815a633b4f90c6eb1a0cb07c3c967f2e00bd7f2e9787a7b931483874b1f70faf62da496a53e7eb89b360f639216f9952574bc509755d43f999a1b18789a517d327455cd7c6d3f53e114b1f933e77f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc5d4b5bb0741edcbfb8d96b5bdc4a3f950a329406f0b44269cae2d3f567270974b006e04af133c0c0b1c9148df0a7cc5900acac2b6465e11296ad7e9c9878ba4326ea1375ae52726489fb6969a7fac3fdfd0f4ff88295abed581e77322b66c845f04cd78b79ed49c8e67a7aade8e77cc59a2a1298c33c2f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15efd2e3a74dd484d959ad40657d2c409cdb1f68105ec29b2aedbe30e9b642ff775402cb033e72beb8e1c3fb3e7fb478503cdd619e324f4b4d446ac527f18b68d07b911c58ec77881f36c2ff251bbf27f4026222c17d305de9270c91da0124951da133b495343c27692efb39065624fb72b8247708e28aa4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9050a553a1f8f9ba81cf75116b41d112245fa70dab84f826d804b54ba7f04b2fede296eba5c7d0ac7953d6012598a376e4d8a36ebdd7a0f1b549eaf25038caee30416202e0bbda3c863abbf4d22cbf96310296fffa581be8cfc7d21155bfd417adc3c4f07ec9a823bd0bd6bc7062de3e1f0898dfc90b99fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17682e9a955afa4822f8dec7b9adb98b885f01542fb6ade276ca868351a3c2ad8c5a7a8761aab6a303e2255307f09018da782510b80544c5aa1c0eb19a2f455e421194776666c31c2f23c5e3076d7f70d9fa678c9ab4f270557c92d9d5e2dd2c8d90856490422b9ee15dd5e50db36a13ac704e83857f4e6e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142eb73440770aa4c8e19ae23d6e60848792b1c8003824aa38eb14a634f64a1a90f46d9c26d4eec11a3237fa200f8bb9a3816bceadaa615c3c9ddbe38b188374426ed1bce5b38bb281d7064481acc2f0e13ac0a4d063d13201a8c338def35e5bfad6d2e6a05ba8c4977c98dbb6c37ae3820686b0f964db09c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17290cce7d4a54a6e205d9c5ee14d618ef62f32b12857319bdc7f1786988e8ecaa0151883872bb847c62cbd0d8a233f5bec6e4b71d029e11c5fdb0c2007de7a9193b33aedbc07f99f2b81b3ab876003f8fee810d0fbc4d17c7cee7ea33afa5735a688d726cb05c2f0d8bc020e9a1fd4386dccae6767458470;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e7167993e31d39dc7fc904703ab4b44035c76d62e94a07678c6baabf70e508695219cb5e18f7b08393f460beb03cb5981c6e5d2f47f6129a6f294eeb5082e15aef553e435a8d6a40ab24504a500e23191bdee9a1adc361ca50ac4c102ac7d9d814a3685a1347568025448616f9e8c20652bd1d18e6445662;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbddb36fbee7f92054fcc5ac741247c3bbd86a345e5a461465594fe20629d5123770aa75fb4a7e062236f972f8eb3b2e91246c474446db41d77e97fb17e89cdb43f1d97035506a56271bdb787cf0a1d488432a661c127861feccc5e43003afdafbfdbbcc3e0375d6d9c7cde80031ed77aedab96ce547c78a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h130e3bb2800af2120010f65147bf7b3ba3bba1b65f6d1d3af51e7f37503e9d4cb983e8c950f2afc8346461b729a9f50689f00c11dbd1042c257520030f85d09cc86af8c8995f8fa610204b590fcd09c150458b76ce4a61580617f0e9828c9a26a1b0772c17140420b98be6bef7e2298628b38545d05036d8f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h53fe24bdc2420b8fa7fa587b7eeff1ff7e069afeb6c03598e07fceacea6d23a2f0a70f9979c156a13711c4633121a30dc3210e78738fb26e5c82db247c2ad50d7a7b5d77d19746dee926f97f0356eda1bc9c410fb46383b08d8e8e28415a20cfa19bb1382688c85b3ed8d96d7b987f1e93872ed43a8c7c10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13d53e4581a3269cb6d378d2719ed9e3f2992b37939df3cbbc75208d22a3177062a6fc8b2b9eec8c103d55ea005cdb9d1399036a9f88b98d07f2382ae53c9e8f9c8c6c751f22493822e8501034775c1b47d0ae46b06a1a09ed6aba8624dcf4615465ace7eaa05a63c6d514c2dfbf732f834e077b07a655768;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd79fdf07dd347a74b779de1a70bd68806cbdc21bc2d96762a5820a813978c69ec4126a1effec9ed9c6140332560ffa961df1b703f3133275706e5dc8b637db96f307c92cd8f42902a87adc40cfdee80e572667acd6d4d9797bc69c594d1d967bf36025936a85c943c2c496437252ffbf41eed00813a1935c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17fecda8dfadbd7ce6a1b5dc447242faf6cf6c9c75ff2523d005229c715d67b13cc08302d534fad1232c4d79dbe8a684bc563d76cf2c828dd203084ca1db36b7e231a3bdb1f0d3aee045b6b21d9383fc4cabbd61bf68c77c61b0dbca024915498b59a5d5c2be352e24eb1bf830a25b15b943d0d8687dcc57d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h171a002154a0479ae270349aeb8e199ef40307d8a0ef6edbfafb277227bbdb5c7cbf0bc1f6f3f928a7de597dbac0d01e575bdd7d79eb1c143eaf310dd1b690e9361786fe90b269b1a4016f0fb6e06da80594a40522699f67a9590d0b69d3a6fb19f9b50b4f7e6ffc11d64ad0548d0cc3b281a455d88b01452;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f5bf899cd959387380525bb1cef43a8bbd0ec44b1a8df06804a37a13a162a4499ea2ce04e15878b7f3f49a633c9e5c80784bec1b081d030d01e1d9019142c83ddde950a105451155da8809437778eee5e312d1cff40813820df809ca3b0589b10fbb8d911f995b0e3f0021c6b309c558de607b71869afa6d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e55e6dd81d079f34a5a48f1ad977aee64e86e3069b0a9a4a7914289755a6096a379c0ee6b257ef45b509de905f786412103500b93a4a47e6c7c7553d1b80ed1a8e0230bd04032301adecb8f042fe0a873be34b2f8a537efb5d5439bd9da0f61329870c34057ac3244ba7b59b0181817075703cc70e169115;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd85c8787449ec53d8beaf5eef1f7433533ccc61c3d3aa65fa8e93812db97392ae12d2bac5ae1f6e4d47ce3fe851fbfa9afac025c7561ba9d7393703d93749caa5e343d3796cb245811fd6b2d57af626bd3660f1fc547b55e61e0a6efbab304bd478916f55b6d57e19e36e88a66eb2dd548fb807725813ab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ca326e15b59340607ab9e4346f2a77ed0fb77f40e9f9eb651e94b126a3fdfca5e5ea53e7c5170740c2d15c85f489f16bbbfa95a71691cd69c128bbad543e245c57396c281ef8f8a13af8d335aff76a737e2977315687c031d91be617233f18214c7e048ecd13f622818d1c8e0c01063c64c75c59d803a379;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h64010b1358ac13306fa8a00854619682b6c71306f6e59e9c87cb9ba588e68ddd6aecae891ddea8a2d07210ad99abcd49d4fd726a46debb7d1a93451b56aaf7dcd3c11dbf646f8475fdf251d95764b0a5bda69d29bcee00075a3e99b6d419ca255be91c611e9eb08b0caf011e77a90bd5d95fb936abadc0a6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c973bf99c75faaf22f2eb5f6c210b85735d55d30626e0dc00aba55298b27cb217240355b11d89b6297ba8a14e30d80c363c5b676704b91fa87effbd622fed65f3cea719591a4a2b314bea70a83175770061cd6fe054de430051155f6871071e27d4d79fd8067c0af67211840c2559a9f85310e39fc52086;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h37df55dd48c591d5657670c147f8427f10b6b539c0f73a919ad53b7bddaa8e6a8c280871014bde308e09fe4d2ad57416f9fd1cc32712cc2efbecf708a41fca9b8efe6626d88c3f6248c3622f936452a9ede3a24c445f73de8a3989874f04e1e2f9519af800f1010328b4123714a45c9541f06281ba0c24fc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b201983c7a51e90592fe8a2ab24950851c657464b0ceef6b9360f661767a31ac2020164f2a376c732f0f9c9f8ffe1053ab42538e2b2b24d1556b976beede5f5c9288c3882386fabdb6f24aa1cb23c43a07556b902f06755a643d75ce7e68ae923da60cfd2356e30ea544885d63530d0c655d10e58283e73b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda230b73046617c4de03ed99a59e41f9c312ad45b7a7d2cb58d98af4a14699445bba6ec77c0f09ea4427071351ffb5c0969e392d73daec2b4ca5087cc8ff0cd9b8059bdea541557e115b2e187d0a5f70576559974aaae3ac6e50dc484148163751395e9abfa5c20485ad58548da5e33b75fafcb63510560a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd860b9cd6ff20228b5f4384233d17d54ca285ba75dafe49d377f396751bdeceee3fa519e0197695be169b8edddbb31fdbf8d894f6d5f808dcc17b636db59aec7a72ab7c501822a098f9f93e921dd643675f079ab23a2c5d16453d2d8a4ef964b64c35b48e608a4f059c49e2de43dfc9ad98ba471be62948;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e989c5a5b3cdb0cd93bd7a3ee3151d87f225fc55d0f7e8b8bd8daa38caff2bd6de3df9c1927ce65df2032c4000ed8316d2c932bbe591ec1560300a16b9c07bd692d3713e0d3c8de348fbe8ef51bee8fab2b3c7ab3ca95909c187819f53cd7862eeefb995edb3ee1f32dfa5440057d73f2675fc1cfc8e54c7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52cdb81641cae31d10c96d74ce0fc69f59dfb7853784b58a80cc69bd0e35756155130a5b31da7cb9e0846835df459f464b0768a0005acf5a445c2de696534b98cfd5bde1fbfea2bf2cbb508701ad0179fb06ac6b4b184953ff8970260b6bec616ad5fd2c74a63d39f3dbf911704104d35c66d1593bf3b807;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17276aa27ef7fd044b8f0253f503856bf567a63d8fbbbcb2cecb294e15389065381d037274a84f218768d939977fa7fb9ab236cf503cf151350d59cdd33e10b24944804d1cc58a8b34b96cbbd10a2b9c4bfc8c60ef08cb90137a069d2463e2ccb0aa46f39e60e0c50a2b8fc783e16dbd35caf361b9929bda7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h190408fc82d24ed7fcc60513fa2d7b68939dc69c043f7a1726df7c196c2e9490d789f174343c91e93da9308869572ecf5211189d8c2b12e28edc8ec53e746be03a286a163d5b6b0e099c8ecd21358224610c52ce76527be73d8169beb777995b8c69b96a6257ebb230e8d9f34acffcbde94a215f105bef1a6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hff6f8a56516905ec96829b7bcb1cda143c4fe6b26f4dcda53cb3580c93366130bdcc48f312c52ece6c91408f901d9e3b7827c34cb0e97085633b0dd748f9f95f53d767f19d2cb941878d8efc322f4cb3c8c05d2f1014a175f3113bcf340a154267237544a228d4a173273b90b92236256a2b2647f7f281a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4451c1a039f8e284858cfac1191e90749185d8ecb713788a14284efba17cdb6bc4022100a2d6cce27febf64c1ffbbb21a18ef0af7519bde0393a8b05befefe58debea7d57b7ff2bd8c48c2ba2d18a9778b2df813b319a4b40a049b7a320a405fe52d99594be3589f62403a6e51861e5f463c7066aca85660;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1abd74a4a4b179815a150a3a29ada5af2380c0cb7a4d25cafd538d352c1b174c6d64cfb0a8ac1bc72e47bedbe010014eb8d466af7aa31b04f0f0db243b44435278f2a8ba63b81995b502ff078d969dbdaf01fe153a6dc91ac4a0944624337ad47f962e0d9c21060bfade7e9597285fe8f4db6b78006e44a00;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9985c669ad0094a27134c27a23245c3775372d48b10bf079c853cc3587de6b611b5ec8b638ace18fefbde901b8c666b9fd1624e0fce58e6c96343bcc6c61f492c8bdee2867fe0b3327031297007b6face7373a462407595a1983ef7bf4be4cdd207eae2d1a929492c9c40a809ed59d904fb4a5c90aa3ad09;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h40e96b1a3de55c1a491ee9742660f10f80fba87279267a7effbefc475c940c16488563d99979e922b8f7992f104ce628b450d75f86e75194686a2c1d283f177f73aeb8dca0f901cb48bb60b4f107bd69e2aab5aad8911424b6b8404112d9ea0559033b390814bc4e81df2f377cc0d09bdd0c5be26fc84089;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hadd9105394ccfa6af84ac7ef3f96514f30383c8418fa91517c6b5a33ebfb22c0fb5e46138e72ebc5f201ae9fb1b58e18c19cc13eb5fb8e3a67476468fb1f93085abb96b72ab5838d05d0da9bd136aa73f5c3c7eb149792a5443ff01dc127724fab57ba1718362878a9fa471ed63cd488e45af4adb14a825e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1006d1532382270ca7663203890dac8dcc3c03f7053bac16cb8be069da00e28a72ac3d579875108c3158bd9b0ec15732dae11d37300362358e65d3935d6d49f506ae52f50401c59414ac1c0b9fd49f0662b88507107b91bb54f51d4cfd87c90f77ec27f6093937e43e56a2fd81459765359198e38473a3655;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151c3d66892811105a020c21908866d5c8fd42bd08e02fd3a3b26cd707a0e8d8be53903f0abdf9665b97ac872d1a4a14cdecc7c6c18c12ddbe624366886c94b230714ee7ba31122229c72526becabcf8f08300379d334bdc8a637baafdd456104b1b2d5fbfad6ce776ff3795a9cd5da3bafb44c07066f0cda;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b095ef04945ab657a4a850d7e344a22cbf2a0c411b3efd11e81a753501219d099fa674e8dece76c4f3d08718aa42822145908bc59cf9d9e33a8d1f0644fc07ae259d1d0f783c138dd218bba1c28689ee81b27e20fa6d9c02145a0024c9eddc0602efcbdce04879d70de7c4b6915ef3572bd98bc5d29cb7af;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e2c3688e383dac5d7f7c0184fddeff17c7356dc9f1e5b2588ccdf2cbf793d9edb1975f5ceb4207aa87b898c465cb837f2cbea96e7bae96a8f8dac0a2afd5eca8b52dee68328679e596d1be971dcbd94801b4855c59e070868b4f328072b76fa7fc2cb1c01246e31427c2213538097544d6fa21b3ffc854cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a0c871905a972ff9447c3e35115bbfb39b807e3e0c9783fbf49f2e770246277df99f9a9bd9aa47bfa6a61e7a313c8772a5850c4568888e7d54efb28cf0a6fc360e61a5370f194a541798dfcfd680ee038c56a0fdf5844a8dc9fd58b58dc870a8e79049af1ad4af5c7718dab0ff19dd12094389273b6f567a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e6a9e69e8b36cbe4b88ea2098941153824c54b59994b7deb18586aa860f82ef8f34bdf3bbdd8591358cac88088dcc72bc1fc38817f5a1b1c73a1c9fc49e860a784c845d3bed66d67fa5592be3cbab8188b0d71e7ebf8f7f126a7f16c5ae51d80e7813480a07d63c860abec713d185959f636bc2e2350244;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5e4dadb15ec9122824541868ca12e1bb42cb006055a8d81ceb4fa38e6051875b758127f01535af1cc2225e4435cfaac1cfaf9354f0b6a71c10dbf1c335d7831e10fea1fa66185200df19aa3d93a75643cd680644b1159aa170934c64b47018faaaef844b991c78db0992431f67987a0a87517622fa6bbbcf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d18601a81a2cc87980cf8112205131e2c9e209800f091af2f52e4519b67fcbc320de5cabcc407cfb03c7ea9ffeab2ce811088de262c702ac6a6658c41c2d5a8e51c6a49acfc2520ef8c1fccfb087065025dcf22c79704efd6cdf1901cb3655f2da3c910b24d72692dd71a4a68df55b06472c52fa178b3cd7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h20f46db9809efa929c3f2d1e1f23ca7cdc5973f4b0b1d122b90823d731ac0efd757e3049a8587e5b3052518ddd175a5bdb8c1f9f25cce470532461fa16881459fcfa396a22e7df99688e7487730c62ecdc287755d939b2f92890e1cc4b21206c2e4d1625041b35b6ad741e1083f71b551e3aad483d569937;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha34284aaba5ae52f83cc429123aa91c23d442f264e4517c364aba23de518777ee84776e72718eab7062f997fb01da58304761351c445cb3455a983fc234aae25c8d67d5e20ebaad3f7092390084c170b6cca8e599b2639ea67170bcc6944e2ab715a0a3b68bf3c1bddd8ec1433df19a376976e399f920235;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9471766a180adc9932b8c66cb277735163ac5693dbad38c288c1eebc19f6566aeb5768b6ad0c20afa1e22f0dced1dc2f71ed173c830e60ae0213195ddd6e7d0167eb1d4f576711efc434c5864caa800000b2aef75652454a99b94c111e39c1534628eda01ee0fc3374955467a428af9c74ab7261965b3877;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h76a499b8c60ca7234de1cc587e8defc5636ad2a68f8aefac0e245214811cb746d5df69a987d283aced5daae745f0b562e61be0523c1074b3e437aa7c07603550de31fc5d4907e9d145a87ec0c6b6083c4a7f81a26ae00e4d69dea7b8a70e75f0a79efa59facd36f686fc5dee654ab61c2881a64748e56579;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1388ac6e89460fd99ee2e21a8c386819dbe0b07f4a586131f4c7c010fc38f63b5efa67da3c111b50530a9736fb549f3e33cd2c77cb58a47acbb3e5ee3a4c021571f60f1dd1702fbfb3d3a7c971decb9fa21e7eb3917c3d60fa70a5ee1c652d02c140aa83e2b32a3e1559251a0724d6e5ad9077737d8bc1e1c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h130002ad15045ea4ff75d54c41d6966c5d376073195d5c7919b2b0538b480d274351b76540c634a0cf0ff114c65fcb410f86fd9087b4a69fab88021483f88486daabf255bace386b84464d29bd766e71c4becf04fd32cec9c33fdc08836b8b1945f94042aa0fd5e39f4b82f362809cf2834e51f985ed262a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h812660ef2e61136f492725ef4c97043510fbfc61249e84e7929d0e1e68bde7d9749bcdd57facfbe5949297c16c8f7d25d250a3e7f26fb643f3f9ab0317904ad57d502799c62414819f8dbcbfaa3ce5eff70a1231a039d6ed7018a6ddc901aceac07e36e13cc1c381c7b53a729fc37b0b22bb035c9b2c5204;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c9eede3308b9f9a223936fe778a713c311c9dbe7317ef223b04cce5471313f0099731f1b8fc3dc10bd1faca66909b66dab00e26485302224173d45512acf49c136c9059fdda2f339d229cb50382958ab0b1b06e1246cddfb6d51b91b7ea87b936ddf5d2e75bb705e52174c283f30247034584f86dbcf8c60;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b9194af7e9d0a2fa750c7b5153df49a3feb892e6943dc0091851d6f0b528c81b2c004a8476d655ff096f56e5d5a01f506fdc61bdb297d55fc9a0f10cbcfde803ff5e0a098ae0c5f3bdae9c3b4811eb145bb6905b311191f1e5dbcf0acf02a9bb5f4cf2613eb99497b688327a1015a1ee3f91bf8eb20fd38;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd9232aaa01dc49c95e8d454db3f7831504c9611f4e87c98c83fff8c9fd77e7adbc751992d29639c2e12f218e5ab1d5b896b03c3a58b7236fb4b41af80e96676376aeec4a42d4944153fcc1b037af01d5e585400dac2a82edeffec94b33fcec7977d046737c153fab2559da293b76f29be9d0f67e51278304;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d727464a378632354a9c1b9efcd0960adfc42d701c301f3626ff8e759a4c21b359033fa48191009e794170d262fcceaddef16527c3f0b99ef1c2144b294aef4cb08a298925e4a198bfa4e5d50a81ce8286333e99b4e515b1815c391c9712be479060ff1d72c88a159b7d8050c1f9893629b0360dad0cf82;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h125188108b95e6c0d87cc46036fc40a965a035bd556acc728d974428631c6b6da8b176e12041b768d688ad23aa354f1d0ca30a16ef56f0331a93636c6d9f121c9d3a26d50d3308994c29c6fd8415c223bede41af106d7e2cfdb4b1320b5a83ba4f04198821864392380117b74aba081ddadf29c371f20fea7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc3531d39678f8c60ed60b17159a47c7698da1a6b088ff347691aa2e0403e35642790b38b5f93d96bf460195e1c308165d7fad4c0806a649819df9d4a09b3f5453cfd4c9028297789b2c91ad303d96b13f97c4b5fc36f7843138b7f80c04e1cafba3cf8107016f247d2ad69c4a4418786bcb18ccad3faecc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h111b5fde0ef7f4baefcfab4418f23dcf483f8c47ec85a6af335e2b06c97c2c4f8bbc50a2a48d9e19e5227645f7c64de694249979945d29375893e6d59c712ffbce97185910f574738b4ce5e71dad15b7a5441a1e5ec6e9a0c6baf9d30437aedf37c736a70497c83ce798e0bbf78f9082d6b8d3baa235d9906;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8910da32e5b382463119b73e3f905728ab9de3bb05012b20dc7456991566257594fe72b6ef25ae1daa65f6a7cb1afb90a776e12d0d6d873cbbddecb8f2ab4351c03b6eb0aef47325ec12357d8403b96a3951ca1546e547dc21b04201563fd45426ccaba0282fc4045962e6e49638093e5eb695965b714fd7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h160fa3368447a888d7674e942b39ae031350eebeb599fa793bd27d8baff099fae00408fab86735d7a344530071848408c2fb926c00ce840c0ac6969776e05cb47df4ba6ba47cbfe8f6c3061bc890a5d6c09ecbfbac716e3f0fafe4ad7067a955be076eb98159f98712c87e9d5d08f71f43b86651032fc8c29;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h121d4e02b6e56a26657d34e6430910a7e78d6fd5d823d1b7af60485b3670e9bab3b8eaba2508fb1068546a6040e0a6a0527fe4e0a9e40cba4313dcb544b162cbe8ea4d5b2d15bc339de03d9203226fb54ac20b42a4cd1282b04c8250529f9d3e10ab19a2a0c393effbce884fba6fc83808f23a35f6cb249b2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc54f1aa5433b2dee30fbd2cb493d98f4712931c55c442b4d2cd0cac9df0d394e98aa214c8df6d807072146ab1309aadbaa75c5ae21bd8ff446ee16535f1422adac7267554205d00460bbf1f18b92c65f2ada6af8bfab270a767a9ddedc1206391d42ac44be8d507a4fc2194ef911e2c7340d22ff279aefc7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3081fefbceca057491c6e4c09067081b73897da2688d3ea7eac0c92cc88740711cd696583da356b153c0034152f4427066305219b873b3c8baa8357a104c2b5ee61baf9803297681cb9c7a87a9f2346bc6cc62c6b0f35046a9fb39925121469aae2a7459d17688e7bb0d55034edf6369e47ea8fbde75d0d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8935cb35f4ecf2bd1244dabae392dc10439233c25fcaa2c5474e9e76f510357450ba1331b4d97cc79c04a0bb8f619b2b2a6919049f7b400b70d8eb8757deda8bd9d829c309b5db5e17aa89ce06c71636c431c2a9ea7d22b15fa5cbbf492a31b8c6712981af376e5d466f7792954841cbf70b434a4e6aceb6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h87b5f6f825ea35f063c3c32108102eab95d68e1a7d70c69ab414d7237f3519aba345033aef0768db94bd9f29c3bcf8543048cae36c4e585322b003de04b319e43e8572047355285ba5bb01f8337d97f8a44bf589e61fd78462c7d72fe989ff0de929b5e5bf2e7be77dad4d3324f724e696862aad9884ffa0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f17294f8f9c8a27d41e80487e7a9cd609e70a1b2f4e6841ed7135a0f8034bdb92747f6ab1dcb3a4961d93ef68e4d6bfa180c3f4af6c7cc43a6431e4ea11ee2c7662f7ff4a137b3f7207a92be8582306e89ef0bcb452152023ca1ea921c38edc2e4ffbdf7bb37b3ee2e921e3b9c516146b9e4ead811c0090b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7011c2e35a0619dfdcfd46c9507705e2a586753b7b8e06f19c94b82abe34f7124892aad631fed64f51d24b772e8499b09301b896d8117d7776d96aeb9779901a03ed5a69c7ff6b75518f27e3c3b7d4c2abfa8590171180210d5b1b00fc945d7e619e770207bc7ebad7e8fa9fa10a3d217d31c7d59beeb8ab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1304d9109c40bdeb4bd6e1368f107b0ebe7ec120a1a2634421e9e40b61347461482ad36d2521312a5612a85fa8c8737367677832bb3265050aace37bba06c6c55a3156faf24503399d441d16119f4acb92148feaec02e4874dc105376ea96f260dba48536adb0c3d5bf7ea2b2842180da2105763b7548fe8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h122eff0703a1b3bebfd2660f38c1f25bece22c2a9753d006e285fc72159524b18797e67715c273b40e3f3c528e9ff5690adb9ff4d3d46aafe3fcc67773ffc185f496b5aede6eff69f6a64ead50f5a9a27ccf996be42e326db14bf4ef622e25be02e6ebb52e2f3abedc8c65e9a92fd0a1a666b7733d1769bce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd8bcb21d49ea444daad3b78bdef5141dacf0c7ca90b93d3e6d9254d1e5d49acb5fd2ba08c1a50e495e1fe2bc9a5bb1843aeb69702fc0c3a56abe22b2fb244ebf5085462e7ecb9e2a68b6b9ab7b930157ac3c82ec92d7490567d5c99c31a1646fecea202cea5e1a026b84818c8a33678fd825907c7968b037;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb5cb2b562dddec3fbc1770a8b80742b98e6d8d10170c1c1ce6a075fc35a706779338223c0822b70b4f759f09e14fcb9be75c68df6a292991f22dcb7c201bcfb2a5bbc5778ad56d9f755686754b0ef2a173897c2aa03ba478b26b3107d818990fcc9b45623e8aaeaa6ab2ce26d62ba8ed8eafc68f05d90a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h135e27c826ed9539d25839bbb63b216c7d43193cf397c679d51715c51d91b93bf23e22c709125a7f1b3fd0a854db3a4176a3ebf9fab837a85d63947116a4eaf924647b10af0c872a8a92eb7323636f6129df4cfe8e3717dbbf065b7e7389e1f7a553f4c530b24416c7dcd7fd28b842b45c186edfee6bccedc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h98b2111f6cf473feb44106fc5ef1e45d783f89fbe762c6524ec640daa584963d214466a1f7869c5fb4d5886bd639274d7d9e13542b448138451b82ab219de56b7dc119b8edc4b9b20d0e28039d3870b72865c1b10ef31badc6c702dd2422fed3833b7610f076f2aa75e8ce23a332243b66dfd395e902eece;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b7024695222384c77859ac3e3523b429ca13f728492e341d4593743617bc581a27b816cde1e2144ac7c0fad3e48176ab951ddd31120a9955842dcf6ee1b04244f37faff6dc9e4d783cc4c325ee3264e9cf79c552117077ed41ba2d01f27202bf3a92db81e3d0e7b9eaf8f2f73d0ff93e9ff376e27ca2dd96;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h272b4d823533529c0111716bd4ed2fa281ee046b5597226d0292325b4bb215645233d9eea94ffa59ec3febee60f75ce1fa1418a112ee9ef046e723723d0d249a21ae541294dc99d92f8532becf3d9c8d92980b5c3d6b1fe19188441638d3b2bfccdc61f511763b70009df6aea8a70d7b79630cf4134eea9e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d7026a20c640f653a89ab6e0fa1df25388f6694c084f9279c8f6cc7fcda6fef478c64dae9da13f5ee81967d894d0fe601aa0e13a15566c57c8257059f6ba6b14925e7ef8506c7fe80c04a002379c70f7edc3f4fbc5222e9207953b4c83433924ab5ffc3231631427cf25168d456ef330b632730ff9de04f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1832db14655b5989f6225d07e70680c3bb142d56587194052a61b8148c292d3511ea9339ff3b785e2f0c13e4460e126d4b654431d52727db409c98a4ef8a4202bc3dc903f6b460e817abfe44226a80e4be7b4f67066ccdb795c307c4fa8d56080a0515ed64cc14455308c3bbf7da7540c9ae9721f4304ae54;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h21b383b6cdccd9c80dda01cc59c2975e32e35e35740c1d122a878909b9488fe43b113df3b7478837b4cac30573eee08b00726bb1b6a354b4ac5a82a4424b12d5e24d55e3cb65aac71607f7e7ca13a01bd6fb5e9b9c6fc505fca43d7e3b660689ea1f25f2614fbadbc672f495f00b0476d5ab6ca82e419a1e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116c8a81978c7dc608434f2b4886442ced850c2f76cfcfaad956cb1e530ba7099ec29e93b5901d7736f92e265603bdb1d8fd4d3bda5337453c237856f48f60733bd576f9fb540f941fae280e2a2f76ebe3a606467035d00f89ebf9a5793e86f2421638789a5b5dbe8007881497646a5c64bf48cefaefdc2f3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82a7530d0c9aedd8c2f1066b4489db13e1fe3f39593fa5094dffe0c4c29909b80ccb9778eae5844dbe6be7b66b1d73249a428df5fcf4b1ceb8b32fbd0614108a3074f354158bd47d15d8919452bbf923273635b8492273680276522dfd2284264a15e2067663c655c713849c51ba7da037167ee6ffdfcda8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f9a4590b78212622717b41a8805d980bea8abe7515cb319c1d972b68ec21f27369efec0d4d3b384cae4ebcd4f3113609754e54042ebe8f07f29436a7474b830ad8d50995db51e63184d413ddcaa96b37983ae93fd01cdad587b400b7963e4d4d6f7819c5e47a1db9128177a022768130a6d66735577d274;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h348bf6869d41870e23997baf3f9bd91dd37680be094de2e6d193d6f5463246c83fe9af57cc3df78b05e44ac79c04dc8536ff4347a8493d29baa8fca4bbdc9c98403c31c3e164aa4495b37e58f8c650d055976af64682e1a7d64ee8aaaff6b28847be5fd2c81830ae5c6ceb2a80581a3254887603e79ce2ce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d5836055a26dc22a9917adaee816b9e4c045d6ec4c6cc92f6edda3f67e27735ad92c8258a26580c8253fe3e97a9397eaf234ec6e71cfff3d39f04d04b3a890460cbb238673f4865a76ef3b224aa2676378870703406a1d2566f2140fdaf02cef24043c4b54c19dac0bf74dfb395c2a446da0b604be991d48;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7bf987ec6ef43fd59077a2b4591119427e34bbf355bd3faecbb54d5d48ed192de9db5591dcd2c08e209efc045b6822cae75778f5eebfa2da00419afcc452af960c590ff9c6e9b0f22a1ec40c6b6655e77615f035ab721e03031332faf6bbd970975c7b45f01293ee44425d60d73b242ec721b1bbd245b0ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c3ad9345e63df58380d96f39b08ffebe448751b4063658f832927d6e43bd0057bff8ce6f4a924cb0f0435e938fe637dd44687b0408d6cf663a0a0098a86eb25358a5958f5afcb91d6f5ea9ee54ce5a573a8886a19bb3492c4e72f8008aa874f413568cb10150cb8825e78efcb6e87fc34f53adac4ab848cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14a659fe15f26b769f838044aae9027ce0f4d69d632edc78480d688e963d09e830d96249e9aee4a61c4c846791e51970d4bddcdc02438f1b4a056232cbf2f4da7a7d8df1debe1da32a784caf28388dc511cb5655a955ce52b612098681c0a1854ef2374144176af413ddb91e9110bdc1ce1b5ad55f5a29653;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h31c771f5f32e62f87606dbbf16f61bde2657f3c604f2c340c0b2514f67a0c8fe30e0795afcccaa58b5d653e4ef340752ca2e84c3326457c1af7f9711461ac4c6dfba522cf89a8cfa8676e5a4937184825347f7a955d8b0492dce2e22c33887343034d50bb145135198340cdd952827ddb54ea50ad0d0ec39;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bcff8261a7b40a1db4acbcf4af3ebb3e768af59e309eae681bd23ab583ec093f95afb1a12ee0a413f5838f0dbf80288c398aa09e550f8c1ca80508f9fae47662b5601ff4c02766f2200f8fbe2c8c7fedd5e07eb62e67968c24e34e8b9c4e81243ee4c225ec145451c228bea8d8565cdcb22af27dee1b547d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8317682927c171066ec681e56e3a0a2f254cee2c0933199187a2f64f652ce00e41df79d45e8563b90693dfa6b2714e0e783f4de67de40f3d9900d0bb4826e0cd4945267c4bb26ce9f9d5dbb3d2717ee183719ca81347e7bd7b03b2e22191bce733c16765983568874979bf4b1124475d1dc56b00eb03bf67;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a0c366a2fef6fe0bdc6f54706373118dc7c0ca441b215fa7b891460b30dafe55df0da6a0112b2a3473f88140db91311d9f99c5787430b6f221247d61479e2d83d8c4dc23bb5a52a88a33fb15345b6a2a3989bc12e0becb07ad979a7bdf87f0e80bccf6da52eb8bfb2aea21f85bb797d343e5bc77a0c5d29e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1669822d098a0329395cb3df3481f51525aeb7a0bf21a0542a32db0dcf92f18115a06e219e956051905533f51778e78ef5d357a221c57e43bc4094bbc95f6ef2c0e4333b49f463fba1cdbe54b85c2224b0969067ecdf89ed67894e2a471ae9647dab043e8b575f5bed4b934e6ee6d1acc82ea710d9a4dfc9f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19bf2783d26adf1a75f18a10df3b282532aab9ade3fccb8a00992dae1a660d23708a2b52e2bee68a814e49ad583134ce56d49e4cb60cecfad62840ac6f11e3238b3485db2bf7ada8e5c68cea6cb8aaf8e312e3e87aabda0347bf2f962738dadb3afe5ecd483cbfeb9160c4ac3bdcc4905e3b5ba4503a1a8ce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h121f7a291536fd4f876517c73a4a5e6d673678e0da2cee3c56ecde8f0362c1c9a161efd18d1821de99ba7c66c280de19b72bd8a28c2dcc82b8ec88abbdb69a345dc95a5a83807f7720b9f0b0bda16228a10cac4c5c33d60cb1a267880a5f0a63ac2d11a8ed9adaa6c29630557b115e12616375d1de66cf680;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15d8be0d852d634a553697562f31853eef4b133d378f5a37011ff6bb33841de94c624ee95d77261886a8dc4fb096545fd322f0248129333724a8053038e28ed962f0d110904385aaa92d00eca34922fd924d863b26792356a3494d6331c5c78fe0043c44db5080f81c883fc88847e5c2871d268af1394b0f7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b432430f09ee94d33054b61770f6a58b63d3da6d089d6f7ef3656f0ed7eac93c3b3852aed3ccc5f212f7f703d1b9b12132e36a7e7da1d90ed4d1e8e31a2094f99c208a45c637cb3083ac7a815ca2229b4a0f38f83c01e063e77d46f08eda68ffa7512ce071ea27204db06df203046602deb93d3ec17d652;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h42924442ee38bb1dd6e75f04148cce8990b85d40e68c0a2bd53ee86e60dc895fa550c9b570568292cfbdda264e432430325b01869e083a26c8739e339657c825d7bb7c634abbb0ead9ece265f252c363babdd76a694daa3ee663fdc8e8eb2ec2240c5dc5f9905d03b039fb3c1257cc07060ae6d2b210904f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h91d472b95974d57ebd6d955a22937aea8a874394c3cf2f9860bec753d00b1dd3d2e5aadb67e2aa8068e6f2b8f14617a9789fd970460e5ad2abbe4fe5279dee5a0768149e4460f4f67d7baedf30fd5879a29a0b3f1600b942bdaaf030fcff09cc6d8682fd92d655751332d677fc2b7a9c62b7ef555b87cd7d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82f548ec7f5011040865d5d3c29b12303b0c66061d74057d68c07d5bb67845d8b861eb66b1c4ff28905ef186a290cab8346d8a721b3503320f62a8bb441afa9e38dd6e47016e486da48a270073b7635e3bf8277852c02598570bfd648d4cbcc397387289f230dca472fe20af3a99fcf30fa2ca40fa3db556;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19dd9ea64f212349fb04472bb1d6fe3559ab9a7060b3622e27ea8123db508f17e5ff7f6c29e3e38abbb38f5b0153608fceff05a625613f5da26808810dd42a75f9cef838cd772d233df1999fbd9d816fbbc3aa7c486a855c61dbce8395dee4ca44b17f883661ca2e3dd9c16c46fd9257154ff16bd993627ca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b9ff2484af6205c31ab94f2b35efdb803c9e527cca7121d3ae968004402bdf696f2b5d40a11ae1da763e0d15d472b8cd6b070329a142de07b8f699b2d344bc0fa7bf0e9f26f1d6d026ff1738c23bde6769d0d1da293195f70e3d84759557f49496c80b639a9ad990106e895cbfb8285b162212849270a96;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h145d01b4d1c14305d8dcc4d532e08ddeba81b6207212a588f837607ec023dde696d196401d5422a3252be4e9afef3b9d06617fc7f8b55830ebcc10f8b15493aceb770ef814fa32e8b7726d56e38f4b349a4feae971264a8350c905c37c8c379e5ca75fdbce936e606b25087133ecbff31f079a4021c1c2450;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ebf5f5954058cf5d69060df4c83007e503aadec80cb45854cb3f61007883ae15f6927242355e517e1c2cffe5e765c68e2c847e5af5a6efdf3ca8f96b25e5c4e74eea7ef49fc7c43f3dda7520d3bc17e6257e578e0518c03779f237f6ea6eb01cbf36bc6ba5f672e4b62932c15a8d8186a7776446183f162c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b52ba20c0a53a3720fd9d7c672ff07c8ffd20eef35dab2d5a1dd93d5569dc7776fd8ef7d53825e13b9421ff578011259bfb0f017ca67591025f05487c49604df312cf34647d5ae5c8dec5e7a052c3a9c498e0d4d06c62e035c2f70070a5d6ed2668efd3267e760e2e9783a3515644512d884cad497453ddd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8faf902f57115e8c7b4a70c46eb6bc420ac74bbee937e97c8f3e19a7621ea1a3597b2754df13a3bb39ce36dadf1d6bf54d976a5ad989a778c14131e812e53b33f30fcfc44298371ef1408944ac04cb21cfbe327a161ef3aeb57703dcc8394b7be5ac834e607cc47b037615250a92afa98115d2643eea811d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a48dfd10ea9aa1d2a8368c20f15c975c6be571f4579a96248f14740c930a86ca69973fe3addfe0372d6fa79b2fc89df751a82363971ca6009ab7c376365be64a028e0fc30c110077a05062e688b25fe652ff2875d16955004590e068ae7e19710aa99b7ed00c4b2e302b68394f5d075b1bb0b1ce45b92fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h217be03b75c2a40d1ce5be8c5ac0a3e9958c340046487338736f684f0d5ef53ac083c8f6b826a0e561984ddd20989e67f3ed157a1fc544f112120782b3842ff115390af03547403b82619cc1ab8861c49f79f9c60d3c44cf0da4fdb8b9ff1c0b3803f58d228ff4a208ab8d4759c56eb58701715b48eb9905;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b9e79bcb62966e657f250fcbf49c060fb79e2a8db0015bbe42dfd3e13d859cfd211e5d4327dd9c3ca3603b16f6eedafb37b6d38d95090c5275952f8e0a360c8270b4320f61919158a5075fad025ec45c5dfca4a33d047eb53ef7eec33343ad879d8e6a712b4ff10f481f574ba3d99854247d8bf7b6ca496;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hff812634d7c02b9888ef54fd1ef90debdde49daff4e8f1c3985d24832675b50b8c467bcec2ade71b20a80052d99f2c160fb8a33bad9a2bad0d30d21690c052c9d7409f32b0ff525c6d81592c4db002b6fdc8e66c71ae01149287f4502fa34d386a28d84875c1ee1e37181af4fd8151ae8313501ee493569a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1971b96f5a2a22cf61ee291114019cdf9688094a3ac470989625790577abcd04904aa0120fe6f5e75a5973ce53460378a4535e0ee56ad6edf3b6152e2c40985c791dfd801576ad0fd76f34dfbd4653907c75bba30d8aa2dccb46094a421568ee179898676d1adf3a1d112d85e41bfc7fdddf541c4af6df179;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h604becb7976a8f785cc9e72160e75b7b5990800bb38707722df67f7ad10175c9c527a995c4af7deb1e9091bb6dc934e14a51d103ab237590a7f8ece80533ef328ac46296f7388b6a809c86a0f68d64aa3ee40ae9d6b8f1a93771ee0aff1b2cc869bc48893010af9c5c0465ef660499631c335b18f96365b9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd22ce6eb307e31c1b2570e44b95637cffa134a4fd534c4deddc485f4d97bf5f1662ef5edbf9484b1a568b339ca21ea4f96333430e1cb0fdffb3f4bb373685d979ae19095233a8613b49c382c24af534e253c4836c0ad1b5b10da99fc4affd2656dccf95a9aa0ac0f18dded775d5769df5cdf02bed10196d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdcc4d5d96aeb14f3eccff7487e1fe91c4c4d05d67b890e4c44edae9e75ded739636f2c8f5e03a01c1437991ec10a197d9c435895e5fd5093ebd018bdea841d5959a1a5bf457f32bb38b748caea0a12b29771d826a207687ce69f9daa3e5fafacd636135ab90c878e915c7244ed759f39bccb50270f1ae83d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b9349ac2552868b52c77037483d188137b3929c412e68c1f5d69df01f682d56092779fbfb773a339755968e62965612aae14f3c7721c36021cb51b313539b8ccc6dd63ad10dd91b107f682fda95a36a18ec86209e846a77b5e876343f02772ec20b913479f6c1d391f9251619ebf5e29ec4560f907a3d566;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d42b1bb98f53113947a4b13f3eaa94fb1cb3b0ff6b4b501ab9235ab351a21775b08ec5d5df1bc0eb89423a136ed05a22156ec893aba7f71f5688378597abd29904fc812706bb11bfa8cad642458f9531b2f4e32aa43b6bf91f5501a2490c8e65e9e57186a8d093086d6452689146481336f2d62890ef3cea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70a4041a07f76e6ff11d06aa7a2cf71f239c967b86f66ea307617a907884d43a924830d953b277db3cde7a158e8f9581ac3b41741e20e70f44f680e6a92ffe768f1bdbdf248a0ba748f1e77607bb708532a9f235059b4a36d69b38d4d5e2d595c1f9acbacfd646a2f5191fd07e2e79272eead73e7457a4d7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h615dd6eb52d1f24324e7e057322ad85cf48bae20fe73b3328fbf319b383eaa1623598528b691f50f18fb3f4cfa2d978918083ff8cfbc481b214ee00f7928e006ac425c6c357cd5487d52adf7ec258d31f082f70fafb458894905589d8a24167235efb68499aa9712c103d2f974410440951495199c2783b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h125b6740d78e2ea0cb5049ab566bc601337720179c87ffcc3ba31fc05a276f5f94c9b5e2e1656c4ed7fd9c0c49fdf592d3a96faa71f69234449c70b36030909d8cc5fd3024dd55638e3f29017d230d865380376effcff0f187426158857b75a9df972105c81c34ede8c4071e9384a40afe2736cce70e3ec48;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha40766137bec46706f246d7ee2ecdf008d21f8c2faf3eeb33766dd396e57ffb6716f7e1111949f022aa782f828ef7669ded3c33c3f2e4c11faa73196c15696351ae9e65b8e207414da4946e98e4e4ca032ab6a990a43f945a016d6249c7c95d7519f3d0bd67facffc8ed944b2a477ebb4a00339e44fc5a03;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf753cdf640c389afac550f3e1f425b28bee1e0cc456c656312b666329a998445b0a933a47ac91cda3fd471d7a97d3bfdda06c5b9abddb5074e6f6df84b83d992f94bd770a85b287887c2a383ffbced6a2916eb06f0d097b28c9d3da72b9b581cdaf0ecfb185fb6c5b0c1c61b7b921509bff531f05079d04a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11b3182ba00d403921bce030094c0d38f86b5b4afa0536ca22b38a851862d5924e98ea02aee1ebd289551e9a4e2beac755bb00dd65a6dd036866a1d02d92b383ec9df44bce64ca9766ddbb7db46075e12c16037afdc012a55503fff0e30a22fca6ccaf0a12d22e51771952373b093e590017a736eba256e76;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h174301b3cc39f28368aa768dda99178e545a4fd5d983948946a19781c76aea217dfdb7c8a9fc6f68b73cc494b0fe07ac78b5d66c3e276c98b6a2715d7c1d241d29587489856d5592e8efd1332cf9a614e69953ee91da3cf7f43cb26eaab05cc66e926f0e4bff6b37c25bf79b5eb10dded8e18f6af660e2a5b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b8ef0147eea2d1f1732c63d49020ba92f38db6a4230fd40a1774bf3621917cb77aafe7ab057857a27dd2e3470867f8f9e44c4c3246c4b7e9e5295c40e95e771daf222a76ab7f6bc11a510dbb8ad742158319dd99b7376ea357c5812d000c3831c872211ce657d4c72cd4f36d5880f1a4aba9762c19c3ac0c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dd1e566da276f690116322e66cd1ae74a50a947cd89ef6580c60e23500695da5551999910381c9f45bdc3876ced7cd0c61138a412634441ac27fe98b708518f50063c15082fd1d70521b6c7bd2d02a5b72a6b8b3794a6c72e7c50b622058331ef83cce494a8cbccc898723fe407e0b16ecb08d12a169dbca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd121293ecbd891212f1f2e6a5588f9e1d5c7b8291323ac29162b7e24f1e3f2f27143523db449d4d0d9449f945456d60b4f91d09cbcd59a20a5ac004f2c6f823f7d425bc960e839188dafc41d133c3f53d64c647526fad53020bd1e69a9847c8648ac1b9849fdce9b4841613a317ac3e9ae4e0a04ba137e60;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c2e3a1b2aef25121b10f8cb4123acd4754bdd352e0da7dc8dd285682d6a99ff21a369e94a34bdb90e1645a64303660581dc8faab2d8affe56c67a6ad6356ed7f6dd2799afdb6cf8513744a45a777f62bd459156120ddd5bc763d16472cbaaaf0d47cac7b1b7c405323c9a68cc9eaaf4e86950d5a06aba15c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heec7b284df56fd10d389a2173ea8f2edd1ca00f063fa32b3e8c560efc6e098dc33aa44a4ba8208258605f8f8dbd39248c280d34a16421b6a4379c99b4275b304f544f647c0af51823a6e8e25f89290231156249f0460c7ff503dfc0725abc1daa2ea458cd624164ff946a18365fcbb35cfbae3705add8861;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h103276c99757deb491acd028ab91b79eddbfc8826fb5246097f3c35a97731b8ff8ff85638443080091689b25580210585466d75b347c866105678a632ea25c4300e9ca5d4003dc52dd6f85c2cb4f1a01fcef329acd6bc49e6ee9b299fb7edb599dcb9e73092dc6c36668ac53cfe28e4bb84f6021519f22a43;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdcb4fba090f83bcf38f47152179e3f7869364e460e123e67e8a13b98873133c983043eeaa66ce51a80604628dc66fd4f9c03cbd2aed1bbb2d1d572d3394ea2392d00c70e111b760c2f84ea770ed755455f7e94fc4d93cee35eab183900f73e0c046587ededd2fcdcc031fb322776fb4cfdc2ce1ce34c26d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10ec53cfa480686f605b7f167879e81d4ad5bb38f64f9270f2fe843a049d588e29ab48dc1a88c483835efd8e24d62a81cdd6817de3973ed18b8d8de72331bddc54305046269ea2eb5ad74b9829f7ddb3f845143c62f970eb2ac8c8e112f4a154f590147c50bec12b70569a4bb63b8fcab4bb6ffe8d8905c43;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf2f78313a63ae8e539a9c93c4527a26ce2a80e04fd6faa54cba706e34755d1e9916d090da327ec11f6fcaedb55a3b51623efd9b735005767744b627102a32920aa3728644e2197b1ea57835eabcfbc2538a252c842c1d98f392c3cd07aabf7005876f57c9e0b3749d37c7fac5d43d813e6d72fd16938f73;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4106411181957164a19f2c71fd809288eec85321a19ec78fc6b117ae472f8621fc770e0902994b8b15cd68d1a989eb0e3fe57e462b3774b48524455f17d970e5768c1d9499eec0a6596fd08567fef40b0f2f48e69cddcd94dd20c32fc4784f91b8a6afb5fa9a97127e9456d8edff4481bd6b08670086fbe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8414020ce313631ad3107506400ade839027865b4d97b7baca82a3cbf6e63bcebfe9e1c4f873686294336a30ad49f61546e380680ff6e9dac3bcd147e771d94be58f485bc896b06562dc009562adb863cebe0c3ded45c91836333fd77a78d9dc7da4dde20566e33231eef9b915cb44afe73d33c3a3e77d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc4520ed929b03c6d23f0e1bf3f40bce4401b3a9373ebb915e3b4183d360fc924bfd517832b9c2c430db5e19b731bf3ce2110330f48b131c805abcb68a78cbd5212172f745ebeb97afb007b6fd0390939247773832b6fdea98565aa183131695274fa407d637319d88b7b77a309b898d095e3e3d848c05ee3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15c4b633434588e9d997b4839c51ec47bea8853dc8abb446cc38dd9917c0c8841d99f002359cda398283c1ab2fe65dca185d67664846409f37c6843ffb120065dd73ac10c4aaaa126e745cb4283b2bfb9ff1e00f5e59fb6ed380e4a6b776cbbdbf2f21ad752c5c6306edd4b0b094ffe8ab15f80d2d191423e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h56b454936656643185940357e947cde2d30fec4dab31f542c3e6422092178ff24d49a7bb4ac5923a0320c59c2b255660e3f93e2de2b3aef78651f18fd6519aabbdd202c71dffccb22cc2571e15d7d30533e0dda0b22ba3798c813140ad3c19d2ed221a1dc7c5b6d1307ac941486e9c185da9bbb966b858ef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcba6f80a9daefc5d85ecd6e3b33e4ec783cb3c7e4c4ea0bfc417f0619d97dae8ed8c9762f8068b3d53a2d67b1aba29184392d3423d2a8163540370963bebd5564faa4ce17971ff7c6be44854d5df9410c817b4283e172d1cc653c4d1bb07f8846121fbd10f3ca8d4326e086b52eee7f56ec14301c6d9fc5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15bf952afd2b94ae28d57f3bcdd6edc60a1c3b33468a11363d0fad7e2b380f0402df3e8cec524f379e4bec1e7f6691ac0a0aef75a6cd909b8aa2cd4e39f76ee46e869459f2d5f6d542b4cd22dba2ad65752a6762bbd915e2feabe548b9cda9112550072b9c3491efcf1b1abaed411e040b0d516e9a6da18ca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he9d6e990e376b23db8cc4908e8ef67dcceed963f1df4beca83a544e8a7ba1e257fd9bbc8a54f7ff744552345a6f8f3ec189443cd95fc1f1f9949c81e4b733a01efa835f8572892edc2b540e2825f0c2e5de086c304242f60aa16234d374b9aa1e86b140a343a10b9491626a9a568384a734acd9fdfab5e4d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h111949aa5a7c1123ac1f6d1616b0cd891bc598b4c3eef0268b34f78970e8aae1d3faa54f80397795535a31d5ea7bd66e0c4898caead2901c93c536fe49043dd789a98931ea1a4474f21e3bc54be1503b55300af10ac8b86829f831a714d7492ddd4f4b21feb55aab5af6482be14a374b369c6d5a179e255c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h165028df9104486a3c5c76b7f6d25f28119ebc669b934d870e4f9ef225a0d369a962acf0c64c17f8c5fade7906746f52c5bae890f97f15175fb7316544959803b5390cc95838fe59bb34b486248bd41a87aaeab92b1317ab05de6b1c23ae0340184d79dc947154348be5551cce429e9ce126674933402b92b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4ac856a3c83526336e91ead3d765b85b46612a8bd078e498ca2e66d15f12e98c158846e05db5893c22cd7d9664c79ca8097752954a8811ba99ef24b148cf61b6d0d834689916cc289fc1b4b05e3d0a2f81c894b8eeb8512a30b1e4344b6e6cd3b3da369817e61b985cb000111ccfaaa04eee7f24f3b4dd15;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a293a3ae446067ba0957454b5fffc24fe7af2afd7b08c41efb96927b600378824a7efef51a6903bc8d67b90135751205e40413f6085d6d0f8aba2b7b8567f0dde4ddab62e799f08024d7b4d5aa339b5f7091d7b3f8b42bc5dc661818e9ce0c91bb878c6ce4205602c5f10e066f2933f292a08886a407cefe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bebc428cd73641d758730d86a9e1230ac89ccd79e6625557a5cacc858a4b9c2afa9b2af91c64763f7f0d8836e7a924b9d53074cfaff4cbb26a295a213786282e498c72638c08e3b7f1739f1f565e5dc179f77c775118acf447593273992e9ef5ff594c873b5a8c5a61def0293b3ab0c858d490da920834ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha670ca5cbd8c72c74c57f9a7a32fb3558c48528528b8638be37c73b566472874a4aa1c8c2a01b2dcb3a02facceb50f0507ea06e794829117be44d776ba7fb37236a31fb9eefa82217ae5cc0e277e441f7cf139bdb22103e6b5670d2c7f3f93aebec0ec60a4e4b07d5a817c7ef8054f006804f13175110d2e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h103a2f6609eba64ea11d452bb1ce2dbf6324c458fd26d3eb56bae963f8bddf4dfe85b6ae5b10ed3147a73e1791d93ccd4f083481f99436a4e4fbbb3b401a0fd078adb15770156931448a46ef5b250c2f859dde41919e2ae37a637bbaab7e9c31545216512ebf63022f9849c4e4955990f9014cc3c0145e5b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bcff6d84994b1fbd745d1b7723a776810a811b4ba589d0c5a0e97f18592df938b650d601395a5c3e3a1743f3cbb76f5be736e19f5eacf60bd589c2834787274070d631e2351126874ff3d826f72be606142685a331d8b669fa134a5951d26f786d648d5664656ac3eb8a3ec0581451b94ab4f12cda3fa471;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1788fe62b9d31f5d317d7a145838db79e6346b97fde54f16cfb60b9415c3ce9c38ae0ec052d3cf87c76abfc993af8d79bb1ae6c7c9ac94a49cae32493769255393a3113872572c881ceecd1e5ea4f4c5cb272074ba053dca66260527fdf49d1ca1f3738c7476c3d28e3bb6dc1df79c8c9017998ccd67ba250;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b6af29794d2fbbcd50cc33181f4eb21b3a535b7d98ebf14268f390039bcd933c294e10b47875c388d692b4388ac3bc437e7d3b80e5913234e5b8ab14e66cdbb7dc4e124214d5c0e0f9bfc536725d72057cba8cefb6d0022038eb2f20828d891a40b6a39a830212b572c677e778a655e77b04135cff615129;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc502343842da4a8c825d879f2e473b86fa3dcdf022babe41b70b96cd55f0c11ddb8ba68525115124d6e5c9353d4441c8877ef0b3306bf5dbbfc522fa0003ac2df7e9beaf57dabdad922e6a2163c9fcd7c2b9390d43ecdec4b88254b9f764c74cc70faa95de3a7bec773a7cabf33ecea7537fd83cd3b864d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h723a0cf42469820cce89cb62fe1f828f0492f772ff846c1d4ff38d6521851dc034cb139ec05150af33218bf669618241b14b8d64265ce996c41f22c195769434159951d0e9395cc454982c991dbe14c59cde1ff42e1f81d6d4d39c2728273c5e54303ef35a4ad01f205805bf931b41870961f4bf82403685;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6d37dcf59b4f064a2f2adc87a8060523401f8791ae5c2940f1e2270c3580bc98a01e15da1f36d9b447a724cfb2f25a986f6c85a1fa18a6f9bcf5a53c016c2e37514518fc01b23f7c5361a9e3cd65829e43abd87487955239cf81c5ed64650f814d6a697f2db330310202e185a8353c1c6cfe2dc75be284c8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da2c884afefcc32ee52671aa2818f800651c9bf6498ebebcc6051a3cfafeecd92523d7ad588f0106fa901b563682561b527a239c9535121628bdb03664646597b8ca0d5f34d2270eb05eff138ccec2b251fa987cdeb3a6d7fa5ecfde2ca0a3b0a94d7866a99bebfb4952a42ce337e3bc76b045434d2ec027;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb03d0e0c40479d100fd816bad404d137815a80ca11d2c721907126880cb87afaeae939bd4817073f08cf17af36de4ec79547db12ca01d43ac113411bc559f53f543ec7674d0aa52cbbafd2e6c918e275a958aa4d893528a3e2d0dafdaf27414df167d6472544dcfb75bcea4129daf3b0f5da06c04fa23175;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16045fc98f2139dca38ea0579c2770259af0276600019db71c0fca499161f2a1d9458cc32ea3bf9a6c7c4a38fdebe1e2bd7b268b8176dddc9c38bfbfac3d6479ebf195d816dc53e1b438c30ddac0301a666c7cee6d945f0fb5e32b3c9960ebbc8a4360dd93a952157c9af72f695023c27b478cf4512e85e1b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h596cd90451f760a007693ac83d5b7d302fe9dcac7fa1e9af96967e550132bc12e52b408f0b891be94bdeed21b1ac11e21a8390f14fb2cd8c8eb3a086dd5a47883f427dfc013194af3884b6489090e99240e9e1d52dac0f0a1de27d5d15359da6efa7d28674a07db9950add8620e3173e7ee72355bb06dce2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b1202d0a47e158d518ca9cffb8451494748d015f9e4b518a6ae4747f8707aed876400621cfde860ed394dfb332b80189d6523d5f6d0bf353d5b741090d00852ab3b552da3f3a0f4c166771836cae3490170584e284a339370c2411239540d25a19537f3925a6e92d6fc592e4a7da99358238b8212a773816;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16004399e8274ff543c786fdfe77ea1bffee4991f0a49426bd183d2b9f244ed5b566245293f4b1af56aceb890be4cfb978d53574c4b3182b1ea59309132d3d596dea6d882285881161d3680c5f150db95e52acd30fabeb374b1acc5e0577e6172a46aa92f5ae2d236c653c68eb99f04ce49e89909a97701b7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3348701307b09e24debe3d42af5660ff619656b0de3481e989e9ac98250e1eeb703dc5414b4bdb37b927bb823358d3f4f5a1ea52aeab137e967242f1b95d8248dcbc19e682d7fe398978227314b9c8cf132f57db261524c16ca8a4eab7bb9aa3812d2a045c42382650e4946149f760cd0a3fe06d8498797e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1328e5d3525e3cc737dda3b0606b53229d7e9f689487ad00f6d877572500b9fce9efc57fd101d2aff4c3d1f58ffa020cc60a1b9fe339db8327af8120b94a1fe1c3145d9a9d97e63a54a52164b1eed7fbdfe45b63e26cbd4e2a3816fd7e65a27220f13b7b93dd0194a058f5f8e4e67dbd7eba32e3ab0639809;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d38d613ebb15ea8509ca3cc3f4858fda22b2278e5d877cd9cb0d33c2bf9d680930da5d67074a510a188d125ff0706c2f00e9429fb62ff749726e17e6ba78e3c703e74fc4668f39d58884f7dcdd70b4e53330d2abf663246754a7169510c592a97ecea970e8fce55ccd25850607a485f4c583de96ed77826f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha1f9cbd9f55918ff76da2520d207392e8c30354c827a4a1866d74968503af45a2645bac06d2bdcf1f3b2462794f82079125b21670bd392e48bec10e2b09475dcc9227679d53f8fbd8c6a443ad6aa170ebbea42d76b7a6f6e03db79f99046dd5c83e5daacfa9076ddeace763b729cd3a5a9a76b6ba3409218;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h198dc63caf57b26016fae0be86241ca6f064c04b4e6e69ea31d40a08d424efd50a7eb540d52e5d2356aaba9a69ed2688f0b0dd70c46949595bfe9d56f750d16d9f201dd1331d8e8c73640053efda960509423a54ce1329eb62f82183e6a28d39512b18ffeea07eaf1f5d6d4181b366b88aab04f9a193bd50a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1831ec1d784a6775ec51638353120e929663a20b1eab0ce2419466801d63531e07597f787828363a0414b00f996bd43c27c54ec7856f828f7bdadecc0a3e27d072d80611f3d4da37164a58529f1d6aa3783686363b15918884cd446248a14151703ec0f4cecf9319dabb81c272e7e1e55e41a85ca8e8ce9bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ff2601bf9401b2d22a55ee6382a7082d3157652fd5d124d052088688455eead06e07cb42bae93fae5ebed8919b007b5bf23f600a46aceb69baad29ea8882a07035a27094674f14d1a6255995d37ef1b82b9310305caa06bc301f79e397d18389d04ccef3a6468f8f406eb1ef18999624ea86b408c5b2282;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bca2002617040c8d3123b3c2591241de1fdc5eaea90b60408bfd109990f235ef8e47446c9a6a6d053b085ece1a780356e26a70f1a9b571a9e14b4688d77f8e6b02f8678709531209ac3ee7f65b69c40b70d357847344efc9b63369078d986f733bbd9ea821f08ee2633e3e85e6329e4daf740caf649cd011;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc7137eaa19a53192f328dc17e44d82c6318a276799453126dd83ca5ee23bc9b801ae7a4c47ef4617aa871350af35be5a9bd44b6cf7daebc8af6a0e3cb35d6dcd223ea6d49d44d48421ae36c2583fa460bf1e45372f0cbcffbf2a39f4607c756df1fc0ec86730d08e6fd7ad06686f15c27f47f5f56de2333;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137967da10fa5131bf05c52a7e2e71bb7bb7f68fde5f861b3358e9daa68707774c5c771705853aef9de2c073dd2110df5ab99844934af12604ee6e5f5de23258cdff0e7346035656d480b11682cd8466d09d6d98a04659258b91216e029001d1a2bf16fac343c9aa20d00d983827b5c75b87a2ce3f196e623;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14968cb37ce525ec73802319521b269f1d084950261fbfd26ee8166c152a8e973ccd857c9b9b8c0913ae35e6f305cda63aebaa086b919aaacb4d9ef3efd76a31fb5e6953806175d786c4aff1017cfc667cca10b402f7a0d63c5f057c652ef28b003d036217208b225f4832806d8e2cf6cff2ac51ceeeafd59;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h360d8ba575617f772fdb3acc85401985999dbae20ff662cfa9331ada9e30d201001c6589422ccb5e9576f1dbad5741b43d41194a412547f4cfbc958157d49e50fac1f387589f212cfa0bb984f13a91ee9d6109e5a687c391019764a4a0fe38a7cb3967cf39165879330ab2efcc5e0ff09c6418eab78d75fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f8547c01cf63f7f80d2428d8a37026769c6811a2bf8c361a0d1376dd279de531265e69a65d119440813209c9cca3ef41f802d6b0e4a97901cb4c93855628fbf8e5d8c79a3aef6b519b2feac149c43fe724adfb78471273df3d15b0dc1351c33d9e8361fdde76906fee5580c42ada759e93588314cb179bd9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h101844f0c38eb9df19ef460cc7997a6ce94cb6d75f2af3d58bff4b86011e993cd4b8b8dd4f692ab409be96f0a33bf54fe55c858945391180a136af4157ed6f659d152e6488e83583b3ca33bfc817a540d2c83e12033d45fe1fdb4d83f80c228b8f567140edf290cd6bc6d9e346fb7723db211b72151c8a0d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17b8e555a6be609a6acbf71301fe684d8c8b567e4444d32c5eb74d66bd96860d25f1187801e30f36a2e0d4d9bf4c90efbea4d48b3d9107e23e321cc52ba500a57f97bc92e53d0dafdd3c7f38ffbba6a546889f08e7a1d2f3e42708de24b1bba3fee287d03caafb1324f272cd652e908ddf2de7dc6b2c61d49;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d515c3791769a8ec78c5798caa9449a6d4d8fa5faa290909d0012b6c273539fbbaefbd8ed3c71991c15c79a93d94c46ba98e378c95d6ea6318479eddd499899d77c1284966c5de4cc8893a0f4c79f4caacade8dbd19cf85a467ffe216b2f20d57a8f5c137b0bed21a750fd20572d983d971d239d9accf48d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc04bc220a271b8191e5c2309c4070404deba2c3e212caa3f53e53c4f82a73a3670f9037913184f3f43a50f569521d86cefdb7eaa6f913121b1021d928ba75be23132edc04a246ffb114f2f8e29fef9b7156fa9a71d955926d151fb041d5db7407594814f3d563d189d1cdb748d9cce141ba6deb70157a3d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8bedf7cf13f90c4b6d6c407e67d61de3ac32dee81b3a91ea9baee41e7e07d4a968a8d8d240c50481c6a5260b891de1eedd52cbacb5a5959f45968a749e9f56ea58e863a1c2998be12b9b72a07b2ad76da076292a70ac7a08efe990617da4566e6bc9f5df1018395461ced58bb3a64d25a28eb223e58c6519;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f761e4b0f241076d599f332cd0a90f4efc914545a4ca8a9955194a48b939e6566987c497993b06d2cdd5cc10c0a4fe2865973cd4653c7ec14a910a4ca26dd7e9d9aa7120cd0134905d052fbfd99384323f4c303c880b046b04a8e22bd2d4488b6a3290eb6d8555c0725a0930f77e670f325d5ba7f1bcffd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h348817d3f3d9bf0a411c683dedd64994232057ae2cccf2785d9833dc86d8bc569b51edf15eeeefad26ea5a2386c8c09e38c94960edadd3180f03ac13f09bd75edda14c7fb6a0f0e462a47917006596c8d04f65cb5c66d2c43b76a17dcf88fcb7795bdbe07ddf1969728e96ca19a9dcc5b002bd4a2f5206e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b2b385f309fbf23eacce20238cdaadb8774519c7cd955085ea261a7778eea72c688929dbe4599a1855e6aa53289937d1847ef4a9149b792b5f459af923f493839cf8ae4e5a48cee8177f7685d034b9278130defbb110795f8a9257584d4c6b889c93edd22e05bc3341e018be73393cb0efd300256c86b45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1777a79bd314c96ce8fe4b04ae058c0fdf38ee79f3aafdd84248b8f3e54dd50407350a6b4b4b10fd6b32dcf85bbcf0e4f1abdb1fe55197f9085c2f82c165dfb08f447bac4db26c813c9145c0e17ac7348d4ddf5e224eec38699e708d23e5a22e5c31a33634066a6c493fa3b969421cbc4b93ecae22c353060;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h268f7aabdc14b0069a2e3d01be3b5a8084db33c36e5e506aebbe3561b17a9f2cdb39b6b279dd94ef811a49d18020f91b480f593b1bbb0ad7d843f8b9fea357f2607385afde09ea1f5ef6e198444447052ea65132aa4b853831c009b13e2b7801863f8af21fab834b075a2abfe3d4f1225299ee75790f4261;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11b9ab05488a67058c73af28d8186838050356807cee64337486e1c1fcf06ef6ecf743648ee038df6d3b006c29da131a971d7bfd04b369e9cb4d59aee88897a177ae5af3688640893e64939ce27f0950177a76558bf596090552e159022d11b9fa129b1f49be6fd2b487cdfb45e773ae1b25bc4f519328a04;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcf610f2c764acc15f88ba72c4f975e8be4066ed2c5b4ef2aef1bbf6a8f896eb170865fe5ba70376000ce719c90e8affd26710f7cec9858bc490b32c1a9897bd7f424cfb3a02e3063f04f959439d5000c7c945c1aacc4ddaae593c149327ebc95f94cb9859645b7a81daf778e202c68fa3965f4a542b9c8aa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104be100f43ac8c27a73abc7dcf2a03379247dacd7591bd20f3dd0f3969f7c8700853195fab79b7615facc47ae841c6fb45ab889448cd66f26243b67029704a76c5337e39b4185f655ae0dffc2d270ad19ed88c5de8394d65239f4600097d54e44c72cadde1db02e5d0bb0d9dfc48f99e4fa458b96eb02b2b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c9c19a2447a3642a5c62085d9d2f6102574f415cd266efef5a3fc76814a7612d25426e9a2065eb3d71da0956b26fc82642dd4e982e70fc83f1c675455cf951d5306dea20a9ca4b97bff9ef3e499d5d758db1a2299d1ffe00600e4f6a578d98d2ee4e80b1ae5201edee325ae4c6a7cca130b5d52e4c5d8210;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6d760ab8a55c0fa3567c5038010fc58b15ad04edacf1d273a3ccb5e95683d3b9eb78b249d2a23b4cb5ad65cafd15961b849750713838135208f0b520bda29ab91e0493ed2f1ac22e49284aee6672d76c02e988a070acf892380e202cede3efef6b21b8861ac73cba0eee7a562aa4a532e6ec770ed6ebb645;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16075899f736cb044491d43cfb8c4fe979303ef032dc149b0211052830f1a54db22dfa74a17088b1b3b9995ff72b41ed1d142f08e06299879e8ec4cd5fb42cf4f6961473ab97c95b15e12b695c6687fc4335296897859aa1246341a297818c91181c6aaeaf5aa670ba3021ee99676cd46ba362d356ec11957;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1880a0dcbb3acc51fb4226d28468020f0bb4e3b9c97cf061194df91b2b1fa2e95d42f760eb824055116114f6afaca7c748d6d53d40f57ddb377d8b0699a74af10eaf885df25de1661ca01c9feb6fb819279acb6c77f683e566f49b38a2a3b84f26252f6b94013adc4c1106943a7fb106bbb2b37fdfcabc0f3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ac747ecc80326a57fc1ecefd900e75b4edbb74b4732ec7c1deaef88225e14b68ab67b4d96803e96652183af341dc39f07f91f97cb4d1ff061bf1491f9a2a7aae94795c8b4bffb97555ac484f441d4379ba7068d1926dd6198d01c81045c6168531d7d7464994d8829864147349c75f720227caf064f35a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c6ce2eda21217b4789630a0cb0a6317beacb807f1c7fd284fac7f68545041faec45cc330474e6d0d275eb5b4282c4feebc177c23da995cd6548efeb002a43736ab66765c29a1b54ff8b236396b1de5732c2c7ae3600325b2aa432e4dc1750d0ec33d3ca7ba68621a51baa2290ec51d6d395431c8de9d4938;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h110c69ead24b7d45559d0dc2369e58d63c9a0152e37c8a9343befcd944e519f123b0c32688ba19ecdb6dbec7b195e3ef77d0fde713e22a48b66e0c72ca3c32b80a8b0fe0c40177e0fd3eef638c85465cc833ee3da84b611f0b8ce4e8c9c795883a2703384355bdf2dd76df47668583ce18e40707edc7bc996;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf4965db5e53504a2f1dc121bd3dcd48e495a6da0710910642760120ea1df933f6d3ef412ebf32da0dc131fac850d904e9fb86a2ce0f236d403502f8456f73d7efa7309aed363945b8f8a9011d2c91e3d4a04350696ade12ad264f5442654e7fa6dd5863a5cbbbeec2a2e46a72d8b0827e4522eb71cce2c30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19010eb0ff1f1ebedf651592b7e366352b810f7a3f4a1e163619f7cfa20b1e600c8e54e153182eb5f7b3cee7883b409490de7b1c7dd4fa7b7314471a02338cb6c910fda231a7874ccf3529a01a3f7798c980b2186e2cfc3b2e3f5a820bc225d7f59fd64b396c3c611f98cd08bbe669101afe25f20a14c971c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1761f297ef25947ad04df3c7a6305dc18250f3859b75ee0a387c314dfe2abac77b9772c1dba9855a962be11551fc066c7cde65ef5c8c323c75a3f8b7318586a9c064de2002d7b95ae09328b3ca65e387816e192b2b076cd3a78d0ca192b830539f45fef948073729ac04fff69b3ba6ee2230bf1e07c5aafaa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he1f27d2e7ebe05ffa7f1ad01f5b222d075bd4c6fbb5157d583ce57856c181901aeb6b23ec20e4da259b177d523d5fadd54e9c491d752c8b454778d952d9b2c968799318a12773bc7378685059bd0566460d926cb122c07007330d94b98fae885044411ff815815bd77181cefb94cf52ce16bc101db67e6b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e3e839dfb109c267caf3232d109b871224f749b68f02ee17b38680e088abc9a24cbbcab83311391c007a4a2882d88be28b212d19f5bc331b7bcc694c6588e10537e5fa48699bcce1b1fa28d837bcda7e067f36794d308503635dfdd51c5574a7906faabe26de027c7718b246d832e056a931c9482a62b13;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11d6bd4e1704fa6679eb5ea2570cfb1f1c5cb7a1723ed0084945a5120063f08616388ade50dbd010c8393066c06196da41bdce455582faaa4ccb095a8e1d11b23496db211b704c12daecad3b30f059b27821875c951679ab0c477f15d50d464c9183b4bf9fc5e768eda1728fddf42dc5e653da18a32a40b49;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13028d2030426aeccd60795e1b2eb959cba9b2a1b1153b7188a198f9316367dc74b733361e727f4d339e32cec00629210e9292999dab9d9800ef83fac2c9c3b5c4803706f36cc5965f8d667a6fb34ba58af9da86e3db6f7b38c983d43a9976c5feb3d13d56e05985cc7917bf26a094c325c9e9e19090f5cb5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3c780b7b3f46247242dc7a595cb115a3bda87560a41152d280aab3b9fa8fc61fa4375ed10301b7dc5bbf8d683d225da52767bc8540984375843e8b8cb9803d5a1a3fb83c9efc782fbbdc85c335e10aec4df80c0aeb2d0dd524dbe3a2e494d701c977210801bb6a7c575e90bfef423fb2b0e095c556b8daf6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e9228d4aa5bae4e658833414b1bb43a1015eb3d1eb7138bac5495436e17f6083c40090f6b3b1827729669baa5f2f8f03781fa417578804e02f3c7e9e256d7d00118b331372a5596b19dc9e7185ac67ba3c3afce0590180abd515761b532e4e3a8e451d367ceb4d89c22c1bbeb72a0ac98ab80f6640fdd68b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1957f119282c3364dec4c71cef3fa612d05a244f9696f85c21a236c850fff888439a3c130188be8e005045837da87255929c424654c939072d3521b8b2b9a0e80f31d5c310b6a832efb9c431254fbd239e70aa3ebd865ab05b7cb2f729dc86ac7c7ee628370ee9446b0303830091974956e22e8c768517497;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb8fee775a543d69bfa0d89dfa75b8f96e30a268886f4b83238a848d318f8d30189dbe0815c6b9a84350fec1419972c94c41148be8249c301f55643a9d90b85441f56abe814de2b69b7076ac0178e69d2a52a093448be127b607f154eb7c530ade693fd474f3720f9e657e2c11c2e84718c4d4467cbd12bb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ac70f12b7600f9e7ae5af134cb56d91c34bf97205b5ca4c5521f7f2d9d46dd8995218f4bbf8b7ef2a6858213ae303b0b8e13c8185e8f44cad3921ca6485b1084ad1e8d298901160771474403fbabe6f02b0809010deff036c0bdcc0aff897f9e12a07f6c61ba3af24f02540f8621c12a1ef0762adbab804;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3b7782ae7e74c83e41cf6da5f3f4633a7bcea3ab3336c6cbe54f8055e8abfa55efdb1f88c822d04ba93c7cbf1102d083454a66033022f6a95a6ae40d9815ad38e1df30cf9f91e39cce09e027c351a58e24044779cc0582b9f50d82bdd58a377558171f21a11ea2d4c42387d47eb7d7881df21aef2699fdc6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heefe88104632bc70e60ecdf08fb07e93cb896ee1e8ec75982d0f52127aa15dcddf124762e49a3a5602e9a46934d59954832bc940612ed9ca101f1482bb816438edbc70e650d5dad993c0180dee77a836af442dfdbab863e0e645f4e865b465a5edf1870411a6d831d7f322cc537b14ecdb6b9836431a6f84;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e586d5df5cc41ff2f769cb295888b8e7f8cfb944ac37a2e12cb53fd8fb7c4b098fd1a71afeecb8849556fe097512ced6d97dc3d77fa902b2b43a2acbc6ccb0b285cd29290a27a70c08a7d45c8691d7c35100842e7959d399d3ca2e18b23a1e9bbb81947ffd967d83fecd29939f05cb163ef5ebdcd36445fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12537b6b8146d3fd32426479a4578425586effc2d49213117ec0ae0a51f64235e40eaa08efa0d444bd43b43cd3a2cb9efaa6d582ea25f13d853b5d3235beeea6a1134c7c0b58394c3d243298aa82ee90a1dc1570d6b504f1748461f22d810a85220c318562d13f742b8051d5d5af829da209d871ce3d4cf60;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa416bf7a9df024d43895920bb7d162878e06604c0e7a76436fa762dae7e79754ddb282cef46bf5eecb40069488ad1e94c59ae40f932a0cdbecb7e74e1744f190326961ece4caefe1f59d7e938519f1b8a6a9294b28c1dcc9d775aaa8448a373c52041d2392b2b5a716c35fddbcc1c0532bcb40d0a7b9121;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a015870570bb6eedb0491a263c7a8f909248118805257c2eb5e0e014f99bca3f8d6497615bb9446a62124d6ff12d20158fc5da66dd170c4259222086a8de4b42615624527e2829b9ed7264899915087dda4803cb3d063b161a6d155cb9e0969dc4ea59431fe51c20119a9005200a1d4400f824da099ec37;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b0f5da167816858844d2b0befc15109956f5e0fc26b4c46d7ef2146bac0c0d3f1aefef4878469babf123143e1822606ae425015b0195774571bf28c7876631a17d5cf4335d01613db8be157d4df163a34f66940d2dcc9949c2f1559aedcf230d36eafa7994d577874130c188a3fa4c1549cbebfe7167377d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fea53d8cbd11e7731bf248e030e7187e2e3e41c3a9b821ae69703bb077fa119e7362a5b2a2424c379b1d3b87709c6e1c76df025af91ea868fb6681254cc5affd296215f660450ccfc07cae5a4992f8165267114fcf36f30d40ff36157a8cb6fbc4ec875efbe7123eca864636e2bc236c096307fd593d45ff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128cada6bb8e77669f9eb054393d156c19c7efd3dcdccd0eca5099f9285c69ecb10e5b36643018fad3ba1dbf63dbd0ef6bfe8a41134dda81eaf8c0ccf89f01d8ed164ec1ea8d13588fb795a68a65b1c1f2ad999efe22308a68929b57b9d738b0178a96aee9ad283607d6779bad13a93d1a4d14f3b0e54c961;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha9f73f319a239eec6755994438c352bc5285c2d41b4bfc245708c74a1a488a27eb2034a700189e4ba7c6deea479ca25a69653d09421a39d8940b40e88cc4b25a1ed552d6fb58e1445ed1e7b1592f7d00138795542ecd78a9cf41153a48f80268b8f6652f7eb9be61de9b0b0a591d570ac08a72c64426eb18;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h195fff03bb7fd6279a7eecf216265ccee83a5be888eac78c3fc49e3e03bd65b80c299c25be601df0dad1151654a6c88e7ba101760313938d42d425bed040a4bbbf82e4ca0a058722d968a45e2ee9037bbf9b838dab77df2abe44af5b193399ebc90f756c384e1daf6934fc679ac8f6d5714e1aabef15fec30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ecd8998b706e1811f57a5cefc612e0d71bdecf8c0747726e06109e903592ca6e4a67f6c992c56fdf922347b2b82988290a922c0612c20bebc7e0af8de861855e3305be103554aa14b94a06780bd9323d337ba2bc2607de97b5b4ad4caeb6ccbed1887c2cf58cf8c7d0c0e6aac179349b758aa5b9dd80904;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16840f8b59990558db56cf828a06cf3ddfe3f4047fc03b49c88474f37c3fcd6b2a3324fa589a04e7555d0df51a18945e08f8e71423a2bda995041ea8f5710e146f45bf57d12273a29936500250eac30e71ba05cf3ee39429e1dc1de409d80b7e52a94207f292fe18f8326d7ee6a84077ac8f665825562b893;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4be6e9d52f4be2f76e321491b133706d28fa3823691935122899c8997a7fb04d61a149547f724da945deef8ef385e06f7d2c5103032ddb78913a8cf1e231bbb6bf2d6cb1293be14a950c4cd13c3058543b09866ad7f3159edac14407cf82923620e05dbfc5e79c0137869c548692b2912943a5fa58490a7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbcb16a817c23a0f570b2fb846555d223acf6b608ef74ac7255e645fa20f2abe3874a1704eea2af6ad889b4e88bfbeb4f8fb6d8923914c684ae2c4d9a7e5ca4082b36d2da2b9cb03a8a813400225a68dd23a4e4a3fdc3a47d5c866f68e19cd4278d53120dc4ca3dc38359657e6da7cd6d0fd8715c2a4d5286;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h105326a25a1e8b0c90a07b6879caeaa88ae0c9e1455ed81c1e09508f9fffca95877f4dda6193b4582d91c4653564dd0105f55ef7e26c4cfb0c033e5f346715f144d3510241653a2daf55f3e7e1c10dea4967305d94d7de0b16f34d11f54b19132cc8b694f8f313c695a6a9b0a366c9f514bc8cd79e783a4fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d158615d9ba9b243705ade30e56cc2f9612a0cd8fff5c49f4ce1ab5f399f0f6b0cdcfe22871040ba25f69bd227a83202fb8cea5452815f265502a25f3468040b722703c82ec9b9f07ce64e7636297d2ecbd692e58c94b90bf22db746e5e1e36589d75c347ed2b174a15f4f15deb25eda8dc48e9a35e3ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf85ac9aeaeb0b326609cfe54e61088b01814c3430722d1c8ef2a44e73726be5344c97fbfc1860016ebd53ec28557bbad9ea2977dd51d8392b7b68df2e3ec6edeb0450166f2acb5c642fc8d41d78f1f3e28fa1e3ee9f8ea54612313baaacac5dc76839fb5f2eef785041ce2a19c73a8f2f62a2a82e611c38;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b46f8c08d059e4ddbc7d66d45e27e55834bd3fe4d5396b9a2b1c221441a5bc97f4081b95f4ab710e47cec927ba88d297564bf85281e97ed3510bcf2d2ec80eafd4ed9effbf7d53267c237e9c325d30b2d472b1f964ac21314f8b04c405b4afd67151b045ade5807bfefd023e178fdeed551156d62461065f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a94900491ebdc11f7da0f27136df57bb4e188d63fdb24f13450a6c4de9548256aa9c3d102131c30dad2e9f689c07cbd31526ffee769b4bc938fe8a52ea70fc7b853769b8c82a255a4865e5d6c353063f2d37791206142521303632d7454c41ad4945dd887e854faf11c1ca975e498d214ca9ba5b6aed4758;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ec44fa5a1b8808b44678d940930163755c0196b8196ddb59bd99e69f8b825b413b92228a63a7c7e8e840da157ac5d2eecf83d201d147325c51d2278be370d1570c54e4064645eb4bfa6dabe17b0c01ccfd71803d19b1bcfadcf78257a0ec3946bcd2bb436d98e4643a0929a7b2bee0ff93f9695b4de22af9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c220d574cee0b9142c93e1972d426265e9dcc267d38e90fe8acf7a244800d2ce9600d3b926a0a5b62bbfaa174a783a48c344852e8b3d12e6678644a8275bd1d84f81d39ba20d97485765dac8bbe55eebe82150eb04a07428cfac0ab3ff476cd29d26e2a859c64462adb53816e7abc718254e71eddb9f127f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h192a6a2477c2624e238aaec8bdb8743e140301ca54dc1b93888d0605d8577df4f7894f98bf883c17481b7e047b599eb11f293e058b66fd6b8a147879a3bd7f2dd23888156ecb7d3db7266b251f263d0307cbccb16273312fd034acbf149359e3b847d770363823a264237cb53ec8c732a873106299e895e43;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1efbd404fe6330e5169ee495991d56c7b65a6d3fad6c5b952962ae05e559e97a6f58c853a0d1d87c0fe6b1639cb6cf0e406296adf4d526cea5d7985d193f19f3b86bf36043c0b5092f5b9c5a766436ce15eb48303d482601d57a40864744c224c046f3f4b0dbfadd2b0d4af71cdc5ffdff6e3af8f0d9b78ff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h27f6b9b679abb85342d2c58fbcf192ac7141662696bccda035c05e565621651c85f58d242c2882a139dee412a2b8a78ce227137a467a7aeef929f759cdf8ff12cff0b05581b5d4c511ab8341125b5fa2df90da9289cfde387869ad977bf3aab645e74e345e6aaf5d61b3b6e53c653bc7f66a37641d4d58a5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h154e94e5af03baa2fcfdf1ea2936135e18cb140232de39e17c386a6940ba3278cdc8f89b969d71d69184ffc672cb227fddbcbcf28574e23659a378f84afd3b884896eeb7139486f9d46040458dea936b5c65c09664d296ed584bb6c826fb8630ff4ff58f77dd040bf925525c15e64d595dd9bd3ca5464c1be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfbb449ff8005555caf32bc9d4885e846c94070de2281404b9753272a11b172351d6d51d4d6420c907d3b2870586366ef414793d7198ef2110958c608b8ada95e45b0af2ae57fd0fd9a39726d9c8622228b1c8b7e1a395fbbea76a5cf8fbf3d70d85101a61bcb2047afb270686dc76de0f4b7e5e271cd06e9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146ba64dda2e7097d267f906870d29ba94ef9e299b9bde4a83f2efbe0f05a97806461457d044ac126c79b74e3d437b45fa4753725899183928b8252278d0e2ae1ee99438f7c171b381d82cbbda659a617a6b74f27e19b9059bc8133cd39dd4e10d251b002e9448a075fe0939378cefe73b209405673fb8c21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h605bf8a112828021c69e1a78b130881015d0f4a0893ef4264d51c89d120977ef24de231170757d5fe833a7f732a2641756931f53be567d2c59786d576fddfcdec52462faca5911930e562b172d33faa4a05481b9d07d1884c5124d2dc45d33d9ec1f8d5f707e9082e4b0f0c38a68844384ef16dba3cbd97a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a880924b9cb7629190f54890cca31715e78a2eb4954a9e06e95a7b63cd3ce49c3de48b95fd49d1963d2c24fe8ba54dfb7747d2d39ac5d4271098efe7edbe3dfb8b4179751298744ae46fe424713dd867b6ebbc406235ac379b518cc2b5eac7b5805668a4573650d50ea5adbb1abc393a35f424557aabc0c5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf196ecfda93a5631d5522189d5aa0d584f508b88c0bdcc0c7a307e63da8367d10eee389f56bf92db0dee8524c93a45d5466ab775b4430d2e059c0020cb5c30c36c882f2ca0266e13ff14b92a1eb669a22e39782162bbe2f05ddac0c4808c684110cc368efb8bcf80080e31e13643360fbbf3ee2fb4e09289;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10ffa57bd298069e41d9c7cd43b45bc776b9927a12af33b9d1d4cc4dad330cdd93e308dde28ef6245b0a7dc300502a8deefd141c88bd7bc4f66275f9aa18aab3ad8d7d255f64ec748b8fcca96d09e8ff5092b9f100c14859a71fcf93225accb1dae4bdcb061e0b23293b998decbc6e1fda8b39c80664226cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4b93fefddfaef1c4836c9bdb8063b4e8186107ed510720cafc26fa0429ec43265b3226fa31e60d080063eeb742851f6de5f3261ec08ac7bc2d10715aaf473401ededf4fd84469978d61fac73b18832545eb63bbc1c7055415666afc4b046f44a3a6ff765699a773ee217e5e6b9c4372166ee91f017b293a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h144672a45d37365312fdd295212285ae0e38db5232100acb95494bd5e44357417902964110596328aa41fb76f0adf2bdaa51688003ff1568fd23748ed23b16e2930c056779438234fec5db6088d8a808ea77973e32986770a011ddc5c0e5091f0b06a164ab957faefe37a4b7f3def4dde1aa1b724805464fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hab031f32661067e89d39856aa54d6afda35651500b6df2bcdd2a47759c7d8a0d2c2cdc8d5742e7f0061cac6b68210b2afbb55d41dd1dc24da20eea49efb373bd8c10286a0e539c30357098744b496826f44bced3c9c72931227185e0331efb0511abfadbd3761dc694006d0f573ade85d2bf36d42b365b05;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de4fb001520683cf5d3339da99826989906ceed0031d96c40862fe14e48fed0c7868b285579881801a41d1e1e78e92d99b58327378bce1b2fc45eb576a328df36f146dfc7b1234f5b1a2e7a76976aec57aff71205b1b71c9835ed93ab17b2f70e8ab7357a75116c79a843d951e74fbedc8a6aadc97cde291;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2d189df54b07cd08a6129f2d5a29f561aee348692501e4b54697aa123e98228a8c7859a2d722c6b3ef699a2f92bc79a0a8a79ed3cd1af4358b16e51da75f33ebd3b11ec8fd9a1b80693f07ff7098904e45ce2ae1e069938836b49bd16e80c432e4338e8c46c58012d383fe256cd73238b0a297c74d1e2978;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f28faa99cc3ed72db6a66dd1eec86b03f1dfff5365d16a4295c81355d9ae5e868967cf4e6fd2d39d53d17268ae04cbf490b1eca88baa9db9920ec310d408c04c5d5bb1c5044883323c0f474eeb9abb5941e2e51c80366da8ac2c455ea32e02358847e7ee919f53062d574635db78b96d6fd232e23919c62c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h321913d03e3976c67ca5f535e37048a74f6698b66f0bc2adb9df2783b9607a347e42af224e5adefb7ac285e9a5c4b5a653e33271a23d44fb260d28efd46ef2605eaa2028ee0e8f1f2fe660b5559a35b445b584ded0fa277a4a7c25fe9c7603781fc6d658c275e1c942b662a3cbb61ad8150625002648df84;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146016c2b8644ce48cdc87e69da8409cb427ecd22467f159ecf9a0ff3676ef1ce0a6b200389349f46008c399f503629a691f7fd33040a0ae5b70f78fbe748196b2e8b5a6e49ddd6ab44cd79466b95a24ff7d8c547456ad02dbbaa2b6c4ff95488fc6be81a41912568af9061609eaaa4a31cf9ab9a7577cfee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147c50350d801c4142164ca2d02ddd69d1117d1b2d7c6f61c2beee278e510659afacb8a70b5150623c38417a80c13c0210d6a2bf4ce762b34ee64556942927500cc143ef6621914e1919b8175cde4f342c5ca540bd1dfc0d22d2dd516d051220856838e011aec5edebe13cc7b745854f67be3ad87e851dfd5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfb9a6fc04223a2e4c146747b4b332172dba1e8fa7223531dc019b39d83f20d1f116128a7496f2e2d3964035ffa21c79acbddb127bbc4ce1a8ccafd1f783420f30912e1e8f83b5867a4edd45b13c13d29d00b75cad905d78b3694df4ea7560012a0479a37e73bd41abe340629b84b72dca65f64bdf83a916e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14dc2c0574c77dd1eee7fc0c3541ef8a2a85842ed1f5ab6609f53de8a27321c9115bdbb618d1af72d77a4687c2c3dd5e25a15633ebc53351c6fe3a793e90615b865bafaa6f960806f0d73873c29396914bc54ddf6daee01d004b6963ecdb43d009566756113b19d82a70b65d90458f6f060787a1fbe311d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he7362e1e14de22650f8ff4a24d3fc9ce186d503e41adff6ce8fb1170085ac6e260b47b2e709ae3f038139a1c11343a8660741f0463468bba2a6244e2bc17061efc6b3e692fb1f4693437d3971d78f5b4300953d824ee9b47bc1becf744ad34d9e9a8108ae8fb550c5d16ace68ec6524f63ec44b8d92c626f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b034b021271f8f4bbb5a61a03fe0974914b6ffab30366f46eba4925bb59277237745e9f9157971c97f40ac656a745b09c270e35f42d2db17c5bb28acd54ecf67271f089c89e482a4e7e7605451d31d7118c15086aaf2ffeb8ed7fdbd5c5d27baa6a66c8da572ebc2ff2042b2ec900bc57cd6a72315a88da2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h150155d39456477537e4b5f51bb557dafbed42af40a3c8f4cba2c4580c0a8dee76c14f28ed4b5c59548b0eb15d0fa5b3913315b5aa822c83b5279c62212f3234710e7a84d9b00a79108ecfa65537b76a7deb4e261f25dcacde6cfa9868363911e751a8eee9c988cab8e5f6920f6e44d2603b48c936c72cd40;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ad3d121c277aaeba61e8a197636ede24ced4f4993a154dddbf1efdb401856b5ca2d3ec5162f69e93a6d37af7c3626798550a48c52c1b6a466470057815c6ff72efd95d8875b836149d753797349393df20970dcff7b0f2587e148d97f913b7b7862f461ef47b7b84b1185234dcd8d012368926dd1966aa9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h245e8fd64c7c18b23385c1d99c91b442e35030839fdb434b2367d44c750b281e050007969fc9befeb022200083850e1c11d1c40f5fcecae584121e15746874e62f6ab6641c3eb066b27030a24166e6a859d63c66d5e1deaf903974599daa15fd9b9b6669feaa021acdf7f5612283c724bbd82a7cdd414563;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a325d066a1315b9cc3a98b295b94d02e87b6a10309cbe88d7d229593ba2e6ac941f45abce28aaae5e26e70740b283bd702a991fe77ba8511be35f0cb7c9a1c543a13eb4f1ea04f78b9c6713271160914f606935f35f528dddc56188ac8417487b894fecbcea529e826692e9b8670ae743803a463ee9cc5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd7906e04bce3b3b2d8624ec0cddc17ce55a21bb0b6bf153e72e1b64693168e5b08ccb615319a64d5a9a538791ca2047dfeda6b965b3cda9b7f07e756b87ce068ea7f3a264761557500843bb80fbb611409b86081a82de2dec5f7ef42e9cf72dcbae1605e9bdf19cc7f8bd8e5a6bbf35d637228dbd7977194;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13247788e901d3be374e8a414b4f669d76a891c1c757d887e338b5d81ba500e60bde57c4318139e118f7a8648599cd2779f56d0b133e2afd24af5f1b82a73cc00fd75606a021cd3ad62fa92dadf36d288de34cc2b5b6345fe7d4a85a90d5e1f956320d6658bd5312bf4b7dca6f7f95a2723bff3f522460d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d28fe899194ebd2b2f8d89b696fda77b7a65bbe6fcebd4e9d15553da574ab34e130d685b9b3c11733e706952f4efaae6ec98ee7bfdac5c88c883bb79893d3a7c89fd683adccc6690987857931006b9729f871aaab4f875c178e501a74820d216863da31b06e24026fe39813610179348616294eec63e8bb2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17b4f7d28b1d032803b6e59d3ad5fb7d799cb3ea91a115758b9a2da66ca577ce8d2a87021c06ba1fbf92e08eabf92c2c17038db3078001f6778104f2e977e87c3a4b4979fd64a0c9abd988a292b58d32834fc00f999cd6e504a5ce66780e45810f15791230edd8e63b10bbcc1583b473a3cb854d427e6c0be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hca7b63b8452f2e01fbe081b7df42d743c830e5940bc06de2a18de761a472358574f52bda704ccf1830dd706b9388df394e32af188dce9145e137caae95a32af7ac6b1232d57184bce36a8e11aa20b1a7252392e3a44e7ff265316e0580924c66b0c9a7985c72213af232915db63e7597d15cd3da01bcb51e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d9a39816bb14414d0bf074ae13a4666c2d7491c966d7b1c2e8d25a8c11804ee302c045e404760a940397ef7d2f105a4edcf3045a347cea765c50849a6585864dd117b2274b3f5b7b2f59ef800497dd2c76f4d399198e3b3aa659d2e45a3fb83775cead701514e1755d73382686cb56ba2a4a6a88dda2f9e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d03610cd0cd569357061592f248369edb92f9ccde52d79a000427b46dec22ea547075ba9a38aec779cae3a31fad21cdd39b634d273c1f6be063ed080b278916a43d97bfd6917e3fc668cd73210b227409146dbe7432139a1dc5354bb01b1422b709ea33d19c9b94b283afaf80c80eaefa78f63193e6cbfb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h172a3a18a3600f9f1096aadff5c9bd2ec1d4359a706efacc19001c02d734a7d7fc80cc19183568d3210aa2e388e2b741bf160d01515c1feb284b94076ee8bdff68cdfbce71a494266fcf02c2d76431dcc2fd5bcb0f2aeeb1abf952daf5bcaef2058682a19ee3067ebd4b1396ba957b01fcdc50f9bd9261be6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ac36d81b2e6f863cc51de0868eeba05df3df640573d001d7ee4c42a50c9523ad5010a2bbc84273225ad0723efc95a07a0ccab65f4916d7ad7fa2838fdd5b3a5516bb5d1dd10c9ef818bc672a8af1778fceab87840b2ffa05cf73fc76b5bfd355a28a513673aca36295e1425ef9e889b89c3d913565d31ea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h525463a323c28b53e03484be3633b7587801d91c43ef201053ab5204d07662ec645e62b363b76ecfc3676e721c9a4d57618eca55509648fd0d7624665e01bf61b09083644092eb4e4f272037e9045e4b5386860b9ee7093f33d67b61763fd62d73b33f47f423515a64d7fde66da7ba7ec89881f1b775b1bb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had92e73de0907804473fa9bcee2b9cca4b6ff38b54806a59e38e219f9010738eefd1c3a0d74f3afa0ddc4219d13800cba8c7aed65a5c7d4bb97041628c41ed06e8c32415be6c3843941b38838d8dec51f4d8898113bc2331ab597ad4638a62708b56ef9e2bc5eba09480afbcafa9ef9f2fcdb5b3bcc65377;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156ecd59511049f4682ed0c82d17624ebbd7c99e2559653d78d7473d1f2d45930ba5b64502a668c29f2211800eef5877972737ed5f68d213d1a7a4d4b5373db482e8d784c9ca2283a6a58d050b0af695171a981e6a7dad93a776a76e6802de531565547ea4796cdfc3744f1ee134aabbce3ce2c233de80f2a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1812f3ae8821f311716601da8352a137784a46bbbb8c3d0716e85599d299e63cad03035896005e17cfd0139c1e2b85b0bea4c4129290fdc61b31329c5cf16aed80969b570a91c5d33debba7fd184ad9ad246ea574a4d3dfe03085d7a9e19bdb67051d87fed321bb3a53f1e7242999e778cb483cba9d9b013;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe445f37d8ef293ba5910a1b9ef5a1a1e4ee53735dfeddf6f78b46e93c42c79e54653569c9973e44c52c78d947715948d036aa8369dbdee5b64420111afe32944fad6efa2b16b7ad8b494ce1ff61cffb5b9692ef41409987d6c4db57ebcced138a04c87c4ecaf0ddc16646069fd41a67b5a019356e30d392;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12189f19446d1db44481ad92963f01650233c9d415ae8cba23c78148f954e3ae82b9ed70934caa7215ea16749159da307acc05872eb6c7889b5994edf16a13184bfe2901158180f95acb74d19b7823fd9bcda081e56a2d96f573cbd73eb55b3797523ebea6ea592ed9b8379d315877a8d14c4df9041c6a665;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5f87345fb187fe3585b867c0b10308fba91a5c1dd713b01ecdbfb21e47664990c39f5c21c111955bacc09aa5500d83952ef202b7d1a2838d73ddf93c8824bc77e715b4fa1db528b62b315e5c247b4f593289952b717d4ee375e137903d400c61a3c65f7f6512a8128264ee94cc60d67959ff144ddd14adfe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14db3a26018779de723642d17f01070969b483fa2cce96f60a7f7944f74350832be7679ff3a7b0b0baf76f65b9d4bb060ab91da3f13e03f4168df6224245f4489be75877843b03afcedceb48c5f54549527b4ce3ffcba61bfa98c011f5995e083b087c0f50c8160832191e3c99bb79e10d789ee7b0cbf7326;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15a8b092328f62e54e8c950dc35ad6a72cc4137f23957e3441aa730bfbf9d33e54a3ac79afbce5596196737efea8aaa7b1ee7edc20c29b5e901f20e8780bc0a18a43011059dd02a3051f5593549c254589de9e37865de5e15f17e1adccb72422ef6a37f723955be78150fba1025866514d23654d352d0ed5c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b06042c77967c9cf3c6209926c5c2161f6938b9e5734866907726271afb7f2873fe490900ef8a0f9356eb6616e100e121e1f45ad50630242567abbf071d0d9d99fc4fae17d21eeaf702e5adbe0c5811d459beb36390186a2c867a97115259d2a0c3c3b66d42a300b38ee9bd8e5214bfefe2dd3810c93646;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151b4bfa21fa8bbea0b7332d135c77e27b36fc6468ef726fcb122c50533a3cff5a5aa4e9cbf4117e8f15f83afbf39b7cc758cb7fc6480a43a8414ee3c40811b2dcaf75f4b941e4b2d957927a96ad891fadbc27eceaafe2531893104195f97ed1b5069d9d603857636bbd3a74711ef23075b3ddf9a68332930;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcde1fdea1d8bcd145046bfff7ac5b61522106e036b6fd3ac38ec207b19f864a8457819178501a1438a26ace78cc3ef8e3a634832e15d29717f5d2afbe4f2e1f68eb9fb32362648625c304591ae75187c59e18202833421d54650672bc70ccf37d18326b4da595a95ecf406392c27cec897fb3c8a6f9ba8ea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0be588748a13810ed7743998e5df7e2df1f4beeecd8e278feaa5d8c4a4bdb0d3030ca25fc90987ec86a3cc7f2593dbe5e0385655e431b12c0750dc002b1ea2c1bf5ef8e174298f2cc2574fb728fea6b1a8a98e3f3d611bf00fd4a6c6167018a5ed8bd39951d5cd1300656be75ce33a6bcd80191bc5d4037;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14573e4f26d4801cf36725df68f7281126b4fba8bb5e8290f85e3a838c8971911d64f853e9fb19cf5eedf8ff916c5dd0ad7aedcf443a08b350b0d1380156338bedddbef072a634e01ca4cdea9d48bdaedaff9cfcd6fe7e7eca8cdf8976bd0b7fea7c45dcfbd54d8c2b90f443132182a70c92d8d52cf30fcfe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88c93a0a6e5867f1f130fc8fdf18777d447ad95a160d7390b73431946159021b9e1d8e9014da13d17da39f84e70d655d3e93b45364838c59f4694f935f302b7610d0f150e2743becdfd34d9dc0910c748d62c6051172f055c6a50233cbc2effdbae49405d546420f10b06363748603415c30d6a2993d071f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1475b56b35b2eb295cb94e5e75e2a3be63084d88a8dcfc85cc5e87862349954550c44e38fa9989c96334c3ad9db019c6466ed4f2c6cb803e4bc86667b753b521685070e763450fc576338e8c805db4eb6d8fec8fed62aa9aec52ea941d873bd175dd1b8e056327be860469d44471751043fc420f09f55fd85;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132c219a2ba8488a678f7aab747061d39fde2412345fe554214e3cc1f5a6b771e7591de1d9e3f96362530c0469a95ca09753946e9f2a0ef3f94cf70cf14859f47149149c257400b322de8fa4b7e8e715ba7f01ebcd1d9d421facc5ec7872ddf99f71be784254c4b1210b71c0271e3cc5806249a7a5668fba3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f77b94938fc1ad2dc0ee259b217069c3150c7bee1670550a6a05053731032fb02dc46a9e82daf1283ace30912ccf3d57229f8d28d79d1ddb64812fc542ae9df9c0686686def70e6d910b2ae682c052f5e4de7812cf957218bec0cb057193083ff142d6ca2afcbb048e1e43eb3151866136d2451414b92a30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14215759285d22939f5782104a31773c70bd54c2fb4eeed4031087db6cb2cccbbb1db65f7ea534d1e809275f34384a0489b9e7a66d656f8af82feaf60234b6de8b1af1644ee062d07a7d8cde7aa49e9018536f37d14db08e3e2680b3d928248cc3a33f6d84ca866b231c11232396ba8c195d46db1404307ae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1767850893fb0a2b6dcf467ada1f325dd901bcc2f3b72cb300f0dd1dda31d6f11b58bfbaa022d159a89fedc49898e42d24fd2dd2479beed917023914c863c9b2124bd0e3d304a042e8b134e3b77aa9feb0779923b56282aa165e51e0e857a2f95a40060b809c7dbdb83633a1689041f51381b754b737af5d3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1946ee89fac3e0c59237edac033513fb43b8a292be4539535ca2c2c82538ccfae90d18787fb6e0b546e4e354815ac271fac03b01cfbd228b6f0bf8a27ed92f59d8f3097f67c80c6f1cde72bdfdedd5e8dc4355e1fec1403391f55b3526ef460363465e540f8eb749d55053c91c4bd08006d0a7f3bcc85e650;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h183f1d49fd78dea40a8627227e9996e4347843c0face890fc1638c016099a7697904203f2c5fdf5532c6b2b8dc5679fca688f8af5be4dff8deb513fb3df664c4882baf6ddef4506f609d02a5431832c23577cd241ca9ddb97d53edf3870476a7124d4ebf2099c78faf7baf55a122a0625ed7d3c422b4cbd3f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b7203bf1b5be29884350d96919e12964b8101c0ac4975d5a78077d152a90b88af9322e7e4c19ea9699ae7314f4ad7a09ace4462074c8c02740a98085c1d9adc3869355313c5286d5954c297f567bd956031bcd7ada6f7af5b21de08f97f149ed10347322be8127ce6efe9510cc501f7755ae750f15592a1a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e919109b3810a1d058160c631d2f9dd170c2b1356ecee9c2c8b36204294140d9563dc9459c905d3d17a95e651c6d20a2a3aec698581103cc078ce5b394971fa32910ccbf994e79e19fd089eb2e47fa787511a7dd25cc95d2b285d5c2585e917df305479460b71bce04c9715d1912f4e7e2a2afac2617c85;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14c9659c5beec248fc03a9b7d813de96bc3be58488c697563773aa8b7b5a1efcb121a53ec2910d4e24119fbf52c1f9c893c401c44a351777d796005e0dd36f1c8629bc67f0ce52d9e0e00caacf30805b825592df937bcd17904c05f1fdbd6e980571cbcc1a6421a84875c0d5157a4d44234c31be631a1d12;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f5c4a967465afb1934246adc60744eab76a39d9bbb959e5f6ab74513dee9cebc3bb8dbf809903bda4bec9c4681b4c09cdd8384c5f7e842bb86c2d1fa401cece42592a81d6d0f54b88fd1852d6685e137effbb6ae205ae3efeefbd711dd4659d4085ef47d06aa5d1354296eff8b451eeee92e15cf7a01eb2f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2106daeaa0003d93e10fbc136b32d35e2203eceba14d23b65aaed643af9d0fe47bf2f9cc61bbcf1de013c8548bb3718a140330aa53b4ecdd6c262f49983baf999cb262832c1831f87f023ec952cbd5bb79722cd4918f4afb462cfcb03e2584817e6890ff0612d3ae2ebf7aeb94a73cf1af765333b3a289fb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h416435d59a741be3e215c898bbcf7d57ecad97531543e78fb494d97da986aaef63e09c7167cdba6ffa0d1d9f2516c7e484ab65a4c83f013d437143fb54d1fa4f3d74d9db63b9c5a06a6c847ae314556c9c02c05c5ed7c6a36319a37d89a7a372623144632079bd39f7baa5cb7ab5a5b05ca01697fdabdb76;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b37c422041087f6bf5e6cf078fd2ed8fab75e8555e126c0b74d7bc463d3b4e83e75e44cfb7e256463b1583a9c68036bc6c5090d03d38162600a8b5d50d6692b644885d4e68b864bfa7e9fb3cf093d65a2e74cce7e2554cebb37415ea46cb79a2462b478383e88cf305bd8efed16fd6370616ba3d95773cf9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h111a691e855c2ce6ddb45d0a7b60e910430d1db21d0679ee23f1dbadaf3dd264ba8730d6b987a3b3bbec5c5e3613d66bb107a4008f737f90c97be92e9b496f529a527a94bdc7123bd9bca3a9fdc1d15213e044e8d0b67480cebde0936cf84c7a97ef44623777563fabc51a33a5be0a28320b1d578f94e9cd2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d91dc6b7767bcc65668b7ddd0ef6bb1ed811ce3915349062bf96209666c59c379149d9af14ff5c64cdb2d803bfb656442f33f097819fd996f5d790d6853429310b73e66d41c2b7969daf43c69a9ac995dbfd3d595246a86e2a5febbcc67f94ac8fbf4c215401757cbd9dd5323906b5595b5b779384808437;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eb57b98f9e3c0a71dff67eb80f42d2b951db7fe04ed540b08bd4f93ce014f2da111dcddd8492cf8a425cbb9c78be4d0b543f69d4fab6b1f8d76b5494b9473524b4d3bd736953e89b175ff9d6c4497f5d625e6dbde7bf49cf8a13a331ae06d0b5ca38795365e9a612a971b62c1aed36d37139bdfc768f0bde;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e6db8c926293591cf8c3e9093b0e8718cb9f3169e6394ce1ce41a4b9800421bb5a23945a877130eba0a9c54d8ee545e8b7923f8711c7d8b69c4e8e90dc20cd491a52f94500488766a5dc416534bd91d182d01996775d0438ad939d9f25bf66d35429446a84fb4d6dd2973025888512f0de17c7a4aa0f7c24;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c14532447ee25f3eb1a222c3de676aed331bafc176b8d853b8e0bba34d35bd03e977c15c790223314c852c2712cd8127b753ae5eb4e395a8ed1e5b82717a1e20eff7cfbbf66fed955114b16b20824789f40bf6f151ee7c37d34f74d2250f70297f4e9ab45a98587a890c1041cc979e819eb45b503b39ddb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c387131c1d4d6e787c40fb2374475c51603e6ee911fd6871e32647ca7af3312a8b5b18f9c91f30a81e00fcf8bf396caa8fd465c164f4faf16da185cbfa9c4d6885b755545ebf17ea6d2ef7749022f48ff865ee93ec02df1bdddf55b7426b535fcb2be0eb688432be9d21c31acd06eff3c7520a75b7ca5858;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1edf2c5d78f501e8487764ed2973bce4bc75b9a362a2d9ad74eee1df72eb01ca0561105d350246be867ba960a7b908f352f169671c7709309d33d80b0efea354738697a29793b8c75232b11c9833a8c856a438430369d4ff0e483f528e534de91fe23b68eb741335d1fd661b4405cc00bc31d9b5bf240d973;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f707baf8e9fb3be28aef25f086028462582b0dda2c77ef485bcd8fc23e221915584fe2fd46f7669d78b9ada5c03984977d47596561d0a51d04ee17d1f9ad944ff34dcbf835146f7326c4eeda2ae5ffffc4b3a50409f2a35956b52bcd86f92fe3b165850f57bda6de5196c3a93801c6b9b04de5bfd6ce395f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14696e2b466ba61c2d079612522fe346107f377fbb0ccb39d33bfd5f3656725301c79b395d393f091273df87ab31469ac8094dbf89aa0492d3aaa01e4657b0d7438ff420fa0e2728cb6a31982573135af90f1c07fc45ccbca7e9adcfbdeae1ab25d8408205915eeb7c7320a840f071fdfe3def7c43c2bcf6a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186d871fcfbd1f51487873c4eef1f3ad741d04ac507594011157dc410e0c35e306b99cc00f621953bec9444242cb3b567a38db479a5d7f21ca34eab12162ce89782d6edea9d5a2f6d5caa8cfca3099b3824fc0fdacf6d0ea6954a94603813101c0da744c7874dc450481f35f9c7789005aea065ab2f377feb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf41a181b911854b5b09587446e6df3dc0cb7adf6a675e36fbdd0353f31d9fd3f95907defa388ec794185996c22c878630d0a5e3994f7e5aa00e6ad63e8e233d4bfb2419385ec381c6ebd2e2ebb380579d265095c59e2f501ce5686466ac44e01c78926e9c933880b3b725d4a405f8b5ea906bea34bafe6f0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d0bc2390d0f2cef12364597d093f1b5836c9062c9f21cbad0fb467ad915fe5a79434be059872262b6dc0ad4b2f944c674cf62e77ebc1028dd3369a35487ac9a7eb6ff7281d7c56570d1e4b3db74e4bff5f02b60715e9fdcfd2772691a67f6b0ef53b97634521e0c55d6fd8b02468826ec2c5c42ddc8b5b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4c4dec02a1d44884b36fd3e4a4ef6b6e8b16a50c20ee6b5296d5f3b8e3133c9bf6821737ddcdaa46596164a235e5d447cecede44b05b53924de86d254314e6b943e6eb4d7d3da8839acfbc90d95df283223e5c31b21443922bd43103d832aca01c7a5d3d900b3ce6bd7c34b82498bde1363046dc548b1524;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha7250259da9c59b273f1767816caa5a2717d3cdd6a975407d9f0f607cd68371694541f1ec47e0b883e3a7c9adf4494bda44054551ba933a3cf975e3805235fddbabc1208746a85db804c2daf12f8e8cd68f770a36c6b264c785aeff0bfb07d00b4068f35408428e803e47be5f0517b3e8151c6b924ffc8b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed791b22d880daee97bedebe545e75e001ca3991dc6589389ab263c1c4858ff815612627f13854c8cc58e789e178cd75e445cde8c0ebfe43567d5eafac7fab6eefcf85743603850a5686caec9ce0ceb513cbb3cc35975bd3e8c599f465705ae408f8b4dd812cabfe845348bdd48bae69828a97303fea4ee4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h34c6ef6ef6712adadc2c7445619d8ba98a05618265dfcf580c5143d304736e69f2a34c98082a36b6b247458db3978bec4503583b79958aad65c6486142cc367b51519a504cffeb0639a5c16b49f7c8a0d7502fd805e7c4f48e16dd3ee2938d5eb596853f37b1607788cf44c23aeeaf2452dbf18585fe7e22;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106df1273ecb55da86077205f705139c470f83ef2e22e5a75b27a7c862b34b3c81e34710b9de79dfb1bee053ac80a217dbff379d272aa61a5046fdac4f9056b7bdc4a10ba66d0975eca9e3554af05b2a11de1784650a9e5481cb5ec478eda8405f4deba7fc967d77069f766eea67c9610fbd8966395fe4399;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f813cf894d83d4d5f505a488a74b8bf9b10ab59ad6b86b35514419377b84e05f03914bfc49d81cfd1cfa9ae56864fb5a8627490c420f655f8c7d54a04cdcb67e1b62846abc9c71caac3859cce700722556501dca499905687c5facd9cff57f637b756f072b904c9cd281acbcd67521945a69a39ad03cfd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b22b4afccca441adfb39a6fb8f3cf82e268efd559fc8f317ee784962e7a52ef90a53e1aa997828728ac66fd50bf2fda3b30581c54210813e994e673cbe1297bf7009c63d818d23aae1b30d7f6e5f39fcbbbb5585d0b6312639ae1734e275cb9c64590f32d95103e1c2381cfe4be6a1ec9304186842c4134;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc31e1b6076db117535db3ee5a3a4930118c9430c16914622dbb3aeb273170d4ae99e3b26d941a48e6d865fe27d187a05e2a7923776b6cd40cf2fb9b3b02eaccbc8c725f2f3726583bcc2a170ae2d38ecddb1130c3586c0237314398b4f1d972d6066460fd9b57abcfdfbfc0d89f89bc5601df28782615cad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d895cb9573b01bc6c2bf6f8ebead3ca94fc587588a0aadf7f02bf1e67aaffe6c3838d220c42746e1d1653ec7e340855d87c91dd85e41a7e8768fc0d9a46ad44ce746fa30da19fde4319c282cd49140578ab9dfb560be2f73ba5b8331eca6757df07ad475c8e111362d165c34d05e9a54e0039ff4a9f2aa33;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab172b9096be59169dcc32f1e895a737d9e23a86a556da4a66d26966a2f4f1a3de0fd294ce77ea1b208011d54af17dc264c2ba444dd4165f4597814016a1ac45869df70b5d1e8228fc6c4519920eff9a9946280c587a1ac46ed41a784c1210700c36f7b976ea38b7a86cfb76e73d1274392af3de1aa23f0b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1adce32bc7e282e3ddd34e75fa1b860f21d89bef9edc88a14b69e3742efb09ca5949869016f7f86bb16a66a1a9d6a1ee3a98b648fed9eb29893196cec83e00481a659e4f42fbec6d919ee0c713dc585bc257a5da0d721a5a3aba8b12136e7ec71dff9beed55ac659c185094deb43b346a1e85cb8965bf3360;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d920dd8a0b32e6b2d4076c7623e188796a2ed6df6ffeb121c2cde2b9c96f60d2b75b29f85efa923df9dca2b6eacb75016bc2561d0f8ef5c10ede0f2ef3cc36f83bb9257cabaa436de4b3acdf4c2118c5c6097769a9a2ffb72c68e40ca580ed0caab56dc6d4221956c36548bfa719ee8b0e1668352a2eb3f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e9fbd535e4bb9bb33367913d3024efef64c824ffa5306000708b4b0e1c576ee8c19a65285297f02d5a8c3fafa92d65e09e4c9e08d4da894406a87de6de308ee58bd96347f3b631b0346f56e60f82d43fdd8a9c16d305c6eed11b3fc747cf3496b67b975a2e1ae7413abac6d70c2c4b0fae68efdead8d293;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc9d6aac17d3fc0f09363087d284053c782bd76e5f9467f30ea45f4b6fc96d6c01b70a1215db256de4f152235a299129b576d6b5575b8dcc0bb898676af6cb04158e958e7323662b0f8d8088910463cc191ed624ccf3b9264fa47e0d6aa520d3bdf421a8ee2eb936cd03ace37ec87a8b94830bc4ac3791581;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc1bed0263aea25fa80888cfd255b13aa88f08471d4b0218c091b5b8ae2eb8f94f094b83eeb8a43fead7ca761ae5eb81becc38eca8d4b58c377c5e841c985fa673c9098f3900cc6e017850a3105caff7926268373a24f12373a550cd07282f56e4037c9f8565741425d29717f9508a075c3a1f3cdd4c7f2f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1811b44d5e9b9e75fd1ee8c34c62f162f4cd2d8d1d0035ef905a470167217ed290ca62a507d4f7d5dfec856a77298aef8104ae889c565e34906dc8bb7e948066d09153dded665deeac5d03b911da3acb5b811edd90312a6442e6fc9d537d6f01eb8b42f00291ab7213544a632d04153c1c246b118462f07;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f113505136e620db7c749ce8579aa36ad30359793a2f4fbb77fca8a6da85011c2c8a39d839ca027dcf14fb8b61687751cb929cd4c3cd61138fb0e3419c1b945c7007022c9fb965ab68d0dec970576b4b51b06854799c5c2e96840172cbd01f438ca26300f30e0139f121944dd8017057648345854161f45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16aa9b6053ec42febc2f0531505a7b1d93fa522cce560031bdef09590220765575abf35e3bf65dd281babaa9011191b2e3cd51c732f9a3458ec73695c9e7075a22d3b1fe40510e9ce74291d64e7bcf07323fa06d1e04afb9e25df5e33a1ee8f06ea4ed03c0b232138dc97c7270347967e542d3e4cd969f744;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c70d76d14f617d01dec0495dd83fe691c4f0be4424964450f68643d44993277d98b5da53fbc5de39d27928ae47cb92b00f364a8094bb07c00ce67ae61b4c02686baf3ef18d2163fe4aa21db46d0d36254446226284f9a5678ad3e7cb57d2568f74a40859d34eb2fa593a6059b3130cbc4266e6c101dec63e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1481a624b9dc8f21cf34f2b4759eb33511a343bc78bb557f27097d645110a1e06e264869c144256ca5b32f85ba156cc52c1d1971ea6fe7ac7a532d5a55ab0b56681484dcce5a1c4bd0ac9c04ee2ae9e455ca588af9d8549415cb812a6cb6f5eff6eae1fdb239303f95a41536e33256ee0b8ed2ed86c271f5a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf64a1a56ac8f6f6566ff2b136bb1d31b08f62b38b1bcd158a86733f1d80b16d537aac79a2f5e8151df2e8354de74d7a26aa4381b536d091f422bdeb67d54c10be5b30e20f423fa4aec14f56bf5cab3dd2d92532776808497d505ca1ae5c6d1ff42a93ed9d856f4d41bf4b08f2664122cd436b5a43794ea99;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd2b680eca8788b90dc823bdb610f2310e1c68042f53014b93d1fcdc8a84a2d0c81067cd942b4b4816c850c9c12bf463f21d7b31233b3642488ec4a553bf6c12ec444fc0db7d3a9dd283960abf1be68a5ac594af4ebcca00d56730b8c1802a2ccaa682e2d9422028986ca89fcd0cd7efe08adfb0b9faf0de;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5a24f71d8c36f49ae6f2c281f54c664a23f56e24a63a332d068c72cb3bb7950f25e0ff571221f074f7286ef1743ad8af1088eaf3acd3a913540ee8683765b86d08bad412360106a3185ac0a8e379abc3418c59929c4b7799167b3dadf0fb70a8557e3f731ae76c7fbd6ed996f7f37edefc0df0b208436726;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h134d3730e4e51f8cd87bfcfae864f5ad10492bd25ef91316114bac31f31ccdfd02e172b8eddde2e9c71357b95b45a372d9270edcaaaf51ac3c1d3fc33689ce721bde08399a49d1f2853dc5493fa501b496b2f0344d759faa9f36dbcda6994d5f830b7fe42a42a19471863ddc4ac6e8fc5e4f4d177d897f8b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128ade4b89d03632c56a0859d604dbab21fc9db8f9d6048335a19ab342b6478ea904e791b011652051fa3ad5fbd747610a1247991d73e8cf722f8b6cbcefe1e845208bf6b3ce3e1ef193f7742a457ad37e8272a35b485c5883e636d6308383aa00fbdcb02c8f614d89a8f8494601509d911d2e0a864d612c0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbee2e798c78b8dd7bfe516130473086153c46d870a01783b63bf2d5953ad49406e9f6b351b4c915af68b320156ff6ce5120c5732a9253bb190aa6d4e1765be58112a17190801a0370296df9bc33e6eb713961dad9738ed5545a936629bce31ad4c9faf054e71b2bd4d65ee5d96e5c1dfcb7c12c5c073e9b3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3279c12ac77a6a44fd8f45211ab300f2e46c0fdc2f7e0e7691198a1ada02c073b1475261f980fb414c98977b765375e9df723483d1856ec1063d35a257c014e72dfe402c6ddf8e1934ece08ebacbc26407ff1213fe866aa6543ac603621907cc211ba8a72c6cb798d3f004b1d32009f5905cf1807c66c008;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168c5e1f51e02925dc8516ca085ff4668b236bb6d6c910dcb88f26b8efe79b8e5f0c14f1854427783db5a085ff4ab741a6bd86754f981cbc41d493c1d1e05e5c914fee56ef72f6974b6bfbe951edc5466a92bd2330f252f36d75c2c5dbfea867da1d717b4640be0bf92eb562ed12c9c83b397f35dba95732d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1807452b75ac483cd1662d2f3edcfc975b49c0d999ffa32fad3af69b1508e97f3b95b96261635faa3056aefde1ed89c8bffc493e5fe9a96fd8181b0c9e94330bd6197476ba66a48f25857a6b6d97ce912b7094d416834e3f522385f9b1064390fab38e4f12bbedf1fa929f2fcb02ebecd24dc6aafa8292b4c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc939b4a594bb6c5982d85a473f5336ff28e6b4961a44e0032572e97cb914c97390e61c5b6b4d68d8432c0366a38bbab80ba243ed65033abf4eb52b833cf0f58ac001d5f3acb7a294acda3489c196b6b3b921858bd0246fa08d245213765d581d90329434b9b6270383237dc44eb87a01672907ded5972f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cc1da1106696ae1bf1a6f658d337a3dfdc30271505789a88316bba2043c5facd090bb404a2972c2501f53e3aa612b4d3c8e172a3acb1b14a0a5cb0eea9f9fff18775dd6ac115c44b3a89cdaa8a5b22168a324eb9ef02c1d2bdce4f30869b8ed3320b521878007351c17e9f5dd736964330306fe4fabda0a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h129fa8f49cd84d19ca8ffffee1c0afe0c9e18fee9f5e4a11292dd27b820e87e8269f1fedb891a9ff22b3331fa39c272d3793bedbd8e81b4a3519b486d11b5fb6962fd51b1d5ed4c53525a83e82bf8a6f419680b994ade7e696f3af7a1d51482bc591105cda8eccfbef9ff7346cde97592cd8acf4fc2fe9f6b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2cfeaa3a06243c2a02716ecbad8257295d62ea173a309db98542b20b704cee28da12e9c94347897033ee19be116280a20b341b8b95a62bbf2a6249f197f42e73c346a9a5fd9ce6467f1d9ee5ab67a8b633ad528f7246aa00914a10d26b0918c6ff4859a9c92fff9adccfeed9d1951c76452fcd28c560768;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d66c31fb66424e7ff03b987f1032c5a04d752a6d2aa4f9b390570492b7d26540deeafa7e4ded38d32c5a12f2344bd37821ad8dbd122ebcbf4c076236ad07dc39c92bb079c47003b2f2848cdf926295e5200669178a772bbad925ed6822f289fd0ca8a291b1d6b811caa718edde8202f4654754c8cd53869;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3e57acc206d35c7ac5078d4afaf903032bc3b7d57056c3fec9e761af44f96925dd689a29ce2cf28b1286ad4223fcdca8e1b396a57cb702134e2e083efeefd547b50ff411e35b8e2280f48b021511d3f5977642f781b279bfa031aa82a1a4ff2989f3edd8bcee1eaf0b551dc20e634387746f7c66b989505;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1822c62a7032972fd78d04e1550413f08f14f43c0c0da4c2edecec7045b5d0df17327f64500dbfa6bd56ca5a519d4fe72c3ba8ef3c023ab1dc6a224291aa7b5aeb3cc12f463886edaebff7f845c8e6025a773b285a02af216701f7e69849c831a4f9727ad8c82f2d58cfb9e55526302ab5a599e48c49d34c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5749c9a5e10a4559477477c85784c846e3e4545076d08284789b4e1f0ce16cb600ed3ab7b0f8071aeae9c6f0273db3d8facf94de5bee9861d645be9d59454aca3fe4183af7eb994a99367e0788f7d8b7301f00f2575d72099cb7988692dc437e5febaf9a927d60b1635612ce913abe38aef7256c454917b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6cbadcf78a0495bc9a22ee9a46cf1878a3521cac67bf37f08eba09e6ab4b7dca84c5ee28993730f9d427404f35ddb3009f82840b6a531ad1246ba3c308d15fcbc879e71f1fee1907c2f752b12146c75388cc1c2d5f5cf4492f64ba77f38a0527c7971f0547b283bb8640ffb62a7621f44dea19319cfe30d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a946d5c9ae0945a51f49bb4cfe552b6717b6c445a1182f2173424e4095118f3bf9fcc947be4f1af6ce0be6ab2894ac11331c79881dc1896f4a89df510a21099ceea58e24f3409b2af52b3d00bc9f8999638655248400548c77afe5885fd009e36e22a391ed14b048254ce78d90914b5e4e3cc2af6123f57;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84961051177a4e7eaa6b576a85e64b6f44da9ce9cc88b3a0a480ea5c081fe27b76c343d176bec61c6106a757e8445d8a9893d54c1d771cedbed6767ad3e741c72059c181544c9081b797dc81b037b58a4875e792e662f7f82a29d56464bf54ed690edea7a4db455ea3d0ca56434a613337c455a250a43c5c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15c58ed59a4466e63ccf67df4d99d24d60cbe51e88cbdb473f21d9e8ff7d058a2fc016667a8d594f3e96805beca46b473b45ee2f72e6fc1c5bd64fa3eedce08a081dd5e1136e83d89d90a90c941d1077f17d6f5a62a9f20add11ec57eca2a47eaa8ada2ffab91e89340cf020a94e0c44597ebdf3009b2eced;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f7cb38bed891b8a0e216e736b892ea7de7e5d9f38e7511e2ab2ec211e2de22c83d7c4968228a202a7a8d2fbbdfce353bffb7e5de157c7263394aa1a19cd717756461202a89c39ac7b5714315cb8581911ae8ecb390c1b4220fb14c9ef226be45ccfbc01bde06d613ad5a7d6b3481731f4af53b173cc30fc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f48f2cdece84fe02f4387deb5c91d1e10405815b50ca89b8887d121c080969f24bf812fae3b99daf1d08a41e38ff1f5ae257ab1462927a656f28a62133704e99a3b09f333bb0e6f4efc213f90f73be5c6132ff5cc1f49daf197c917969e8a799b29846be3f7f6e65f08ba6a6029f2945ad3a59255804b387;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1df7d9d2071fc9f9086474d85b71521afcfbe6c5d4202b18bd1830b366c8486faebfa8a8443e05cbb0474d7adb9dbffc91bdaf213ae0b1404c285a8667634ec96db077d847c5b42f067982bf9bc5ad58e5d3bebfafe396ad6fb892856e60255837ed58f226c1458774d3ebc0e8f83b369f1c268e650b61373;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5da87d4ba46d0ace29192ef2d0336b99cdc7008b87a6319b26c7d371cce634c370145c9e7ffb94cee353c1cf9808a382f638b95c6e35996f358d7216de2f1cdb507efffa74d56722813ce61566be3f545c358516026623effe327fa6dc2598d4b191ff7289db284bc9bd9bc6235f56b2c2c3e5d0d948e0c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h133bde21a7daf7271b790df7de96a0bba6762b79b74b38417408a9766f1673303f917bbfaf93527d22f0f961a8a8cb948e6683c6209eb9bcc618e4d8c96d07a00c402d323b41f6d89d2ff9b3dc0a4666dfe2201bec6f664753ac7ccca9142004ce968deec9c8f90235eb7fe3c83d5029d4e35e9f76de647d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181d3dbec0bfd225910953bf4d51953e47299bdb7b9203c3f6ae0630cb008d13cec4be36a15df42b6e309153c23d62ca4b814168fe81dc59173acec96605327580e9109399aa1c1ed0895beb1e60ccb7c1396f9d2b24b080bacb17b256939e9d48081a820b1efb6e4543771705ad0ba480dab2be3ccf21239;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9a0b254a17e8721bbf9e45510e54ee953857080c8abccb7e02032559ef7817fcbdf8e96f9ba4847f8e377a106e150ad1320f060f1049ae500114f9d440fabccc73a20331805d864f00b38e4cf48985f6cd5cf04923e7e25a37d92b06aec9c53937518e544149ef11186f21e091cb9aa2c09f82c6a9f00eda;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9566dae82ea6ffc1440fbe4548d345402a49cbe1bb28d1329719fd65bb652cdb51973366c9811ab8bdb3de079bf98db2f76d9c475df3744d01975f50d6355550c0381188df8369e760e10d9e8aeb1d9270f864db112808447cb23adbc106d4566652f2c0b7a2469951954b0dceccc4de74a02bc8164459f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa9ba3aff1befa5286a3c9a7726e214c2452eda3468c62249747df78078de5cc81e629ddcc87cc548e4aafec4be7aa75ba900fd54813254e5d60eee11b8e88f8f98376efe8bc242b40d302093cff93ca3d2208b68ab0778150f6f5de9905b692255ad43e22735eeb3f08903e96cc145bf38de60702987e41;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h163ea0dd6735f60122b2d5e19d30d6841a90559e158c7d2dc0aad674375e71289672ad419736461d81d23114d796f9612f3e7908f577951c0a3768a3cf633a82d3dd6eb3af6e133577b114ea71df4e695c88b14734563f20240a34db710b81c1f81588ef09e95897f7bbe5ab7e5fd4fcecf5ec6ad4193b331;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fd839799e4e3ff701aa23312f81942db2cf50fa94fe6fbf1ee7512e6ce226158d400cf7ef3894c43b2c7c077db0fbf91d057e4a156d74e5eac2f2ebbd24a39f33347f2d4272cd59fe09342f309807190dc46b02217e61aca8c098ca50470b08753bc5d198d0e570759daf3916045c4a15de97f075ec65731;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hba3bcfe1306c6f0a67b0c2e3bce82155ca1f5cd0f041f3868dde3aa0b930d131f03eb405649b835a275fd7e39dadeb6431190da50a6ed24c842cc0aa1951bfc6b398e1d84f639329e74757d1787065ac723930c956045541462519a5b1b91bc9f25dee39558c0a962699507f30a93bb2efed9e703f2aabee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h508f5a4b043e5604776e855d3f5ee44389bed4018b780a68bd062948c06b51cabd5fef1b3a89471020f676b42d14c9dd1cb759c70e18f49b1ec573a1717eed2730bbe922ea3f9dc6ea4b98a8c5c3995724580d4e75d915ffeeb6c1f97a6d453aa65123365594ec46248bdebfaffa3297400316682bdd90fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c694a6a0ccc2c65a57fe5538ee00231181423c10bb3fb03aef3dc207d772743c029e0130ea1bc0187d26b8c915c426662fabd55b2fe3a302600e7fc1e533faac8e3cc94aaefa25bf683a505b5a81cb08a094c814fd428fcbceabb6b4939ba7b2389792299f42fc529fbd5c7a1cc2378b86d8a50c15eb447c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1939f2a54e4d89bbcdc4494f29412a67b76fb22ab0db5fa73bf8dfd3793f5e85234957f2d57222d9fa4be81afe2a533ee19d2780f408be1b5acb13a3bcea126f9b6f8ba9fb4571163c0b3cade984913108c1db6d97b53a7449d69334ef2c29ffe548191695e2e32ce49e0e100d6c974ba8da5b461b4b042d7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hca21ddc6ea06401326df976882b98156d2c01dd43d29b68b4d359a678a20b331fe1e487335feda06b8ecc8592b19321c9759497c45e7b174fed8167be94dc0476c577a375dbe7946cf0feb4a3175ce37e681cc67da6b0047f652433e458867175b982977184f480104cc60210aa08e084b214c7b68e6660f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d63b1c7524eaf18d9bee8d345ed9499b0749cfbad2b5e934cf50454258afb135cba4679cd339aca32be8139de18fee91df4ded0b7eaeffc5aa50f7c0c6f85e30a5cab67e895486fe090a88924267115b5ab83f5a3c475cb9a893489d74d17956136ebfd092162b2ba1b6e3251229c10a918229054e11abc0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h26a1067b5612b76fcbeaf91cf9115320ae94901e985a69742baef2e60957d03aec6f3b1820e42a1507fde4ffea23a9ad45baea989c50cbf922445e3ba36d084354cf433e8f3e9177de4aa6c18985439cfbc09362ec08994aaf00b61a73425cc5904f6f9af4de9dac68f27facb475d24be6d7344bd60c3020;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88616a602ec21bc5a3e78848cbf34f80ba635aa415a3f83241382cbe53910054c80d559c6d4511ea3333ed5d96ba6723d2b3467b1d4f7c9179593eb4e8bae7e9a30e0d31b90ecd8563f724e2d6a7b384508ee8fe8da33724d5cdbe229010832b450a532ba5d9d91f6dc982db483d306753c5ede82a093d72;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4604862722badac59328d06de54fc6800282f345e624b16708e516bcfbc3e5505098bfdb6f7bd1a74ace498190ebebeb270ae9ebeedb1c33e67d1c23c94178469d4ce4ef886795b8ea50479574289b08e1a2fc4f9635670f6637b8f6a2ba21818a7e6ca7c32e422ba3436aafb2a57989f4fe7685faa0c982;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1823c91e5723deb2ba013f898a799d1edca1b448d2af88625303e7defa6db0bffa463cb44f0e8b25c4a3fbf6e3ef86cf25392afb2c13b12bded4a5d303af721a07fd653dd797fd2926299739c1967dcb8e66a22a821185eee8504a888ed490ecea1a2521df8f8d9b2e6997684dce6c70f9211264831717027;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bed9152d0d62aa1bbc4fc4d76b32960b1cb01389d9cd3815487fe3af952d9982b9e63269f73fdf1b58eabcc4a243b7ff5f68fe0b6316fb336896c37b82baa23cfdfec91ecf58bf7a7db3f1fd0a05032befacb819109d05347ed4d98e5efcc5009ee8e401cac6881fe89e4277e506594cfb045269987bf265;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f67604df8401ccbc946cc7bb7d01afb63025a7d2d6a6eacffe6597e4514cf74443fd6a34a2ee9563b731a3cc6edf4f643b0f2d52a8ee711e958c3e61efe5e977fdf99ea41d4d39ed2b112b103edeea6e5427ccd3ad8b580d430192e42338e062a83d2050706f836c410f8cc5e2f3d9afee159f7b9e44636c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b82363089917ec929347fe98bdbd5d0684862001c189fca1cccfa0e0092056bd6407dc4be7b9fe2f93eff2624d38b50b743ea382b821ca47f72afbcc843d213648b065ffbcc958a1e3777506cb9abd1174ce2e55629406e9d3f80b609cd68246bb916684fdfdc972857a1b4b174da9beea21ddc3afb2842;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5173393845a951549605b58e5b96adb938d56f4adcf89d47ad2e88eed97ed8ebb2fa10e1d145f895b30b79dec2762052dfe7fa934acffd2ae5463fa189ea90cc8b6ba00fdbbcbc956754f7c5625056b20c64979f918e4b36dcdb91e85ebc47ebfd1077f55e91e81c111a47687930ec792975e166710b8ca1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d9621114f6459bd3c0a5f7e9ad441ba230937ea3db70b90e8bc8f2a1af077de88d7e35e1f42a2729a7bfbfc00ef9214d574758c1aaf21a7b7255a863f41cfcc25704c21a4f5b36d1744b77b4bbe41632fb023e3eea7923f96a436b7246854446b305bd429afba38b5c88ac57969cf0c53643c6a88175d744;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4db71c3a56fd457fdba382dc773b13ea8d75ac9067a7bbbf9e37958f942e28bbe21ab7099b8a4332435ceb5a92a96666960b5261d775d4d8b5e067244ac8ce3134846ab7c354412125e9b17e273e30bc67a08839ace8a43208bf847ac761212abb71e074032888ae4595ff5d240ea1626061b4b14bada591;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1118d6035b7a592ad32d829d42f70fcdc25d7cf2164433e74365f86a91a7845cc79963aa7fa12bc7ec511ba0b451b9176f2a49bd89287f71264ad25a0d23371f4b84c19e7160b4251d37037310684681d06c10061e743aec27d6e938967fda9f7afb010e2bc1afe15d87c9d98af447b1b5be6b1362f1b3757;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h543d7a12fb33996273356282684363427e8f00fcacf9852aed5eaddc07f00b386b0e8601689763064f953b1a3ec6f6467697cf71487c3f5d7dfa7a085df2336a5c139260b350f520800a94ef05eb094498c1ff21c1d16b27485accfbf92878195b5dce40185adf15a7619073823e3f2d0e3886acc996a9ff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he4f33f3f89e8cd81693ca8e0f50acc1065f48982e9a20a6decc44c924b8438a1e0c8d4926867581aa7cad4c369994e99fb5b1b06f8f260fecd6df436c78abf321dd1b43b2353931bc7fe1b10ecf616c2217b99f7e150ec88b7691f203ac29bf91a50a63bcf1a342686aca10c2dd5b9b77902ab83b32f351d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec6ca7f6a544234ae03358daee3f0c38b981b73102033c7b4cad28d8e7aaa63eaf0834836afffd1c85120f2846f0c5edaf023051344871bbc059347758020fca903ea3289f386cacb380fb001ddd403f06c99fee344842eabe3c3512712bbb7c4bdb0a6e0cfadfe8e1aae8942f1b86cee79003345d359f58;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h827f486ead28c92d361cd592232df900e5c676ebda4085e78b889c8b6106eb1a1f94240eeb28ffdd061b187fdb9f09045e7771257f1114fc6a61f4bc6ea1a43d4f018758be03c12d92be1846c75469e5b25b1f924c25d063073191788b451271172d82dbb32eee83bc00bfe7139b3f631c7b65bb5c4d7b24;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha265702516c6729a5c9668510fef145115a369f182e88f5440302b352b20a59522dfc6c4b9d2e82eb3d1911a016af134f101431aa2ff3a4b6e1733688b1412d88b9d0a74c110fe2d6c699b1ebed4d78aba4de2fd9633a6f6a0d25f17da8cc5061a6a41fd9eba313bdde1236e56c6467b525eeff9f0622da0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcfd5d51f8bd08ae2334f1625519ce12ddfab23153e9afc9f1fef97d94b1ec517f027525a413fd3439a4b72448dfaa11ad0b696ee65c475a13f9dabf1dfe21358634dc8edda1fe6cedcdb57552dc08df056c64314bf25149b5629a635e364cb6c89809d20ea69378ca995528b37e097b42340d58a54ea7d26;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142bb3127ae363412525e37b40e261c096c2be0180e05a916c0bf891c418a3c3eec4412132049c904ef55b4a15a2d493fc7f90c3c286d0bd3cd305dc7567e38856bf88cc39765ed0adbfe40340a16de4b53f3c16d83ef22d6c074e0483218fdd6e58120e7fbb92cab002aebb939b4cd3c5f4e3427d293086e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h97503b0ad33bb4fb023df864e0d278aa0192104eac8e9f4cdc404f923b1557eea18c946379f68cbd8ea22c6fa05bffa69b8ff4b92a8309fbb29d53a9d5d8d903b4c60e2aecce2e56780b31ec3a944ea2931017a4a4ad33d71c59a483822ab19405b83ac6cda7dae1c44372d9e4a01b7d1ece7eeb9a3a6297;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h93985a45a0ed2f51886839c4a6c7e41e3d6e47514e969d1a3f0e8b2cc4a3123864e928a8277dca1bad1b0260ddab6179eff07b89119fc6392362737d788071461b19539e4ddfc3a063d17cea2056eb9e56db36470ecb389c2a11bf2f1e9afae0e5cc44278a5db5fc1ccb95b762345697aa53f961c50fb5dc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1225041f94d024273dcdf98c9e1381e62b0bf527a29d03141a33ad0eb001b273d2c43a13add48bd62bc674ded2c8749acf228c4ad23d98e424ddb00a72e4c562f92316113a53ce0aa1693015fd2e0a32eb5b92447568475ec6e4aa04f48a3d03f0f7f1b22850b2f380d6dc544df397fe579e06da1f879ca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1505ee7da5766b9c95118244ab95c8168eafd896ceaee2ba6054aac6c464c073c4c4bbd4384fbfc55265a60887fd494258a26026262f9ab92889f5db8fa02c538ca14ed66d67fa5d7c9064349ad0738a725e07274f1f68bf4528c0ddeca31af985f63f729638f66fda65964226adb6deeb01a4ce9975e463b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1751298629b421c372cc74fd2ae4c1baa4209e2891da80515da82c34f71a6fbbea7541146a4f54d353bc984bd4152ccfdc736b3d0e0b2f4b4d4f4793e73305840370d79882d0b79b893b0d98c1523ad252591cbc74979cc47b381f77718697ec771002ef8040e3f6b0bc0ce1b9aeb0abf7ea6aef47b1ca195;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2fdcdfd87594d47733cff59a6c9ec36ef1913837ef2fc59f78061b9d8bd8d6a3671c2a23e7eb06051160400b130836c1f44283c4b9a85c38b30670bc346ec25c73639712b668f263fb181ab6a5e63690378aef9bcfddfa8e8362fd948a015a4c8a71924afec704ba97bd881e5603b7535b569a77802595c5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b9294ac62f69256dd3ade6e510f7261fb4458464af8a2190553e4c6c8f536bbd0444e097d569c7db394f88877e96ef31199a54f9d70a08a862839247590e0d6cdd4b869cf404b2d41c31267328b64295cd5dbe02ec5ecce2d3170cc1dfa2a185026735cdd245735615c4531154a02e9e26d4e2f8a489a86;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h121a88eefd684d3b83b0a8295d03423258a5bb99f3ccfd5dea17391a2b6c94c1784b10a874df0dfb1bf44e7f8f69e928d7363ade2def01e82e99542de386c006bd7012c741fdb580f007b63a3de4b8328e81a072c2c41b06d9e62dd4121929f07d7c8e7d367b6e2b4ddf1487dc63fb73535bc0455a048565e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1278671c4728b7047a2536a14ce91a8fcba4c5fceb3e49ea3c0e37030660937a60b37519124585d6eaea2dbcbf03e75803b2a596d1ff9a8e9bb4608b3b73cef81d13dcb6ab506eac51763230f2706ab46060891f965ba65001c10cf549b6acf2c6f61c0e510517e6896f3ab45c563abce796fc66d29ce1c03;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b609e9bd04b183ce984ac9bff68f33aef6a0abe5be29c79c97718a4f81d986eff2ca1bda6553a14c1810d6b898b9e7f0f734c7bea730af589dad4c98b3528400a2fc80146bc939ab85b0fe3760880e904426900767194178eadd3f79e83bdc3fd3765bb7a053000b647f720cc49fd4437b78de2740e9f337;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h125cb0a12b963fecbac9c276f73bc2d90795cabb4f3ac0c2e6d62fb37c8066ab89a4c5c56f076e9af1956ab0191fdd996eeb6222a333a93a3d7ef289384cf0bb893038158f59630a83cd5d481ca096a1712ebb30bb979b29f0d9210ae2050a97ec9ccfb1836d26ced84000281c55fe8dfb8d0f6a578a53046;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9410f4a6b6e85e263fb0187b52a55af76ee0c74357e363037eb7edd10f65f84e61629d9725b89c48d8dfdac6744fd122be65ca2afd45677addd823d151d29a7fd3c0bd1cbcc2693b6904dc8bd2fecd682cef5fc8f6b7c53cfa76b263a484cc4e5f7c5336a0cf3ac39d17f28aab98950926cc3b43212b07e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h40ff44a58c0c771ff6b6b243669789c7aa7c1b17af903b6132a063d00ce71bb10418e973618ed12542d53035fd312538a548a40553674af151087a27cc2ef590d2f545d70b6d5d65b387070b901cfb1fd4174b31abfd4d869538d774d67959e60d2217fc71fc5dca2cda63aedbf86b64ce66f70010073b1d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175f5a33e3f4641a4da645bc3c5f389c6f18edd9db0c7c71e71345450fe003f7cf8d1c666c666735612edb1b9a717736f295123a44cdd269fb483752ca2b1fa82da1704791d07fc15c9397cdf348af53da48e9461feada79bcd998dfebde9134f66e8e0e9db35bf37169b699c14001c9a8420f2c3ba2a2fde;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6bbcc9e99feb83675093ba607132c2e102e56097ae78189801147a3736a07fe439e27dbcb28d57c186b9c02fb75b16247d9c1168fa4e2afeeeec16c0d526c35ff594be377a15c558a87b78517af14227f281ac7f764140dfa97944b5b0da69f8b4ae976e746140436bd9b1604d1e309a8a88847eabc2fd6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h605d6044e801c006b678908367df988203a2844e859d765e89368e33522670b7a6138bd6cd01590a0fe100b0d28d2a326c74cd513344c175aa7892ad5d41502cb4fa102475f88fb6ca4f1089d4c189592bbe2e279b285f586dbc158b2e1a55ec37b562298978d566fe410f64aef941d71d811c0e2c67849c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h139530327532c5f39b423320e93798725eb95f89cdd9ff77bf830b7d2c70ab0e71dc7b0e22b79c9165e8a59a695d2d9a55e61f1687f7b22b86bd592577f41221e2e728da05bf83a3c695baad57dd249e8701ef065c96a21df08d6853d9c0063cff78f321ab325af7209d18af3b43ce0e6b1c266e0e67bd2f8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52f0eeba2f4a60db9d37a9116974c8d79c2d07eb262364ceaeea4a86cbb3f902ce24ca48266e432a0cfb1d31bc90a3e213661d3f8b0c13ce33a7e3d70da734b2daf1c109198cbf4d7d789fb994629a2d56355c284dbf0f8c37112308c7cd69932a3e2237f0b31db84a501f9a232613b43e718dbd6fcf3806;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17d5c7d38ca235ef7513da2e0aa19961275838fb608a47812b7df7559ddc7e86f96c5179c3003ec054678d2372180b848c5d60fa63fbaf34bad36770ebbc9486e4f47f5efdb65711b2f20b9594614a7713a927b731e250a6fdc142b725ea3ef07631943e00acdfba8afa65d47cd0852347d662bbd81adeb64;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h152117052f05d0458564cbf3174ef9ccd579a473d876dda8e9f7d3b4c2886813e57896189334f9e3df5dfb0374a153fa3b8f20a5735f6f291a4854d43068b1b39fd108fbff35b8bcbd999ad5078ab6e38d55074c52ff1c656570088460af57a51da4f61669f28d20cfda98b7a65f02de461f50f4da883f542;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd29039341eda83ea5b9d0421b78a64b2b21f88fef9ec0be91099f53c79e7aba641696a85c110278c2721bcb50c4975438eeebf8bc0b7953804d4fd70763ab7e2ef20459214644bacef4a04f5b9d4ac3faa43a2578d991a65ee7cc8758d1d94d3288bb1c380ad39d991aa5d755395bc652201e690706090d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h390a5ca8c7b3f0c4246f8819d47a715e733fb8aaf4a1f65dbb5e3a17a0aa04bc9c0b17abaf06f6e75e21392f3943cc4b72f642d6d178faec2fabf4d9437062aac01a6d8b17c9bf3b60e868e58466a78d2f2b6a45d25b6c729913cd8873dcd8cd0e889ddbd7dd16152e6309f54ccb15c8c1d7f3529636101b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h152c329c66f64e187d00d194a00a6b632bdafbe5c1f9e315eb6e79b1b0d5fb7e0667d241d078ce9bbe27e4ff8fb8425ff9e8d2fa0067f1af6e3b8edf4c9d29221250dc1103e9e79eef44bf402ef2548872ef62b5a90d6ac6e85f0712b9d9415ee01853520ef2b98b2d2c9b1f10cf17da2d5117694d85217ab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1535f40578f2d5d756983d023632e4c27c13062ddf29573d5eb20ceae4a5de9b899b1156f0fffa016caa1e3be86ef5f7b18c439d76e76a9748ff665c517facfa83d6bfface3723a59f67b57f328234387deac99e59b00ad6b69869756b61e3c026df749f581c057d39984c66a5852a52b387489fb217345f7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9cee63e86f42e886d19674e55f0e6c110f1bfcafae91d1dcbef9cd7709391bb0bbf7fe13c95069a5c1e3e22143134d0525954286409180af141238d6618fd0e39afed5c52ee05ce3d9eb25428f8030263750c14e868f71d933146f4391be03c140e9fce073922d29af53fc7ca085b9eadc02259a3c2a1f24;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c05cc4b4b9162cc92218c053fdd00b8ad80647fee301360de006bc151e25be920cb69266262602db880ea7cb37cc7f76d186e2d198063253ec7cd26ee0f88c614cd2165772817f960049e1cf956b54aaaac637b96a1a50b01747a01bed05c44a787eca85e42467242dd4e17b486225df0b7c39cd557a408f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142f37c506b70da86109929551195287aba385729461f1e78f12ebc51a3152ead778429cdeabfdc4fcb924631e9dd144cd4a493e996ad6e235e1b3c6a02bc37c89949f56421a24c7ada86e90e0f96703c23d4bb8aed3ac0da78730697e910b277294fe475a1bbb827ad269b72125704b94eb613828da7b4c6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h124906f3211a74e2110eaa237fcdf1508edd70bf5950b282c958c8ba175a7a93456e843b5785f4778132e5552641a6b43899fc81aee825852986320e50799250a4d98fcfe51410e82ee7dd8e498f4e40a80e7920b9247581e9739f61b40f517bae10a336e821b36bfc04cd398e495c87292d91278780f9794;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61d7f05eb4f61f48a9ae5cbae956f6923684ba4f38b38ebb2ed2dd35a3a896519a9b7a3f36646800417be5626435d47938e17677cc4cbec2cac0cd06bb819cb675440e875d64599fa1dfae6312f6a61dc8d3e42e1c26ce6a1d06be56eaa4906c7bf47348080861a54a472785cd5ca57da3db4f967f2e325;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6cf138f3e8be7ccb01b7b6027c2cc3992d95c10d819a9cce2d98821c4751ff0990d8e3084b9bc1c42c33d33bf8876071c02c5c784c64ba8247553dcac4bbcc81c4a44b8c006224219c4ec40ecf8846feaf7fa2080d4cd521813b5d7e6ceb8f447c9f50cd9b8c213468dd09b95d31107ea0ca99de7d6805ee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1823ce26aa1c80afccff351b240cc5adacd4325baff36a6d77fac39d96c071b9bb184616fcb6e2e472267a09b0bf555cd2292ed8376f2fadc76cfa4757ff7a2ece51a3883b3ec30f80654126568aef5f61b96f9758015df3370a72179a224e6f2971421c0071ee42e7f6d32b2ffc14a10b8caf35881c8ce86;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he8f4e1be509f1d5da6fef127b35ab03a8e46780f44cd7ae0a1cf5ebec8dfef5ce2dc6905a496e0bf20221a6366d9d61061b6bfc0e7af0eaf9597681b2a40cb9f3376e71e8e3394500d4163614da3f7c68a34654b8d039de5a69e220ab7a00b0298e53b83e9a191a09a6d46f6116e4e19e6a63dd8a010896a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2dcb1ab4eaf538a69d4f263c6c75158110dbe3559071c42af43673fc6188bd3d95733ffd1640ad3fd1769a004d40d50dd2d40dcfe31d785f1d750e9866bad3fd9a657380665406014e0b861c2a89e3cf231d99e764671b8a3e333c6a4ca6e55f68799980879b116ea922bccecb500f62aab7c56c8a23eaf9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he3e296b0ea84687683da07175a8d1657f2517980c3aba44061386f053cd557b1e6a1399165a79d9251717727d377f48327d263283179fd7a74b088274601340a9a46413e70c3974aa93c70814d2308f4936f02365ba32afd175035f722837c9ce045e04e0e915c424ca2bffa13f8e7f12c31efad30bc3602;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cd1485b5e6ab75d40ae0703f3a9d573551c92144d23c8077d47728df5ba547e131382af896d2253fc5821dc23c74e0cb0e4b21b57edca2ff6ae4dcb1db8dd83c41ea95bb18f9066e9ac05045500519704b10e9abdefeceeedef48b38d34f2248ab4734c86eb352b6304e24d1dbac71edb2d7ea6d2ecbf0c5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17dacffd63014ace7d59588a4e0fd042e5019ee96e0f8758d7888415e7aa84eae2ca283ef6cde7da27def3f10996049c0a5e7d5344432ec85b254deef6b31f261db58a91f344893473c362a32bce605dc28108dc7de375ccf3ae07508cfc48a4c2e7fd825c5ba16f9d57d956cbee538c31c5d77f60281fe3b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58509232b1a113c002c52bda7344ca4848a386a7a2699c49d56c02713b0d0d348cd2ff60cb14f4c3a955f90df729c29f6fd26d8ebc5cefc36c7c4ea2d4a104b181fc7b886c8bbe7e4e85a5292eeb0932df0eebd815b06cb45b64cda69d79080d3aea4172c1b20eb376db28cdbe2d1445518a72d7147dab09;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h90572693ce4014b2b5f9df45a0593ca70732bad89a24b0908d7d97ffa51a7736e446b7a7e1b273709da4f84482bdf19446f34986e8c424a3a24cf2bb9c8d62423eaecae591c48d6b91c85cbc4b75e1c20b67cbd135b4110bbc8fe47b16ab01a4d8a4a53dd7a6ff207ac12a4e4e46ff746007a689870b0131;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha183fc340675e3339a7dafc306465566254d0533b257c192ea9e8d99df1e2d10200b321a9b2d715f4710c27ff0fb78ce24947223b9d0cd65976aed2ba880d8d75018442503c4d95de3f3e4d17024963ccf1feaf2226f433ae7cfbd2561c6ffb357106b72ba2002119d755052309a421572a9df0b83410571;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd817d131f86f7fb2ad35264291ee508ea59ed1dde7802244c1fb14dfcf01f1383aa7b0dee8a6fb3c10155da01f906f1e8c76d4bbdbb230ee164dd960a47509402e0c302f7c29b538b524763504574c6e0e0e7c77a659e5b19aff666340df4b7b9d50239dcb2c91d15d197d028522fb6a70d04b1f2c2dc866;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc172458768a974b597f77178d7ad91ccc884d678db9209d86a8200b9cf1c0c16280831e81d5bf150adfe771347129fcb9fdfd158bf64e17ea52d896611d21bace57dfaf394507d3ae9a10acc1b8697cb37c028e8d19c3c38d9577e45c4b447426ca962c4da10f75693d2504430cebde6922d4631ea1859b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d60573c0beba8c2e344c805aba6f6c8e061fd1f4be6335e58598c26b0ff2af6d48f0c71f1206023631429f9d99921fb570d3973888a7255154d7a082fddccfa022423570d7f8f6bb3c1877d9ab64275848fc04c03ef15adb221639301776f856c69b5582f518168360e03f5cd6febb2692faac219f7f6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b23b921f00fb195bd3f8b2890174512871a01b81cc1b6694cf523221bb0a4075bd9471ecf51c74d2b9c8ed1652ba6f266c7f0abf279fb6ffb1d6166d31827e22d728f82015807bb8d2ee2ab82ea1248edabec9769c4761ec83ebf686de2570ee39969a234d0f3f734d869ba11dd4ce29c05d9d927ea81e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dbe0afe7b4a8b05ce557f1bddf8ca84299d48aed44973e579cbb4f261a944c3d7612f7608dc8920692b25bfaaaf3a4e614d2dbff0444b79de3708c6dd607f2d627d4766e892a78e9f8c6a30c26fde6edf6903435970e0b8e71633ba15a6dc7ea158d1e4852e176bb545e6efd15f159b300f1845a7baa0b09;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82d4cd2a0e0cfb4c080780852cd5d22ec3f2f5d524dad5965e9715b2d37f23474674d91eccfb728a8546cb16ef6536371953bf550f35034c926453224338ed4737c24e30b8d14226b2ff72ba8fdcfad42ca32d3010ee8d1e09242dd758e71aad6f50c51c926170f4dd2cc64cbf08513040a49708ba2d9adc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e8f951c8d55c197181853b5fbfba570ffe33959587347b1abf6968ee529ec9cc06368c88a3bec1f63ab9cd0aae92021387097a24fe37a2eeaceedc56f660001409599bae476bc3d2b9217db89366d6935efa3b14ca3665d21a97471e9b3caada6c31526cd927306a583b1e19a034a1a974f360c505e138ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52f7404ef389214e819f6c5d84193121931ad7803755062ad52e2ffc76317b92b50c11ff4e3aa03ae2d3e8022d7e001bc17108c435ff5033e1607865f74b2b738585cbd47e1d84fc9aa4ae0acb0ba87e40f56f034ea453b31bea060013e6ec210033c255f800ba86bb34553bd5d42512c328533b342ebdd3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1773314258e1ce543e8d7e3560e4265aac74b27930b5e83a66d0b39ec01cc0f5b4bbecb90e153eaa7b98ca0382f07a15b2ad906527df9c7c486be606988ce77e824be6cc19449b6cae349bc1bce57b233457776387684e21534060b929e9955886bfd522236c77236ca3663fa94e606c9e0ce17b8b3084bc1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15551497c1f46c66d5c06bbff8d6c564842c88fe8a37325aa8c6ba4e6cefbd16cc7ff408ee772b04c71b9e93f8f1760d1cc77be5f2daddb0cb777316a673016a17ece966c84c42011bc95bce31b15c01eb3cf86de0f1f3104a30560de91b17c2386805713181d6ce2b736c6b3b4d6819472aff9b27eaf98dc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8eec87ffea3d6ba4df0d46789c95a48347ec81802f61ce6db72b345c5084e1c7175f131151b694142f9c16312ebfb6df3a1e5d39cb41b9c8216b54db366e8043ad1f438833bb4603142e36525cf771d7fa3e6acd71b51f3535c31bac7615a021936c1decf1611e823845c9a34e50785af5ecfe2397cc1be;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd79954a560e7157141c263430c8f4d6c5e08371f4a0f3d03c9c59e793019383d9eeaf024319fdc858b5b9f5b62ec38549fd5e564766761434d958aa55e10a39e0da2af6ae8ef262aa102b94d3e2b4b8c4c60cc6ecba80096c64801dfaf691fd4c705ffac78494ad41dddb8cf1a12f5e7da7559a5ebb057c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h92a7dc93217670db53c80e258126bc90901d963e97e963ffcb6a67cc880553e2f9a38041cf4ba80274e727514a74646eea1dcfc27d2ceb328bbe6a444e6ad759de9af3d8e1362f6ef3821d740e1bfcb9510c3949a453485ca0449799137157f47138b532e41b9456a3c0223171b457c5db8b58726feca97c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb822865d494e5b933307129a7bacbf0e7874ed66d4585efa6a1e5e827c138f8edecb8e4a1699aaf46575337082ceb0241414a6d7b6f8241115bec155bb7e1f31ac25116fed0300edf4f420bf0142f5689a4c6c7d70fbe893e4bf934165292516c6f96e87f00ceb26641ee11aea497b0889038714765974b5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f9de22eb365d78eea28e63110e6fd9dc4a8c2486a0bad3d5008ecbef2342932fcd98275eb00aec821483a9d29b1ec2325a6f673839c2a1b79b2ebb1cf78797e748066b1e92ecf8a8f1a9c54d7027b668a74075ea2cc5d62ca928d8035c400442b6552180e0f7e653c6e3b45ec92260a30c6ddec3b3dc750;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h665c3b3d6255d884238ccc195bf3308bf79ba1de8f1e51191484367ece5ed8eb54fb9ca9b4432af24f05f362059be841879a5df584fe5f77fcdd52f631c4d5b97c222f7efa6ebecb5713e955eb0e2a6ca135d8801ff76c5e289fc83e09ee00b7b451eedbc97348377b5ffedf6e264f96573313029a1a4844;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1594c0af542a902f3126f2dea250e61a7586d8a84c7bcb88ec25e807ca7ad4ee362df578397dc199febe6a93abd9a0cd88e7a8655ed0bb6cae841e80ca99925512f1970e50e2e677c34fe9f4885a16e64edb1f2a8b446b9f00671b08b0e3633a5bca156f2300cb6cac1a102260a2392d20c27925836e9609e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ebd938edd2f9795d85bc1947c5c263f1da97f39825bc8f09c079ca8af49ee2fa066095793c4b269eaa3136a7a40612084602df07c730d7a889439ff7ae49484cc8e8f9320c410676d44e987e349f1790ed2d27e761538169a319ea7118cb35263d609b011e372c2f305efad10908ff8365a0d5b1277e0c48;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1abce8e7ce5c23ecebe05a797d8137248b1ca93f1bd0f167b6d064feb266d7dd011353d6d064a0b27526e6e7b68034ec5e59250847ede424386ddbc708ef13ba84a2245127fcdac83745c01aef5c39748097d232f9539cc96bffaa5eca4a3dc77f2343d244b891f9c701c042a24dfe68335f2effd66631724;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6845dcb19fd56c748622f1de30d1c29e64ca4143caf9b665e75fd0365c784e673177862288e34586d1d80b4cc436085e9b5af74c22388685ca5413dd121c933d2a9314414449a8095220fef8d19ff1d0eb1a3123bfc9b986273f650479295bac315ccd3aac6eeaa40d8e89b1e37516f5619c01e5150a3da;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfd98b74457e605f79f7979390b5e930f005c2bb5f152260bd8d027a1e57ad0ee5891e7d43d1a5e3afb19f2ea4a33e2f744871156c064f7ab7ab8a20857b14bf1763b6578759f9ebbcb1032783aa3dcf96a42cc2b8fe25b8008f6526222cf958583e3296015a129a3792faab946b4d3be20ad187f829aa089;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha94c1261c85e23a2f65a2ebf990d818a9fa6d9415e25dc532bb709241ea044a1910bfb05a75fda69373ebcaf94d9d7747747b7d1d4c3b086bdd9c5be559be9e76acf18c85867eaa205ed45cb996c52b9e269b1f6354f2b3d305627605b6965fb6b8bb21a4b7d30cdd1a027dcbdf1ce51b917376603334cd5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h726ffdb8e6f3bfc2622ad7db32b8a670c654cb62c361caf92553f309216c3df34b187fba2f5b09c88ddced9159d5172cd6d1b5e464a202d2038b7e1d4502ab397438dfc4e3d1896554dc90b1219605afda5fc72a570ffa6e82fa161d4c44b5b9e63f4980e0b45df06769dd8aefa9d3e1b185436c67c01572;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h63f20318a21c70705720acf035da6a2d58ca3805d4a330da0e9f2fb8c306c568b6e2102b9a9f2b109548b45a9f9b4e74162c65a86c6254df50e3df587de2f81974d3d346e18816b3aac10a3172a369e607fdf10162cb0e53ece9dabbd2d780479f1e628ef97b65617c26a1f1620838cdcc3d6d0bcb76bcff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b00f14596fe362945ba94e21a74201106f0290fd8f10aa7b65f848d53d7ab3dae18020e1858ff8f12ed6fe58e4ced3ec7db37468b40e17a887dd982a0d7c8a7c821f9f69120547fc685c8f9f42888e5588143aee96f8cddb9506139942f83f593f4e7077bd0056e942ea0f516554513edc9dcfd999d4229f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e9985fce53672a3c962446e36127f41e959dc59b61b6fc8cd9226c18ab5cc9877bfbdcc80ee08614533285b8608aac24ec304452f28dfc91cc96b6a63d5a7d96f04c164c8edb37b9f210e172746515605f68247b918ea0e4207799a9d3651d0cac7ddd6490c28350198623c3706175add7cacb8164c6ac1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc2a632efa5f6c43e7ad9b1635c3f4525eaaf5a868b94dfbdea4530f0dd651bdbbb5dd14508073a135b3e19109e629ed56221baf76503f0655bdeeefeb07d0c1133e7c65174dce5ebd78dac2c0d280eda83032ea706a19b5a2287548e832fcf6b2286e11cc7450a7008049e487044dd945d9ada6de28ae1b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h148c9a676db2af4069247aab27d8fb8d5696af652fbf595ba647b4ebc92cf1d34f0d0fc2449b410b9833d38aefa7cc459f3fac71aef8fe139fc283fe6abfd3be88b1bf2e5f66c957fbd79ed453e882b78e304a581e27308675e53f1cabc669650346af44c0e75c584a388a4bd83add4bdc3a8ad02e5630074;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b259e9049814af69882cea4d8235a898ba05471ab23dc15b908d1ba057e74567139a414f3d8a198e7111deceae0e093be6be4b96dfe43efdaee9fa8b21567cdf8e87320db3c3da8cf9e3f7abc5001ed67aafa69aa073753f615c2d34f04ed7102c54d65654cf3ff71d131065caa07e3b57364ad420274ea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3421ce90d7b8cd5ca2fe36a8d3d890dd9091cc8d094a6259f31d07401dfc1910e74a861b4740b5bff8b4771e3adbd8f443097a526aeeba312a171090ac2b56999adfc276763b9751dcc52fadc260188122f17a68cb11781cc613da4223257144706c0f69d4134efead3c8f296a6c1a07c6a83149375165dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc4e1a7f1177de1d3554c7240b81a3dc64ee87255510e961e714cdc9ec8cb0b511617e8a26d639803c0ee79bf8a95061ea148fa5cc3034742e26b18f1e9019e59eb18f0070530dfa66ca1227a6309f2dacd93a3e72ecd87de2c30fa1c3f7a1fc9ca5cd201e60d6ec5fb4dbe2c825c0834392aba89577c3302;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc45f4174490fa40d0a508ec4ebe9d65989fa517cc60faa1e6676f0c880839c8c3f8eafef67516fc1b788c7f539e63a81bc79f14ce99dfbf9c8a2d01d6ca8e951d0e6729dd4d6dc26ff15c1bd39a7c45c1dff57f529fbaae636b9008d37150ee54a7e26e21fc6ba7bf5ea45730318642bcec280146e840c3a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h99a4c958e9807f421be29288db0e235b346f2c5be4fca003722afd8380e10b7889b82a249ba66710073b5679fd067cef4744c1060e058ec2066af0908a0f21fc9cbfc1b1370818eb71ac14d1d30d987f876f828241a34574e9af68577792d9ff7b6d0b3cbdc04e7edc72967017b89f50bd9ed29533fd3e1d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h918694dbc6fc7f571af67529f7da8a3734b26666422e326e0f401492a3bf191e0cbf43cb76cb824efe0bfd2da4567566d4d38be71bf5da05fd6dd378ce3c4cc8bc98b56300a4a1fdd51583b490865624d6bd360b31b31e2541bafc842cbc7595314dfbaf7c8809e8c6c3835db919683adfdbbb77016afa22;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e60c5b808cc71dc651c5a24ea709cbaa6a49d4f18673c63047a5f807d0fc119dc2a32b000003f1803273f11d8b4aa6df1f0e62550c1b9dab9b13c6733dfd5e9249b8b288f4b96c749d3f949c55faa393b07e9a1d1f12dec04374e7c14715d1381202aa518d9f641cac3c9b7628a0f960142ddd933b3e78e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e2ffe95a0964d09590f9305adac34451f810aef6449412cc950d9e10d43b3253e8882b350172adcaa9823f7aa4db690321ecd7a822ce107a71ed971078c3c074dc8e00809b4ca79a8cfc4cd7d28589b78100c98dd11e08aa5b68c73acb4f9de2465729f3a8338fc84a0a7a97d54d782aaf1f5c6b906619d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1852aa488a97b99bf3ce19adb15656a6e747ec3a87ca33a6639a78a7ec5b74d74b3364a75bc47908c197f73d8b670826519e3e1621b2383cb6a383b131b5f5554cc4b6ad8aeaaa829da81fc58f799a257b7bd128ad6345d114f6d43ef7667ea9513cce5c5bcf5753657a5c34416ac943ea6a924266f520ff9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h192075a89dedc0186d2fa9a47621bc31ed4696372fc085007ddf6e1fd14c030091f1ef185e2645434f9090e628cacf3f93dc333db66b5a30487eda1a6f7eb5df3baa5b51874729b8c23552e8d02250ea7e7613ad4bd6c3fe90ad947caf21997c2f06ce74348bb661ab2d086c1f936662abe63df8c89bbba2d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12deb04280eb58509d286c37ee451b55d810ae26188707e3b3c9a3d1be6b6f277b18bc8725f3319358c1a6ca647a0d13e8c115c70520fd4e64a89f672ed371d41521c272f53f109030d0f9fa3ed90ab2a55b8f42ddb5128cdbccf24a9abb3735b316245c1b8faf638d640c315ed4bca0d34eaedc11304657f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8b828159912ab116c053c88f9cb7564a0c731f61a5f17682cc27362e73f290c70b3bcee671ae8076ab1c91378cb0963ce49ba71952b1b6ec9771b85eb92032bb3958103cb53abce27d5cce62c509392889891cc27feae85e30d81a857e67e20d3c42914f7af65772fecad542038c813a4b01519a128bf5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19ad6fdfc06a0aa5bb5d478487537eacbde0d32721160a240900ad6031a7f87454aaf7a4218c9b60dbe609091ef6ee7058b033770ce2891b520ee925da69186d61b18e291d51201ee373778d6d41cefcafb04ba12baa4d65fc77fe9428a859927258a6cc47c0e8f6b38030039b3f4f3b3a03406ec9d8ebb30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha93f36544f5fd11cc9ed80865e59d17e66b6d7ea7041a3d28eda7d6dd6032151278594f0e468c390ef264d2ddd21eaa7279105288a6200bfa88acd311bd233d1b23bd1fd6a978be06f72538182279e4a3bbd9854700bb22bbc091162dc30957e6547600fd6b1c50b9983e47f3dba369c4ac1c143b7dc1eab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h653f991e64b3a6999167b50ad5b4f818845d6c12d88dd82d5eb421eca4d601699a3521bb777af290495e17558e244c1c62a7c2a3857af6a9295a6096e13b6939a3fc4f717f1c3f4c981017ca756cfc0ad08aa7dd5b39ad41ee2c1d2feff1274701bd917ff540fbef1be6970010b29db6f70898c8f313c5e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1abb5465a71605d0556be6f5c9b855d7af7ab394f55742fd491520696805a77ff30096bb9780f601a9755d86e4f6fb59a36518db231c0a4b0f9207adb09fb586cb9f3b6741cab4333a5f9b5d2da43314d5727dd88c34704509f93d22c591f6a06913d9b6448257e838fb77795904a93b4f0a4fa246a3ce74;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6202a89b0186be245093c2b3ef99ab5b5bbb16c489394729e8bc44f6dec32d5008017ca7098ebaeaa8f2d9e7b29d81df01bfe4baead5881f401f74a099406f44cc566bfd4a392b32c4090ead05b2ed6c64b3993f00a163df3c2392bf5559ca75a2cc5a1d53f8b6c565da9bc5b68acf69ca7e2560ee742921;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc6c975f1c720e6fcb77b8d8a3853ff6a74b2008d8d6c78958006433d4847834e909215fe4562eb788ab91cbba94546431e661b49a294de979132675f26a299d9986f6c43ca4d90883b29059eab5e9fbab8acb259326f14581cb3bf72dcdcc89fb48a1047fb1e5db7cd0847ccc5c46020ff82bc93f7aee732;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h370eee0dd37e3942ff27d91133de5716f9333c6142e950e505c7fa208e3ac3b5c3c33da9a02cc272236ed29b346e368a1e97f4861b608847ccdec55d83f63c5faadcf3c56e88c936f4544ec278b6f9b1fc73df13a209866b1de5315f807192228ea88d28e5fc118f732e9e6478c64a30b256a64fc5cbdbe1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc7fffe9d86f07fbba5b18d9479242595c8a62e8d939895285f637e06d9e6d0b130bbbcfce3ae87d2e8287889f76570b86392e3f7cf864802553a8c54bed46b09873fd0854a122cb49577bafab7a0c66df4078051359729c1a112e2b07907921164da8551b95da5f76950020b0ebd279eb3c53e9505e550b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde2dc86230323d7c0ec64b4209bec11d0070861105f5bf2fbd1a1657756f855b9254bc5b2ee4af6d988f9d7249b1ee6f2e07f14fc6cbbe759762bc2ff6ddb49c284bb1452b3bb6b772b5d46cc294cf28c5b3f7d46708c089c3e0375eae0bbfd2ce92373de5960a01f864ad4749456947f5f8f4b722d54909;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18c470b146f9be153c11ce007eaa73b2d6a3d7e1dd13a5bae126a3cab10cf3ac5dab02c654347060623d51d6af816123e943c7844aca0f0cac4cef55abb13ee09cb81178baf8167216f92fb033826be8d2b3763d9b8d6bf94bd2327add784424a18e802b4e07220dd498566e495570a0d2b4afed2c1b2f9af;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cd80b844e7e3032cbcfc09479c13caaa2731a8d17c012d91c8185837ddd1dc52e336896d355171622b830266ca345e68a934b542fa539c3e52e10f59a4113335ef49bb574198811ece4d70812257bf6f81e445a2b091924118196abef6d4b84cab70cfe408ba619fc7db0c129a6f6001fb4eb019af70897f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cda98e8da15223144c1815c7ffc93ed7ee73f7554fa4fee54b4af9d801e1919d838f738cfd32f40a580105ca663fd5ca5c7aef6cc2cbbe7b7b3707cb40044b45e404c46f4c4adcb57df668f7357ee483314bf945474dc3a7ea7590ccb9ae12d1f106692fc264669401401bf9e4f8712c9ef6fdfb5e20c2b2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a06e5705a39043592bccf494e79011bea6bbc0edbebeaf6479a61a12a0038f73c4be952a793871dc19c86d1258acfe3a0902a6f2c539aa38608539e45142e53262f841002f2a5b5ae3449503e00cb5493c82715de76de3e352f56bf101b43c24286e4da06329ab2f96ea180406da60d16642d0fcb4ae3fb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haeab4b8f6601b3604fe2931e1b50b2be60cf1fec852902a9b8aa1df1e39e53a58ae988050d674bb21a53f8fff5362606b29058d002f81697aeff438da237dfce9122adfe40dfacbcc14706cc014413942a64d186ab0b131bbb66eeaa1be82133ecb108e879290bf00e4d2568aeaad4af52b9006f4544f8cc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h122716d53110dc4933c893eb4e4c3e050ff0f84e0690c6b1e5446144bf9ade828c40fde2761b9b526cc5dee4ffe4b2dcb99da24b58e0e156ee59dcc0967e0823eafd1f6fb6c4faaf92d4b6150a9fb652b9b6557b2a6be010a0a3b04eb5fffdd81e460060c79a49df8df031666df1f30ca14480cae6644fad1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h155175bdacfec6476abe5967416094954ba063bd8d1e6431b19a64b0a136b880c677036d613eb77d94197ee15f2979de9f8ac2b00ab566ab50f81901d3649d3269bd3417b0604adf374437e9db85d000474027b071d3ed16fbe69e39dc7dfe6334acc3fd05c04306d2734bfcf6224c47c6168d15246a0a24f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha6c786cd3e0600c32fb5221c7e66cdcd2cd1ab1294a8aa47455687b03184c0b7e769e8ef2ca2f00cc2fbd255aa5fdaa2199f9bcec79c48a1668e3b9ea6b9aba6b9faf8862912c2e904a6825f5dd8568addf35f5fccfe5aa82cbf58278cec9330359374472c802657d99294d75e1da267b4d29d0cbde91c70;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdddd68c02099d7d302d11a25dfba50e10d8518ca574389b73d55d87ba2ecf07f95199b3bc207df136981cbc0b420bd5f89287fc590fd84468345afddb129adcf02fe33b3f002b86292f39aa672f4eceb4f9d33cf3e7f1d91db5a0b37d5d74c749b20f5e853650b5ed237b4593c276712f6c6192f4c860b04;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3feac501747affd2b19376bf4562b4293d8eeb2c3bac18324d023f2d0d14b571019e59370f0973b44f1060b277f191a82a7137bd3bd0e60caaa964a0e91c7498de292d8373b7e4db621c0456b905d5dda788f8d50e8cc1b2175bdb80af41f35887d30f12dc81142d43229b849f96f29f3ee34b1a5f78c380;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15eb23687cc153122b4e8c5b1e0f27eff6225a74c8184b730f6eefbfd81c1db3275af0788824ca28cacf160af001c62871bcedbb29571a9884bf768a8a90cb223dda9d70bf8f9453e05ecf8fda29be93c469c2c62423c50a2bf192675371c9d4d97af94aa5d8606a709d8cd0e8778a52f74cd10e67bd13b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16631643028659aab7fb31f4db8964e3be71da7e9142d629ae8055f62ed20562659106f496a317537af02ba364ca4af0e7da9ed3a43d6b4b5787b73815465082e2a6d0f5512040205ada97d203fcba6a46a94c7131dabedbc5422f8209425d9b354ec540f7a2d714c77f17bababc796e692bded8dca95ce68;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h111344dc5463275627142fb49cf951128d1463dda3853f1fac114445c1d1aff3268ee08968b00583765a8e06f59d2bbdcd15f07c6fb344e32b8f2f720badf43f9597c645619931362b664fa7c207ced312b311964669dc5ec993d234b4f3f7faa4944e08ca959f6d38ccc8a4390bf0da54ef006b1ebb096fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hed969daaf1b436d6572216b666bbf39fd0ae662894e641db9972ce270c5ac5271685b34b9eaa3321936c98aa8c50e6ee5b61742558ebf887f7ad4afe9a6ca4d7f7c92a55ae94c79f75f81eeb671efaf05db1ed67d4e5f93a7ff8155d51a815d61a766a50b25fd3be514e88e0fcff7702cd5d71b60b17a66c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcadd56ad551e5f393537d7ce10ade93c5983f5eea7110d895a948dc13b30aa49d6176990f298d691f0abd3a2ae48160f71dc8996ee54b7224df40ca1a6f4d0dec28449c8fdc783b4c188b53016146841c2d34b23d7e8ad7630eb68abca9d9a29cc8e26831cef30183d92b0332c985d0b0ffeceb183cafa8e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h30d1297219d10f0241bd7a9829ae2f4f27526ae370466afd060c57a0df1c8befc918d96047517c6a7b3ac14e1d144ea4b61e29859f39817a8413c045a752f39230146df1023d7cede7d6388c39869d97a2329ac51adc7a2f371f446d00a9aab8e98e2d80e4a6e242a09da5bb458d12f00ecd9849027c90e7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf7fb33943fdad71b44d9dc4ab51fce9cb6bf2bf139f22ef75aa1f29842ba4cca85873a96bd54bd86d84adc09108b0d7be9d8a286bbdd6f4a56406ff80cddff70721f4737d150240801eb8f814e0d8eb0616f91b3204fee9722f5d0230f8a81555d390635ded0ad6d068e33ddf876bf3f667fde60541ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h194267118aa00b3373812d4296e81d380f555e380868f206258b6c767a590d7044696a2d1d6f5aa7cccb206e8fbb9cee3922075027c36105e25638bf9396d65bc9cca0179a24b7c031608187d5b59dbf75fd3fbaf023d1d78f9bf7e620bd85a0967295588c620470fc7f7552c6783a80a5240828312031b98;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bea83f1ec05646b4cedf0798af0ded51ecd5da0eec707c421b00cf442d0b27bb4ef5bf9e40df3768f14766cbeb5556c82ac955760da1ee5c4ec664268a8c83fcaa9c339773d1e651bdbca918cdfad9e2b80b8c87100d533a68e72b4c6ce82120171a193b1b30c1615db5aa216916b760696a43fb00804f72;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b8ed6d6f76a099989292ea1fd3d31237fec98f40a422f75d21ebdba326aa642c54d938e392f615698fefea56bcc1fc5924e3dcb3e4a525c2a35f145187411cd5ea3b2bb524af60a13f04e30344f650f8520848183673de88036a940d82a832035a67d03fad2d2ddec0a5bb2b745eeaa96564d21b4c7f2c62;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h72ee290349ae3aa35f7b9d01ac27eb9b474fc0d7b53b3d0f3cca804edd2a6b0e687abc24266c6d08f14cfc17efbbbf5a47ef8578415965bd23b48499f6c213e01448e0a7d619258e8697276b680a249e4e695daa8d792788d200f3f54da459bda87b9ff712c450495296471b82b40bee388d46f6f57c7bf5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfd528ed18d3f8116fdfe92b922eac175b149cfef5bcdc5850e37abe90e7d94f64c7cc23154293965c1c9f95f129795bc62503fe062dae04893ad42ba204f52a70b59399ec5dbd4d3e3a8244201b566eed91d5115801afc573091e1219f0cddf10bf8028886f08efe8729d98a8436a61f331dcf194b6c1e71;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5925f0b0b46fd9b96cf878ec1d40fb537871891f8836b60467df29f23cff6562dba2dd2d75abdb82a6472290ef11ae998130b2d88233c8fe7d9fb9a332ad9b1a554abc1b4bfb2710c01e5e8321982a1ac1ac7c8abb3634f53c154a3bf11edb0a90809eedf3dfb86802d7e24b5c5f0d130e3f44c43200390;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1833e8fd5043726c7a93a653bf6abc17b8f6a566423e97763993aa930603ee5174e3a9d10e4d55791453065ddad146801c0fb27293e7d7be2d4805885ed55e22b94388c24d17b17800139d12821d25be4da0f9c608d5c8b30e5a47ca27362ae1c188eee33ab66b2bab4b6501c91f2f503c5ad5f52f7c73f43;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10105a672cf40a98d5395fc98d95ba0b5fd18f7681e3d5520275f59dc26dfc521af8f21a4280eb77f760110c92a2df48311baf05d37286b571eec5c063151b92f4125eb68b10072942d523684659b825709e5fb8ccb84f2385256a6c42c5197ed4f03b0fb0acbd64e0bf4cf22090622250b1a2b84cab6c1c6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a663390e6db31b9b3209214b4bca4b871bce6a6c6048652e103aa06ea7d129d730c5f75043499d9ff0f97ad1dd043f194c5ec9261b9fb5178688970f75f7fcddba30718d5ace7f44f0b22f8814523140307854043808c56fad90a62904981c45270b38096db68b2e3fc0aeda80d53f4de87fefd19b5f2b2d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h64d7312ba93ec4633d4d60be976301483e41bab5bcc741412220957dfc22207e74f17182fb41115edcd3a7a7fbd9a136e1453fff4f511dad5579bb703fe88ca018358972d103023d7c616abeddcb908c0df8581a8b013ac6470f328fbdf842a2477953c390beac17a217d1f5ad460a4283f9876e52436238;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1012a82ee5dc54597789e571bcde72d92d3483adefffece04e72a895dca097cee732d63f4e356d1574575b7755cbe3ed1609f9ef51b415f552f91344b8c4306f63a8a7ee12768f61639ae35b21bfb2b6409c1fa0dde112597ce83dffe979d178055fd3b7c1e61bda4d4a453a3150efc6d90a695f61feb9e14;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hae1c5431ffb9cd9c74b917bfcd34b898bfed2b2fb111c95ebb48ee7334b1da702ed8141d44bdb87724b5225e12aed39f0155612b592528cf5a0d5c09204a1e27cdd1c9c7974d2d0faf99f85a0f9e5a128fee62143f637c45fcfe482d711b42a2e89c2a51ea707c5cd6d24779a46551579f1bad78b6355d99;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf8dfb725c30c518915eb4174c5c18683f097ef94262fe02600e60d770f6ea40cad9d25827a7c23588b4a2d3eafb500ae145c46c622e050c1ef51b70f0bfb5cab5348d3401800594fafaf600fddf4b1a1151c5f60fded516873a0bafc16f477dd5f253dbdcc13f3f21c1d32c6b5b364142d1cb96a81d0534;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4151d598bc1ea8a9d6f4aea0396870a85be514406e559843df802eaa2bad7a5577e5de265abe11760b67d20b4f86e1321d01433e1fc64f6114d465dc425349232ed08d39de384c15c62c0a00d892318cee43eaed54da93c478b844ff4250f5102d25fb420bb3f0f822cc8230b12339131d94014a44baaaeb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6193a97ec875daf5f63f000e96c6ccad54c1f9307fecdf14e74636e5229708540c65288e96fdc5fa88320bba4f781ddcd5f46b781b242d4d17e7b022352672d959d533fd83efeb01b8417289902fb81d541e163b714c64ad0536082e5940922771a4dbed645d938c20e333c958f69a5d06900c59a0621e9f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1793202cde8f9c578224674e369d8273a64e5d084fbb4f01c8dc40e8552e32e65fd5e282d3968dd1460a4bb9e5a5329f894650a73422a46a75eda76d365f6bd7c48db9a6f85c09fb91c1a8f81b847231652659dd077f5987cd98a0e2a2e10e2bec71446cc65874d7e34533ec8ac97c233529dc71a484d4e88;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h592dd12328036ee08f71a0219caf711cc3ad9ffd21b6ec72aeb65f0bd2cd5d58890daaa2ab2d2d423bc6ac4a0d8860b723eeda9abc5eff75cd7d3a9cd066f5505b3d0f52ab61f6d3d0e0b7f15455918ef6209b4b456eef003b07dd728e72f24c4641cfcbe3768022d40358e0ae27bb22f39ea53595747547;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ac836b5da38461facef30f61a56c4e6c46387cf2a8537864532155272a05408017588a34387fb0a019f8603454d3a94e1255fa84152149a77b0db84123440daab793e0970e60d1bae43bdda1d2551eb314182e5654477ecd9501d50ffc8831ec947bdba336319ff69a74fe8e2c435b6362fada35e4241d33;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fccd0e231ad7b598cb8e4f5350ebafb34e957f826d3940b9628f39fe2244370eb35062eed1f54e4466991f8473bbc4c15390b7dd1ba0255a48bbb97fe5bfbf8696a8120915b412eb772db0824615ec1e4a5e23cf853b8b6988a839b69c8459353002439cf99642db3652b5a4b260eeda3943b8aabb91db17;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h745ab58d4ffb8962b4c99a4cd46f061ba862808cf01ab681e7e121c028a993696a7d8e32404ac49a65e435a49a688b2f0216a47eddf9707a1e4e45bddd1891c4e75589ce7f7504690e2e872246c5362fbf1febb07d71b73bbb76a039b77c4bdb1988f91c05abd84bb0e16fc20b053fab8127b75fd36abe1b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71fe229b4b3ecd236ea548515e7ff4830611186075bc81f922eb369f3f0dec88dc2ff89335fca5f9068ff4e350cb85e08f33318db6ca98dc078a6dfa9e6de7aeca63342ed2359c6379650192539f26c21b1f9bc6f12518d5a383d9badf14a31de3ad37fcb7435e8ccb6eeb312029ccfe8ee2c4230e4bf7bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h103b28396a81481b7b01f28215578c20a0f42594c715567f9d8dc8f10ba211a92472702b1ca2e8333931a770a20b269b77ab510802988e03073ad247c17628b488d4e7e25aff8ece0b61704c7e8d1d8ec8a164b939e7492c32fb1259412ac0ceaf99cf1a7637dc3309db8efcdb78630ef95c74fedd9f7a0a3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1635718f8e3a1b5835a3018ca5e41ad58522d2693d7319719474be799fd80436bb6ab293e2287a2e209840e2ba408d444a0a2dd046b1aaa85a1622c702d5138e973f7197113cfa7d1003552ec464ca1c558184a871afb4b780e076543c43e091183a063f792468ae7b38b87afbe469a97fd5193c57941c3db;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2a300b339736ea1ff0d29563321176b7fe1bf64e6f69f2ce98f863984f109deca50db456cd6483e060d1495ff74d78961f365997ce045217714bc5c68dfcd1d0811fec74352e543335fabc1f2dbad14651d64bad21f8ccbe4d414b6f32481fd8d7fb26fdc83ff73ec8be9272bd1b7a59053c093ad3e592d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h20a816986378d2c477e33a0ab5964b8e0983c76ed3d543a1b0926375de5a47b1e63ce22c7df107e407c4e22b928190b013dc650574dcae29fe27235108641964c8fd3af31e5b942e3c7099ed56d92ea9920c1b15cc6dfef0ae77ed43089e87872dd93211f786b7b197109bdb05393e6a133ab202ca9a371;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd30e4d5c1fda42a383c9671d3f4401373c185adc2bb0910c5a79b7d61fd3834b53f6e6de62cd5c4f29c7efb1c7781ae38d6370a74ed129c472c99cac82fc4d2c93fdbefd1fa9273c0b140b097ede85a6eaa413823f8598d29f523123e5fa061fb51fc91e6e5291195355381223113ef8734b579058dcb1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e1f6ecb05eebec42dd8bcd9b48954b8126baf1acd560eac5baead616d45342baaf0f1de437413ea718b847ae17ef4bad0acba5d0c28a13837c766c0c3bdc5ae3a6e953729589f44e2cae30839169683d59b410f60358587321a3c6c2bb2306c2f4c41e3011219543f8b8f8775cd7191f6b5c555c382ee828;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e653fd5ab7994a34160bbb3db5e6d28d0f6df3fb32301cb2c234f759efdbea434d9b0b2cc1f9d9506eb6f26ea48d56db95b68fff5fce71ef67035ae37b55c785bb01e9e828ab8240ddbc0442a202a0ded0c750d92967c3e3198120b83eadb4ef176ebce478609704cdfe53544c12be250f81c87e4f5ec37e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h46729c98c5e47fc620307ca3590dcc552f7969f127b429acbcf61844464790afde6dc7435f8b2e9ca602d9e3ba4ebc2ec43a514055d3714451aab437e345348b5354f44355a0d25d9a1d41e19652d53785fbbfb340faf5d8cfd757801aa1e81674adbadb91f70142f593e5f6a85ba96be22047ce1580d3c5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16375cc117bf2d792b11e80eab6fc0c50591c209a2ecc1152cbd7b970755ce089ada64ad002ae996dabe5259bc3e7c3ae1b9e6cbbb845126abe80606e86ab61cfee5f96c9c25a66c87b7881264e1312089b4a49638b4f96499212f48c4ee595992d0716cda9ca287fb792c90de60aecb8b76e952993502e32;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h34d71664dc34b4c776a239bb8fd51dffe6c5fc6e95621150bfe75a701585321a2035291818e02fa323dc145d6f61ce0795a343f9df6ca7dd4582de1dfb690f746ab959a96d1274326a66be90b39cf46339645b964e8bd846a0034db29ea61c612f58821e2fe867e3c604b0e7b66e4781a2568113c98cdaea;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h652de983737db14642d2a82e9f7d3cacbab43b334d647f19b9b21ae73ad41b8946f73ad498192c93b7d1886ff003099071ed2c9bd2c8d88fdf9fefc860b1a1057f4e78576acf5e737bf58b4573ede93e333df2ee5021cd2d591d06e8e33f2fc20b0faeea85986b42a67f50a040800dd3c805714fe0fb7333;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d9b985218c693d9d84cefd4055965ca6b86d5775c7f10e71de091d9100a76a1b5c89d2c365e9bbdf74723d87ced9b21080885a12e8669f74704d62a683f95ba7f08ff949e7d42a9acc747cd1506ea922842a8358963ba1196a826c826eb192fe778f0e1e02e5fc01b9bb411ca580d6550999e78d8aa8484a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h23ba2986719c516fb9f6bdc5b78bda1868db8d1d0653fc565f2440b8946cdfd5495b2708c258c9b5e18606ffd9744d9eceefc4a4e8495411cb326097d7bfb3c52f622f667c10ab3872eabe4febea5d0909fc7ce71c47b2ec08aef1cbdc7a818215fea1811c5d745a0cc5d50070d735c529fce4f763bc05fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11fdc4c5d68a9bd704937aa098cdc03fb105e3aad1f14944e369e2d525211f00bf4ff279de637e689784157257dc939c3fc2d9dfa9121db6f28a491dc00a3b6e9955932d33ef9857fbc2a6236018cfef47311c96233045ed27ad5b7b73a1b7f0cc86ed4cf5916e67a107d4f473bde405c071f313e53b81f64;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14cc4d6eacc803f68f9324611829ca19b0c195cce7e89b4708d0212c8931b5c0ddc572a09be8abcf0b899495fe37f3ff1ec6e369f4f72dd378157d130759d92a6c2907f3ac2c25ad0825fb3750875e1db0c26ce825b6bee7c57f5811c6aeb3ea10c8d8f260bc2144ff866df8b934abded47ccdc390d61b65d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h29c621d245e7b743f41014104dd72c932a8800119714cbd609cd41da70c814be547a1ea8fcb7e2fce78671cdaeb8e512940fc5afdbb5ebf3ae0df93acdeef908b12e3e18c755a32a4a2b3a526a053d054e1198a7b15a89f3912741419df4cd85e841f8da8026d281a23f8234b3a01945e83d4919b5e8725a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de0de7702589d867a5d1e27f4ed53f88b62c11a0a10f29b79f276a91b6f1b4bbe451e5419a37b3b16d48a8e1bf0baceefe8de94823187870ef72b7aaf2a96f726ecee8b8ab3c8d840d06a2b80b4f13f65cd75c3a5c84be3d21e22282147af475beda9144a421814c8af35e8225268d69c2b2b79882eb802c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b61e8d8ef02cb86c8205aafe657ac91eedbe5441cc457cf37c2b7944b2dc30f0a9efc0cdd27c147d49b6f4773a8eca331b794adf33870a48699f61f1bea101ed93f4dbc4a91ca36e56aeca4ca116c00f97364eab416b1fd040f7381aeedcde92e17dfb3c0fe45632376f14c5fdb61339793af1c78de8a2df;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h89c323d923878d96a3be84c331b4f1230f688af094381dcdf31828787550f0b37b007fe53f397acbe4a8b51dca38554700bf08a2c42b78ff9f9f9a21047cd5658d2fc5fc874362cd5c07cb7ecbbc632e1b8da36c0899e57040b3edf0d52d03bfd190d421a02410aaf7a7f5e099a7bcd9fd604b64f56f234c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h44c9d3182d3e75d9fdd1555574b601017c67f65810df12cff440976a672fd3a6ec8ccf45ded87f8c8ae2c7c9f947f40c189d9ad4ead28d530fba52ed1002f717411777b0be0ad486e001525b730f1cf11773643f88f6110e4ac23ef822fb7007c574ff968e253829bc8d4bd4cc477f90d8912283dd2ddbe5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dd0ba59dab6cb1103452f27f66b5bb598c2c740c4ad60657ae25a2588a7114ab21640b244478f75685088db7f0b5cca0c6424ef8460ccda6e32962d8fd853f41e0ee2f6f7b134427fc12a08acbe1261a3670d1400c72a87877065aab52a5df6ea0bcf334fb73bc46e8a90d1079751b143550cef07cba2c7c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd785ba79001ab2fc5b389fc800bae243211c80bc3a1722174f37f03df70c499a88bec3cc8a1a28a326d8439fc61a1f06634705d8759d4566029656ac80beeb86d1592b522021acf05d54119f55ac96620fd3dbc54c60ade42d78ccb153a53e7121f24d9fb0d2d74867f0dd47b4de188f29fff8b3c94e0b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h122c36aae0f18d33a8181576cbeca65921ae198fea0949c9fa4c1bdaaaab92eed4ad79f8db73ff90dc21bdcdad0978991ea8b36469a24265601a65706085e91b890ca7d9ef308632665a9bb2c686bc96e5496625d5cb985f4f3c05a937bea00b6295a92693754f03f7ab7d01e5ef937ce72dd2819731e5734;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1371aa933c4f0c15911393ea51b0cc8401fb782b6fa396316cdbf2f6d8835708ff98578b0a0e45f4a1ad26d415be6ef036fd3c661b7f6c01a6d1951e8b024695b0dda19bf4ee47307572d3dd46fa9cdd032b1b8fda8d3fa789207a298ed2e8d605119984a5ec87ebe75b2cfa4731119a4c80ee718ad8db93f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10eb5c7ba02012c49a557bca36630a351efeb997e5610960bfa2022b6ddb2d0fbae5e0b9d5a15db8f6680ee10983cd0cf581bf16eb2e94bc855020eab9830837b0883c915eb11205feac8f6951c257fa655208cd901703b83222e4ac647990b0ae8094cf40b4d095725fa978e32de939351df330b113a88e2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1ad1744df9f2ccac72bf9c38a2d2d9fc311b86910b9ed7cf66d037932be36c2627381a4f1034ba1fb4b8348f49e75db74ec87f47a54a21428068fafad241c010eae6798231ac641323c0d7f253a760dedfd00d400bc2547d1ad992b7a2e60e3737bf4e4da541cf82c56a62f5625a5a323345abc39b47d26;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f98fa1accc001f5d97a60948884dc2ebe7e993e74ed8ae844cbc6b9a65dcbbcb6941cf8073f804035042b68adb6878a22180c3ba7b793db937ccd71ecad01042de0d2732b90f865b7fe3128748b9d3f85feb0438a41d5bb695e82bb865ab51a1eb3ccd31cd757b8ec46e5ea11cefd6a9a4bb9eea5b2f1b50;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17287fa14a82d8236f3997d85c9c3e015b6b528c7499bc0ff06ab0fc4c67de380bbf9e60480442794c38bc5f33a904af06a388e554ebd5c43df66e1ab49020d4b7449d08b8e7acdcbc96535b2160c16aa590993752f76e8c65f55db9a4c4d71252ea70f149163128c7912cd3d824f4fc328ee6ae9347e4055;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cbf5560d821d9e65fd1f2bd67b7d1b4c718de3f8f14e911a9e8db96970b4e9541a1aaf1871668a8e2eb33a660cf6e64db942f2e24d3d6880b1b4191ddf49afae72c6870cc880f9a2538c2a67d964caf406b2fbd6b435c3cc5194de2b1df65a44335f3ce872ff0fc2b8fce21f346ac6466715ee4a3275e4f6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9a57174b59b410aded684db862ffdafce845eba90cbed27638368e730e1088580c8ed23b5d19d1de4e35ecab30fae3fef65d1a9a670b5773bf42ef41033f63f0d7123685853359c8f3fd762cff107b18e7d59c47c8afb64629b9b14a3920c67edc4feba2931124da2a148cd47b48d0731b4b47d4770d3acf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f895d33f96fd7c11489785225b232fcbce914f0a80ecc9fee7667260951397a6fd4ddd630325fdff0bebcd31b6974bc2467ea70da8cf7a8aa4205c80903fd969c6bdd55791fdbbab660322a0e28a68beda5eb0971aef755fd65b59f1c741217a57de4411423d59f0ee9a8656675484f074c0991f082088fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he5e217cf03e25ead5b5b13b897a4812fca8ad0cb3be019362d30be6af345ee4b8244ec31307dc94bb9fb0108ac654d38bab095c544e7d86ca5dbbd25f6df7479aa04dc94988470e3423f174e1942dee1de70a3beeefad9a4f82883f2af49cf1e067200f90906af3991f6dc20df551adea94001bfad018a95;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d7d1fbdb10b674f480478ac2c3dbdf195014f2194899fa9c90a88df88a559b7c99d74c3c35b287e57657c10588265594bb993ddcff31c14f00f230f5233a762f1a55324fbf21eb9a62c26502e2934756875c8047274809a5486b22bc4a55d2e27b068c2e4fbcf814cd3271d6ab2b297d0d5834e87be2450d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d039eff921b679cfd73bfa0126c9e588a9bec9a8c64a4da6c52464b0ed914af08fced0ff406ffae9578ae26866019855e2c38d3b74b7dcf364fe19d5eb73398d0a955cb3f277ffdbd17f19249b91d8e8fa7a99f696111fe9dd1c9da1c90bb44df259467e81542b66db1fe1b6d05f16107fca1538d38b16a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a27d102a617166227d05d148873c9a223f17bfe0f548f400f2352928f560049e73df0248aa77ae8be950f076f6b721a90cb2f570cd4d1c0feabb880115b301a5b6a99a9686c1d9ae491e731c9d62d56440e72f6ecfd62672125ba407235285ceb851c782be98933950e961d38fddf426fbb39e8c12f0b5e1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1241977c52976d1dac1d05159e0a73568f8f0342093122ac1cf268f1dfc97c6398a0c2ddca09defee1134477d3914463a66f32fc4ddc1fbcc2c767c424870974f542cfabdb9c01a45449789ade57bf7f434f65065bf86b6eb6b3e4b4c5e79c159f5a1366c2d1b046ed2320381b38b08f0c024214b86ac37cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1af6620642bc6479ff82a8530752ee946cb9591820707c72939189664155343920076bd87aa38ecbdc82849475dcb4d4ce9aa608816a53f2af776d6edd697eebd8ba46646b50fdfcbeba48b9ff56c264d6e8cf59453f8c9dda89706bf00bd8a6adccd593641ce3b012eea93a35e9f95f846f8c28302d6424d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h31aaf131e6f017dbf9b1990eacad39907dfeb9f4f91c5827d242efed3c44535650a40ce6a099df29a988a47d6f5d017b5556f0395f6464bd2201c1cdb38f714472c18e1740d150fa2c7c33e6a3448935c4c95061f947f8c66735a790d2e44a24b5a2a4c81e6bf352b7e408c7a3e498fd2a0dacf932fd5680;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3917066425da5ace1cf51cb442880d0c8dfa449bc77cd838699bd5b2dfe4091f5b9c126e0e3b6bda6254be72b16907e521103173f013a0913cc77befe6fac8bb460794139b583c99c0576b619601e766e8a50b6fc4c01e37afe9ee90b41ae51dc1a3172ee7be528841a302594f4402ad5ada631af321b779;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b058a0e86afa1bc5a8fb7335fdc4bfc0702653dd804edad1dcd1f4fd099cbe7473d00b3cded00553c13af4fb2219d9522286733e89b368c914b96a8d39a12df8d9eccfa78b8bd879742e07178282f42845ff3cd1f2a177ce3eca696b72ec5f13a4153efa5bed1ddf6cd610645bd8010749e2d720d6288b1a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1448aef022505b1a801bc9c7dec89f87ce1d7342894f24a286a8db159cae5ff9bbebd4270589b02569cd1626676151b5dd4bb4d1a079b0934b0bec75041cbe5cc0f39ae7de7b04cca63d6ee41b94e131a795c10f15b4d4749640a1f4fd4dff07d27c2eaf27f2675c9f18a9016729f286ef2f115d328bf07d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha39eed007cbb104da7ef0a95d7b58fc8a5a1b3074c42128ce30e46b92a172a7dfd28c403f9bbcf3beea3ecd443394e1e00de65b81af3f511b6a8c51609136b1ed0fe0906094dfdd26da533ca4232c36a1a0526aee1ae112039354d3c9cef7fbaaa0c5c83a45154076a7327478efe6cb6a77d4e8cffa6c73b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha1d7c37e537fa40ac2482a913907623e172d358a8043e40d8ff14ff4955d1df4983c74967674e236ea95127a08af5215978df3889e2943359a1ea80abfc3179dbc2cf737860b7781d6af58c50e300330ba0a5b2589cd5373e7a1aa0b4742a9f87bccd32f71952169a728a4eab0334b5cf54212cafd8c49d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16313b01a8d5a55da13d75f1b9102be53e399680c0003aea561af24cde090a7cbd54884bd39a113646ca928867d7d16c4f61cef89bdbc62061317e7a0de7bf785d768db6d426fdae8d627b913a3b69a41adddb13772f1a252b9acfdaa635c7149ca2d28f407e1472e4c2ea0ed40332a3793fc78c78c52ec74;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h36400c72fbf4f061248bc7ba3c9c38e3ffeceba3aa0e6007737c278c2867e1710a6b76af8a1acd11e2b9c94dbcda3a53cb9db594e3914901d4a33a64519d2d1b5da9bba4fdc843b5eddebf35abf32ca350754cf382d2f498f02329b65bf89a1f42b43c01eef3f9f2c45d22386d6e9b5118365af2de5ff5a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3426b42577352cfd6f944e62876a446231e3e0589d1ed5d316ff0697e0068fb7a575e25f8ec86a269d0a595dc391272c9b4164377e291a08ec17d6f5b0e1875d85b4f297c72f13294f5b7fb8e1fc0ada4b1721e6d55596d26ef2d9f3fc14c32f65791d689ad1a60e93f9eb0cf793d383334d50405c526d75;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a36ed7e808a0c7ab3caca2e51150b7788c24c94d3c10185619f49c3630d6d81fe6cdbfc1bc4253f48e0848ed198980069d0af077a6c2256745ae61ed340738190609bbbee3da6ced541195b3324457f42bf9bfcbc48ed862d7d6620bde17366c657b01f53394be2576fb3c7f735191a68412c03a03567876;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h891ecbc53864e5ae24b8560700680caeab42cb36bb1477c21989f65b51ac219000fa3473db72e73f667eba52277778b3485aaf02461de1f6363bc165c5fba960ac60df1b3c27759961c741a735be57e4b53b908f2b8a5f4ae38c43e2231968d2571f47d5fb92c4a7e62a3d8ba1880fb9a71f4e71eb910762;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1725c5e9049f5ee4a44e78b6dc3d7f2f9fa9db6c982803480b3febb4c88bb652366560e2f2cbe1262a39624debaa5dfcdb504de394e8b56c31331e29159e894a570fa83197acdc68e0501ee1d0b21459fe72321477f25b7c98556d8b93d14a843202a45d3117430c2d984ef001744ee40fd3ec93d2ea562de;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he08b4c5c367a9e376603b5c3de8883f07e55da731833f79eca1bd146e97b245627dcfcaa9976defda041c505aff96a3431802b84dc46ae2abbbd93a4b9ebec08f6ee07662f464fb209d76d4868f23267932ffdd6ca58b69817efb9130affd30761460e09f4fba269a6a5d29a278e49848186fb66936eed18;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed26b4f7103f3630df03919bf3233d8366e807a707100f910becada03b610622336be962ded40b7c95f6751899143e93adf81e116fd0a56ad5f4a3537b8157f79a94e1feea667f09962389f6d070b6ac953c3e57c8b378f0483d7cf30cf1caf8928e6edc60765332559b2d6069a47e1c7a1f056106348f53;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157268d2760a15e8e72c8269dc1fca1e67ab79aac083df3e27b28fc1087793956adcb36954744eef41db02ed1518e43d2b508b11b7ead6027b3f144bf3d09780398ef9d1d384619e7f4aec7cad366e982de7f003f0c900eeee5f232826545d80bad87adf15af6cf65aa737d6c32d3e272fd48a41f4a535aa4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18477d974600e1d90b090ba921445b684e819a56e17568aee801de783722972096bb36ed94f20f2d1e95447052e76fac3899eeeef926a2409d89ec47ec3534d93aec337ebee80bcaf2e33999bf1ac5dad691b52587c6bfa4fc3aa055fc22df5185abbafb32cec59725d467524959267e7b4caddad3fbad497;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb9ee5c090c6622fad0160422fd6b07664f6cfcb956eee9f885b87d61a225c85be2ceb232bdfbe36d097f82e33dbfd1c7891e090d34e45371d698f3a24c84428a27ffd06f905eb402ee388bcda1684427da019cae97b018384d91f78d6f17a67f62e66ea86431dfd23ac4080c1ece6da7ac975b44bfd6801b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc18a7f07422a1253bc7bb3d00d9509d2e65fd3d072bf16a7dc1c9b1e48a94b094b01f99330eec564104168146b12a08760b061023b70b3e4c35d5f8299e515a6e4a8ad275f526ec2e8e81d040621344974371a03d3587dcfb96116a81722784a99a6c08acc288b134e25df4c729e8882f3cf613b955c41c6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1242b1d932a45be73a883edf3384eb9536a022ba7f02995336e871d35dd7295cc35e35f62dedb3ef78ecf35593cdeb7d9a97bdb2632ceb3bb8bfd97529429958e2a9bcdcc9f56b876f77efefe0e74e144b6692dd33f6727c8fd3cef02dd91f8712b332a883257aa8825aec736d00c724357061b1614f3197a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he3f31a55b9f3b7e9513035451b7eba57405f89ce1ac00082833769ce2985a71cc85da980c39fc05bc62fca1cfffd679c562e0e9e103b635d1f9584f69aee463ad8a663000d6e2ed40eeac9db44aacbf711e15e7b7a16d9ba6419397b64ef6fda4e8535f8d16a4dc4bfdc6c969f48f51fd577ba31b4b7435e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4e34397dadfe16ca2df4ebedf9368b94e2a93b399685c9788011ee8fb777b27e7cdbdce7ae2694fd6bc8eb0fae028907d8b3204b34fcba8b053c34d96aaef565b76e8ac8b4e132ea46dcee7761aefa8f4840646109bf07205c7d50fd1669b1155ccaf6ee39191d928c3c090d9f9fb2ba4c2372d38a37149;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3dfa3bb316b8568a7f4148143bfedb44b6b0bb9f426b15e0c4482596aae60094bfc717eedd15c66b5f3e0d1d750280ee4db21a6dc8d43136b8be29ad3bb2f40c6f81a62a52b3f4b909e70e8394bd7fb4e9f0ee103b6e86dbc6ae705ac9ba318bc291435cd3cbeb111a2c71b759513ba86237788a18b532b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef0f8efd3f96ccf54c6c410eed2108b27fa213ff6f2574a6f600e9b0c8f65931a276329990cc415532aba3bd46b278f64c871bacdc3749c292ee1813869957afa7ec9f3e6170435fd9a52fcb82457ddf744479eab29bf25a5558ce9605bf57e508df79cd18223b6cc744acc9eadcdee28960c620759ac195;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb88aacb7ef44c698cb816d5bccb0e0d8061a4360aff95133ea89cca9a4b0a19201873d0a8e2b50dc31882c41937a92edde6b21026506417bb68b2739d9443df945042f2db8333eef04fea9dc5abb514b15c6f4a19c6c6c806a96f310831482679dd8a884e549b8ed168b46ff918b9dfcc1d39c50a774dd7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc0d0e465ec41fea9e94d4f0191835aeef323ec9d7c9f2021c4a965fddde9404a7cd23b30e7d4d3527f79f620023d7e3032800a5ce97399921cfdbfc9e6f706e6fdf24aedd2bdd4f715de1ba59c886dc2dd892464a48bdd74a0496f6e6d492b77ebaef4f65859e2a118d5a6d118f0301ba91227c8d7a69901;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e84bbe7cb3e973dda019ce82411533fee772a36c02705921a0dbc26f319f70ce9dc78bd83a0e916efdd1f3f203c27055409fc212ddbbd0f4d087f810a04f9c6f70824b79ab5050cd5cb3c6c6bcf303efc73de18f466ee0d0ddcf96c46c9b0b7576f2970933d506cc776c0eb3a62102652f2854422ad8b75b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h191dec7087144a6cfbb3ec99a112eefbda2430d98965c59c0fce8a7797e5a56eee0ab0b3aacf0a76ff3bb2108f40c4fdb6a33b5f7fec9d99457ad19aaac925a228d8579632216add00059e79cf60cd847baf6f8c84d82dd8fa97e260f7c6b43b797136ded630dd69c90aa5a275c93e05844a738eb44632030;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ec919dd648dcd9c16b56f4447da856f74a2a451c1f5fcc5dee2414862c7d15dbb904fb0b36571ff67f0d6381706b255b155a1e9802e8b6ddd9bbac269c2199918d5a538220d930ad4920fad32f03d7ed5dd9bb9a6148657de7cfb80b38f44cefbeb620d3b80e651f4d057954a9b459b2ddaeecd1370c4cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61f137e3342a7f4ed0c9aa826e6df086e147798be88216d545c1583b8ac3a7ac5ab5eae227a096afd421683ed265b58ddf2c504452a36b63b0b9dcaa64b5eea16ec9de2738adac7be0d988bf45914cdbc20b927b7382eaab1b2cd5ea16ffbacba937a499326a089c4ce5c17d217eee9c3426ffacc9b57c35;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3ed3706118dcb88b120ced83780ed7414e1574d8a7ba8a9c7a9e1c8bd232de143938134a200ea4edfc8816f12b8572fe9fc3d9e22f06c12f709ec1f25bdcbfed8e58955206335f891e0515e87816b0356f4c2de5a513cde03a28d4dadcf52bb52bac56d6373c30b8a874d9643baa06848cf6ff0b268a391c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b84c9058044a3a0cb3d5fb16bc4475afd02eee464c5c7a9536ef208725b3cfe02087c42616bf84a39e7893e1d2abc2fb35ee6c66797f4057389992b19ae090df27f0a525bb523bbe89c75b3efbf907e7d452d78f5be90df81e84c0fd109847eaf29d885dfaa4f7ae52c1f9bc767f7e1b155bc43b5db6f5c7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1618a8fe910fc57dfdedfeb273e5c2c5c6c100294ccc3e6ffebae42a9ca74385eb91866e8fd48a7970da46304d666ce033258e491c1bfd9657b8128c0a3b3dd143a9dd43ee980c77609fe7ffda02e8da56190c4bba1086c3114a75143b860b0999179b23a9a62f13f945e56c191c61ea2cbec95ea6ba4743a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd8ce45fbd2262bb6ca83613a978155846fa6645169cc21395229385d8b98f0adeb7d23a2b62cc5f27ce7ce4b3a38c77d5624dbf26368d701f49a04b603f5a7fd748a78ebdc1bd0390e7ccca10dacf978debe08253060aa3d5eedb5c69680912d7876bdfa7a65a08cd00bb64071d19888cecf402bb60f7199;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h554aa82258d659be015f89ceabe3d7d7d66b60e7a6d20258e28621c73cb4e0b16e3982576f5baf6b9816b8ded9e5b8522eba4db3033a14eaf64067f1e364aa4289c9d30d2b68c82988338d78d0111285cada17fc2527d85312f902a82e49a07687fe15021a1a03e2884616bd56ebbff8440f5881a709ca0f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ff945c1aec8b4bd869d1b1eaf73f555e90c705627f94a30cc63bc9b9a94ba6a195355984a9e255d569c3d65ee0cc16b2ae0d2b24484cd2e5df394075d2c0531288da877d03e5353ae19e0d7a591bddac748533677cabcee902b5a1d7a4fffd565a967c02b724911f89ebd038918b9660992f2276bd3074f8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11d65e6a80fb1f83edcfdc7aa4bf1efb91de045e405a0ab8cb912473763c42de7bc2e8aae5cb93587a4b0bea31b5bca6fce28eeab7279b745051c6c23da1f49e63a69d5f28e8dcde1d3c301ccde2842dde01a59cafca3db37f32b020999f0bd388d30de50f5cde0b8c4d97d6bf32706d9c99c8467be979467;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ced94a2830eea287bdc879ec3927efd2b880b0bc692fda134630d49066f1b8677ea66e9920a3abe0258db40e0a2235cfcce5cd458e4fb92057c00f8d7ab54f6258477c0291c74364911bce1b9c92134c263b743e253042fe2b61b01fa8df1f836143dc7310d80990e8609ec37416671129ae120e2ca4dcf7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116b7dca4280ec43d65da09affaf958cde12979669d245dc14713d3ad9e3d37c38cc93429d843677ed334249d15ac152e7675c6e33c87c364b4577c5181010d10b693794d630fca45dc42ef76fa3670bf7f681c3f809d578340251b01c0292d0a4b377345ca7875ece057a46a0e7c7604acf37830ceb569f7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h182e02526050aaf9565d1407cfae72de586373353c8b9c51f30201a645b0c179b44ba55d9533b4cd854b9e91ebe795156372f8720de122ca6dd655b695066d930774e411ec5c1a89c655b73bdb3cf59b884ba0db3f8ccfe40b8679c77efd1557e39de6d84fc08abeea2105707a2b41ca3e59ae752e4178dfe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a417e2bdd8657ff03f538a7e321c87b67572ada286302f76f1617ef3583f3711a88c2aa22187191d451b76f588bc79639010b5e86f908c7fb8c07b189079127d4b9206d1b63ca66965a389748deda904dfa97717f457f70534a07531fcfa991d8be9640144347d84bb34e9397b23d5eb7d47309dfb96305;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1666eef57cda25211c31247de8a36196586254d1eb6f48ab75d8be5dc6f313d137fa43a5237d0317ca37bd849bc5735fbd9103abcc6deb64075c347df3f50970e037e64bbaa2cab2f11a375d00bd167fb7b5a257a85768ebc676ae3b59a957f934f514af52db6e1e58a16f37d97214d2c35eb46ab5d83cc8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1539faeb3ec391b12006d5cb409ab2b318dd2f8e42a1fa36def8ed5c290be3003ae8b1eb2cd70d750d3d48747b7629b2de02b3c53878d7d2b9a1408ba2c1fd6f798f4cdff9de9836a0fb366adfcc5f83a1a6b4e5382a15b09a76dd0a3d650a7e142418398e17961aaae43bef6681efca01a4e73034f7167e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19929a98038a6718405f15f5f47c1737290eb71a47a1431d3c1654426e6721fa1f9c59561618153ed330d7caa356a62e973b92569b2a180b2036b376c022cf04f3c3a007e3203f6fc4db5b0055ea1dd7e87e2bde389ca4f94d95f25316bc093086338f4e26d9a2594e05158495f91f5015640199129b97909;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h108d378b3ae541002eb2b9612fde16d340f4e251511b43db03f169e5d2928834383a248fbd7c51be4e4c65cd8715cad115e542c1f79b813257f6fe75c09c0c9f08b8ce3382a3257fc448873b3b950e159f9bb6b167041cc012aa3724db0f1671630e224fe607c6433f919991403f0be5fa2337c2018b23eef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h150bb79ae918fa9b141b3943cb8e431cbbfe2dea8e0ad72ca1a22d3da37dcbab49ea3b09b3ac722787e1a163501b2ecaac75e86364d746415d0a68dd67435838fb4b34df5dab612053c221bef53fa9189c6be3f4323a09ab8f8e0dd732945c91ad3301141c98162ee630eada04ad03679a0a0c8cd5c5c400d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc16f0335ec21e8a80183c44bc6e21eb21895cd8703aabf10bf762b75eb417b33b8073cc5dcd67aca9c60ebebbf0087d306e07d699b45d7db6b8a4ea2b9f6019e2cb8b77cb5d3be57bd304d7f6443903083f14e0e25772f406858041882b3eb3c5b104904bbaacda2dfc4c0b5f21ee92ce87265f91fdbfd71;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heec7370d0b1fd5bd9e1fa434349a809a45d7051b53cbddee50e1cd420664bf04a9d9f10d6e452c5e346ae1b44d0f9040a858902ef2b713aca450d7b43ad8258b66d501064d99ab662d363c3d8b7b1b244c524254806ab651d83296417cd8d4945192817e78821075610ccfc428397559a94323fe80a07995;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b0a87b2f82e770a008ea61e3766db4e3c002ccf53bcbd6be1cfa0e31d6ea7d6b2df1eb5c29d38a5f24e545e115e49264bc9ea248c6a4718970313902454ceb08dade9aab2f4f1d9f83607f8eb289ec0cf46d5010f1830b2ef2fd5023ae7c3655fe655a2aeb9b9071eb09a4f5dc9aad3a3da825f0a0f6de5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h100cf95fc409f81c10f6dc982c17a83680083a85eafc7821c8e9beda7863c84e3befe65ce2589d0e37c76261a774acf6fb5b9b7b0ae258eb9f0fa1fc1675dc91cd6cf3800923a91755f289565fcf408e6193db4b77e1fefdd7d0f5f4ce46886fe8dde193a3e2d2f8b0feec13bcf8281f599ebcca7591bbed3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde0135f987ab60995e13c65d4441d6cd20aee52200f0a46d4059d7c492eac177b63577077fd8e1a9ba490fc6dbb34ec1962f30d099c235107f19f4ba97ee6365ea0d465e9271c93f5825cfcf2a70753620470e11f9d38db8dae659ad47f14a0087c3ede9b7f122dc8a3227f2a3fa6c0092c98fe9b1a5abd2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1447f36d3ba4534d7ee14d08f2b1dabbf56099aaa3b59212db1a1cd456647bb4131f1eb2100ff40902045468a18ebd47754cc1bd7a3cecac272fcf9f5da4157e1e62bcdbb99212fae0bf0cc50f5e39047d1209418c7835ca68e63309d5d7b98c0c7f9cdd880874b07095d790260f26d2ff30699910f997ef6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h51c30b151a3a15af9f699fc15826666f0989dd3e0fa23eba4cde31705b95699b9c9b9a4f57873ddfa617269506a690d102d7640632af13022a9290d346e793af6a93551e8a4811148ea4da7e4b743d295f22a4edde96c71d44d778a69dcaa8d51c449fd2b32cb6f54ef844568c51e5765a2cce04b1ffce66;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7d420e22fde4c307470fe0aaac68f6ae7e6f2cfbc25d52d12fb059e5129f9c6b51a19ffaa2c4f72d4be83b1f64d1a12c73f8ef2794eb77ac937768dbccfb322a2c9d6d66be6bf7cd44557d6c8a0a2a9d3efaf189b3b4eb25e880a12888840e48e5f7a73cdf1b8180b091286b2fab91b54d8d48d7c562cbd3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b8666dd93050e9790f950a3c0c63917818eb84970a7eb4959020621e49e7b416ab56f52aae0922d03d474a1d89a4d2fa20777fec67999b78748ff5c73fd810449d4ce214f0344ee65e41a19c1323b222b77ad8ad3bc92731b857245337d6432873ef155ce189db5c94c7376b03e5a99037cd90e260190a5d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h296bf856153f499c7e38788fcbd40c4b8d03fdee0fe1e99596af1a95a6bf8062e1151188d6d242b7f85eeaa35258b59576123b473dfc3af0a5a63dcb4fa7ea43171cf236d1d772ca375f182949a9cc1ea73721e60e997e72ec1ab217ea87c519a6cd4688161d93c75356096833658f7a4899afc849c6b57d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa928ceb91a0ba92233e3c3a55aebf59ddbdc394809a7b20a60a568514d89594069f475789e3f0d41f311baca7d849afd9287803935340e6019f2542fdfe6523ef699f6b0eadc632412b30887a76505fa61c7ecb4b1a5fc57c0d33481b28b12ba13f529d6ebe344a57d2f844d5b72ca6adfd673b3e6df77f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h323924ad8dfaf10e6715f2d3f219479d0229ccaa65c7160a962e87cf0a78cf886d19712029e4149f25fc8a69dca5e3697322c607de4c4d6367f7b7abcff9e5c856dbd46306a45e7c0fc952ab0e6461b973d8c050de57d64dc6c9fada9bef50bba0daa2139048416da77192720e9c6817a05107bd5ede3ffa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cd39edca0a9ff2ed5755019d0da520b41d3f6d34f04dcb035c7b8f9cf83aaadb743dd09cc63728aeb0872218f9e952c54c810d1666dbf24c0c15bf05742ea24ebbee10378656e309053d2de2c03069e549e163612cdf1b712966b3ba2375f63c52bd50a0caaad9357c9b136813713b81527d0e73901ba3f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f3e4b7f7dc780a02c0dc25d4ec9aee4e6aab35d1eadeda0ddf06b94bd569a6313f69f176db3d986fd27d922a61842114b221ceab78a751d1f095348c35a5722485921c133b28c1f57b1db88c1a64952bf9807ee48b8c8715dfe780f377c187d96e081b90700725b7a13509d16a3d25bcd1ef229e3fd57294;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d10d0c9773cc889460e7f73496a2625999560c4c71c9868c0f4893cfa83050ff937ffa3782505e16c5aa0a0411526aa41d6533ea29bc5c46519ba9f16063e994998dcf48febb1376c3d05be714441f31038acb41d15f999e5b15a086dea7906a33fa4f07a0b407614174bbbba37061cc66eab29b17566c5e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18fa43fd35c0183f70cb52041fd79e0cb3d87511af3b097d9ff79047c60ee7ada47d69dd75b013b4e11a63042e204708b7a9b9393ed375bd8fda9213a60af953a233d8ae6b34c94e053efb6ff62b4342ea53ac32ad20c3cdd90fd7dd7020c34669544cd76e026a02fd3d51e733545528a8809d1f4523d6396;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h91710ffa80b871763b55f811fda24313026845b278ca23971d808c6bb8425b6092f23a37383609ee20850c76c8dbca1c009ee4fc3e6128742b2cd2ae7fd09de2fd8738baf8a7f5e1221d2213bf044aaff17451c62af7f0106cd4818d7842b933d9029bf21ce50793ba245845963b1f014c3edd78034637a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c66e07702d633bc9954f8822767a9913b4d45d163ac550569a3a21b6bea2bd6ad321d8bcb79d77614021cbbadedfa60431d3477bb942dd8a16f5bbab2f436bc1069d7869f968459a60a4287d692e85504bbf79214547eb9b9dba87ec2089b4e5b39a6a41ab5ccd450ea7d0409b1397439fba6037ed6cc141;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb34cf25afbb00d5c5ae7093bcca03c1f0f691b5adbe1b91d8b5f7caeab8fb332d857a58911d69e797514f43a9b1e75f3e51dd6c17b56b728ddf502aa2448a6162ba585389000432cf944afcda12da60d0ea4f2bd1dd592a6a56a26566445f5ecd2d7e24c616af103441aaa08e41fbde58809990d0cc5ac7d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d482fbdd2c3e833824175ce5c76598040168fd0afdbcf48b937ffb6005821a41b7eca5059a4b1fa0e3b0914955b6ac510701c04f5a0ff3d5a14dc3f93796364a9df5ccb351ad217bda82c5247b5c2dc70cca36a5efe365d4876954229fec83c5297f142a0b884feb0aad3f993e8b5fdc741579558464e013;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2f374fd09a452170a0d58f6f3e60bd144ae924341cd825274b702d03aa84581dc43d27f22f0a8daa8a0bd26235957f114ccb7d23ccbe5c013b91d54c021a360d0dbc330120fe6a2275dfeecf380ef840f414053dfe23e57415248dd56f9043b7f72a446b6b91d3af6c37b10b577f64039ef978533f1a4da;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h114d13f0174ce5438630aded6d98a4a31fd17d9a7e39c005d0d173af7bde774ee99a154fc258015e70e23eb3a2a1165c788c7a158ab9b41c760792a9ead417eb9923477670d7b27af6da8afb8efcbe8ed629e16db026fa51caff202e148d037d42721ff4acfe810560db9a5ee84c86c93902634976ad04787;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8bbc13533c0be10328ef6027ce3ddc67acdd75a93f6a0a20eb65d918e8224aebc6e525c6f85f945937f3c94575f74fb2f48d634e22380d8112152cefbcacf8b57fa3df66f8bca9cd47c7ebdfa0e9870751b4094eb8307adf096c157dd0813a0ae71c5c19184447bea5b02ced7fedfb64ec629cf663570a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9717569e8faec035ca0673a6de119c437f4c8b119e6e81df500d2c09d3eec88f2109562b49420c52d7693bf31b4b50889528609d633931128e1893cd7b1d995e8146386cebafa14c17679e4171f8742dc8edb5454c840bc02a07a63505c6a6ec3bb1b3b904b3fd0ab2fb7fa5db48de9d5f821f45bf70a87c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h136a22381744b31ddff7041e1f03a03294fe328317240dbfae8f54b63b7a5f2f174af37a607e75b9b50f799276db9429ba0f59a72687f2a4074ab956f268c5be1513dfb120685cfeb0817cec339a3754f0e34375fc742264f7731a2559708e6270c75081d81b3ce7f116dc78f6efafe8bf1a9e24f0773dc7e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18015ecaa2746900ff3ba99ffbf79a060e91d992c09c6b538d3cda4bacbe41fc7ca0034903acd6e3a22ce9ab07ceb2fd7ba29401492442ab2ce78d4724af1721356a7a344f3c0be0707d1890b22ecf9cd759ce0664eaa35719ccc185b2d568b07f6dd5e90e0641ef7510fe36c9428c52c2de2d113f8e77d89;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a1a4a53cdd3e83ec722aea33f70fe4727d193af42a9353c32f9febaa64c2a166746ae0c9ea01e7e57a06a2186a7f5be3f793171c5c973a9fa4592d341dae5425152389d239d7d1d7f132d34ac2b721038ceb2cb19537ddd722d74d548a30232550f6ec22e8d5bfc5d17226d98f9eee4687cebf98679ac0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1092c80a2560803c80a341f56992d0b5fb5a75208e5f7c05a897c3db3c6961c2b95b2f524f70e789ffeb2386eb36f933ec2f50f22999345655038981a135f0ab5e9db9f1cbeaf5f80cd1768bbceee280e2dcea2c1fb9b54d223208d13be7cbca466a60139ecd90419328c1824d483829227d96287bf5c5d6f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19ae3eaf6f907cc2ca06f693aa2461e740c3b1e80812f628853b31fd8c59bcbddc95d344c99ff4219f3e0fd2f14e028b192eda2e50e1eb959b70361df9696ad475366c7aba092daee9cb2dc428c12cbea08b099c2edbf00627f1f289a7265432cec7a39e0fa24d4e80555b120a5163ee0d6c39dc9ac863fbd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13b42aecff3dde8a30a9027953ba5645ba80e63f8a021708732de39769f4e22dad11aa4906e5c50b3d8813de571fcfe2dfc1acb3008e1cd858fb7dc19ec09b1b847fb1b966771f8ba15cf2dc292c0269d64210eeb9b60d424f80aea170da2398d1726286091cf4968fc2efab21204d0d223fb5e873edc4ca7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ec773d906352dd8850cc8cc649af6425d7eddac2fb7f704711d2de2d811a8aea008bd5ba4c98aaeb946467661fd68001140b738d57a0b5718e9c63f0417aecdc1d09417b602916d99dcf8d879fbe78b58362a704bb245e0d1c062020827017e91324becfc3cecc661d5c2d090e047e48999a149a2d068c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f76afc47bb5ce0611ff170818ca1841b51b0b2e6dd2b0bdcee11c63a4e97f7b4c768237382f35c3c18a6199ee2051ade2df48012e1b2a475f4695b5486510920e7da41970cf0a3c4973f8d810df14b7a7d148fbb5732997b587a4f7d6626fd57af454fd9d38b9dc45f9ec42a0119687d43cf80217537a23c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h861b708cc74ed8487547476f83d899f0b902a8e6259a7e8157b83ade6491f934b8178ad83ff9a3c48d4a56cd27cc2fbedf04b9c7b92a2cd3b06715a12d5f247ac65cd5bdfd01551c4627f2ca9db924ff84cecaa3a1fd3c173650df9dc6d71bf8182c24b64d4013372e2b314aa363678d93ecf19ca320e9c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1072fbd8f9db7968399ed6f52a34e22e2fd0d9fe31986a969823b2385c45fcb349cddb765f5839fb44684350042dec8e1458efad0cd1bd2427434d4bae33557cff99b2ac635598a800efb53892ba2f5210a7213497d6c16f051c8b05364588d5157236951dfc94eac1f9d89779c59661ca15f22649bc00806;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6eb7a220e62c3962b1ffe039d14a14122cde40ac44c7f92936d10ee17c7cd930c5a88d42f656265e0e4c84d0e5bb2d4beb035edafac3f753d45eb59b6d1945092639b9a976c25ef5729d403dcfbdc0c9520dbb6aec0d97dbde51ffd5ac19f002cd64c4b365b3dea5aacc065ae6ec0bf02cd7977abe89095;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hea7fddf159e73fc56440288586d0054035044ed7374a1d9fb6c70cf56d8911e166c45a667d3c21b2750033da5aea01d1aad7f33e15967e8f1020bcb32a0f76b3d9c46410ab706db357060fa0f78a378ebcbc86a020c29c3c6f1f893715c247da4d4c7b72b77891cf9e0c9dd7bb75e3c7918e1d662b866f69;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd711884c121939cbd98089dd349e50bc3ff75191c67a9d5d1696ddc1dbcc5aea77ac65df0018558053139a2ada033fbb6bd61b286b5a3969ce5b61420d26d106ee44a37145736cd1505fc6ef11c26f4487d0329f80c56d184d1419d153f6b878add09e5c19169f1c45c11b0179cb9bc24211c5e3e95a7af2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1708caa271e284f63bc221e9382cc5b0abb90c269bab2b3c06525259e7ee7c9a52fddeeebd15c5a5256e50bc1c4b139facf5674ad697006e2d3e19a5bc8d44115ad16204f920ee81b208aabf0a2b2abff8e8a7e610b5282f767567833e31e31f49c1a9b2f5b3fa9b02f67b86c387b5e3c27710195d927d616;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196c0379f88f54cba3e4b333bab114183c2cb7b80f604308a648eddf0e53f8aa826343c0f450c65a74d0311efeb0796347720d3c9906563321579ce4433d2dc5a6008ea1bbd26b5f8a41f5189576f3000a1f63fdba0af0d0076845aa60f71a08b47d7f6966dd808e9f8fed311d239c8305a249e67d64659b2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13cebfab600c8a115bcedf28d5ddcec3a3211ef399fb08fd45e64372ba5cae00ef326d52aa1fa6282bb7ebdea018dc7b659d99f21701317ac43ab82749e0678b8745f39e24b2be936e3313243deedc49440c0233dcea1e1651baad28882507c61e37d500803112238f47a6e6f7cc297b651e314f802643c2e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6d576fcee028ef661730381d19970c620c1a59976e74a168328d717f55c92562aa367512f41dc8e35760d03f4d6a08194696d2529c41411c9652ac12dfd7e89f9a61cab13d714b722ebf7910deb904ddde4f9e88bafd61f26a690055a73d91ac303a06c8b35ff8c3b870ebdd78d52838cb6ed34287b09d9e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2fc7662e66eda7f7a1e6f8a7834ab45c70bba8b21d0792351d0ead4847622ba3086ec660acf587356ee00fd5029c24865f37dbc30f7d30e36843552277bf99c1f312892e53195fd00124d8c7f6c508b46d89c6a350d4a4c9fa55dab2c4e2bb4c8db6e45c4772ec8743496c45c36e8c700a42f6202b35ebeb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b8050b97fd89a901a9a4fb628176566d7bab12f537a1a789c2220974a2d9b3e537079406cf65876bf9c6d7a3759d3205208e58405b5359b765fac1d366f650e4b483b4f95390ad37eca21e55e324dc71e79319692e99de3bcca11c265cbaa75109d53f24d1140dd0b1cbe729cbc1259d1ec311034fcaf21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6cb6ddff0cd5d4f5b26bcd33d6dddc255e5da5791cbf0c10e8d0007b21fe9e4b2753d0ff9f44cbf78924a114bb282718892adfecc53a6a1a296e76f718005d822bae9ea93ca8118350c59e22829a35173f81d2564c2b2c03e5520b0546ac29291a1625c04fd4bc8780ac0df77eb06385ac962ca3ad7c4ab9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h190019b6ea05eab75dfc77b493d15988d52728d62efb210db0e4c9caf3d0ed48aebe4f3e3e77142b968f585b013b7b74cabbdf4764b2a96736bcbd0f1fd6ea6f7a8a28dacee099073a5573449b8f2fb57a3363bcbecd807a3bad520930f53430127185086124d9aecdc4c18a660814fcc9a96762fcd0f6def;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c88a0c8eab648ad6439af07dea8bd643077d8851ebbb293dd4f29dc84685c8fd580f8478c4eb43d18bd595980df28c204cdce13a49a3b98a9bd7c0c408701e249197dbbc82c9908d34879f0da08b4bf8771a97ba600c2d1331b9788beeee97bb5848b18260eec4ea696594c76b0b4a0d0b92da7df613e41;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f6902b622d715566220f9b325cd6890d1bcd614b80a795eb01f04d092b08eb13cfbd1eb052e48025d60b8d6c6f1a5054e2a936fe051882403d07e950c975017105f74ba7fb7b7475ca004d3078ba67c43aacca17c1079e50d33486d10bb5e3ffee4171c19f19accfd447e671947dd3301ff8ed3e7814918;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he9ce915a54fc8728ffc0b55f66128ac3b23ca4b8eae95ac76de8309a6443acf108f332ef931491274d5647c2a95406c35cb87ea7854d0a1e11bc3cd8b7d105d3223f0c8279ded3a957bdfac2df88f68ed3fc86a8aed96f1fc9b7a547c7605803317d6e75c6ffea61e0c697822e85dee4d299deabd7fbadc8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha8bc8ed32a39e777ebba7d81a3c8dfcb7ab7faf2a0280c643930a2bf76bcf3bc044df4db836989ec0618206ea8690b9168575540b6305203e5745e3ecde238c5c8b7f4cebf63d37c8fa0fa80aa44b8c0a3bd4deb2d50bcf8e2f8d3031102eadbac8c36abbaa51df864683511012b37b612f88001e17913c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1374af595d874ab081536c74d147e46499d2e79966c3ce9ca787a15ca1361dca6a27b475cc148c6212d06839161c7965b1a7daefe5217a06d2d96961321c16aef2577b5019a5269ae7eb96337725c45bb9aba7e4b880f2881bad6c5956d71c40be33f1b021a7d2ee825b47a8b48912ce893a216851dde746e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e3751f8330ce76a148f7001ac184c092aa7df0ad1543b508b785decdd367edf086f0a89bf874074fb0978f730be0a98995b8700e09e45a603d9e89c827a4ab885ca28138b10749a60886efe36ebd0f1cb7be342ae84da67dc06ecdf8bf1ce2e2965d036c65c35e80a78dd94e05ad805d1404185f850f28f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f9f7bbbc37d05322f1c800e525c2306c8372a769a5a435f1ae43d825204035dca2a0f11bbb79abbe22f236c0d309046e2f8da324e30f4eba19b248bced63771ec40c10b6dc854cbff7088af72f78b96fb524b210d97c398565c0067c794db42da2a194fb29b702a474c0a73e584a7b8bd1aa5f08b14094;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a9a456b04f85fe0a643584410471a6cd039e48a708c65dbb03d084a242249ace752e53e213ead1c6c4ff5209497cf5ddfa9e1e76c3734efeddb75b3ec1e7d4d181b6a50ab7b1f0c9196147412d7133ced237b31bdafda9049687bc68e82595b7515f8178dc98d007a81bb535f97be04de8086bd61c2686d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ba4113eaf9d45d8df3a8069de211879d41ed16a8eacc97d9b965c75a59509fd23a15d327336e75392393f2b422117101611ba1beaa5f7360e7cc31e621ab182f0709dabfb251fecbc95cc538c5b6af0a9ab541b31ed092f387feb1d3736c7c28f4d9bc94d220b0afa6e654459536f81c6ec3d8a22166cbf7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h144b9dcfe0cb86df337fd4dc10ebb4ee812530ab1e81d0984a0a6ebe6ca629c05da5b3a669d0a693d3d27fa4fbd84e7fc91bc820eb54ea8a591d6d5e59efe3b48d455006bf0168192d925fbe0bfeb718b265965c4f59b69ca829cb1cdefb06f94c458ada28ddd88260923c188772dbe130cdf6f687aba898d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f2d8a92cc64c465f650c92bcba7ba18c71ad682a5466a4e149dd9d83c4a809bf13f8202117beebc969aeb6f25d037c35ec62ecfc05d5d4a23ce974eb3d7cb2c74da4d9b7aa396d66ff792be47481a04121632109d252d7d886f9174f89f9255fab1e212e38410126a0653623977fbb329ed4d9388be79f5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c88c9c210d87b53709a164577fa79c3f6766c5f5fbac5d3195ee56262a0b5d554c468aef8b00e9cda52a6bac56a47c5ca3c46d32917ee9a9dc216b1aa133aaac8fcf5215a420453ef47ba71833c549f9cc102a9e20a0e6ffcd46fb1e43996808417c5e171778574667d6f69c37f2e4c32cabac6bf6699343;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a798a7fa121d8ade8cef8e942e2acd11758926c8fbe583b107fb73a1be780879fd2b98d19388bdbdd915807cb0db775f68abeb79053cd8fe2ee858b34e656a6ebee6893cc3f8820610cb2abb581514c8771ad119fb97c3effe162591fd093f60eea0b1bd8f150382c48d9f7c93459f5dee1cf1cbf7949705;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f1d69c88afaf503d829cb038c8fc532fb88111265549a1f7d574aadada094e20181371ed35ff2e9c50ec64790534ef74ffa341446483bad6259b88a5e040dc8572befbecfd67e9fa7a1ae289c24c0fd36133d772c75f59a676733ed456ab8e12c4e65ffbdcefd3af1a7e01421b5d216e18c0bd2f7809fb7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbbf615a0f35148dc77c199142ee4f884fd70fcae26b94e2b4024727c847c028951ee834bfc21923e9c348a922e52ba3baf15c5f3d675387f0b1fe8c62cf63ee327d6d76e79f3bcd552901afe8711e5932ddfb48c6ef1207aee04276cd023cb79151af1841887b5248462cb523123502fd2de5b259ad57352;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc94457a07e2cb43e4b06d337e0f61d0f2a0fe62c68c4ea52fa5ab912db26c469f2aa22fb83f9328bbd8414c9876ec78863b78354eaae379958bda9ddd2314107a024aa3cbe4905852cf4ec85dd2a532714a39e949a982e7f48ba18065b5216518f92b28ddf7a447c4edd6036da127f40fa51793ac618fe44;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5258024b3ee140ba9d21d06f322ecb8e5620f502354df597858914e19955a27c9c313b660ed2cf0a152eaa49dfd69a473b812e833b748c42c52176c60916efe4583f62c58f70ff0e46c442f38ba1be1e931e2b888ead91b64cc0dd11a2fb48205927040c0467968421726abf7d098b44982a99c3d867d195;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b30ae78bd86e82d6d9978eafe9095c315bca0246d1bf1574361cd1d46e4f25e7f9202964092b6c78349f78f30c3053069cd371967c055a90376f310a6d13d20bff3c29a04cca544f0b63d874bf273dd032e1dd744e911b86e804772dc74410a2a338e1913d782697ca0e70f2a395c156aafa4496af5e31b0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1083c6f3db49d1c7672afac3bf7f2031d0fb371eacf1d44358a3065e1b7ec7340367b33cf4d9ed16e9ac30a780c63d7777c5eab9bf1d88998a631d6f7f8c583e2ce68d9086013494fa713eedffbfc210dcf09e54b64ae5791f3e3ce1385cb19e718596eeb4756df401f86e76582ae2b34acc5c8dcfad9e0c4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17313d66a6e3aaa7796a2f6e90020ec2fb166902d593c04046e6ef66c34adfd82dff247da2782300fd599373dd2e4c238a4e5a51a02afedd7def7c6f540b64d143dca73c99d8c8da923a2febc88e0bd98da0ddf7fab45572b2c64710f08da3acd9645f83c4e7b68266518de845d231dda03a9fc534b8acd41;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f41ef0dcb43c5226661ff191d3395ae37e62deeb4b9bfee9e8b2597edda729977eb6149b308ed750b58fe4ac55498b0c3e21b6845b97b250e030aa000ec8f7a41dac30381a05875b2caead4d49e3646db7bbc4d23152c97aab23fb7c292c0225b9dbe7c8a5c8e6adaa663efbf6754b4995ca91ce7d158c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12da9c5725b350427dcdf6fa0f2423809000bccd910534b0a2ef68ceaf22a4796cbcfc0947f3cad2a9f31073b97ffd9de4ed732b2b8e79fb4f375296d7bb73553602e2c89109a1b9a1beb53b1809fae1fc9e05bd5bbf0760e0e706a139a408779e9211b9d8cd5b239546a7969d8b0e5b4706d140e5890eda8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a342f5ef4ef3c62069b1e32d0b9c69042b1dd4974c7860a1ed76ae5d33df0d31dd6e2ae0fa63350ac8c56c2c8dd872cb653fab467161a1f77d4f4e67cb4c5c9c691ea0f535504bd893ec227e8a4f18b9b1cec9168c042a707109704b77cc67caac5a444619b061ecb685668742db4d5e4822249546d72497;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h171c981ccb354e226e0cf838769cb3cd771f3eb77f78f56943071dbaf2143bdf747386b5b029ba4af9394604466cc4221da2c0fa936943c50ee4d7ddae58a591c19cb64f9ad11386474c42598720efd1aa42b73d6179c8897fedbf4e3c20b6ee10991651078588eb3fad697be4e6a27e9613791e94983d6b7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2184dd735362d7bc1a2388731d0c273b8cf3d9036d325173c20ef3da5489cb5541d0f648b2c6ed4efcc3bd063e7af3d0035f607704b7d218530aa83b7051e3398b76ab9ae5eb15afc0d5e23b216a2e6a279e2c950f2e835c73079f994150143ac11dcb2aa54ca82b5969e9eac0fde57ff969f57db4cd9f2b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbcc8984fd43944884d84223f30405067c771be54788b3104cef7badd910cc9d7d312d65dc301fe215f75e351055d817037b6a20fcd0db7e0f5b39f10b0edb4d563c110529af0259e021824dd68dd0ed77cce7206a399896d5e1b3789aa9dd65434990b5252814e77dbfbab52b03aef95c7751a8e515504fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1db07dd329b3b1f44002e25376734e5d28e88ba5855cc6604a6a7b4ca0fea904e74e5057ad7f290cebdb993d0b8385313b439d006cfa4faf910256ceab7aa0951210d04f36dbae6bb4d4811981edac57cb9db78a254ba0009897a69d07bab9503fdfeea1b09e99b399371da60780157391d933ef72d19a470;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18ec8fad951ff1761105ae63cbcd555da3dd9397f7811053c02f142fabbaae2aea46d304eb487d4010a6708a356a1325a58faeb3e5ac1cfe083be2fe6b1dd12f280ab2df648f32acbfd6306f1d0aa87929ef01d98627545cb5e1f99864f025e6d8193afcb1c695e8fbcbb24370b66d07e574df912926cd93;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a494f1a31322dfdc3dcb4ed605df88ab30a232eb69c0a7cb6aa2fd3fe6960fd3d59dcfec3febaa1bbaa8ed50d23f3e303d6d19644a00f15008fda7accae9a2ddfcf1b889e6847507e3fcaa00494b1a9582fcc6e718328addcfc2b9a764db6ab32ac84147a814e21a846cabd60809fd96f26a2ce587cd80e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a52edaf7dc550fb1cfcb8e20c983397cbb33af2dc6d9d779693986e1e9bc4a60cdc0c4dc9a63493e237b469cc2e7124f82378aabea7042ef45cf1a2b0c7b0bcd30ec37a7d6ae1d34b6cc0d3d83eb04ae554448d7fb9742c92656a8fb66f6134d532ba1f4d617b2455d28aecc1557308633a6c77a17f17daf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e3a8340e6294f59bb6aab706f697d7ae02515f0b6b518e0202a5b25273e4603111ea56609f7f6786795a480328a452a6e5befa9fb6d7ccfd27013a3ec8a84d2d94798abe7045addf4174061e1199343e29931b0ac2fa7f2469af76b21dc6c339751dd30339d82a5a19bb8718732bd8c8d5db77b254d7ce0d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dbffa9e1ecb2c5f604201edb30f8d9fec6985a98696ec8336f8c941bbad9265450c914586b7cbe5f9fc46e7924999b0544918176cbfd3017b353f9c210150e1efe5fe0facb04c99f6c9b931e4a641aee6c2c5e2aa9425c34c652fa7e7080aa5ab0bf807e1aed68d5b24aaaf51c3ae49d6c420fe7885e8dc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h178704e07f54416e55954bdacd6e3693e462d8c4ccd164a3413d3913241b3b5e43f7f1df7adda20cc5d71991b5c3b7b02f53a0b072cb0230c44ce04871ecd11d0c28310a818c5b692b7b24d8927347513a316b166098570cf223b8af6c63a5f205f9cb0e2de42927dc8e798909311047221701e0599cfd5b7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1feba2f11647b3445939bd0d66286cd1a75e0152c6cef4bafd06ef39cbd71ee419c36b6eb93f1dd784e99b93106bc6ba64fe661f1f3a3a0e5d6321ca748290070791a8ade96caa7b0ca6be755f88eea32b1e49ba231b0fdb965d96ac48c51fe94710d159302cc1541b18579e83978852baef089aca38918bf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h92c1ad1f409b992aca1b4951ac5fc75b254de72f11d9354246e6aa0042ce651c4ae352c681f575c889ac2715b75f0f64b6c1d333ad5daaf4a122846deac34e4001a3ba4470fa1c304db4679aa6dca8d25d31fca7497421795993bdb04a7a0d32566779f3c01cc0a037067c5b62db1d4c9ee3278bdee8a98d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f69b74a0f6f9c74b2db9779e307ceb7c9ca35a01c68951b21b9df2abbe8ea76ccbbaa9da627ec6750aa42779e735e9194764a22c3083635135d36c163b38942d05028f43204c6455c173cdd2ea97a02c4f53c231f0e035f0cfc329cd3dcf08d04717fd209b82f5e8c9faa8e3103005451eb08d3b4d4cee45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h243851225bb943fa7486fab0baf461bc4b3273842eb76bb6ab29f3cf6e0a663dddc3cb071f03c87e92d7cd3bf16f309bea958577d3c20f210980194177c8b7e44e90bba81b3ee157b22f5e73718f51680530efb5b39325278fb3c3ae4675530208d6524c40f871fbd542338f556ae1242b97abd759038e6f;
        #1
        $finish();
    end
endmodule
