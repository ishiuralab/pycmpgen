module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20);
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    compressor_CLA486_12 compressor_CLA486_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20));
    initial begin
        src0 <= 486'h0;
        src1 <= 486'h0;
        src2 <= 486'h0;
        src3 <= 486'h0;
        src4 <= 486'h0;
        src5 <= 486'h0;
        src6 <= 486'h0;
        src7 <= 486'h0;
        src8 <= 486'h0;
        src9 <= 486'h0;
        src10 <= 486'h0;
        src11 <= 486'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA486_12(
    input [485:0]src0,
    input [485:0]src1,
    input [485:0]src2,
    input [485:0]src3,
    input [485:0]src4,
    input [485:0]src5,
    input [485:0]src6,
    input [485:0]src7,
    input [485:0]src8,
    input [485:0]src9,
    input [485:0]src10,
    input [485:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [0:0] comp_out19;
    wire [1:0] comp_out20;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out20[1], 1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], 1'h0}),
        .dst({dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [485:0] src0,
      input wire [485:0] src1,
      input wire [485:0] src2,
      input wire [485:0] src3,
      input wire [485:0] src4,
      input wire [485:0] src5,
      input wire [485:0] src6,
      input wire [485:0] src7,
      input wire [485:0] src8,
      input wire [485:0] src9,
      input wire [485:0] src10,
      input wire [485:0] src11,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [0:0] dst19,
      output wire [1:0] dst20);

   wire [485:0] stage0_0;
   wire [485:0] stage0_1;
   wire [485:0] stage0_2;
   wire [485:0] stage0_3;
   wire [485:0] stage0_4;
   wire [485:0] stage0_5;
   wire [485:0] stage0_6;
   wire [485:0] stage0_7;
   wire [485:0] stage0_8;
   wire [485:0] stage0_9;
   wire [485:0] stage0_10;
   wire [485:0] stage0_11;
   wire [85:0] stage1_0;
   wire [154:0] stage1_1;
   wire [197:0] stage1_2;
   wire [195:0] stage1_3;
   wire [240:0] stage1_4;
   wire [229:0] stage1_5;
   wire [169:0] stage1_6;
   wire [161:0] stage1_7;
   wire [238:0] stage1_8;
   wire [240:0] stage1_9;
   wire [179:0] stage1_10;
   wire [170:0] stage1_11;
   wire [156:0] stage1_12;
   wire [78:0] stage1_13;
   wire [30:0] stage2_0;
   wire [57:0] stage2_1;
   wire [53:0] stage2_2;
   wire [83:0] stage2_3;
   wire [88:0] stage2_4;
   wire [74:0] stage2_5;
   wire [97:0] stage2_6;
   wire [88:0] stage2_7;
   wire [70:0] stage2_8;
   wire [91:0] stage2_9;
   wire [98:0] stage2_10;
   wire [81:0] stage2_11;
   wire [111:0] stage2_12;
   wire [51:0] stage2_13;
   wire [26:0] stage2_14;
   wire [11:0] stage2_15;
   wire [13:0] stage3_0;
   wire [25:0] stage3_1;
   wire [16:0] stage3_2;
   wire [24:0] stage3_3;
   wire [33:0] stage3_4;
   wire [31:0] stage3_5;
   wire [44:0] stage3_6;
   wire [37:0] stage3_7;
   wire [30:0] stage3_8;
   wire [42:0] stage3_9;
   wire [37:0] stage3_10;
   wire [53:0] stage3_11;
   wire [46:0] stage3_12;
   wire [33:0] stage3_13;
   wire [25:0] stage3_14;
   wire [17:0] stage3_15;
   wire [4:0] stage3_16;
   wire [0:0] stage3_17;
   wire [8:0] stage4_0;
   wire [11:0] stage4_1;
   wire [6:0] stage4_2;
   wire [6:0] stage4_3;
   wire [12:0] stage4_4;
   wire [14:0] stage4_5;
   wire [15:0] stage4_6;
   wire [18:0] stage4_7;
   wire [12:0] stage4_8;
   wire [16:0] stage4_9;
   wire [18:0] stage4_10;
   wire [15:0] stage4_11;
   wire [17:0] stage4_12;
   wire [22:0] stage4_13;
   wire [16:0] stage4_14;
   wire [7:0] stage4_15;
   wire [11:0] stage4_16;
   wire [3:0] stage4_17;
   wire [6:0] stage5_0;
   wire [6:0] stage5_1;
   wire [4:0] stage5_2;
   wire [5:0] stage5_3;
   wire [3:0] stage5_4;
   wire [4:0] stage5_5;
   wire [6:0] stage5_6;
   wire [5:0] stage5_7;
   wire [11:0] stage5_8;
   wire [6:0] stage5_9;
   wire [7:0] stage5_10;
   wire [7:0] stage5_11;
   wire [6:0] stage5_12;
   wire [10:0] stage5_13;
   wire [7:0] stage5_14;
   wire [6:0] stage5_15;
   wire [3:0] stage5_16;
   wire [6:0] stage5_17;
   wire [1:0] stage5_18;
   wire [0:0] stage6_0;
   wire [6:0] stage6_1;
   wire [4:0] stage6_2;
   wire [6:0] stage6_3;
   wire [3:0] stage6_4;
   wire [0:0] stage6_5;
   wire [2:0] stage6_6;
   wire [2:0] stage6_7;
   wire [6:0] stage6_8;
   wire [2:0] stage6_9;
   wire [3:0] stage6_10;
   wire [3:0] stage6_11;
   wire [1:0] stage6_12;
   wire [5:0] stage6_13;
   wire [4:0] stage6_14;
   wire [1:0] stage6_15;
   wire [2:0] stage6_16;
   wire [3:0] stage6_17;
   wire [1:0] stage6_18;
   wire [0:0] stage6_19;
   wire [0:0] stage6_20;
   wire [0:0] stage7_0;
   wire [1:0] stage7_1;
   wire [1:0] stage7_2;
   wire [1:0] stage7_3;
   wire [1:0] stage7_4;
   wire [1:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [0:0] stage7_19;
   wire [1:0] stage7_20;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[10]},
      {stage0_3[20]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[11]},
      {stage0_3[21]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[56], stage0_0[57], stage0_0[58]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[12]},
      {stage0_3[22]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[59], stage0_0[60], stage0_0[61]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[13]},
      {stage0_3[23]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[62], stage0_0[63], stage0_0[64]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[14]},
      {stage0_3[24]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[65], stage0_0[66], stage0_0[67]},
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_2[15]},
      {stage0_3[25]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[68], stage0_0[69], stage0_0[70]},
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_2[16]},
      {stage0_3[26]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc207_4 gpc17 (
      {stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77]},
      {stage0_2[17], stage0_2[18]},
      {stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[17],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[18],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[19],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[20],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[21],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[22],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[114], stage0_0[115], stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[23],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[120], stage0_0[121], stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[24],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[126], stage0_0[127], stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[25],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[26],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[27],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[144], stage0_0[145], stage0_0[146], stage0_0[147], stage0_0[148], stage0_0[149]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[28],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153], stage0_0[154], stage0_0[155]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[29],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[156], stage0_0[157], stage0_0[158], stage0_0[159], stage0_0[160], stage0_0[161]},
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage1_4[30],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[162], stage0_0[163], stage0_0[164], stage0_0[165], stage0_0[166], stage0_0[167]},
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage1_4[31],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_0[168], stage0_0[169], stage0_0[170], stage0_0[171], stage0_0[172], stage0_0[173]},
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage1_4[32],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_0[174], stage0_0[175], stage0_0[176], stage0_0[177], stage0_0[178], stage0_0[179]},
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage1_4[33],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc606_5 gpc35 (
      {stage0_0[180], stage0_0[181], stage0_0[182], stage0_0[183], stage0_0[184], stage0_0[185]},
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126]},
      {stage1_4[34],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc606_5 gpc36 (
      {stage0_0[186], stage0_0[187], stage0_0[188], stage0_0[189], stage0_0[190], stage0_0[191]},
      {stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132]},
      {stage1_4[35],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195], stage0_0[196], stage0_0[197]},
      {stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138]},
      {stage1_4[36],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203]},
      {stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144]},
      {stage1_4[37],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209]},
      {stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150]},
      {stage1_4[38],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214], stage0_0[215]},
      {stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage1_4[39],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220], stage0_0[221]},
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162]},
      {stage1_4[40],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226], stage0_0[227]},
      {stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168]},
      {stage1_4[41],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232], stage0_0[233]},
      {stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174]},
      {stage1_4[42],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237], stage0_0[238], stage0_0[239]},
      {stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180]},
      {stage1_4[43],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243], stage0_0[244], stage0_0[245]},
      {stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186]},
      {stage1_4[44],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249], stage0_0[250], stage0_0[251]},
      {stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192]},
      {stage1_4[45],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255], stage0_0[256], stage0_0[257]},
      {stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198]},
      {stage1_4[46],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261], stage0_0[262], stage0_0[263]},
      {stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204]},
      {stage1_4[47],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267], stage0_0[268], stage0_0[269]},
      {stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210]},
      {stage1_4[48],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[270], stage0_0[271], stage0_0[272], stage0_0[273], stage0_0[274], stage0_0[275]},
      {stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216]},
      {stage1_4[49],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[276], stage0_0[277], stage0_0[278], stage0_0[279], stage0_0[280], stage0_0[281]},
      {stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222]},
      {stage1_4[50],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[282], stage0_0[283], stage0_0[284], stage0_0[285], stage0_0[286], stage0_0[287]},
      {stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228]},
      {stage1_4[51],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291], stage0_0[292], stage0_0[293]},
      {stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234]},
      {stage1_4[52],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297], stage0_0[298], stage0_0[299]},
      {stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240]},
      {stage1_4[53],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[300], stage0_0[301], stage0_0[302], stage0_0[303], stage0_0[304], stage0_0[305]},
      {stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246]},
      {stage1_4[54],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[306], stage0_0[307], stage0_0[308], stage0_0[309], stage0_0[310], stage0_0[311]},
      {stage0_2[247], stage0_2[248], stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252]},
      {stage1_4[55],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[312], stage0_0[313], stage0_0[314], stage0_0[315], stage0_0[316], stage0_0[317]},
      {stage0_2[253], stage0_2[254], stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258]},
      {stage1_4[56],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321], stage0_0[322], stage0_0[323]},
      {stage0_2[259], stage0_2[260], stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264]},
      {stage1_4[57],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327], stage0_0[328], stage0_0[329]},
      {stage0_2[265], stage0_2[266], stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270]},
      {stage1_4[58],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[330], stage0_0[331], stage0_0[332], stage0_0[333], stage0_0[334], stage0_0[335]},
      {stage0_2[271], stage0_2[272], stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276]},
      {stage1_4[59],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[336], stage0_0[337], stage0_0[338], stage0_0[339], stage0_0[340], stage0_0[341]},
      {stage0_2[277], stage0_2[278], stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282]},
      {stage1_4[60],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[342], stage0_0[343], stage0_0[344], stage0_0[345], stage0_0[346], stage0_0[347]},
      {stage0_2[283], stage0_2[284], stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288]},
      {stage1_4[61],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351], stage0_0[352], stage0_0[353]},
      {stage0_2[289], stage0_2[290], stage0_2[291], stage0_2[292], stage0_2[293], stage0_2[294]},
      {stage1_4[62],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357], stage0_0[358], stage0_0[359]},
      {stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299], stage0_2[300]},
      {stage1_4[63],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[360], stage0_0[361], stage0_0[362], stage0_0[363], stage0_0[364], stage0_0[365]},
      {stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305], stage0_2[306]},
      {stage1_4[64],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[366], stage0_0[367], stage0_0[368], stage0_0[369], stage0_0[370], stage0_0[371]},
      {stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311], stage0_2[312]},
      {stage1_4[65],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[372], stage0_0[373], stage0_0[374], stage0_0[375], stage0_0[376], stage0_0[377]},
      {stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317], stage0_2[318]},
      {stage1_4[66],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381], stage0_0[382], stage0_0[383]},
      {stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323], stage0_2[324]},
      {stage1_4[67],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387], stage0_0[388], stage0_0[389]},
      {stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329], stage0_2[330]},
      {stage1_4[68],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[390], stage0_0[391], stage0_0[392], stage0_0[393], stage0_0[394], stage0_0[395]},
      {stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335], stage0_2[336]},
      {stage1_4[69],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[396], stage0_0[397], stage0_0[398], stage0_0[399], stage0_0[400], stage0_0[401]},
      {stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341], stage0_2[342]},
      {stage1_4[70],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[402], stage0_0[403], stage0_0[404], stage0_0[405], stage0_0[406], stage0_0[407]},
      {stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347], stage0_2[348]},
      {stage1_4[71],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411], stage0_0[412], stage0_0[413]},
      {stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353], stage0_2[354]},
      {stage1_4[72],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417], stage0_0[418], stage0_0[419]},
      {stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358], stage0_2[359], stage0_2[360]},
      {stage1_4[73],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[420], stage0_0[421], stage0_0[422], stage0_0[423], stage0_0[424], stage0_0[425]},
      {stage0_2[361], stage0_2[362], stage0_2[363], stage0_2[364], stage0_2[365], stage0_2[366]},
      {stage1_4[74],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[426], stage0_0[427], stage0_0[428], stage0_0[429], stage0_0[430], stage0_0[431]},
      {stage0_2[367], stage0_2[368], stage0_2[369], stage0_2[370], stage0_2[371], stage0_2[372]},
      {stage1_4[75],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[432], stage0_0[433], stage0_0[434], stage0_0[435], stage0_0[436], stage0_0[437]},
      {stage0_2[373], stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377], stage0_2[378]},
      {stage1_4[76],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441], stage0_0[442], stage0_0[443]},
      {stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383], stage0_2[384]},
      {stage1_4[77],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447], stage0_0[448], stage0_0[449]},
      {stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388], stage0_2[389], stage0_2[390]},
      {stage1_4[78],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[450], stage0_0[451], stage0_0[452], stage0_0[453], stage0_0[454], stage0_0[455]},
      {stage0_2[391], stage0_2[392], stage0_2[393], stage0_2[394], stage0_2[395], stage0_2[396]},
      {stage1_4[79],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[456], stage0_0[457], stage0_0[458], stage0_0[459], stage0_0[460], stage0_0[461]},
      {stage0_2[397], stage0_2[398], stage0_2[399], stage0_2[400], stage0_2[401], stage0_2[402]},
      {stage1_4[80],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[462], stage0_0[463], stage0_0[464], stage0_0[465], stage0_0[466], stage0_0[467]},
      {stage0_2[403], stage0_2[404], stage0_2[405], stage0_2[406], stage0_2[407], stage0_2[408]},
      {stage1_4[81],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[468], stage0_0[469], stage0_0[470], stage0_0[471], stage0_0[472], stage0_0[473]},
      {stage0_2[409], stage0_2[410], stage0_2[411], stage0_2[412], stage0_2[413], stage0_2[414]},
      {stage1_4[82],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[474], stage0_0[475], stage0_0[476], stage0_0[477], stage0_0[478], stage0_0[479]},
      {stage0_2[415], stage0_2[416], stage0_2[417], stage0_2[418], stage0_2[419], stage0_2[420]},
      {stage1_4[83],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_0[480], stage0_0[481], stage0_0[482], stage0_0[483], stage0_0[484], stage0_0[485]},
      {stage0_2[421], stage0_2[422], stage0_2[423], stage0_2[424], stage0_2[425], stage0_2[426]},
      {stage1_4[84],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc606_5 gpc86 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[0],stage1_4[85],stage1_3[86],stage1_2[86],stage1_1[86]}
   );
   gpc606_5 gpc87 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[1],stage1_4[86],stage1_3[87],stage1_2[87],stage1_1[87]}
   );
   gpc606_5 gpc88 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[2],stage1_4[87],stage1_3[88],stage1_2[88],stage1_1[88]}
   );
   gpc606_5 gpc89 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[3],stage1_4[88],stage1_3[89],stage1_2[89],stage1_1[89]}
   );
   gpc606_5 gpc90 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[4],stage1_4[89],stage1_3[90],stage1_2[90],stage1_1[90]}
   );
   gpc606_5 gpc91 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[5],stage1_4[90],stage1_3[91],stage1_2[91],stage1_1[91]}
   );
   gpc606_5 gpc92 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[6],stage1_4[91],stage1_3[92],stage1_2[92],stage1_1[92]}
   );
   gpc606_5 gpc93 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[7],stage1_4[92],stage1_3[93],stage1_2[93],stage1_1[93]}
   );
   gpc606_5 gpc94 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[8],stage1_4[93],stage1_3[94],stage1_2[94],stage1_1[94]}
   );
   gpc606_5 gpc95 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[9],stage1_4[94],stage1_3[95],stage1_2[95],stage1_1[95]}
   );
   gpc606_5 gpc96 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[10],stage1_4[95],stage1_3[96],stage1_2[96],stage1_1[96]}
   );
   gpc606_5 gpc97 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98]},
      {stage1_5[11],stage1_4[96],stage1_3[97],stage1_2[97],stage1_1[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage1_5[12],stage1_4[97],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110]},
      {stage1_5[13],stage1_4[98],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage1_5[14],stage1_4[99],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122]},
      {stage1_5[15],stage1_4[100],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128]},
      {stage1_5[16],stage1_4[101],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[174], stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179]},
      {stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134]},
      {stage1_5[17],stage1_4[102],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185]},
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140]},
      {stage1_5[18],stage1_4[103],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191]},
      {stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146]},
      {stage1_5[19],stage1_4[104],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197]},
      {stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152]},
      {stage1_5[20],stage1_4[105],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203]},
      {stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158]},
      {stage1_5[21],stage1_4[106],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209]},
      {stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164]},
      {stage1_5[22],stage1_4[107],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215]},
      {stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170]},
      {stage1_5[23],stage1_4[108],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221]},
      {stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176]},
      {stage1_5[24],stage1_4[109],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227]},
      {stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182]},
      {stage1_5[25],stage1_4[110],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233]},
      {stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188]},
      {stage1_5[26],stage1_4[111],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[234], stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239]},
      {stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194]},
      {stage1_5[27],stage1_4[112],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[240], stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245]},
      {stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200]},
      {stage1_5[28],stage1_4[113],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[246], stage0_1[247], stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251]},
      {stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage1_5[29],stage1_4[114],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[252], stage0_1[253], stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257]},
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212]},
      {stage1_5[30],stage1_4[115],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[258], stage0_1[259], stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263]},
      {stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218]},
      {stage1_5[31],stage1_4[116],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[264], stage0_1[265], stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269]},
      {stage0_3[219], stage0_3[220], stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224]},
      {stage1_5[32],stage1_4[117],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[270], stage0_1[271], stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275]},
      {stage0_3[225], stage0_3[226], stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230]},
      {stage1_5[33],stage1_4[118],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[276], stage0_1[277], stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281]},
      {stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236]},
      {stage1_5[34],stage1_4[119],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[282], stage0_1[283], stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287]},
      {stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242]},
      {stage1_5[35],stage1_4[120],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[288], stage0_1[289], stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293]},
      {stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246], stage0_3[247], stage0_3[248]},
      {stage1_5[36],stage1_4[121],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[294], stage0_1[295], stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299]},
      {stage0_3[249], stage0_3[250], stage0_3[251], stage0_3[252], stage0_3[253], stage0_3[254]},
      {stage1_5[37],stage1_4[122],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[300], stage0_1[301], stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305]},
      {stage0_3[255], stage0_3[256], stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260]},
      {stage1_5[38],stage1_4[123],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[306], stage0_1[307], stage0_1[308], stage0_1[309], stage0_1[310], stage0_1[311]},
      {stage0_3[261], stage0_3[262], stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266]},
      {stage1_5[39],stage1_4[124],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[312], stage0_1[313], stage0_1[314], stage0_1[315], stage0_1[316], stage0_1[317]},
      {stage0_3[267], stage0_3[268], stage0_3[269], stage0_3[270], stage0_3[271], stage0_3[272]},
      {stage1_5[40],stage1_4[125],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[318], stage0_1[319], stage0_1[320], stage0_1[321], stage0_1[322], stage0_1[323]},
      {stage0_3[273], stage0_3[274], stage0_3[275], stage0_3[276], stage0_3[277], stage0_3[278]},
      {stage1_5[41],stage1_4[126],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[324], stage0_1[325], stage0_1[326], stage0_1[327], stage0_1[328], stage0_1[329]},
      {stage0_3[279], stage0_3[280], stage0_3[281], stage0_3[282], stage0_3[283], stage0_3[284]},
      {stage1_5[42],stage1_4[127],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[330], stage0_1[331], stage0_1[332], stage0_1[333], stage0_1[334], stage0_1[335]},
      {stage0_3[285], stage0_3[286], stage0_3[287], stage0_3[288], stage0_3[289], stage0_3[290]},
      {stage1_5[43],stage1_4[128],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[336], stage0_1[337], stage0_1[338], stage0_1[339], stage0_1[340], stage0_1[341]},
      {stage0_3[291], stage0_3[292], stage0_3[293], stage0_3[294], stage0_3[295], stage0_3[296]},
      {stage1_5[44],stage1_4[129],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[342], stage0_1[343], stage0_1[344], stage0_1[345], stage0_1[346], stage0_1[347]},
      {stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300], stage0_3[301], stage0_3[302]},
      {stage1_5[45],stage1_4[130],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[348], stage0_1[349], stage0_1[350], stage0_1[351], stage0_1[352], stage0_1[353]},
      {stage0_3[303], stage0_3[304], stage0_3[305], stage0_3[306], stage0_3[307], stage0_3[308]},
      {stage1_5[46],stage1_4[131],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[354], stage0_1[355], stage0_1[356], stage0_1[357], stage0_1[358], stage0_1[359]},
      {stage0_3[309], stage0_3[310], stage0_3[311], stage0_3[312], stage0_3[313], stage0_3[314]},
      {stage1_5[47],stage1_4[132],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[360], stage0_1[361], stage0_1[362], stage0_1[363], stage0_1[364], stage0_1[365]},
      {stage0_3[315], stage0_3[316], stage0_3[317], stage0_3[318], stage0_3[319], stage0_3[320]},
      {stage1_5[48],stage1_4[133],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[366], stage0_1[367], stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371]},
      {stage0_3[321], stage0_3[322], stage0_3[323], stage0_3[324], stage0_3[325], stage0_3[326]},
      {stage1_5[49],stage1_4[134],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_1[372], stage0_1[373], stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377]},
      {stage0_3[327], stage0_3[328], stage0_3[329], stage0_3[330], stage0_3[331], stage0_3[332]},
      {stage1_5[50],stage1_4[135],stage1_3[136],stage1_2[136],stage1_1[136]}
   );
   gpc606_5 gpc137 (
      {stage0_1[378], stage0_1[379], stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383]},
      {stage0_3[333], stage0_3[334], stage0_3[335], stage0_3[336], stage0_3[337], stage0_3[338]},
      {stage1_5[51],stage1_4[136],stage1_3[137],stage1_2[137],stage1_1[137]}
   );
   gpc606_5 gpc138 (
      {stage0_1[384], stage0_1[385], stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389]},
      {stage0_3[339], stage0_3[340], stage0_3[341], stage0_3[342], stage0_3[343], stage0_3[344]},
      {stage1_5[52],stage1_4[137],stage1_3[138],stage1_2[138],stage1_1[138]}
   );
   gpc606_5 gpc139 (
      {stage0_1[390], stage0_1[391], stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395]},
      {stage0_3[345], stage0_3[346], stage0_3[347], stage0_3[348], stage0_3[349], stage0_3[350]},
      {stage1_5[53],stage1_4[138],stage1_3[139],stage1_2[139],stage1_1[139]}
   );
   gpc606_5 gpc140 (
      {stage0_1[396], stage0_1[397], stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401]},
      {stage0_3[351], stage0_3[352], stage0_3[353], stage0_3[354], stage0_3[355], stage0_3[356]},
      {stage1_5[54],stage1_4[139],stage1_3[140],stage1_2[140],stage1_1[140]}
   );
   gpc606_5 gpc141 (
      {stage0_1[402], stage0_1[403], stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407]},
      {stage0_3[357], stage0_3[358], stage0_3[359], stage0_3[360], stage0_3[361], stage0_3[362]},
      {stage1_5[55],stage1_4[140],stage1_3[141],stage1_2[141],stage1_1[141]}
   );
   gpc606_5 gpc142 (
      {stage0_1[408], stage0_1[409], stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413]},
      {stage0_3[363], stage0_3[364], stage0_3[365], stage0_3[366], stage0_3[367], stage0_3[368]},
      {stage1_5[56],stage1_4[141],stage1_3[142],stage1_2[142],stage1_1[142]}
   );
   gpc606_5 gpc143 (
      {stage0_1[414], stage0_1[415], stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419]},
      {stage0_3[369], stage0_3[370], stage0_3[371], stage0_3[372], stage0_3[373], stage0_3[374]},
      {stage1_5[57],stage1_4[142],stage1_3[143],stage1_2[143],stage1_1[143]}
   );
   gpc606_5 gpc144 (
      {stage0_1[420], stage0_1[421], stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425]},
      {stage0_3[375], stage0_3[376], stage0_3[377], stage0_3[378], stage0_3[379], stage0_3[380]},
      {stage1_5[58],stage1_4[143],stage1_3[144],stage1_2[144],stage1_1[144]}
   );
   gpc606_5 gpc145 (
      {stage0_1[426], stage0_1[427], stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431]},
      {stage0_3[381], stage0_3[382], stage0_3[383], stage0_3[384], stage0_3[385], stage0_3[386]},
      {stage1_5[59],stage1_4[144],stage1_3[145],stage1_2[145],stage1_1[145]}
   );
   gpc606_5 gpc146 (
      {stage0_1[432], stage0_1[433], stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437]},
      {stage0_3[387], stage0_3[388], stage0_3[389], stage0_3[390], stage0_3[391], stage0_3[392]},
      {stage1_5[60],stage1_4[145],stage1_3[146],stage1_2[146],stage1_1[146]}
   );
   gpc606_5 gpc147 (
      {stage0_1[438], stage0_1[439], stage0_1[440], stage0_1[441], stage0_1[442], stage0_1[443]},
      {stage0_3[393], stage0_3[394], stage0_3[395], stage0_3[396], stage0_3[397], stage0_3[398]},
      {stage1_5[61],stage1_4[146],stage1_3[147],stage1_2[147],stage1_1[147]}
   );
   gpc606_5 gpc148 (
      {stage0_1[444], stage0_1[445], stage0_1[446], stage0_1[447], stage0_1[448], stage0_1[449]},
      {stage0_3[399], stage0_3[400], stage0_3[401], stage0_3[402], stage0_3[403], stage0_3[404]},
      {stage1_5[62],stage1_4[147],stage1_3[148],stage1_2[148],stage1_1[148]}
   );
   gpc606_5 gpc149 (
      {stage0_1[450], stage0_1[451], stage0_1[452], stage0_1[453], stage0_1[454], stage0_1[455]},
      {stage0_3[405], stage0_3[406], stage0_3[407], stage0_3[408], stage0_3[409], stage0_3[410]},
      {stage1_5[63],stage1_4[148],stage1_3[149],stage1_2[149],stage1_1[149]}
   );
   gpc606_5 gpc150 (
      {stage0_1[456], stage0_1[457], stage0_1[458], stage0_1[459], stage0_1[460], stage0_1[461]},
      {stage0_3[411], stage0_3[412], stage0_3[413], stage0_3[414], stage0_3[415], stage0_3[416]},
      {stage1_5[64],stage1_4[149],stage1_3[150],stage1_2[150],stage1_1[150]}
   );
   gpc606_5 gpc151 (
      {stage0_1[462], stage0_1[463], stage0_1[464], stage0_1[465], stage0_1[466], stage0_1[467]},
      {stage0_3[417], stage0_3[418], stage0_3[419], stage0_3[420], stage0_3[421], stage0_3[422]},
      {stage1_5[65],stage1_4[150],stage1_3[151],stage1_2[151],stage1_1[151]}
   );
   gpc606_5 gpc152 (
      {stage0_1[468], stage0_1[469], stage0_1[470], stage0_1[471], stage0_1[472], stage0_1[473]},
      {stage0_3[423], stage0_3[424], stage0_3[425], stage0_3[426], stage0_3[427], stage0_3[428]},
      {stage1_5[66],stage1_4[151],stage1_3[152],stage1_2[152],stage1_1[152]}
   );
   gpc606_5 gpc153 (
      {stage0_1[474], stage0_1[475], stage0_1[476], stage0_1[477], stage0_1[478], stage0_1[479]},
      {stage0_3[429], stage0_3[430], stage0_3[431], stage0_3[432], stage0_3[433], stage0_3[434]},
      {stage1_5[67],stage1_4[152],stage1_3[153],stage1_2[153],stage1_1[153]}
   );
   gpc606_5 gpc154 (
      {stage0_1[480], stage0_1[481], stage0_1[482], stage0_1[483], stage0_1[484], stage0_1[485]},
      {stage0_3[435], stage0_3[436], stage0_3[437], stage0_3[438], stage0_3[439], stage0_3[440]},
      {stage1_5[68],stage1_4[153],stage1_3[154],stage1_2[154],stage1_1[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[427], stage0_2[428], stage0_2[429], stage0_2[430], stage0_2[431]},
      {stage0_3[441]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[69],stage1_4[154],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[432], stage0_2[433], stage0_2[434], stage0_2[435], stage0_2[436]},
      {stage0_3[442]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[70],stage1_4[155],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_2[437], stage0_2[438], stage0_2[439], stage0_2[440], stage0_2[441]},
      {stage0_3[443]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[71],stage1_4[156],stage1_3[157],stage1_2[157]}
   );
   gpc615_5 gpc158 (
      {stage0_2[442], stage0_2[443], stage0_2[444], stage0_2[445], stage0_2[446]},
      {stage0_3[444]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[72],stage1_4[157],stage1_3[158],stage1_2[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[445], stage0_3[446], stage0_3[447], stage0_3[448], stage0_3[449]},
      {stage0_4[24]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[4],stage1_5[73],stage1_4[158],stage1_3[159]}
   );
   gpc606_5 gpc160 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[5],stage1_5[74],stage1_4[159]}
   );
   gpc606_5 gpc161 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[6],stage1_5[75],stage1_4[160]}
   );
   gpc606_5 gpc162 (
      {stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[7],stage1_5[76],stage1_4[161]}
   );
   gpc606_5 gpc163 (
      {stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[8],stage1_5[77],stage1_4[162]}
   );
   gpc606_5 gpc164 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[9],stage1_5[78],stage1_4[163]}
   );
   gpc606_5 gpc165 (
      {stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[10],stage1_5[79],stage1_4[164]}
   );
   gpc606_5 gpc166 (
      {stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[11],stage1_5[80],stage1_4[165]}
   );
   gpc606_5 gpc167 (
      {stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[12],stage1_5[81],stage1_4[166]}
   );
   gpc606_5 gpc168 (
      {stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[9],stage1_6[13],stage1_5[82],stage1_4[167]}
   );
   gpc606_5 gpc169 (
      {stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[10],stage1_6[14],stage1_5[83],stage1_4[168]}
   );
   gpc606_5 gpc170 (
      {stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[11],stage1_6[15],stage1_5[84],stage1_4[169]}
   );
   gpc606_5 gpc171 (
      {stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[12],stage1_6[16],stage1_5[85],stage1_4[170]}
   );
   gpc606_5 gpc172 (
      {stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[13],stage1_6[17],stage1_5[86],stage1_4[171]}
   );
   gpc606_5 gpc173 (
      {stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[14],stage1_6[18],stage1_5[87],stage1_4[172]}
   );
   gpc606_5 gpc174 (
      {stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[15],stage1_6[19],stage1_5[88],stage1_4[173]}
   );
   gpc606_5 gpc175 (
      {stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[16],stage1_6[20],stage1_5[89],stage1_4[174]}
   );
   gpc606_5 gpc176 (
      {stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[17],stage1_6[21],stage1_5[90],stage1_4[175]}
   );
   gpc606_5 gpc177 (
      {stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[18],stage1_6[22],stage1_5[91],stage1_4[176]}
   );
   gpc606_5 gpc178 (
      {stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[19],stage1_6[23],stage1_5[92],stage1_4[177]}
   );
   gpc606_5 gpc179 (
      {stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[20],stage1_6[24],stage1_5[93],stage1_4[178]}
   );
   gpc606_5 gpc180 (
      {stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[21],stage1_6[25],stage1_5[94],stage1_4[179]}
   );
   gpc606_5 gpc181 (
      {stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[22],stage1_6[26],stage1_5[95],stage1_4[180]}
   );
   gpc606_5 gpc182 (
      {stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161], stage0_4[162]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[23],stage1_6[27],stage1_5[96],stage1_4[181]}
   );
   gpc606_5 gpc183 (
      {stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167], stage0_4[168]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[24],stage1_6[28],stage1_5[97],stage1_4[182]}
   );
   gpc606_5 gpc184 (
      {stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173], stage0_4[174]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[25],stage1_6[29],stage1_5[98],stage1_4[183]}
   );
   gpc606_5 gpc185 (
      {stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178], stage0_4[179], stage0_4[180]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[26],stage1_6[30],stage1_5[99],stage1_4[184]}
   );
   gpc606_5 gpc186 (
      {stage0_4[181], stage0_4[182], stage0_4[183], stage0_4[184], stage0_4[185], stage0_4[186]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[27],stage1_6[31],stage1_5[100],stage1_4[185]}
   );
   gpc606_5 gpc187 (
      {stage0_4[187], stage0_4[188], stage0_4[189], stage0_4[190], stage0_4[191], stage0_4[192]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[28],stage1_6[32],stage1_5[101],stage1_4[186]}
   );
   gpc606_5 gpc188 (
      {stage0_4[193], stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[29],stage1_6[33],stage1_5[102],stage1_4[187]}
   );
   gpc606_5 gpc189 (
      {stage0_4[199], stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[30],stage1_6[34],stage1_5[103],stage1_4[188]}
   );
   gpc606_5 gpc190 (
      {stage0_4[205], stage0_4[206], stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[31],stage1_6[35],stage1_5[104],stage1_4[189]}
   );
   gpc606_5 gpc191 (
      {stage0_4[211], stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[32],stage1_6[36],stage1_5[105],stage1_4[190]}
   );
   gpc606_5 gpc192 (
      {stage0_4[217], stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[33],stage1_6[37],stage1_5[106],stage1_4[191]}
   );
   gpc606_5 gpc193 (
      {stage0_4[223], stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[34],stage1_6[38],stage1_5[107],stage1_4[192]}
   );
   gpc606_5 gpc194 (
      {stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[35],stage1_6[39],stage1_5[108],stage1_4[193]}
   );
   gpc606_5 gpc195 (
      {stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[36],stage1_6[40],stage1_5[109],stage1_4[194]}
   );
   gpc606_5 gpc196 (
      {stage0_4[241], stage0_4[242], stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[37],stage1_6[41],stage1_5[110],stage1_4[195]}
   );
   gpc606_5 gpc197 (
      {stage0_4[247], stage0_4[248], stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[38],stage1_6[42],stage1_5[111],stage1_4[196]}
   );
   gpc606_5 gpc198 (
      {stage0_4[253], stage0_4[254], stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[39],stage1_6[43],stage1_5[112],stage1_4[197]}
   );
   gpc606_5 gpc199 (
      {stage0_4[259], stage0_4[260], stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[40],stage1_6[44],stage1_5[113],stage1_4[198]}
   );
   gpc606_5 gpc200 (
      {stage0_4[265], stage0_4[266], stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[41],stage1_6[45],stage1_5[114],stage1_4[199]}
   );
   gpc606_5 gpc201 (
      {stage0_4[271], stage0_4[272], stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[42],stage1_6[46],stage1_5[115],stage1_4[200]}
   );
   gpc606_5 gpc202 (
      {stage0_4[277], stage0_4[278], stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[43],stage1_6[47],stage1_5[116],stage1_4[201]}
   );
   gpc606_5 gpc203 (
      {stage0_4[283], stage0_4[284], stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[44],stage1_6[48],stage1_5[117],stage1_4[202]}
   );
   gpc606_5 gpc204 (
      {stage0_4[289], stage0_4[290], stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[45],stage1_6[49],stage1_5[118],stage1_4[203]}
   );
   gpc606_5 gpc205 (
      {stage0_4[295], stage0_4[296], stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[46],stage1_6[50],stage1_5[119],stage1_4[204]}
   );
   gpc606_5 gpc206 (
      {stage0_4[301], stage0_4[302], stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[47],stage1_6[51],stage1_5[120],stage1_4[205]}
   );
   gpc606_5 gpc207 (
      {stage0_4[307], stage0_4[308], stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[48],stage1_6[52],stage1_5[121],stage1_4[206]}
   );
   gpc606_5 gpc208 (
      {stage0_4[313], stage0_4[314], stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[49],stage1_6[53],stage1_5[122],stage1_4[207]}
   );
   gpc606_5 gpc209 (
      {stage0_4[319], stage0_4[320], stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[50],stage1_6[54],stage1_5[123],stage1_4[208]}
   );
   gpc606_5 gpc210 (
      {stage0_4[325], stage0_4[326], stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[51],stage1_6[55],stage1_5[124],stage1_4[209]}
   );
   gpc606_5 gpc211 (
      {stage0_4[331], stage0_4[332], stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[52],stage1_6[56],stage1_5[125],stage1_4[210]}
   );
   gpc606_5 gpc212 (
      {stage0_4[337], stage0_4[338], stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[53],stage1_6[57],stage1_5[126],stage1_4[211]}
   );
   gpc606_5 gpc213 (
      {stage0_4[343], stage0_4[344], stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[54],stage1_6[58],stage1_5[127],stage1_4[212]}
   );
   gpc606_5 gpc214 (
      {stage0_4[349], stage0_4[350], stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[55],stage1_6[59],stage1_5[128],stage1_4[213]}
   );
   gpc606_5 gpc215 (
      {stage0_4[355], stage0_4[356], stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360]},
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335]},
      {stage1_8[55],stage1_7[56],stage1_6[60],stage1_5[129],stage1_4[214]}
   );
   gpc606_5 gpc216 (
      {stage0_4[361], stage0_4[362], stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366]},
      {stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340], stage0_6[341]},
      {stage1_8[56],stage1_7[57],stage1_6[61],stage1_5[130],stage1_4[215]}
   );
   gpc606_5 gpc217 (
      {stage0_4[367], stage0_4[368], stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372]},
      {stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345], stage0_6[346], stage0_6[347]},
      {stage1_8[57],stage1_7[58],stage1_6[62],stage1_5[131],stage1_4[216]}
   );
   gpc606_5 gpc218 (
      {stage0_4[373], stage0_4[374], stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378]},
      {stage0_6[348], stage0_6[349], stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353]},
      {stage1_8[58],stage1_7[59],stage1_6[63],stage1_5[132],stage1_4[217]}
   );
   gpc606_5 gpc219 (
      {stage0_4[379], stage0_4[380], stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384]},
      {stage0_6[354], stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage1_8[59],stage1_7[60],stage1_6[64],stage1_5[133],stage1_4[218]}
   );
   gpc606_5 gpc220 (
      {stage0_4[385], stage0_4[386], stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390]},
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365]},
      {stage1_8[60],stage1_7[61],stage1_6[65],stage1_5[134],stage1_4[219]}
   );
   gpc606_5 gpc221 (
      {stage0_4[391], stage0_4[392], stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396]},
      {stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370], stage0_6[371]},
      {stage1_8[61],stage1_7[62],stage1_6[66],stage1_5[135],stage1_4[220]}
   );
   gpc606_5 gpc222 (
      {stage0_4[397], stage0_4[398], stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402]},
      {stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375], stage0_6[376], stage0_6[377]},
      {stage1_8[62],stage1_7[63],stage1_6[67],stage1_5[136],stage1_4[221]}
   );
   gpc606_5 gpc223 (
      {stage0_4[403], stage0_4[404], stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408]},
      {stage0_6[378], stage0_6[379], stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383]},
      {stage1_8[63],stage1_7[64],stage1_6[68],stage1_5[137],stage1_4[222]}
   );
   gpc606_5 gpc224 (
      {stage0_4[409], stage0_4[410], stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414]},
      {stage0_6[384], stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage1_8[64],stage1_7[65],stage1_6[69],stage1_5[138],stage1_4[223]}
   );
   gpc606_5 gpc225 (
      {stage0_4[415], stage0_4[416], stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420]},
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395]},
      {stage1_8[65],stage1_7[66],stage1_6[70],stage1_5[139],stage1_4[224]}
   );
   gpc606_5 gpc226 (
      {stage0_4[421], stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426]},
      {stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400], stage0_6[401]},
      {stage1_8[66],stage1_7[67],stage1_6[71],stage1_5[140],stage1_4[225]}
   );
   gpc606_5 gpc227 (
      {stage0_4[427], stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431], stage0_4[432]},
      {stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405], stage0_6[406], stage0_6[407]},
      {stage1_8[67],stage1_7[68],stage1_6[72],stage1_5[141],stage1_4[226]}
   );
   gpc606_5 gpc228 (
      {stage0_4[433], stage0_4[434], stage0_4[435], stage0_4[436], stage0_4[437], stage0_4[438]},
      {stage0_6[408], stage0_6[409], stage0_6[410], stage0_6[411], stage0_6[412], stage0_6[413]},
      {stage1_8[68],stage1_7[69],stage1_6[73],stage1_5[142],stage1_4[227]}
   );
   gpc606_5 gpc229 (
      {stage0_4[439], stage0_4[440], stage0_4[441], stage0_4[442], stage0_4[443], stage0_4[444]},
      {stage0_6[414], stage0_6[415], stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419]},
      {stage1_8[69],stage1_7[70],stage1_6[74],stage1_5[143],stage1_4[228]}
   );
   gpc606_5 gpc230 (
      {stage0_4[445], stage0_4[446], stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450]},
      {stage0_6[420], stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425]},
      {stage1_8[70],stage1_7[71],stage1_6[75],stage1_5[144],stage1_4[229]}
   );
   gpc615_5 gpc231 (
      {stage0_4[451], stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455]},
      {stage0_5[6]},
      {stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430], stage0_6[431]},
      {stage1_8[71],stage1_7[72],stage1_6[76],stage1_5[145],stage1_4[230]}
   );
   gpc615_5 gpc232 (
      {stage0_4[456], stage0_4[457], stage0_4[458], stage0_4[459], stage0_4[460]},
      {stage0_5[7]},
      {stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435], stage0_6[436], stage0_6[437]},
      {stage1_8[72],stage1_7[73],stage1_6[77],stage1_5[146],stage1_4[231]}
   );
   gpc615_5 gpc233 (
      {stage0_4[461], stage0_4[462], stage0_4[463], stage0_4[464], stage0_4[465]},
      {stage0_5[8]},
      {stage0_6[438], stage0_6[439], stage0_6[440], stage0_6[441], stage0_6[442], stage0_6[443]},
      {stage1_8[73],stage1_7[74],stage1_6[78],stage1_5[147],stage1_4[232]}
   );
   gpc615_5 gpc234 (
      {stage0_4[466], stage0_4[467], stage0_4[468], stage0_4[469], stage0_4[470]},
      {stage0_5[9]},
      {stage0_6[444], stage0_6[445], stage0_6[446], stage0_6[447], stage0_6[448], stage0_6[449]},
      {stage1_8[74],stage1_7[75],stage1_6[79],stage1_5[148],stage1_4[233]}
   );
   gpc615_5 gpc235 (
      {stage0_4[471], stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475]},
      {stage0_5[10]},
      {stage0_6[450], stage0_6[451], stage0_6[452], stage0_6[453], stage0_6[454], stage0_6[455]},
      {stage1_8[75],stage1_7[76],stage1_6[80],stage1_5[149],stage1_4[234]}
   );
   gpc615_5 gpc236 (
      {stage0_4[476], stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480]},
      {stage0_5[11]},
      {stage0_6[456], stage0_6[457], stage0_6[458], stage0_6[459], stage0_6[460], stage0_6[461]},
      {stage1_8[76],stage1_7[77],stage1_6[81],stage1_5[150],stage1_4[235]}
   );
   gpc606_5 gpc237 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[77],stage1_7[78],stage1_6[82],stage1_5[151]}
   );
   gpc606_5 gpc238 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[78],stage1_7[79],stage1_6[83],stage1_5[152]}
   );
   gpc606_5 gpc239 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[79],stage1_7[80],stage1_6[84],stage1_5[153]}
   );
   gpc606_5 gpc240 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[80],stage1_7[81],stage1_6[85],stage1_5[154]}
   );
   gpc606_5 gpc241 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[81],stage1_7[82],stage1_6[86],stage1_5[155]}
   );
   gpc606_5 gpc242 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[82],stage1_7[83],stage1_6[87],stage1_5[156]}
   );
   gpc606_5 gpc243 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[83],stage1_7[84],stage1_6[88],stage1_5[157]}
   );
   gpc606_5 gpc244 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[84],stage1_7[85],stage1_6[89],stage1_5[158]}
   );
   gpc606_5 gpc245 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[85],stage1_7[86],stage1_6[90],stage1_5[159]}
   );
   gpc606_5 gpc246 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[86],stage1_7[87],stage1_6[91],stage1_5[160]}
   );
   gpc606_5 gpc247 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[87],stage1_7[88],stage1_6[92],stage1_5[161]}
   );
   gpc606_5 gpc248 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[88],stage1_7[89],stage1_6[93],stage1_5[162]}
   );
   gpc606_5 gpc249 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[89],stage1_7[90],stage1_6[94],stage1_5[163]}
   );
   gpc606_5 gpc250 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[90],stage1_7[91],stage1_6[95],stage1_5[164]}
   );
   gpc606_5 gpc251 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[91],stage1_7[92],stage1_6[96],stage1_5[165]}
   );
   gpc606_5 gpc252 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[92],stage1_7[93],stage1_6[97],stage1_5[166]}
   );
   gpc606_5 gpc253 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[93],stage1_7[94],stage1_6[98],stage1_5[167]}
   );
   gpc606_5 gpc254 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[94],stage1_7[95],stage1_6[99],stage1_5[168]}
   );
   gpc606_5 gpc255 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[95],stage1_7[96],stage1_6[100],stage1_5[169]}
   );
   gpc606_5 gpc256 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[96],stage1_7[97],stage1_6[101],stage1_5[170]}
   );
   gpc606_5 gpc257 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[97],stage1_7[98],stage1_6[102],stage1_5[171]}
   );
   gpc606_5 gpc258 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[98],stage1_7[99],stage1_6[103],stage1_5[172]}
   );
   gpc606_5 gpc259 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[99],stage1_7[100],stage1_6[104],stage1_5[173]}
   );
   gpc606_5 gpc260 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[100],stage1_7[101],stage1_6[105],stage1_5[174]}
   );
   gpc606_5 gpc261 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[101],stage1_7[102],stage1_6[106],stage1_5[175]}
   );
   gpc606_5 gpc262 (
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[102],stage1_7[103],stage1_6[107],stage1_5[176]}
   );
   gpc606_5 gpc263 (
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[103],stage1_7[104],stage1_6[108],stage1_5[177]}
   );
   gpc606_5 gpc264 (
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[104],stage1_7[105],stage1_6[109],stage1_5[178]}
   );
   gpc606_5 gpc265 (
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[105],stage1_7[106],stage1_6[110],stage1_5[179]}
   );
   gpc606_5 gpc266 (
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[106],stage1_7[107],stage1_6[111],stage1_5[180]}
   );
   gpc606_5 gpc267 (
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[107],stage1_7[108],stage1_6[112],stage1_5[181]}
   );
   gpc606_5 gpc268 (
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[108],stage1_7[109],stage1_6[113],stage1_5[182]}
   );
   gpc606_5 gpc269 (
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[109],stage1_7[110],stage1_6[114],stage1_5[183]}
   );
   gpc606_5 gpc270 (
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[110],stage1_7[111],stage1_6[115],stage1_5[184]}
   );
   gpc606_5 gpc271 (
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[111],stage1_7[112],stage1_6[116],stage1_5[185]}
   );
   gpc606_5 gpc272 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[112],stage1_7[113],stage1_6[117],stage1_5[186]}
   );
   gpc606_5 gpc273 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[113],stage1_7[114],stage1_6[118],stage1_5[187]}
   );
   gpc606_5 gpc274 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[114],stage1_7[115],stage1_6[119],stage1_5[188]}
   );
   gpc606_5 gpc275 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[115],stage1_7[116],stage1_6[120],stage1_5[189]}
   );
   gpc606_5 gpc276 (
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[116],stage1_7[117],stage1_6[121],stage1_5[190]}
   );
   gpc606_5 gpc277 (
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[117],stage1_7[118],stage1_6[122],stage1_5[191]}
   );
   gpc606_5 gpc278 (
      {stage0_5[258], stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[118],stage1_7[119],stage1_6[123],stage1_5[192]}
   );
   gpc606_5 gpc279 (
      {stage0_5[264], stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[119],stage1_7[120],stage1_6[124],stage1_5[193]}
   );
   gpc606_5 gpc280 (
      {stage0_5[270], stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[120],stage1_7[121],stage1_6[125],stage1_5[194]}
   );
   gpc606_5 gpc281 (
      {stage0_5[276], stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[121],stage1_7[122],stage1_6[126],stage1_5[195]}
   );
   gpc606_5 gpc282 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[122],stage1_7[123],stage1_6[127],stage1_5[196]}
   );
   gpc606_5 gpc283 (
      {stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[123],stage1_7[124],stage1_6[128],stage1_5[197]}
   );
   gpc606_5 gpc284 (
      {stage0_5[294], stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[124],stage1_7[125],stage1_6[129],stage1_5[198]}
   );
   gpc606_5 gpc285 (
      {stage0_5[300], stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[125],stage1_7[126],stage1_6[130],stage1_5[199]}
   );
   gpc606_5 gpc286 (
      {stage0_5[306], stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[126],stage1_7[127],stage1_6[131],stage1_5[200]}
   );
   gpc606_5 gpc287 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317]},
      {stage0_7[300], stage0_7[301], stage0_7[302], stage0_7[303], stage0_7[304], stage0_7[305]},
      {stage1_9[50],stage1_8[127],stage1_7[128],stage1_6[132],stage1_5[201]}
   );
   gpc606_5 gpc288 (
      {stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323]},
      {stage0_7[306], stage0_7[307], stage0_7[308], stage0_7[309], stage0_7[310], stage0_7[311]},
      {stage1_9[51],stage1_8[128],stage1_7[129],stage1_6[133],stage1_5[202]}
   );
   gpc606_5 gpc289 (
      {stage0_5[324], stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329]},
      {stage0_7[312], stage0_7[313], stage0_7[314], stage0_7[315], stage0_7[316], stage0_7[317]},
      {stage1_9[52],stage1_8[129],stage1_7[130],stage1_6[134],stage1_5[203]}
   );
   gpc606_5 gpc290 (
      {stage0_5[330], stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335]},
      {stage0_7[318], stage0_7[319], stage0_7[320], stage0_7[321], stage0_7[322], stage0_7[323]},
      {stage1_9[53],stage1_8[130],stage1_7[131],stage1_6[135],stage1_5[204]}
   );
   gpc606_5 gpc291 (
      {stage0_5[336], stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341]},
      {stage0_7[324], stage0_7[325], stage0_7[326], stage0_7[327], stage0_7[328], stage0_7[329]},
      {stage1_9[54],stage1_8[131],stage1_7[132],stage1_6[136],stage1_5[205]}
   );
   gpc606_5 gpc292 (
      {stage0_5[342], stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347]},
      {stage0_7[330], stage0_7[331], stage0_7[332], stage0_7[333], stage0_7[334], stage0_7[335]},
      {stage1_9[55],stage1_8[132],stage1_7[133],stage1_6[137],stage1_5[206]}
   );
   gpc606_5 gpc293 (
      {stage0_5[348], stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353]},
      {stage0_7[336], stage0_7[337], stage0_7[338], stage0_7[339], stage0_7[340], stage0_7[341]},
      {stage1_9[56],stage1_8[133],stage1_7[134],stage1_6[138],stage1_5[207]}
   );
   gpc606_5 gpc294 (
      {stage0_5[354], stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359]},
      {stage0_7[342], stage0_7[343], stage0_7[344], stage0_7[345], stage0_7[346], stage0_7[347]},
      {stage1_9[57],stage1_8[134],stage1_7[135],stage1_6[139],stage1_5[208]}
   );
   gpc606_5 gpc295 (
      {stage0_5[360], stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365]},
      {stage0_7[348], stage0_7[349], stage0_7[350], stage0_7[351], stage0_7[352], stage0_7[353]},
      {stage1_9[58],stage1_8[135],stage1_7[136],stage1_6[140],stage1_5[209]}
   );
   gpc606_5 gpc296 (
      {stage0_5[366], stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371]},
      {stage0_7[354], stage0_7[355], stage0_7[356], stage0_7[357], stage0_7[358], stage0_7[359]},
      {stage1_9[59],stage1_8[136],stage1_7[137],stage1_6[141],stage1_5[210]}
   );
   gpc606_5 gpc297 (
      {stage0_5[372], stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377]},
      {stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364], stage0_7[365]},
      {stage1_9[60],stage1_8[137],stage1_7[138],stage1_6[142],stage1_5[211]}
   );
   gpc606_5 gpc298 (
      {stage0_5[378], stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383]},
      {stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370], stage0_7[371]},
      {stage1_9[61],stage1_8[138],stage1_7[139],stage1_6[143],stage1_5[212]}
   );
   gpc606_5 gpc299 (
      {stage0_5[384], stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389]},
      {stage0_7[372], stage0_7[373], stage0_7[374], stage0_7[375], stage0_7[376], stage0_7[377]},
      {stage1_9[62],stage1_8[139],stage1_7[140],stage1_6[144],stage1_5[213]}
   );
   gpc606_5 gpc300 (
      {stage0_5[390], stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395]},
      {stage0_7[378], stage0_7[379], stage0_7[380], stage0_7[381], stage0_7[382], stage0_7[383]},
      {stage1_9[63],stage1_8[140],stage1_7[141],stage1_6[145],stage1_5[214]}
   );
   gpc606_5 gpc301 (
      {stage0_5[396], stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401]},
      {stage0_7[384], stage0_7[385], stage0_7[386], stage0_7[387], stage0_7[388], stage0_7[389]},
      {stage1_9[64],stage1_8[141],stage1_7[142],stage1_6[146],stage1_5[215]}
   );
   gpc606_5 gpc302 (
      {stage0_5[402], stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407]},
      {stage0_7[390], stage0_7[391], stage0_7[392], stage0_7[393], stage0_7[394], stage0_7[395]},
      {stage1_9[65],stage1_8[142],stage1_7[143],stage1_6[147],stage1_5[216]}
   );
   gpc606_5 gpc303 (
      {stage0_5[408], stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413]},
      {stage0_7[396], stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400], stage0_7[401]},
      {stage1_9[66],stage1_8[143],stage1_7[144],stage1_6[148],stage1_5[217]}
   );
   gpc606_5 gpc304 (
      {stage0_5[414], stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419]},
      {stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405], stage0_7[406], stage0_7[407]},
      {stage1_9[67],stage1_8[144],stage1_7[145],stage1_6[149],stage1_5[218]}
   );
   gpc606_5 gpc305 (
      {stage0_5[420], stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425]},
      {stage0_7[408], stage0_7[409], stage0_7[410], stage0_7[411], stage0_7[412], stage0_7[413]},
      {stage1_9[68],stage1_8[145],stage1_7[146],stage1_6[150],stage1_5[219]}
   );
   gpc606_5 gpc306 (
      {stage0_5[426], stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431]},
      {stage0_7[414], stage0_7[415], stage0_7[416], stage0_7[417], stage0_7[418], stage0_7[419]},
      {stage1_9[69],stage1_8[146],stage1_7[147],stage1_6[151],stage1_5[220]}
   );
   gpc606_5 gpc307 (
      {stage0_5[432], stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437]},
      {stage0_7[420], stage0_7[421], stage0_7[422], stage0_7[423], stage0_7[424], stage0_7[425]},
      {stage1_9[70],stage1_8[147],stage1_7[148],stage1_6[152],stage1_5[221]}
   );
   gpc606_5 gpc308 (
      {stage0_5[438], stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443]},
      {stage0_7[426], stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430], stage0_7[431]},
      {stage1_9[71],stage1_8[148],stage1_7[149],stage1_6[153],stage1_5[222]}
   );
   gpc606_5 gpc309 (
      {stage0_5[444], stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449]},
      {stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435], stage0_7[436], stage0_7[437]},
      {stage1_9[72],stage1_8[149],stage1_7[150],stage1_6[154],stage1_5[223]}
   );
   gpc606_5 gpc310 (
      {stage0_5[450], stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455]},
      {stage0_7[438], stage0_7[439], stage0_7[440], stage0_7[441], stage0_7[442], stage0_7[443]},
      {stage1_9[73],stage1_8[150],stage1_7[151],stage1_6[155],stage1_5[224]}
   );
   gpc606_5 gpc311 (
      {stage0_5[456], stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461]},
      {stage0_7[444], stage0_7[445], stage0_7[446], stage0_7[447], stage0_7[448], stage0_7[449]},
      {stage1_9[74],stage1_8[151],stage1_7[152],stage1_6[156],stage1_5[225]}
   );
   gpc606_5 gpc312 (
      {stage0_5[462], stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467]},
      {stage0_7[450], stage0_7[451], stage0_7[452], stage0_7[453], stage0_7[454], stage0_7[455]},
      {stage1_9[75],stage1_8[152],stage1_7[153],stage1_6[157],stage1_5[226]}
   );
   gpc606_5 gpc313 (
      {stage0_5[468], stage0_5[469], stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473]},
      {stage0_7[456], stage0_7[457], stage0_7[458], stage0_7[459], stage0_7[460], stage0_7[461]},
      {stage1_9[76],stage1_8[153],stage1_7[154],stage1_6[158],stage1_5[227]}
   );
   gpc606_5 gpc314 (
      {stage0_5[474], stage0_5[475], stage0_5[476], stage0_5[477], stage0_5[478], stage0_5[479]},
      {stage0_7[462], stage0_7[463], stage0_7[464], stage0_7[465], stage0_7[466], stage0_7[467]},
      {stage1_9[77],stage1_8[154],stage1_7[155],stage1_6[159],stage1_5[228]}
   );
   gpc606_5 gpc315 (
      {stage0_5[480], stage0_5[481], stage0_5[482], stage0_5[483], stage0_5[484], stage0_5[485]},
      {stage0_7[468], stage0_7[469], stage0_7[470], stage0_7[471], stage0_7[472], stage0_7[473]},
      {stage1_9[78],stage1_8[155],stage1_7[156],stage1_6[160],stage1_5[229]}
   );
   gpc606_5 gpc316 (
      {stage0_6[462], stage0_6[463], stage0_6[464], stage0_6[465], stage0_6[466], stage0_6[467]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[79],stage1_8[156],stage1_7[157],stage1_6[161]}
   );
   gpc606_5 gpc317 (
      {stage0_6[468], stage0_6[469], stage0_6[470], stage0_6[471], stage0_6[472], stage0_6[473]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[80],stage1_8[157],stage1_7[158],stage1_6[162]}
   );
   gpc606_5 gpc318 (
      {stage0_6[474], stage0_6[475], stage0_6[476], stage0_6[477], stage0_6[478], stage0_6[479]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[81],stage1_8[158],stage1_7[159],stage1_6[163]}
   );
   gpc606_5 gpc319 (
      {stage0_7[474], stage0_7[475], stage0_7[476], stage0_7[477], stage0_7[478], stage0_7[479]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[82],stage1_8[159],stage1_7[160]}
   );
   gpc606_5 gpc320 (
      {stage0_7[480], stage0_7[481], stage0_7[482], stage0_7[483], stage0_7[484], stage0_7[485]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[4],stage1_9[83],stage1_8[160],stage1_7[161]}
   );
   gpc606_5 gpc321 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[2],stage1_10[5],stage1_9[84],stage1_8[161]}
   );
   gpc606_5 gpc322 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[3],stage1_10[6],stage1_9[85],stage1_8[162]}
   );
   gpc606_5 gpc323 (
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[4],stage1_10[7],stage1_9[86],stage1_8[163]}
   );
   gpc606_5 gpc324 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[5],stage1_10[8],stage1_9[87],stage1_8[164]}
   );
   gpc606_5 gpc325 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[6],stage1_10[9],stage1_9[88],stage1_8[165]}
   );
   gpc606_5 gpc326 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[7],stage1_10[10],stage1_9[89],stage1_8[166]}
   );
   gpc606_5 gpc327 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[8],stage1_10[11],stage1_9[90],stage1_8[167]}
   );
   gpc606_5 gpc328 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[9],stage1_10[12],stage1_9[91],stage1_8[168]}
   );
   gpc606_5 gpc329 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[10],stage1_10[13],stage1_9[92],stage1_8[169]}
   );
   gpc606_5 gpc330 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[11],stage1_10[14],stage1_9[93],stage1_8[170]}
   );
   gpc606_5 gpc331 (
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[12],stage1_10[15],stage1_9[94],stage1_8[171]}
   );
   gpc606_5 gpc332 (
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[13],stage1_10[16],stage1_9[95],stage1_8[172]}
   );
   gpc606_5 gpc333 (
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[14],stage1_10[17],stage1_9[96],stage1_8[173]}
   );
   gpc606_5 gpc334 (
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[15],stage1_10[18],stage1_9[97],stage1_8[174]}
   );
   gpc606_5 gpc335 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[16],stage1_10[19],stage1_9[98],stage1_8[175]}
   );
   gpc606_5 gpc336 (
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[17],stage1_10[20],stage1_9[99],stage1_8[176]}
   );
   gpc606_5 gpc337 (
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[18],stage1_10[21],stage1_9[100],stage1_8[177]}
   );
   gpc606_5 gpc338 (
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[19],stage1_10[22],stage1_9[101],stage1_8[178]}
   );
   gpc606_5 gpc339 (
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[20],stage1_10[23],stage1_9[102],stage1_8[179]}
   );
   gpc606_5 gpc340 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[21],stage1_10[24],stage1_9[103],stage1_8[180]}
   );
   gpc606_5 gpc341 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[22],stage1_10[25],stage1_9[104],stage1_8[181]}
   );
   gpc606_5 gpc342 (
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[23],stage1_10[26],stage1_9[105],stage1_8[182]}
   );
   gpc606_5 gpc343 (
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[24],stage1_10[27],stage1_9[106],stage1_8[183]}
   );
   gpc606_5 gpc344 (
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[25],stage1_10[28],stage1_9[107],stage1_8[184]}
   );
   gpc606_5 gpc345 (
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[26],stage1_10[29],stage1_9[108],stage1_8[185]}
   );
   gpc606_5 gpc346 (
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[27],stage1_10[30],stage1_9[109],stage1_8[186]}
   );
   gpc606_5 gpc347 (
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[28],stage1_10[31],stage1_9[110],stage1_8[187]}
   );
   gpc606_5 gpc348 (
      {stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[29],stage1_10[32],stage1_9[111],stage1_8[188]}
   );
   gpc606_5 gpc349 (
      {stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[30],stage1_10[33],stage1_9[112],stage1_8[189]}
   );
   gpc606_5 gpc350 (
      {stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[31],stage1_10[34],stage1_9[113],stage1_8[190]}
   );
   gpc606_5 gpc351 (
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[32],stage1_10[35],stage1_9[114],stage1_8[191]}
   );
   gpc606_5 gpc352 (
      {stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[33],stage1_10[36],stage1_9[115],stage1_8[192]}
   );
   gpc606_5 gpc353 (
      {stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[34],stage1_10[37],stage1_9[116],stage1_8[193]}
   );
   gpc606_5 gpc354 (
      {stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[35],stage1_10[38],stage1_9[117],stage1_8[194]}
   );
   gpc606_5 gpc355 (
      {stage0_8[222], stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[36],stage1_10[39],stage1_9[118],stage1_8[195]}
   );
   gpc606_5 gpc356 (
      {stage0_8[228], stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[37],stage1_10[40],stage1_9[119],stage1_8[196]}
   );
   gpc606_5 gpc357 (
      {stage0_8[234], stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[38],stage1_10[41],stage1_9[120],stage1_8[197]}
   );
   gpc606_5 gpc358 (
      {stage0_8[240], stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[39],stage1_10[42],stage1_9[121],stage1_8[198]}
   );
   gpc606_5 gpc359 (
      {stage0_8[246], stage0_8[247], stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[40],stage1_10[43],stage1_9[122],stage1_8[199]}
   );
   gpc606_5 gpc360 (
      {stage0_8[252], stage0_8[253], stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[41],stage1_10[44],stage1_9[123],stage1_8[200]}
   );
   gpc606_5 gpc361 (
      {stage0_8[258], stage0_8[259], stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[42],stage1_10[45],stage1_9[124],stage1_8[201]}
   );
   gpc606_5 gpc362 (
      {stage0_8[264], stage0_8[265], stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[43],stage1_10[46],stage1_9[125],stage1_8[202]}
   );
   gpc606_5 gpc363 (
      {stage0_8[270], stage0_8[271], stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[44],stage1_10[47],stage1_9[126],stage1_8[203]}
   );
   gpc606_5 gpc364 (
      {stage0_8[276], stage0_8[277], stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[45],stage1_10[48],stage1_9[127],stage1_8[204]}
   );
   gpc606_5 gpc365 (
      {stage0_8[282], stage0_8[283], stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[46],stage1_10[49],stage1_9[128],stage1_8[205]}
   );
   gpc606_5 gpc366 (
      {stage0_8[288], stage0_8[289], stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[47],stage1_10[50],stage1_9[129],stage1_8[206]}
   );
   gpc606_5 gpc367 (
      {stage0_8[294], stage0_8[295], stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[48],stage1_10[51],stage1_9[130],stage1_8[207]}
   );
   gpc606_5 gpc368 (
      {stage0_8[300], stage0_8[301], stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[49],stage1_10[52],stage1_9[131],stage1_8[208]}
   );
   gpc606_5 gpc369 (
      {stage0_8[306], stage0_8[307], stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[50],stage1_10[53],stage1_9[132],stage1_8[209]}
   );
   gpc606_5 gpc370 (
      {stage0_8[312], stage0_8[313], stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317]},
      {stage0_10[294], stage0_10[295], stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299]},
      {stage1_12[49],stage1_11[51],stage1_10[54],stage1_9[133],stage1_8[210]}
   );
   gpc606_5 gpc371 (
      {stage0_8[318], stage0_8[319], stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323]},
      {stage0_10[300], stage0_10[301], stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305]},
      {stage1_12[50],stage1_11[52],stage1_10[55],stage1_9[134],stage1_8[211]}
   );
   gpc606_5 gpc372 (
      {stage0_8[324], stage0_8[325], stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329]},
      {stage0_10[306], stage0_10[307], stage0_10[308], stage0_10[309], stage0_10[310], stage0_10[311]},
      {stage1_12[51],stage1_11[53],stage1_10[56],stage1_9[135],stage1_8[212]}
   );
   gpc606_5 gpc373 (
      {stage0_8[330], stage0_8[331], stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335]},
      {stage0_10[312], stage0_10[313], stage0_10[314], stage0_10[315], stage0_10[316], stage0_10[317]},
      {stage1_12[52],stage1_11[54],stage1_10[57],stage1_9[136],stage1_8[213]}
   );
   gpc606_5 gpc374 (
      {stage0_8[336], stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341]},
      {stage0_10[318], stage0_10[319], stage0_10[320], stage0_10[321], stage0_10[322], stage0_10[323]},
      {stage1_12[53],stage1_11[55],stage1_10[58],stage1_9[137],stage1_8[214]}
   );
   gpc606_5 gpc375 (
      {stage0_8[342], stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347]},
      {stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327], stage0_10[328], stage0_10[329]},
      {stage1_12[54],stage1_11[56],stage1_10[59],stage1_9[138],stage1_8[215]}
   );
   gpc606_5 gpc376 (
      {stage0_8[348], stage0_8[349], stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353]},
      {stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333], stage0_10[334], stage0_10[335]},
      {stage1_12[55],stage1_11[57],stage1_10[60],stage1_9[139],stage1_8[216]}
   );
   gpc606_5 gpc377 (
      {stage0_8[354], stage0_8[355], stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359]},
      {stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339], stage0_10[340], stage0_10[341]},
      {stage1_12[56],stage1_11[58],stage1_10[61],stage1_9[140],stage1_8[217]}
   );
   gpc606_5 gpc378 (
      {stage0_8[360], stage0_8[361], stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365]},
      {stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345], stage0_10[346], stage0_10[347]},
      {stage1_12[57],stage1_11[59],stage1_10[62],stage1_9[141],stage1_8[218]}
   );
   gpc606_5 gpc379 (
      {stage0_8[366], stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371]},
      {stage0_10[348], stage0_10[349], stage0_10[350], stage0_10[351], stage0_10[352], stage0_10[353]},
      {stage1_12[58],stage1_11[60],stage1_10[63],stage1_9[142],stage1_8[219]}
   );
   gpc606_5 gpc380 (
      {stage0_8[372], stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377]},
      {stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357], stage0_10[358], stage0_10[359]},
      {stage1_12[59],stage1_11[61],stage1_10[64],stage1_9[143],stage1_8[220]}
   );
   gpc606_5 gpc381 (
      {stage0_8[378], stage0_8[379], stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383]},
      {stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363], stage0_10[364], stage0_10[365]},
      {stage1_12[60],stage1_11[62],stage1_10[65],stage1_9[144],stage1_8[221]}
   );
   gpc606_5 gpc382 (
      {stage0_8[384], stage0_8[385], stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389]},
      {stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369], stage0_10[370], stage0_10[371]},
      {stage1_12[61],stage1_11[63],stage1_10[66],stage1_9[145],stage1_8[222]}
   );
   gpc606_5 gpc383 (
      {stage0_8[390], stage0_8[391], stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395]},
      {stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375], stage0_10[376], stage0_10[377]},
      {stage1_12[62],stage1_11[64],stage1_10[67],stage1_9[146],stage1_8[223]}
   );
   gpc606_5 gpc384 (
      {stage0_8[396], stage0_8[397], stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401]},
      {stage0_10[378], stage0_10[379], stage0_10[380], stage0_10[381], stage0_10[382], stage0_10[383]},
      {stage1_12[63],stage1_11[65],stage1_10[68],stage1_9[147],stage1_8[224]}
   );
   gpc606_5 gpc385 (
      {stage0_8[402], stage0_8[403], stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407]},
      {stage0_10[384], stage0_10[385], stage0_10[386], stage0_10[387], stage0_10[388], stage0_10[389]},
      {stage1_12[64],stage1_11[66],stage1_10[69],stage1_9[148],stage1_8[225]}
   );
   gpc606_5 gpc386 (
      {stage0_8[408], stage0_8[409], stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413]},
      {stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393], stage0_10[394], stage0_10[395]},
      {stage1_12[65],stage1_11[67],stage1_10[70],stage1_9[149],stage1_8[226]}
   );
   gpc606_5 gpc387 (
      {stage0_8[414], stage0_8[415], stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419]},
      {stage0_10[396], stage0_10[397], stage0_10[398], stage0_10[399], stage0_10[400], stage0_10[401]},
      {stage1_12[66],stage1_11[68],stage1_10[71],stage1_9[150],stage1_8[227]}
   );
   gpc606_5 gpc388 (
      {stage0_8[420], stage0_8[421], stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425]},
      {stage0_10[402], stage0_10[403], stage0_10[404], stage0_10[405], stage0_10[406], stage0_10[407]},
      {stage1_12[67],stage1_11[69],stage1_10[72],stage1_9[151],stage1_8[228]}
   );
   gpc606_5 gpc389 (
      {stage0_8[426], stage0_8[427], stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431]},
      {stage0_10[408], stage0_10[409], stage0_10[410], stage0_10[411], stage0_10[412], stage0_10[413]},
      {stage1_12[68],stage1_11[70],stage1_10[73],stage1_9[152],stage1_8[229]}
   );
   gpc606_5 gpc390 (
      {stage0_8[432], stage0_8[433], stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437]},
      {stage0_10[414], stage0_10[415], stage0_10[416], stage0_10[417], stage0_10[418], stage0_10[419]},
      {stage1_12[69],stage1_11[71],stage1_10[74],stage1_9[153],stage1_8[230]}
   );
   gpc606_5 gpc391 (
      {stage0_8[438], stage0_8[439], stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443]},
      {stage0_10[420], stage0_10[421], stage0_10[422], stage0_10[423], stage0_10[424], stage0_10[425]},
      {stage1_12[70],stage1_11[72],stage1_10[75],stage1_9[154],stage1_8[231]}
   );
   gpc606_5 gpc392 (
      {stage0_8[444], stage0_8[445], stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449]},
      {stage0_10[426], stage0_10[427], stage0_10[428], stage0_10[429], stage0_10[430], stage0_10[431]},
      {stage1_12[71],stage1_11[73],stage1_10[76],stage1_9[155],stage1_8[232]}
   );
   gpc606_5 gpc393 (
      {stage0_8[450], stage0_8[451], stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455]},
      {stage0_10[432], stage0_10[433], stage0_10[434], stage0_10[435], stage0_10[436], stage0_10[437]},
      {stage1_12[72],stage1_11[74],stage1_10[77],stage1_9[156],stage1_8[233]}
   );
   gpc606_5 gpc394 (
      {stage0_8[456], stage0_8[457], stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461]},
      {stage0_10[438], stage0_10[439], stage0_10[440], stage0_10[441], stage0_10[442], stage0_10[443]},
      {stage1_12[73],stage1_11[75],stage1_10[78],stage1_9[157],stage1_8[234]}
   );
   gpc606_5 gpc395 (
      {stage0_8[462], stage0_8[463], stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467]},
      {stage0_10[444], stage0_10[445], stage0_10[446], stage0_10[447], stage0_10[448], stage0_10[449]},
      {stage1_12[74],stage1_11[76],stage1_10[79],stage1_9[158],stage1_8[235]}
   );
   gpc606_5 gpc396 (
      {stage0_8[468], stage0_8[469], stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473]},
      {stage0_10[450], stage0_10[451], stage0_10[452], stage0_10[453], stage0_10[454], stage0_10[455]},
      {stage1_12[75],stage1_11[77],stage1_10[80],stage1_9[159],stage1_8[236]}
   );
   gpc606_5 gpc397 (
      {stage0_8[474], stage0_8[475], stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479]},
      {stage0_10[456], stage0_10[457], stage0_10[458], stage0_10[459], stage0_10[460], stage0_10[461]},
      {stage1_12[76],stage1_11[78],stage1_10[81],stage1_9[160],stage1_8[237]}
   );
   gpc606_5 gpc398 (
      {stage0_8[480], stage0_8[481], stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485]},
      {stage0_10[462], stage0_10[463], stage0_10[464], stage0_10[465], stage0_10[466], stage0_10[467]},
      {stage1_12[77],stage1_11[79],stage1_10[82],stage1_9[161],stage1_8[238]}
   );
   gpc606_5 gpc399 (
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[78],stage1_11[80],stage1_10[83],stage1_9[162]}
   );
   gpc606_5 gpc400 (
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[79],stage1_11[81],stage1_10[84],stage1_9[163]}
   );
   gpc606_5 gpc401 (
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[80],stage1_11[82],stage1_10[85],stage1_9[164]}
   );
   gpc606_5 gpc402 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[81],stage1_11[83],stage1_10[86],stage1_9[165]}
   );
   gpc606_5 gpc403 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[82],stage1_11[84],stage1_10[87],stage1_9[166]}
   );
   gpc606_5 gpc404 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[83],stage1_11[85],stage1_10[88],stage1_9[167]}
   );
   gpc606_5 gpc405 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[84],stage1_11[86],stage1_10[89],stage1_9[168]}
   );
   gpc606_5 gpc406 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[85],stage1_11[87],stage1_10[90],stage1_9[169]}
   );
   gpc606_5 gpc407 (
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[86],stage1_11[88],stage1_10[91],stage1_9[170]}
   );
   gpc606_5 gpc408 (
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[87],stage1_11[89],stage1_10[92],stage1_9[171]}
   );
   gpc606_5 gpc409 (
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[88],stage1_11[90],stage1_10[93],stage1_9[172]}
   );
   gpc606_5 gpc410 (
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[89],stage1_11[91],stage1_10[94],stage1_9[173]}
   );
   gpc606_5 gpc411 (
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[90],stage1_11[92],stage1_10[95],stage1_9[174]}
   );
   gpc606_5 gpc412 (
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[91],stage1_11[93],stage1_10[96],stage1_9[175]}
   );
   gpc606_5 gpc413 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[92],stage1_11[94],stage1_10[97],stage1_9[176]}
   );
   gpc606_5 gpc414 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[93],stage1_11[95],stage1_10[98],stage1_9[177]}
   );
   gpc606_5 gpc415 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[94],stage1_11[96],stage1_10[99],stage1_9[178]}
   );
   gpc606_5 gpc416 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[95],stage1_11[97],stage1_10[100],stage1_9[179]}
   );
   gpc606_5 gpc417 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[96],stage1_11[98],stage1_10[101],stage1_9[180]}
   );
   gpc606_5 gpc418 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[97],stage1_11[99],stage1_10[102],stage1_9[181]}
   );
   gpc606_5 gpc419 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[98],stage1_11[100],stage1_10[103],stage1_9[182]}
   );
   gpc606_5 gpc420 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[99],stage1_11[101],stage1_10[104],stage1_9[183]}
   );
   gpc606_5 gpc421 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[100],stage1_11[102],stage1_10[105],stage1_9[184]}
   );
   gpc606_5 gpc422 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[101],stage1_11[103],stage1_10[106],stage1_9[185]}
   );
   gpc606_5 gpc423 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[102],stage1_11[104],stage1_10[107],stage1_9[186]}
   );
   gpc606_5 gpc424 (
      {stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[103],stage1_11[105],stage1_10[108],stage1_9[187]}
   );
   gpc606_5 gpc425 (
      {stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[104],stage1_11[106],stage1_10[109],stage1_9[188]}
   );
   gpc606_5 gpc426 (
      {stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[105],stage1_11[107],stage1_10[110],stage1_9[189]}
   );
   gpc606_5 gpc427 (
      {stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[106],stage1_11[108],stage1_10[111],stage1_9[190]}
   );
   gpc606_5 gpc428 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[107],stage1_11[109],stage1_10[112],stage1_9[191]}
   );
   gpc606_5 gpc429 (
      {stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[108],stage1_11[110],stage1_10[113],stage1_9[192]}
   );
   gpc606_5 gpc430 (
      {stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[109],stage1_11[111],stage1_10[114],stage1_9[193]}
   );
   gpc606_5 gpc431 (
      {stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[110],stage1_11[112],stage1_10[115],stage1_9[194]}
   );
   gpc606_5 gpc432 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[111],stage1_11[113],stage1_10[116],stage1_9[195]}
   );
   gpc606_5 gpc433 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220], stage0_9[221]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[112],stage1_11[114],stage1_10[117],stage1_9[196]}
   );
   gpc606_5 gpc434 (
      {stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225], stage0_9[226], stage0_9[227]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[113],stage1_11[115],stage1_10[118],stage1_9[197]}
   );
   gpc606_5 gpc435 (
      {stage0_9[228], stage0_9[229], stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[114],stage1_11[116],stage1_10[119],stage1_9[198]}
   );
   gpc606_5 gpc436 (
      {stage0_9[234], stage0_9[235], stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[115],stage1_11[117],stage1_10[120],stage1_9[199]}
   );
   gpc606_5 gpc437 (
      {stage0_9[240], stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[116],stage1_11[118],stage1_10[121],stage1_9[200]}
   );
   gpc606_5 gpc438 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250], stage0_9[251]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[117],stage1_11[119],stage1_10[122],stage1_9[201]}
   );
   gpc606_5 gpc439 (
      {stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255], stage0_9[256], stage0_9[257]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[118],stage1_11[120],stage1_10[123],stage1_9[202]}
   );
   gpc606_5 gpc440 (
      {stage0_9[258], stage0_9[259], stage0_9[260], stage0_9[261], stage0_9[262], stage0_9[263]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[119],stage1_11[121],stage1_10[124],stage1_9[203]}
   );
   gpc606_5 gpc441 (
      {stage0_9[264], stage0_9[265], stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[120],stage1_11[122],stage1_10[125],stage1_9[204]}
   );
   gpc606_5 gpc442 (
      {stage0_9[270], stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[121],stage1_11[123],stage1_10[126],stage1_9[205]}
   );
   gpc606_5 gpc443 (
      {stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280], stage0_9[281]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[122],stage1_11[124],stage1_10[127],stage1_9[206]}
   );
   gpc606_5 gpc444 (
      {stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285], stage0_9[286], stage0_9[287]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[123],stage1_11[125],stage1_10[128],stage1_9[207]}
   );
   gpc606_5 gpc445 (
      {stage0_9[288], stage0_9[289], stage0_9[290], stage0_9[291], stage0_9[292], stage0_9[293]},
      {stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage1_13[46],stage1_12[124],stage1_11[126],stage1_10[129],stage1_9[208]}
   );
   gpc606_5 gpc446 (
      {stage0_9[294], stage0_9[295], stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299]},
      {stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage1_13[47],stage1_12[125],stage1_11[127],stage1_10[130],stage1_9[209]}
   );
   gpc606_5 gpc447 (
      {stage0_9[300], stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305]},
      {stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293]},
      {stage1_13[48],stage1_12[126],stage1_11[128],stage1_10[131],stage1_9[210]}
   );
   gpc606_5 gpc448 (
      {stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310], stage0_9[311]},
      {stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage1_13[49],stage1_12[127],stage1_11[129],stage1_10[132],stage1_9[211]}
   );
   gpc606_5 gpc449 (
      {stage0_9[312], stage0_9[313], stage0_9[314], stage0_9[315], stage0_9[316], stage0_9[317]},
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305]},
      {stage1_13[50],stage1_12[128],stage1_11[130],stage1_10[133],stage1_9[212]}
   );
   gpc606_5 gpc450 (
      {stage0_9[318], stage0_9[319], stage0_9[320], stage0_9[321], stage0_9[322], stage0_9[323]},
      {stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage1_13[51],stage1_12[129],stage1_11[131],stage1_10[134],stage1_9[213]}
   );
   gpc606_5 gpc451 (
      {stage0_9[324], stage0_9[325], stage0_9[326], stage0_9[327], stage0_9[328], stage0_9[329]},
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316], stage0_11[317]},
      {stage1_13[52],stage1_12[130],stage1_11[132],stage1_10[135],stage1_9[214]}
   );
   gpc606_5 gpc452 (
      {stage0_9[330], stage0_9[331], stage0_9[332], stage0_9[333], stage0_9[334], stage0_9[335]},
      {stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323]},
      {stage1_13[53],stage1_12[131],stage1_11[133],stage1_10[136],stage1_9[215]}
   );
   gpc606_5 gpc453 (
      {stage0_9[336], stage0_9[337], stage0_9[338], stage0_9[339], stage0_9[340], stage0_9[341]},
      {stage0_11[324], stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage1_13[54],stage1_12[132],stage1_11[134],stage1_10[137],stage1_9[216]}
   );
   gpc606_5 gpc454 (
      {stage0_9[342], stage0_9[343], stage0_9[344], stage0_9[345], stage0_9[346], stage0_9[347]},
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage1_13[55],stage1_12[133],stage1_11[135],stage1_10[138],stage1_9[217]}
   );
   gpc606_5 gpc455 (
      {stage0_9[348], stage0_9[349], stage0_9[350], stage0_9[351], stage0_9[352], stage0_9[353]},
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage1_13[56],stage1_12[134],stage1_11[136],stage1_10[139],stage1_9[218]}
   );
   gpc606_5 gpc456 (
      {stage0_9[354], stage0_9[355], stage0_9[356], stage0_9[357], stage0_9[358], stage0_9[359]},
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346], stage0_11[347]},
      {stage1_13[57],stage1_12[135],stage1_11[137],stage1_10[140],stage1_9[219]}
   );
   gpc606_5 gpc457 (
      {stage0_9[360], stage0_9[361], stage0_9[362], stage0_9[363], stage0_9[364], stage0_9[365]},
      {stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353]},
      {stage1_13[58],stage1_12[136],stage1_11[138],stage1_10[141],stage1_9[220]}
   );
   gpc606_5 gpc458 (
      {stage0_9[366], stage0_9[367], stage0_9[368], stage0_9[369], stage0_9[370], stage0_9[371]},
      {stage0_11[354], stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage1_13[59],stage1_12[137],stage1_11[139],stage1_10[142],stage1_9[221]}
   );
   gpc606_5 gpc459 (
      {stage0_9[372], stage0_9[373], stage0_9[374], stage0_9[375], stage0_9[376], stage0_9[377]},
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage1_13[60],stage1_12[138],stage1_11[140],stage1_10[143],stage1_9[222]}
   );
   gpc606_5 gpc460 (
      {stage0_9[378], stage0_9[379], stage0_9[380], stage0_9[381], stage0_9[382], stage0_9[383]},
      {stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369], stage0_11[370], stage0_11[371]},
      {stage1_13[61],stage1_12[139],stage1_11[141],stage1_10[144],stage1_9[223]}
   );
   gpc606_5 gpc461 (
      {stage0_9[384], stage0_9[385], stage0_9[386], stage0_9[387], stage0_9[388], stage0_9[389]},
      {stage0_11[372], stage0_11[373], stage0_11[374], stage0_11[375], stage0_11[376], stage0_11[377]},
      {stage1_13[62],stage1_12[140],stage1_11[142],stage1_10[145],stage1_9[224]}
   );
   gpc606_5 gpc462 (
      {stage0_9[390], stage0_9[391], stage0_9[392], stage0_9[393], stage0_9[394], stage0_9[395]},
      {stage0_11[378], stage0_11[379], stage0_11[380], stage0_11[381], stage0_11[382], stage0_11[383]},
      {stage1_13[63],stage1_12[141],stage1_11[143],stage1_10[146],stage1_9[225]}
   );
   gpc606_5 gpc463 (
      {stage0_9[396], stage0_9[397], stage0_9[398], stage0_9[399], stage0_9[400], stage0_9[401]},
      {stage0_11[384], stage0_11[385], stage0_11[386], stage0_11[387], stage0_11[388], stage0_11[389]},
      {stage1_13[64],stage1_12[142],stage1_11[144],stage1_10[147],stage1_9[226]}
   );
   gpc606_5 gpc464 (
      {stage0_9[402], stage0_9[403], stage0_9[404], stage0_9[405], stage0_9[406], stage0_9[407]},
      {stage0_11[390], stage0_11[391], stage0_11[392], stage0_11[393], stage0_11[394], stage0_11[395]},
      {stage1_13[65],stage1_12[143],stage1_11[145],stage1_10[148],stage1_9[227]}
   );
   gpc606_5 gpc465 (
      {stage0_9[408], stage0_9[409], stage0_9[410], stage0_9[411], stage0_9[412], stage0_9[413]},
      {stage0_11[396], stage0_11[397], stage0_11[398], stage0_11[399], stage0_11[400], stage0_11[401]},
      {stage1_13[66],stage1_12[144],stage1_11[146],stage1_10[149],stage1_9[228]}
   );
   gpc606_5 gpc466 (
      {stage0_9[414], stage0_9[415], stage0_9[416], stage0_9[417], stage0_9[418], stage0_9[419]},
      {stage0_11[402], stage0_11[403], stage0_11[404], stage0_11[405], stage0_11[406], stage0_11[407]},
      {stage1_13[67],stage1_12[145],stage1_11[147],stage1_10[150],stage1_9[229]}
   );
   gpc606_5 gpc467 (
      {stage0_9[420], stage0_9[421], stage0_9[422], stage0_9[423], stage0_9[424], stage0_9[425]},
      {stage0_11[408], stage0_11[409], stage0_11[410], stage0_11[411], stage0_11[412], stage0_11[413]},
      {stage1_13[68],stage1_12[146],stage1_11[148],stage1_10[151],stage1_9[230]}
   );
   gpc606_5 gpc468 (
      {stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429], stage0_9[430], stage0_9[431]},
      {stage0_11[414], stage0_11[415], stage0_11[416], stage0_11[417], stage0_11[418], stage0_11[419]},
      {stage1_13[69],stage1_12[147],stage1_11[149],stage1_10[152],stage1_9[231]}
   );
   gpc606_5 gpc469 (
      {stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435], stage0_9[436], stage0_9[437]},
      {stage0_11[420], stage0_11[421], stage0_11[422], stage0_11[423], stage0_11[424], stage0_11[425]},
      {stage1_13[70],stage1_12[148],stage1_11[150],stage1_10[153],stage1_9[232]}
   );
   gpc606_5 gpc470 (
      {stage0_9[438], stage0_9[439], stage0_9[440], stage0_9[441], stage0_9[442], stage0_9[443]},
      {stage0_11[426], stage0_11[427], stage0_11[428], stage0_11[429], stage0_11[430], stage0_11[431]},
      {stage1_13[71],stage1_12[149],stage1_11[151],stage1_10[154],stage1_9[233]}
   );
   gpc606_5 gpc471 (
      {stage0_9[444], stage0_9[445], stage0_9[446], stage0_9[447], stage0_9[448], stage0_9[449]},
      {stage0_11[432], stage0_11[433], stage0_11[434], stage0_11[435], stage0_11[436], stage0_11[437]},
      {stage1_13[72],stage1_12[150],stage1_11[152],stage1_10[155],stage1_9[234]}
   );
   gpc606_5 gpc472 (
      {stage0_9[450], stage0_9[451], stage0_9[452], stage0_9[453], stage0_9[454], stage0_9[455]},
      {stage0_11[438], stage0_11[439], stage0_11[440], stage0_11[441], stage0_11[442], stage0_11[443]},
      {stage1_13[73],stage1_12[151],stage1_11[153],stage1_10[156],stage1_9[235]}
   );
   gpc606_5 gpc473 (
      {stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459], stage0_9[460], stage0_9[461]},
      {stage0_11[444], stage0_11[445], stage0_11[446], stage0_11[447], stage0_11[448], stage0_11[449]},
      {stage1_13[74],stage1_12[152],stage1_11[154],stage1_10[157],stage1_9[236]}
   );
   gpc606_5 gpc474 (
      {stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465], stage0_9[466], stage0_9[467]},
      {stage0_11[450], stage0_11[451], stage0_11[452], stage0_11[453], stage0_11[454], stage0_11[455]},
      {stage1_13[75],stage1_12[153],stage1_11[155],stage1_10[158],stage1_9[237]}
   );
   gpc606_5 gpc475 (
      {stage0_9[468], stage0_9[469], stage0_9[470], stage0_9[471], stage0_9[472], stage0_9[473]},
      {stage0_11[456], stage0_11[457], stage0_11[458], stage0_11[459], stage0_11[460], stage0_11[461]},
      {stage1_13[76],stage1_12[154],stage1_11[156],stage1_10[159],stage1_9[238]}
   );
   gpc606_5 gpc476 (
      {stage0_9[474], stage0_9[475], stage0_9[476], stage0_9[477], stage0_9[478], stage0_9[479]},
      {stage0_11[462], stage0_11[463], stage0_11[464], stage0_11[465], stage0_11[466], stage0_11[467]},
      {stage1_13[77],stage1_12[155],stage1_11[157],stage1_10[160],stage1_9[239]}
   );
   gpc606_5 gpc477 (
      {stage0_9[480], stage0_9[481], stage0_9[482], stage0_9[483], stage0_9[484], stage0_9[485]},
      {stage0_11[468], stage0_11[469], stage0_11[470], stage0_11[471], stage0_11[472], stage0_11[473]},
      {stage1_13[78],stage1_12[156],stage1_11[158],stage1_10[161],stage1_9[240]}
   );
   gpc1_1 gpc478 (
      {stage0_2[447]},
      {stage1_2[159]}
   );
   gpc1_1 gpc479 (
      {stage0_2[448]},
      {stage1_2[160]}
   );
   gpc1_1 gpc480 (
      {stage0_2[449]},
      {stage1_2[161]}
   );
   gpc1_1 gpc481 (
      {stage0_2[450]},
      {stage1_2[162]}
   );
   gpc1_1 gpc482 (
      {stage0_2[451]},
      {stage1_2[163]}
   );
   gpc1_1 gpc483 (
      {stage0_2[452]},
      {stage1_2[164]}
   );
   gpc1_1 gpc484 (
      {stage0_2[453]},
      {stage1_2[165]}
   );
   gpc1_1 gpc485 (
      {stage0_2[454]},
      {stage1_2[166]}
   );
   gpc1_1 gpc486 (
      {stage0_2[455]},
      {stage1_2[167]}
   );
   gpc1_1 gpc487 (
      {stage0_2[456]},
      {stage1_2[168]}
   );
   gpc1_1 gpc488 (
      {stage0_2[457]},
      {stage1_2[169]}
   );
   gpc1_1 gpc489 (
      {stage0_2[458]},
      {stage1_2[170]}
   );
   gpc1_1 gpc490 (
      {stage0_2[459]},
      {stage1_2[171]}
   );
   gpc1_1 gpc491 (
      {stage0_2[460]},
      {stage1_2[172]}
   );
   gpc1_1 gpc492 (
      {stage0_2[461]},
      {stage1_2[173]}
   );
   gpc1_1 gpc493 (
      {stage0_2[462]},
      {stage1_2[174]}
   );
   gpc1_1 gpc494 (
      {stage0_2[463]},
      {stage1_2[175]}
   );
   gpc1_1 gpc495 (
      {stage0_2[464]},
      {stage1_2[176]}
   );
   gpc1_1 gpc496 (
      {stage0_2[465]},
      {stage1_2[177]}
   );
   gpc1_1 gpc497 (
      {stage0_2[466]},
      {stage1_2[178]}
   );
   gpc1_1 gpc498 (
      {stage0_2[467]},
      {stage1_2[179]}
   );
   gpc1_1 gpc499 (
      {stage0_2[468]},
      {stage1_2[180]}
   );
   gpc1_1 gpc500 (
      {stage0_2[469]},
      {stage1_2[181]}
   );
   gpc1_1 gpc501 (
      {stage0_2[470]},
      {stage1_2[182]}
   );
   gpc1_1 gpc502 (
      {stage0_2[471]},
      {stage1_2[183]}
   );
   gpc1_1 gpc503 (
      {stage0_2[472]},
      {stage1_2[184]}
   );
   gpc1_1 gpc504 (
      {stage0_2[473]},
      {stage1_2[185]}
   );
   gpc1_1 gpc505 (
      {stage0_2[474]},
      {stage1_2[186]}
   );
   gpc1_1 gpc506 (
      {stage0_2[475]},
      {stage1_2[187]}
   );
   gpc1_1 gpc507 (
      {stage0_2[476]},
      {stage1_2[188]}
   );
   gpc1_1 gpc508 (
      {stage0_2[477]},
      {stage1_2[189]}
   );
   gpc1_1 gpc509 (
      {stage0_2[478]},
      {stage1_2[190]}
   );
   gpc1_1 gpc510 (
      {stage0_2[479]},
      {stage1_2[191]}
   );
   gpc1_1 gpc511 (
      {stage0_2[480]},
      {stage1_2[192]}
   );
   gpc1_1 gpc512 (
      {stage0_2[481]},
      {stage1_2[193]}
   );
   gpc1_1 gpc513 (
      {stage0_2[482]},
      {stage1_2[194]}
   );
   gpc1_1 gpc514 (
      {stage0_2[483]},
      {stage1_2[195]}
   );
   gpc1_1 gpc515 (
      {stage0_2[484]},
      {stage1_2[196]}
   );
   gpc1_1 gpc516 (
      {stage0_2[485]},
      {stage1_2[197]}
   );
   gpc1_1 gpc517 (
      {stage0_3[450]},
      {stage1_3[160]}
   );
   gpc1_1 gpc518 (
      {stage0_3[451]},
      {stage1_3[161]}
   );
   gpc1_1 gpc519 (
      {stage0_3[452]},
      {stage1_3[162]}
   );
   gpc1_1 gpc520 (
      {stage0_3[453]},
      {stage1_3[163]}
   );
   gpc1_1 gpc521 (
      {stage0_3[454]},
      {stage1_3[164]}
   );
   gpc1_1 gpc522 (
      {stage0_3[455]},
      {stage1_3[165]}
   );
   gpc1_1 gpc523 (
      {stage0_3[456]},
      {stage1_3[166]}
   );
   gpc1_1 gpc524 (
      {stage0_3[457]},
      {stage1_3[167]}
   );
   gpc1_1 gpc525 (
      {stage0_3[458]},
      {stage1_3[168]}
   );
   gpc1_1 gpc526 (
      {stage0_3[459]},
      {stage1_3[169]}
   );
   gpc1_1 gpc527 (
      {stage0_3[460]},
      {stage1_3[170]}
   );
   gpc1_1 gpc528 (
      {stage0_3[461]},
      {stage1_3[171]}
   );
   gpc1_1 gpc529 (
      {stage0_3[462]},
      {stage1_3[172]}
   );
   gpc1_1 gpc530 (
      {stage0_3[463]},
      {stage1_3[173]}
   );
   gpc1_1 gpc531 (
      {stage0_3[464]},
      {stage1_3[174]}
   );
   gpc1_1 gpc532 (
      {stage0_3[465]},
      {stage1_3[175]}
   );
   gpc1_1 gpc533 (
      {stage0_3[466]},
      {stage1_3[176]}
   );
   gpc1_1 gpc534 (
      {stage0_3[467]},
      {stage1_3[177]}
   );
   gpc1_1 gpc535 (
      {stage0_3[468]},
      {stage1_3[178]}
   );
   gpc1_1 gpc536 (
      {stage0_3[469]},
      {stage1_3[179]}
   );
   gpc1_1 gpc537 (
      {stage0_3[470]},
      {stage1_3[180]}
   );
   gpc1_1 gpc538 (
      {stage0_3[471]},
      {stage1_3[181]}
   );
   gpc1_1 gpc539 (
      {stage0_3[472]},
      {stage1_3[182]}
   );
   gpc1_1 gpc540 (
      {stage0_3[473]},
      {stage1_3[183]}
   );
   gpc1_1 gpc541 (
      {stage0_3[474]},
      {stage1_3[184]}
   );
   gpc1_1 gpc542 (
      {stage0_3[475]},
      {stage1_3[185]}
   );
   gpc1_1 gpc543 (
      {stage0_3[476]},
      {stage1_3[186]}
   );
   gpc1_1 gpc544 (
      {stage0_3[477]},
      {stage1_3[187]}
   );
   gpc1_1 gpc545 (
      {stage0_3[478]},
      {stage1_3[188]}
   );
   gpc1_1 gpc546 (
      {stage0_3[479]},
      {stage1_3[189]}
   );
   gpc1_1 gpc547 (
      {stage0_3[480]},
      {stage1_3[190]}
   );
   gpc1_1 gpc548 (
      {stage0_3[481]},
      {stage1_3[191]}
   );
   gpc1_1 gpc549 (
      {stage0_3[482]},
      {stage1_3[192]}
   );
   gpc1_1 gpc550 (
      {stage0_3[483]},
      {stage1_3[193]}
   );
   gpc1_1 gpc551 (
      {stage0_3[484]},
      {stage1_3[194]}
   );
   gpc1_1 gpc552 (
      {stage0_3[485]},
      {stage1_3[195]}
   );
   gpc1_1 gpc553 (
      {stage0_4[481]},
      {stage1_4[236]}
   );
   gpc1_1 gpc554 (
      {stage0_4[482]},
      {stage1_4[237]}
   );
   gpc1_1 gpc555 (
      {stage0_4[483]},
      {stage1_4[238]}
   );
   gpc1_1 gpc556 (
      {stage0_4[484]},
      {stage1_4[239]}
   );
   gpc1_1 gpc557 (
      {stage0_4[485]},
      {stage1_4[240]}
   );
   gpc1_1 gpc558 (
      {stage0_6[480]},
      {stage1_6[164]}
   );
   gpc1_1 gpc559 (
      {stage0_6[481]},
      {stage1_6[165]}
   );
   gpc1_1 gpc560 (
      {stage0_6[482]},
      {stage1_6[166]}
   );
   gpc1_1 gpc561 (
      {stage0_6[483]},
      {stage1_6[167]}
   );
   gpc1_1 gpc562 (
      {stage0_6[484]},
      {stage1_6[168]}
   );
   gpc1_1 gpc563 (
      {stage0_6[485]},
      {stage1_6[169]}
   );
   gpc1_1 gpc564 (
      {stage0_10[468]},
      {stage1_10[162]}
   );
   gpc1_1 gpc565 (
      {stage0_10[469]},
      {stage1_10[163]}
   );
   gpc1_1 gpc566 (
      {stage0_10[470]},
      {stage1_10[164]}
   );
   gpc1_1 gpc567 (
      {stage0_10[471]},
      {stage1_10[165]}
   );
   gpc1_1 gpc568 (
      {stage0_10[472]},
      {stage1_10[166]}
   );
   gpc1_1 gpc569 (
      {stage0_10[473]},
      {stage1_10[167]}
   );
   gpc1_1 gpc570 (
      {stage0_10[474]},
      {stage1_10[168]}
   );
   gpc1_1 gpc571 (
      {stage0_10[475]},
      {stage1_10[169]}
   );
   gpc1_1 gpc572 (
      {stage0_10[476]},
      {stage1_10[170]}
   );
   gpc1_1 gpc573 (
      {stage0_10[477]},
      {stage1_10[171]}
   );
   gpc1_1 gpc574 (
      {stage0_10[478]},
      {stage1_10[172]}
   );
   gpc1_1 gpc575 (
      {stage0_10[479]},
      {stage1_10[173]}
   );
   gpc1_1 gpc576 (
      {stage0_10[480]},
      {stage1_10[174]}
   );
   gpc1_1 gpc577 (
      {stage0_10[481]},
      {stage1_10[175]}
   );
   gpc1_1 gpc578 (
      {stage0_10[482]},
      {stage1_10[176]}
   );
   gpc1_1 gpc579 (
      {stage0_10[483]},
      {stage1_10[177]}
   );
   gpc1_1 gpc580 (
      {stage0_10[484]},
      {stage1_10[178]}
   );
   gpc1_1 gpc581 (
      {stage0_10[485]},
      {stage1_10[179]}
   );
   gpc1_1 gpc582 (
      {stage0_11[474]},
      {stage1_11[159]}
   );
   gpc1_1 gpc583 (
      {stage0_11[475]},
      {stage1_11[160]}
   );
   gpc1_1 gpc584 (
      {stage0_11[476]},
      {stage1_11[161]}
   );
   gpc1_1 gpc585 (
      {stage0_11[477]},
      {stage1_11[162]}
   );
   gpc1_1 gpc586 (
      {stage0_11[478]},
      {stage1_11[163]}
   );
   gpc1_1 gpc587 (
      {stage0_11[479]},
      {stage1_11[164]}
   );
   gpc1_1 gpc588 (
      {stage0_11[480]},
      {stage1_11[165]}
   );
   gpc1_1 gpc589 (
      {stage0_11[481]},
      {stage1_11[166]}
   );
   gpc1_1 gpc590 (
      {stage0_11[482]},
      {stage1_11[167]}
   );
   gpc1_1 gpc591 (
      {stage0_11[483]},
      {stage1_11[168]}
   );
   gpc1_1 gpc592 (
      {stage0_11[484]},
      {stage1_11[169]}
   );
   gpc1_1 gpc593 (
      {stage0_11[485]},
      {stage1_11[170]}
   );
   gpc1163_5 gpc594 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc595 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc596 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc597 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc598 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc599 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc600 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc601 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc602 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc603 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc604 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc605 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc1163_5 gpc606 (
      {stage1_0[36], stage1_0[37], stage1_0[38]},
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_2[12]},
      {stage1_3[12]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc1163_5 gpc607 (
      {stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_2[13]},
      {stage1_3[13]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc1163_5 gpc608 (
      {stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_2[14]},
      {stage1_3[14]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc1163_5 gpc609 (
      {stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_2[15]},
      {stage1_3[15]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc1163_5 gpc610 (
      {stage1_0[48], stage1_0[49], stage1_0[50]},
      {stage1_1[96], stage1_1[97], stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101]},
      {stage1_2[16]},
      {stage1_3[16]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc1163_5 gpc611 (
      {stage1_0[51], stage1_0[52], stage1_0[53]},
      {stage1_1[102], stage1_1[103], stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107]},
      {stage1_2[17]},
      {stage1_3[17]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc1163_5 gpc612 (
      {stage1_0[54], stage1_0[55], stage1_0[56]},
      {stage1_1[108], stage1_1[109], stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113]},
      {stage1_2[18]},
      {stage1_3[18]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc1163_5 gpc613 (
      {stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_1[114], stage1_1[115], stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119]},
      {stage1_2[19]},
      {stage1_3[19]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc606_5 gpc614 (
      {stage1_0[60], stage1_0[61], stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65]},
      {stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc615 (
      {stage1_0[66], stage1_0[67], stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71]},
      {stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc606_5 gpc616 (
      {stage1_0[72], stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37]},
      {stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22],stage2_0[22]}
   );
   gpc606_5 gpc617 (
      {stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[23],stage2_3[23],stage2_2[23]}
   );
   gpc606_5 gpc618 (
      {stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[24],stage2_3[24],stage2_2[24]}
   );
   gpc606_5 gpc619 (
      {stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[25],stage2_3[25],stage2_2[25]}
   );
   gpc606_5 gpc620 (
      {stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59], stage1_2[60], stage1_2[61]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[26],stage2_3[26],stage2_2[26]}
   );
   gpc606_5 gpc621 (
      {stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65], stage1_2[66], stage1_2[67]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[4],stage2_4[27],stage2_3[27],stage2_2[27]}
   );
   gpc615_5 gpc622 (
      {stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71], stage1_2[72]},
      {stage1_3[20]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[5],stage2_4[28],stage2_3[28],stage2_2[28]}
   );
   gpc615_5 gpc623 (
      {stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77]},
      {stage1_3[21]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[6],stage2_4[29],stage2_3[29],stage2_2[29]}
   );
   gpc615_5 gpc624 (
      {stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82]},
      {stage1_3[22]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[7],stage2_4[30],stage2_3[30],stage2_2[30]}
   );
   gpc615_5 gpc625 (
      {stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87]},
      {stage1_3[23]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[8],stage2_4[31],stage2_3[31],stage2_2[31]}
   );
   gpc615_5 gpc626 (
      {stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91], stage1_2[92]},
      {stage1_3[24]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[9],stage2_4[32],stage2_3[32],stage2_2[32]}
   );
   gpc615_5 gpc627 (
      {stage1_2[93], stage1_2[94], stage1_2[95], stage1_2[96], stage1_2[97]},
      {stage1_3[25]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[10],stage2_4[33],stage2_3[33],stage2_2[33]}
   );
   gpc615_5 gpc628 (
      {stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101], stage1_2[102]},
      {stage1_3[26]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[11],stage2_4[34],stage2_3[34],stage2_2[34]}
   );
   gpc615_5 gpc629 (
      {stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106], stage1_2[107]},
      {stage1_3[27]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[12],stage2_4[35],stage2_3[35],stage2_2[35]}
   );
   gpc615_5 gpc630 (
      {stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111], stage1_2[112]},
      {stage1_3[28]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[13],stage2_4[36],stage2_3[36],stage2_2[36]}
   );
   gpc615_5 gpc631 (
      {stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117]},
      {stage1_3[29]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[14],stage2_4[37],stage2_3[37],stage2_2[37]}
   );
   gpc615_5 gpc632 (
      {stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121], stage1_2[122]},
      {stage1_3[30]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[15],stage2_4[38],stage2_3[38],stage2_2[38]}
   );
   gpc615_5 gpc633 (
      {stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126], stage1_2[127]},
      {stage1_3[31]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[16],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc615_5 gpc634 (
      {stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131], stage1_2[132]},
      {stage1_3[32]},
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage2_6[17],stage2_5[17],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc615_5 gpc635 (
      {stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137]},
      {stage1_3[33]},
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113]},
      {stage2_6[18],stage2_5[18],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc615_5 gpc636 (
      {stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142]},
      {stage1_3[34]},
      {stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119]},
      {stage2_6[19],stage2_5[19],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc615_5 gpc637 (
      {stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146], stage1_2[147]},
      {stage1_3[35]},
      {stage1_4[120], stage1_4[121], stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125]},
      {stage2_6[20],stage2_5[20],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc638 (
      {stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151], stage1_2[152]},
      {stage1_3[36]},
      {stage1_4[126], stage1_4[127], stage1_4[128], stage1_4[129], stage1_4[130], stage1_4[131]},
      {stage2_6[21],stage2_5[21],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc615_5 gpc639 (
      {stage1_2[153], stage1_2[154], stage1_2[155], stage1_2[156], stage1_2[157]},
      {stage1_3[37]},
      {stage1_4[132], stage1_4[133], stage1_4[134], stage1_4[135], stage1_4[136], stage1_4[137]},
      {stage2_6[22],stage2_5[22],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc615_5 gpc640 (
      {stage1_2[158], stage1_2[159], stage1_2[160], stage1_2[161], stage1_2[162]},
      {stage1_3[38]},
      {stage1_4[138], stage1_4[139], stage1_4[140], stage1_4[141], stage1_4[142], stage1_4[143]},
      {stage2_6[23],stage2_5[23],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc615_5 gpc641 (
      {stage1_2[163], stage1_2[164], stage1_2[165], stage1_2[166], stage1_2[167]},
      {stage1_3[39]},
      {stage1_4[144], stage1_4[145], stage1_4[146], stage1_4[147], stage1_4[148], stage1_4[149]},
      {stage2_6[24],stage2_5[24],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc615_5 gpc642 (
      {stage1_2[168], stage1_2[169], stage1_2[170], stage1_2[171], stage1_2[172]},
      {stage1_3[40]},
      {stage1_4[150], stage1_4[151], stage1_4[152], stage1_4[153], stage1_4[154], stage1_4[155]},
      {stage2_6[25],stage2_5[25],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc615_5 gpc643 (
      {stage1_2[173], stage1_2[174], stage1_2[175], stage1_2[176], stage1_2[177]},
      {stage1_3[41]},
      {stage1_4[156], stage1_4[157], stage1_4[158], stage1_4[159], stage1_4[160], stage1_4[161]},
      {stage2_6[26],stage2_5[26],stage2_4[49],stage2_3[49],stage2_2[49]}
   );
   gpc615_5 gpc644 (
      {stage1_2[178], stage1_2[179], stage1_2[180], stage1_2[181], stage1_2[182]},
      {stage1_3[42]},
      {stage1_4[162], stage1_4[163], stage1_4[164], stage1_4[165], stage1_4[166], stage1_4[167]},
      {stage2_6[27],stage2_5[27],stage2_4[50],stage2_3[50],stage2_2[50]}
   );
   gpc615_5 gpc645 (
      {stage1_2[183], stage1_2[184], stage1_2[185], stage1_2[186], stage1_2[187]},
      {stage1_3[43]},
      {stage1_4[168], stage1_4[169], stage1_4[170], stage1_4[171], stage1_4[172], stage1_4[173]},
      {stage2_6[28],stage2_5[28],stage2_4[51],stage2_3[51],stage2_2[51]}
   );
   gpc615_5 gpc646 (
      {stage1_2[188], stage1_2[189], stage1_2[190], stage1_2[191], stage1_2[192]},
      {stage1_3[44]},
      {stage1_4[174], stage1_4[175], stage1_4[176], stage1_4[177], stage1_4[178], stage1_4[179]},
      {stage2_6[29],stage2_5[29],stage2_4[52],stage2_3[52],stage2_2[52]}
   );
   gpc615_5 gpc647 (
      {stage1_2[193], stage1_2[194], stage1_2[195], stage1_2[196], stage1_2[197]},
      {stage1_3[45]},
      {stage1_4[180], stage1_4[181], stage1_4[182], stage1_4[183], stage1_4[184], stage1_4[185]},
      {stage2_6[30],stage2_5[30],stage2_4[53],stage2_3[53],stage2_2[53]}
   );
   gpc615_5 gpc648 (
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50]},
      {stage1_4[186]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[31],stage2_5[31],stage2_4[54],stage2_3[54]}
   );
   gpc615_5 gpc649 (
      {stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55]},
      {stage1_4[187]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[32],stage2_5[32],stage2_4[55],stage2_3[55]}
   );
   gpc615_5 gpc650 (
      {stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60]},
      {stage1_4[188]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[33],stage2_5[33],stage2_4[56],stage2_3[56]}
   );
   gpc615_5 gpc651 (
      {stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage1_4[189]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[34],stage2_5[34],stage2_4[57],stage2_3[57]}
   );
   gpc615_5 gpc652 (
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70]},
      {stage1_4[190]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[35],stage2_5[35],stage2_4[58],stage2_3[58]}
   );
   gpc615_5 gpc653 (
      {stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75]},
      {stage1_4[191]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[36],stage2_5[36],stage2_4[59],stage2_3[59]}
   );
   gpc615_5 gpc654 (
      {stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80]},
      {stage1_4[192]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[37],stage2_5[37],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc655 (
      {stage1_3[81], stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85]},
      {stage1_4[193]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[38],stage2_5[38],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc656 (
      {stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90]},
      {stage1_4[194]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[39],stage2_5[39],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc657 (
      {stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage1_4[195]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[40],stage2_5[40],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc658 (
      {stage1_3[96], stage1_3[97], stage1_3[98], stage1_3[99], stage1_3[100]},
      {stage1_4[196]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[41],stage2_5[41],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc659 (
      {stage1_3[101], stage1_3[102], stage1_3[103], stage1_3[104], stage1_3[105]},
      {stage1_4[197]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[42],stage2_5[42],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc660 (
      {stage1_3[106], stage1_3[107], stage1_3[108], stage1_3[109], stage1_3[110]},
      {stage1_4[198]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[43],stage2_5[43],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc661 (
      {stage1_3[111], stage1_3[112], stage1_3[113], stage1_3[114], stage1_3[115]},
      {stage1_4[199]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[44],stage2_5[44],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc662 (
      {stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119], stage1_3[120]},
      {stage1_4[200]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[45],stage2_5[45],stage2_4[68],stage2_3[68]}
   );
   gpc615_5 gpc663 (
      {stage1_3[121], stage1_3[122], stage1_3[123], stage1_3[124], stage1_3[125]},
      {stage1_4[201]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[46],stage2_5[46],stage2_4[69],stage2_3[69]}
   );
   gpc615_5 gpc664 (
      {stage1_3[126], stage1_3[127], stage1_3[128], stage1_3[129], stage1_3[130]},
      {stage1_4[202]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[47],stage2_5[47],stage2_4[70],stage2_3[70]}
   );
   gpc615_5 gpc665 (
      {stage1_3[131], stage1_3[132], stage1_3[133], stage1_3[134], stage1_3[135]},
      {stage1_4[203]},
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage2_7[17],stage2_6[48],stage2_5[48],stage2_4[71],stage2_3[71]}
   );
   gpc615_5 gpc666 (
      {stage1_3[136], stage1_3[137], stage1_3[138], stage1_3[139], stage1_3[140]},
      {stage1_4[204]},
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage2_7[18],stage2_6[49],stage2_5[49],stage2_4[72],stage2_3[72]}
   );
   gpc615_5 gpc667 (
      {stage1_3[141], stage1_3[142], stage1_3[143], stage1_3[144], stage1_3[145]},
      {stage1_4[205]},
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage2_7[19],stage2_6[50],stage2_5[50],stage2_4[73],stage2_3[73]}
   );
   gpc615_5 gpc668 (
      {stage1_3[146], stage1_3[147], stage1_3[148], stage1_3[149], stage1_3[150]},
      {stage1_4[206]},
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage2_7[20],stage2_6[51],stage2_5[51],stage2_4[74],stage2_3[74]}
   );
   gpc615_5 gpc669 (
      {stage1_3[151], stage1_3[152], stage1_3[153], stage1_3[154], stage1_3[155]},
      {stage1_4[207]},
      {stage1_5[126], stage1_5[127], stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131]},
      {stage2_7[21],stage2_6[52],stage2_5[52],stage2_4[75],stage2_3[75]}
   );
   gpc615_5 gpc670 (
      {stage1_3[156], stage1_3[157], stage1_3[158], stage1_3[159], stage1_3[160]},
      {stage1_4[208]},
      {stage1_5[132], stage1_5[133], stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137]},
      {stage2_7[22],stage2_6[53],stage2_5[53],stage2_4[76],stage2_3[76]}
   );
   gpc615_5 gpc671 (
      {stage1_3[161], stage1_3[162], stage1_3[163], stage1_3[164], stage1_3[165]},
      {stage1_4[209]},
      {stage1_5[138], stage1_5[139], stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143]},
      {stage2_7[23],stage2_6[54],stage2_5[54],stage2_4[77],stage2_3[77]}
   );
   gpc615_5 gpc672 (
      {stage1_3[166], stage1_3[167], stage1_3[168], stage1_3[169], stage1_3[170]},
      {stage1_4[210]},
      {stage1_5[144], stage1_5[145], stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149]},
      {stage2_7[24],stage2_6[55],stage2_5[55],stage2_4[78],stage2_3[78]}
   );
   gpc615_5 gpc673 (
      {stage1_3[171], stage1_3[172], stage1_3[173], stage1_3[174], stage1_3[175]},
      {stage1_4[211]},
      {stage1_5[150], stage1_5[151], stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155]},
      {stage2_7[25],stage2_6[56],stage2_5[56],stage2_4[79],stage2_3[79]}
   );
   gpc615_5 gpc674 (
      {stage1_3[176], stage1_3[177], stage1_3[178], stage1_3[179], stage1_3[180]},
      {stage1_4[212]},
      {stage1_5[156], stage1_5[157], stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161]},
      {stage2_7[26],stage2_6[57],stage2_5[57],stage2_4[80],stage2_3[80]}
   );
   gpc615_5 gpc675 (
      {stage1_3[181], stage1_3[182], stage1_3[183], stage1_3[184], stage1_3[185]},
      {stage1_4[213]},
      {stage1_5[162], stage1_5[163], stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167]},
      {stage2_7[27],stage2_6[58],stage2_5[58],stage2_4[81],stage2_3[81]}
   );
   gpc615_5 gpc676 (
      {stage1_3[186], stage1_3[187], stage1_3[188], stage1_3[189], stage1_3[190]},
      {stage1_4[214]},
      {stage1_5[168], stage1_5[169], stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173]},
      {stage2_7[28],stage2_6[59],stage2_5[59],stage2_4[82],stage2_3[82]}
   );
   gpc615_5 gpc677 (
      {stage1_3[191], stage1_3[192], stage1_3[193], stage1_3[194], stage1_3[195]},
      {stage1_4[215]},
      {stage1_5[174], stage1_5[175], stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179]},
      {stage2_7[29],stage2_6[60],stage2_5[60],stage2_4[83],stage2_3[83]}
   );
   gpc606_5 gpc678 (
      {stage1_4[216], stage1_4[217], stage1_4[218], stage1_4[219], stage1_4[220], stage1_4[221]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[30],stage2_6[61],stage2_5[61],stage2_4[84]}
   );
   gpc606_5 gpc679 (
      {stage1_4[222], stage1_4[223], stage1_4[224], stage1_4[225], stage1_4[226], stage1_4[227]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[31],stage2_6[62],stage2_5[62],stage2_4[85]}
   );
   gpc606_5 gpc680 (
      {stage1_4[228], stage1_4[229], stage1_4[230], stage1_4[231], stage1_4[232], stage1_4[233]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[32],stage2_6[63],stage2_5[63],stage2_4[86]}
   );
   gpc606_5 gpc681 (
      {stage1_4[234], stage1_4[235], stage1_4[236], stage1_4[237], stage1_4[238], stage1_4[239]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[33],stage2_6[64],stage2_5[64],stage2_4[87]}
   );
   gpc606_5 gpc682 (
      {stage1_5[180], stage1_5[181], stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[4],stage2_7[34],stage2_6[65],stage2_5[65]}
   );
   gpc606_5 gpc683 (
      {stage1_5[186], stage1_5[187], stage1_5[188], stage1_5[189], stage1_5[190], stage1_5[191]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[5],stage2_7[35],stage2_6[66],stage2_5[66]}
   );
   gpc606_5 gpc684 (
      {stage1_5[192], stage1_5[193], stage1_5[194], stage1_5[195], stage1_5[196], stage1_5[197]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[6],stage2_7[36],stage2_6[67],stage2_5[67]}
   );
   gpc606_5 gpc685 (
      {stage1_5[198], stage1_5[199], stage1_5[200], stage1_5[201], stage1_5[202], stage1_5[203]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[7],stage2_7[37],stage2_6[68],stage2_5[68]}
   );
   gpc606_5 gpc686 (
      {stage1_5[204], stage1_5[205], stage1_5[206], stage1_5[207], stage1_5[208], stage1_5[209]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[8],stage2_7[38],stage2_6[69],stage2_5[69]}
   );
   gpc606_5 gpc687 (
      {stage1_5[210], stage1_5[211], stage1_5[212], stage1_5[213], stage1_5[214], stage1_5[215]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[9],stage2_7[39],stage2_6[70],stage2_5[70]}
   );
   gpc606_5 gpc688 (
      {stage1_5[216], stage1_5[217], stage1_5[218], stage1_5[219], stage1_5[220], stage1_5[221]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[10],stage2_7[40],stage2_6[71],stage2_5[71]}
   );
   gpc606_5 gpc689 (
      {stage1_5[222], stage1_5[223], stage1_5[224], stage1_5[225], stage1_5[226], stage1_5[227]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[11],stage2_7[41],stage2_6[72],stage2_5[72]}
   );
   gpc606_5 gpc690 (
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[8],stage2_8[12],stage2_7[42],stage2_6[73]}
   );
   gpc606_5 gpc691 (
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[9],stage2_8[13],stage2_7[43],stage2_6[74]}
   );
   gpc606_5 gpc692 (
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[10],stage2_8[14],stage2_7[44],stage2_6[75]}
   );
   gpc606_5 gpc693 (
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[11],stage2_8[15],stage2_7[45],stage2_6[76]}
   );
   gpc606_5 gpc694 (
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[12],stage2_8[16],stage2_7[46],stage2_6[77]}
   );
   gpc606_5 gpc695 (
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[13],stage2_8[17],stage2_7[47],stage2_6[78]}
   );
   gpc606_5 gpc696 (
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[14],stage2_8[18],stage2_7[48],stage2_6[79]}
   );
   gpc606_5 gpc697 (
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[15],stage2_8[19],stage2_7[49],stage2_6[80]}
   );
   gpc606_5 gpc698 (
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[16],stage2_8[20],stage2_7[50],stage2_6[81]}
   );
   gpc606_5 gpc699 (
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[17],stage2_8[21],stage2_7[51],stage2_6[82]}
   );
   gpc606_5 gpc700 (
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[18],stage2_8[22],stage2_7[52],stage2_6[83]}
   );
   gpc606_5 gpc701 (
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[19],stage2_8[23],stage2_7[53],stage2_6[84]}
   );
   gpc606_5 gpc702 (
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[20],stage2_8[24],stage2_7[54],stage2_6[85]}
   );
   gpc606_5 gpc703 (
      {stage1_6[102], stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[21],stage2_8[25],stage2_7[55],stage2_6[86]}
   );
   gpc606_5 gpc704 (
      {stage1_6[108], stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[22],stage2_8[26],stage2_7[56],stage2_6[87]}
   );
   gpc606_5 gpc705 (
      {stage1_6[114], stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[23],stage2_8[27],stage2_7[57],stage2_6[88]}
   );
   gpc606_5 gpc706 (
      {stage1_6[120], stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125]},
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage2_10[16],stage2_9[24],stage2_8[28],stage2_7[58],stage2_6[89]}
   );
   gpc606_5 gpc707 (
      {stage1_6[126], stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131]},
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage2_10[17],stage2_9[25],stage2_8[29],stage2_7[59],stage2_6[90]}
   );
   gpc606_5 gpc708 (
      {stage1_6[132], stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137]},
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage2_10[18],stage2_9[26],stage2_8[30],stage2_7[60],stage2_6[91]}
   );
   gpc606_5 gpc709 (
      {stage1_6[138], stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143]},
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage2_10[19],stage2_9[27],stage2_8[31],stage2_7[61],stage2_6[92]}
   );
   gpc606_5 gpc710 (
      {stage1_6[144], stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149]},
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage2_10[20],stage2_9[28],stage2_8[32],stage2_7[62],stage2_6[93]}
   );
   gpc615_5 gpc711 (
      {stage1_6[150], stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154]},
      {stage1_7[48]},
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage2_10[21],stage2_9[29],stage2_8[33],stage2_7[63],stage2_6[94]}
   );
   gpc615_5 gpc712 (
      {stage1_6[155], stage1_6[156], stage1_6[157], stage1_6[158], stage1_6[159]},
      {stage1_7[49]},
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage2_10[22],stage2_9[30],stage2_8[34],stage2_7[64],stage2_6[95]}
   );
   gpc615_5 gpc713 (
      {stage1_6[160], stage1_6[161], stage1_6[162], stage1_6[163], stage1_6[164]},
      {stage1_7[50]},
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage2_10[23],stage2_9[31],stage2_8[35],stage2_7[65],stage2_6[96]}
   );
   gpc615_5 gpc714 (
      {stage1_6[165], stage1_6[166], stage1_6[167], stage1_6[168], stage1_6[169]},
      {stage1_7[51]},
      {stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147], stage1_8[148], stage1_8[149]},
      {stage2_10[24],stage2_9[32],stage2_8[36],stage2_7[66],stage2_6[97]}
   );
   gpc615_5 gpc715 (
      {stage1_7[52], stage1_7[53], stage1_7[54], stage1_7[55], stage1_7[56]},
      {stage1_8[150]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[25],stage2_9[33],stage2_8[37],stage2_7[67]}
   );
   gpc615_5 gpc716 (
      {stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60], stage1_7[61]},
      {stage1_8[151]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[26],stage2_9[34],stage2_8[38],stage2_7[68]}
   );
   gpc615_5 gpc717 (
      {stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66]},
      {stage1_8[152]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[27],stage2_9[35],stage2_8[39],stage2_7[69]}
   );
   gpc615_5 gpc718 (
      {stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage1_8[153]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[28],stage2_9[36],stage2_8[40],stage2_7[70]}
   );
   gpc615_5 gpc719 (
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76]},
      {stage1_8[154]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[29],stage2_9[37],stage2_8[41],stage2_7[71]}
   );
   gpc615_5 gpc720 (
      {stage1_7[77], stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81]},
      {stage1_8[155]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[30],stage2_9[38],stage2_8[42],stage2_7[72]}
   );
   gpc615_5 gpc721 (
      {stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85], stage1_7[86]},
      {stage1_8[156]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[31],stage2_9[39],stage2_8[43],stage2_7[73]}
   );
   gpc615_5 gpc722 (
      {stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], stage1_7[91]},
      {stage1_8[157]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[32],stage2_9[40],stage2_8[44],stage2_7[74]}
   );
   gpc615_5 gpc723 (
      {stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95], stage1_7[96]},
      {stage1_8[158]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[33],stage2_9[41],stage2_8[45],stage2_7[75]}
   );
   gpc615_5 gpc724 (
      {stage1_7[97], stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101]},
      {stage1_8[159]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[34],stage2_9[42],stage2_8[46],stage2_7[76]}
   );
   gpc615_5 gpc725 (
      {stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105], stage1_7[106]},
      {stage1_8[160]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[35],stage2_9[43],stage2_8[47],stage2_7[77]}
   );
   gpc615_5 gpc726 (
      {stage1_7[107], stage1_7[108], stage1_7[109], stage1_7[110], stage1_7[111]},
      {stage1_8[161]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[36],stage2_9[44],stage2_8[48],stage2_7[78]}
   );
   gpc615_5 gpc727 (
      {stage1_7[112], stage1_7[113], stage1_7[114], stage1_7[115], stage1_7[116]},
      {stage1_8[162]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[37],stage2_9[45],stage2_8[49],stage2_7[79]}
   );
   gpc615_5 gpc728 (
      {stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120], stage1_7[121]},
      {stage1_8[163]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[38],stage2_9[46],stage2_8[50],stage2_7[80]}
   );
   gpc615_5 gpc729 (
      {stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125], stage1_7[126]},
      {stage1_8[164]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[39],stage2_9[47],stage2_8[51],stage2_7[81]}
   );
   gpc615_5 gpc730 (
      {stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130], stage1_7[131]},
      {stage1_8[165]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[40],stage2_9[48],stage2_8[52],stage2_7[82]}
   );
   gpc615_5 gpc731 (
      {stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135], stage1_7[136]},
      {stage1_8[166]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[41],stage2_9[49],stage2_8[53],stage2_7[83]}
   );
   gpc615_5 gpc732 (
      {stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140], stage1_7[141]},
      {stage1_8[167]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[42],stage2_9[50],stage2_8[54],stage2_7[84]}
   );
   gpc615_5 gpc733 (
      {stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145], stage1_7[146]},
      {stage1_8[168]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[43],stage2_9[51],stage2_8[55],stage2_7[85]}
   );
   gpc615_5 gpc734 (
      {stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150], stage1_7[151]},
      {stage1_8[169]},
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage2_11[19],stage2_10[44],stage2_9[52],stage2_8[56],stage2_7[86]}
   );
   gpc615_5 gpc735 (
      {stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155], stage1_7[156]},
      {stage1_8[170]},
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage2_11[20],stage2_10[45],stage2_9[53],stage2_8[57],stage2_7[87]}
   );
   gpc615_5 gpc736 (
      {stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160], stage1_7[161]},
      {stage1_8[171]},
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage2_11[21],stage2_10[46],stage2_9[54],stage2_8[58],stage2_7[88]}
   );
   gpc606_5 gpc737 (
      {stage1_8[172], stage1_8[173], stage1_8[174], stage1_8[175], stage1_8[176], stage1_8[177]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[22],stage2_10[47],stage2_9[55],stage2_8[59]}
   );
   gpc606_5 gpc738 (
      {stage1_8[178], stage1_8[179], stage1_8[180], stage1_8[181], stage1_8[182], stage1_8[183]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[23],stage2_10[48],stage2_9[56],stage2_8[60]}
   );
   gpc606_5 gpc739 (
      {stage1_8[184], stage1_8[185], stage1_8[186], stage1_8[187], stage1_8[188], stage1_8[189]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[24],stage2_10[49],stage2_9[57],stage2_8[61]}
   );
   gpc606_5 gpc740 (
      {stage1_8[190], stage1_8[191], stage1_8[192], stage1_8[193], stage1_8[194], stage1_8[195]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[25],stage2_10[50],stage2_9[58],stage2_8[62]}
   );
   gpc606_5 gpc741 (
      {stage1_8[196], stage1_8[197], stage1_8[198], stage1_8[199], stage1_8[200], stage1_8[201]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[26],stage2_10[51],stage2_9[59],stage2_8[63]}
   );
   gpc606_5 gpc742 (
      {stage1_8[202], stage1_8[203], stage1_8[204], stage1_8[205], stage1_8[206], stage1_8[207]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[27],stage2_10[52],stage2_9[60],stage2_8[64]}
   );
   gpc606_5 gpc743 (
      {stage1_8[208], stage1_8[209], stage1_8[210], stage1_8[211], stage1_8[212], stage1_8[213]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[28],stage2_10[53],stage2_9[61],stage2_8[65]}
   );
   gpc615_5 gpc744 (
      {stage1_8[214], stage1_8[215], stage1_8[216], stage1_8[217], stage1_8[218]},
      {stage1_9[132]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[29],stage2_10[54],stage2_9[62],stage2_8[66]}
   );
   gpc615_5 gpc745 (
      {stage1_8[219], stage1_8[220], stage1_8[221], stage1_8[222], stage1_8[223]},
      {stage1_9[133]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[30],stage2_10[55],stage2_9[63],stage2_8[67]}
   );
   gpc615_5 gpc746 (
      {stage1_8[224], stage1_8[225], stage1_8[226], stage1_8[227], stage1_8[228]},
      {stage1_9[134]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[31],stage2_10[56],stage2_9[64],stage2_8[68]}
   );
   gpc615_5 gpc747 (
      {stage1_8[229], stage1_8[230], stage1_8[231], stage1_8[232], stage1_8[233]},
      {stage1_9[135]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[32],stage2_10[57],stage2_9[65],stage2_8[69]}
   );
   gpc615_5 gpc748 (
      {stage1_8[234], stage1_8[235], stage1_8[236], stage1_8[237], stage1_8[238]},
      {stage1_9[136]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[33],stage2_10[58],stage2_9[66],stage2_8[70]}
   );
   gpc606_5 gpc749 (
      {stage1_9[137], stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[12],stage2_11[34],stage2_10[59],stage2_9[67]}
   );
   gpc606_5 gpc750 (
      {stage1_9[143], stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[13],stage2_11[35],stage2_10[60],stage2_9[68]}
   );
   gpc606_5 gpc751 (
      {stage1_9[149], stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[14],stage2_11[36],stage2_10[61],stage2_9[69]}
   );
   gpc606_5 gpc752 (
      {stage1_9[155], stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[15],stage2_11[37],stage2_10[62],stage2_9[70]}
   );
   gpc606_5 gpc753 (
      {stage1_9[161], stage1_9[162], stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[16],stage2_11[38],stage2_10[63],stage2_9[71]}
   );
   gpc606_5 gpc754 (
      {stage1_9[167], stage1_9[168], stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[17],stage2_11[39],stage2_10[64],stage2_9[72]}
   );
   gpc606_5 gpc755 (
      {stage1_9[173], stage1_9[174], stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[18],stage2_11[40],stage2_10[65],stage2_9[73]}
   );
   gpc615_5 gpc756 (
      {stage1_9[179], stage1_9[180], stage1_9[181], stage1_9[182], stage1_9[183]},
      {stage1_10[72]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[19],stage2_11[41],stage2_10[66],stage2_9[74]}
   );
   gpc615_5 gpc757 (
      {stage1_9[184], stage1_9[185], stage1_9[186], stage1_9[187], stage1_9[188]},
      {stage1_10[73]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[20],stage2_11[42],stage2_10[67],stage2_9[75]}
   );
   gpc615_5 gpc758 (
      {stage1_9[189], stage1_9[190], stage1_9[191], stage1_9[192], stage1_9[193]},
      {stage1_10[74]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[21],stage2_11[43],stage2_10[68],stage2_9[76]}
   );
   gpc615_5 gpc759 (
      {stage1_9[194], stage1_9[195], stage1_9[196], stage1_9[197], stage1_9[198]},
      {stage1_10[75]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[22],stage2_11[44],stage2_10[69],stage2_9[77]}
   );
   gpc615_5 gpc760 (
      {stage1_9[199], stage1_9[200], stage1_9[201], stage1_9[202], stage1_9[203]},
      {stage1_10[76]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[23],stage2_11[45],stage2_10[70],stage2_9[78]}
   );
   gpc615_5 gpc761 (
      {stage1_9[204], stage1_9[205], stage1_9[206], stage1_9[207], stage1_9[208]},
      {stage1_10[77]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[24],stage2_11[46],stage2_10[71],stage2_9[79]}
   );
   gpc615_5 gpc762 (
      {stage1_9[209], stage1_9[210], stage1_9[211], stage1_9[212], stage1_9[213]},
      {stage1_10[78]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[25],stage2_11[47],stage2_10[72],stage2_9[80]}
   );
   gpc615_5 gpc763 (
      {stage1_9[214], stage1_9[215], stage1_9[216], stage1_9[217], stage1_9[218]},
      {stage1_10[79]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[26],stage2_11[48],stage2_10[73],stage2_9[81]}
   );
   gpc615_5 gpc764 (
      {stage1_9[219], stage1_9[220], stage1_9[221], stage1_9[222], stage1_9[223]},
      {stage1_10[80]},
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95]},
      {stage2_13[15],stage2_12[27],stage2_11[49],stage2_10[74],stage2_9[82]}
   );
   gpc615_5 gpc765 (
      {stage1_9[224], stage1_9[225], stage1_9[226], stage1_9[227], stage1_9[228]},
      {stage1_10[81]},
      {stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage2_13[16],stage2_12[28],stage2_11[50],stage2_10[75],stage2_9[83]}
   );
   gpc615_5 gpc766 (
      {stage1_9[229], stage1_9[230], stage1_9[231], stage1_9[232], stage1_9[233]},
      {stage1_10[82]},
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107]},
      {stage2_13[17],stage2_12[29],stage2_11[51],stage2_10[76],stage2_9[84]}
   );
   gpc606_5 gpc767 (
      {stage1_10[83], stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[18],stage2_12[30],stage2_11[52],stage2_10[77]}
   );
   gpc606_5 gpc768 (
      {stage1_10[89], stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[19],stage2_12[31],stage2_11[53],stage2_10[78]}
   );
   gpc606_5 gpc769 (
      {stage1_10[95], stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[20],stage2_12[32],stage2_11[54],stage2_10[79]}
   );
   gpc606_5 gpc770 (
      {stage1_10[101], stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[21],stage2_12[33],stage2_11[55],stage2_10[80]}
   );
   gpc606_5 gpc771 (
      {stage1_10[107], stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[22],stage2_12[34],stage2_11[56],stage2_10[81]}
   );
   gpc606_5 gpc772 (
      {stage1_10[113], stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[23],stage2_12[35],stage2_11[57],stage2_10[82]}
   );
   gpc606_5 gpc773 (
      {stage1_10[119], stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[24],stage2_12[36],stage2_11[58],stage2_10[83]}
   );
   gpc606_5 gpc774 (
      {stage1_10[125], stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[25],stage2_12[37],stage2_11[59],stage2_10[84]}
   );
   gpc606_5 gpc775 (
      {stage1_10[131], stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[26],stage2_12[38],stage2_11[60],stage2_10[85]}
   );
   gpc606_5 gpc776 (
      {stage1_10[137], stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141], stage1_10[142]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[27],stage2_12[39],stage2_11[61],stage2_10[86]}
   );
   gpc606_5 gpc777 (
      {stage1_10[143], stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[28],stage2_12[40],stage2_11[62],stage2_10[87]}
   );
   gpc606_5 gpc778 (
      {stage1_10[149], stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[29],stage2_12[41],stage2_11[63],stage2_10[88]}
   );
   gpc606_5 gpc779 (
      {stage1_10[155], stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[30],stage2_12[42],stage2_11[64],stage2_10[89]}
   );
   gpc606_5 gpc780 (
      {stage1_10[161], stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[31],stage2_12[43],stage2_11[65],stage2_10[90]}
   );
   gpc606_5 gpc781 (
      {stage1_10[167], stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171], stage1_10[172]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[32],stage2_12[44],stage2_11[66],stage2_10[91]}
   );
   gpc615_5 gpc782 (
      {stage1_11[108], stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112]},
      {stage1_12[90]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[15],stage2_13[33],stage2_12[45],stage2_11[67]}
   );
   gpc615_5 gpc783 (
      {stage1_11[113], stage1_11[114], stage1_11[115], stage1_11[116], stage1_11[117]},
      {stage1_12[91]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[16],stage2_13[34],stage2_12[46],stage2_11[68]}
   );
   gpc615_5 gpc784 (
      {stage1_11[118], stage1_11[119], stage1_11[120], stage1_11[121], stage1_11[122]},
      {stage1_12[92]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[17],stage2_13[35],stage2_12[47],stage2_11[69]}
   );
   gpc615_5 gpc785 (
      {stage1_11[123], stage1_11[124], stage1_11[125], stage1_11[126], stage1_11[127]},
      {stage1_12[93]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[18],stage2_13[36],stage2_12[48],stage2_11[70]}
   );
   gpc615_5 gpc786 (
      {stage1_11[128], stage1_11[129], stage1_11[130], stage1_11[131], stage1_11[132]},
      {stage1_12[94]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[19],stage2_13[37],stage2_12[49],stage2_11[71]}
   );
   gpc615_5 gpc787 (
      {stage1_11[133], stage1_11[134], stage1_11[135], stage1_11[136], stage1_11[137]},
      {stage1_12[95]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[20],stage2_13[38],stage2_12[50],stage2_11[72]}
   );
   gpc615_5 gpc788 (
      {stage1_11[138], stage1_11[139], stage1_11[140], stage1_11[141], stage1_11[142]},
      {stage1_12[96]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[21],stage2_13[39],stage2_12[51],stage2_11[73]}
   );
   gpc615_5 gpc789 (
      {stage1_11[143], stage1_11[144], stage1_11[145], stage1_11[146], stage1_11[147]},
      {stage1_12[97]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[22],stage2_13[40],stage2_12[52],stage2_11[74]}
   );
   gpc615_5 gpc790 (
      {stage1_11[148], stage1_11[149], stage1_11[150], stage1_11[151], stage1_11[152]},
      {stage1_12[98]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[23],stage2_13[41],stage2_12[53],stage2_11[75]}
   );
   gpc615_5 gpc791 (
      {stage1_11[153], stage1_11[154], stage1_11[155], stage1_11[156], stage1_11[157]},
      {stage1_12[99]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[24],stage2_13[42],stage2_12[54],stage2_11[76]}
   );
   gpc615_5 gpc792 (
      {stage1_11[158], stage1_11[159], stage1_11[160], stage1_11[161], stage1_11[162]},
      {stage1_12[100]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[25],stage2_13[43],stage2_12[55],stage2_11[77]}
   );
   gpc615_5 gpc793 (
      {stage1_11[163], stage1_11[164], stage1_11[165], stage1_11[166], stage1_11[167]},
      {stage1_12[101]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[26],stage2_13[44],stage2_12[56],stage2_11[78]}
   );
   gpc1_1 gpc794 (
      {stage1_0[78]},
      {stage2_0[23]}
   );
   gpc1_1 gpc795 (
      {stage1_0[79]},
      {stage2_0[24]}
   );
   gpc1_1 gpc796 (
      {stage1_0[80]},
      {stage2_0[25]}
   );
   gpc1_1 gpc797 (
      {stage1_0[81]},
      {stage2_0[26]}
   );
   gpc1_1 gpc798 (
      {stage1_0[82]},
      {stage2_0[27]}
   );
   gpc1_1 gpc799 (
      {stage1_0[83]},
      {stage2_0[28]}
   );
   gpc1_1 gpc800 (
      {stage1_0[84]},
      {stage2_0[29]}
   );
   gpc1_1 gpc801 (
      {stage1_0[85]},
      {stage2_0[30]}
   );
   gpc1_1 gpc802 (
      {stage1_1[120]},
      {stage2_1[23]}
   );
   gpc1_1 gpc803 (
      {stage1_1[121]},
      {stage2_1[24]}
   );
   gpc1_1 gpc804 (
      {stage1_1[122]},
      {stage2_1[25]}
   );
   gpc1_1 gpc805 (
      {stage1_1[123]},
      {stage2_1[26]}
   );
   gpc1_1 gpc806 (
      {stage1_1[124]},
      {stage2_1[27]}
   );
   gpc1_1 gpc807 (
      {stage1_1[125]},
      {stage2_1[28]}
   );
   gpc1_1 gpc808 (
      {stage1_1[126]},
      {stage2_1[29]}
   );
   gpc1_1 gpc809 (
      {stage1_1[127]},
      {stage2_1[30]}
   );
   gpc1_1 gpc810 (
      {stage1_1[128]},
      {stage2_1[31]}
   );
   gpc1_1 gpc811 (
      {stage1_1[129]},
      {stage2_1[32]}
   );
   gpc1_1 gpc812 (
      {stage1_1[130]},
      {stage2_1[33]}
   );
   gpc1_1 gpc813 (
      {stage1_1[131]},
      {stage2_1[34]}
   );
   gpc1_1 gpc814 (
      {stage1_1[132]},
      {stage2_1[35]}
   );
   gpc1_1 gpc815 (
      {stage1_1[133]},
      {stage2_1[36]}
   );
   gpc1_1 gpc816 (
      {stage1_1[134]},
      {stage2_1[37]}
   );
   gpc1_1 gpc817 (
      {stage1_1[135]},
      {stage2_1[38]}
   );
   gpc1_1 gpc818 (
      {stage1_1[136]},
      {stage2_1[39]}
   );
   gpc1_1 gpc819 (
      {stage1_1[137]},
      {stage2_1[40]}
   );
   gpc1_1 gpc820 (
      {stage1_1[138]},
      {stage2_1[41]}
   );
   gpc1_1 gpc821 (
      {stage1_1[139]},
      {stage2_1[42]}
   );
   gpc1_1 gpc822 (
      {stage1_1[140]},
      {stage2_1[43]}
   );
   gpc1_1 gpc823 (
      {stage1_1[141]},
      {stage2_1[44]}
   );
   gpc1_1 gpc824 (
      {stage1_1[142]},
      {stage2_1[45]}
   );
   gpc1_1 gpc825 (
      {stage1_1[143]},
      {stage2_1[46]}
   );
   gpc1_1 gpc826 (
      {stage1_1[144]},
      {stage2_1[47]}
   );
   gpc1_1 gpc827 (
      {stage1_1[145]},
      {stage2_1[48]}
   );
   gpc1_1 gpc828 (
      {stage1_1[146]},
      {stage2_1[49]}
   );
   gpc1_1 gpc829 (
      {stage1_1[147]},
      {stage2_1[50]}
   );
   gpc1_1 gpc830 (
      {stage1_1[148]},
      {stage2_1[51]}
   );
   gpc1_1 gpc831 (
      {stage1_1[149]},
      {stage2_1[52]}
   );
   gpc1_1 gpc832 (
      {stage1_1[150]},
      {stage2_1[53]}
   );
   gpc1_1 gpc833 (
      {stage1_1[151]},
      {stage2_1[54]}
   );
   gpc1_1 gpc834 (
      {stage1_1[152]},
      {stage2_1[55]}
   );
   gpc1_1 gpc835 (
      {stage1_1[153]},
      {stage2_1[56]}
   );
   gpc1_1 gpc836 (
      {stage1_1[154]},
      {stage2_1[57]}
   );
   gpc1_1 gpc837 (
      {stage1_4[240]},
      {stage2_4[88]}
   );
   gpc1_1 gpc838 (
      {stage1_5[228]},
      {stage2_5[73]}
   );
   gpc1_1 gpc839 (
      {stage1_5[229]},
      {stage2_5[74]}
   );
   gpc1_1 gpc840 (
      {stage1_9[234]},
      {stage2_9[85]}
   );
   gpc1_1 gpc841 (
      {stage1_9[235]},
      {stage2_9[86]}
   );
   gpc1_1 gpc842 (
      {stage1_9[236]},
      {stage2_9[87]}
   );
   gpc1_1 gpc843 (
      {stage1_9[237]},
      {stage2_9[88]}
   );
   gpc1_1 gpc844 (
      {stage1_9[238]},
      {stage2_9[89]}
   );
   gpc1_1 gpc845 (
      {stage1_9[239]},
      {stage2_9[90]}
   );
   gpc1_1 gpc846 (
      {stage1_9[240]},
      {stage2_9[91]}
   );
   gpc1_1 gpc847 (
      {stage1_10[173]},
      {stage2_10[92]}
   );
   gpc1_1 gpc848 (
      {stage1_10[174]},
      {stage2_10[93]}
   );
   gpc1_1 gpc849 (
      {stage1_10[175]},
      {stage2_10[94]}
   );
   gpc1_1 gpc850 (
      {stage1_10[176]},
      {stage2_10[95]}
   );
   gpc1_1 gpc851 (
      {stage1_10[177]},
      {stage2_10[96]}
   );
   gpc1_1 gpc852 (
      {stage1_10[178]},
      {stage2_10[97]}
   );
   gpc1_1 gpc853 (
      {stage1_10[179]},
      {stage2_10[98]}
   );
   gpc1_1 gpc854 (
      {stage1_11[168]},
      {stage2_11[79]}
   );
   gpc1_1 gpc855 (
      {stage1_11[169]},
      {stage2_11[80]}
   );
   gpc1_1 gpc856 (
      {stage1_11[170]},
      {stage2_11[81]}
   );
   gpc1_1 gpc857 (
      {stage1_12[102]},
      {stage2_12[57]}
   );
   gpc1_1 gpc858 (
      {stage1_12[103]},
      {stage2_12[58]}
   );
   gpc1_1 gpc859 (
      {stage1_12[104]},
      {stage2_12[59]}
   );
   gpc1_1 gpc860 (
      {stage1_12[105]},
      {stage2_12[60]}
   );
   gpc1_1 gpc861 (
      {stage1_12[106]},
      {stage2_12[61]}
   );
   gpc1_1 gpc862 (
      {stage1_12[107]},
      {stage2_12[62]}
   );
   gpc1_1 gpc863 (
      {stage1_12[108]},
      {stage2_12[63]}
   );
   gpc1_1 gpc864 (
      {stage1_12[109]},
      {stage2_12[64]}
   );
   gpc1_1 gpc865 (
      {stage1_12[110]},
      {stage2_12[65]}
   );
   gpc1_1 gpc866 (
      {stage1_12[111]},
      {stage2_12[66]}
   );
   gpc1_1 gpc867 (
      {stage1_12[112]},
      {stage2_12[67]}
   );
   gpc1_1 gpc868 (
      {stage1_12[113]},
      {stage2_12[68]}
   );
   gpc1_1 gpc869 (
      {stage1_12[114]},
      {stage2_12[69]}
   );
   gpc1_1 gpc870 (
      {stage1_12[115]},
      {stage2_12[70]}
   );
   gpc1_1 gpc871 (
      {stage1_12[116]},
      {stage2_12[71]}
   );
   gpc1_1 gpc872 (
      {stage1_12[117]},
      {stage2_12[72]}
   );
   gpc1_1 gpc873 (
      {stage1_12[118]},
      {stage2_12[73]}
   );
   gpc1_1 gpc874 (
      {stage1_12[119]},
      {stage2_12[74]}
   );
   gpc1_1 gpc875 (
      {stage1_12[120]},
      {stage2_12[75]}
   );
   gpc1_1 gpc876 (
      {stage1_12[121]},
      {stage2_12[76]}
   );
   gpc1_1 gpc877 (
      {stage1_12[122]},
      {stage2_12[77]}
   );
   gpc1_1 gpc878 (
      {stage1_12[123]},
      {stage2_12[78]}
   );
   gpc1_1 gpc879 (
      {stage1_12[124]},
      {stage2_12[79]}
   );
   gpc1_1 gpc880 (
      {stage1_12[125]},
      {stage2_12[80]}
   );
   gpc1_1 gpc881 (
      {stage1_12[126]},
      {stage2_12[81]}
   );
   gpc1_1 gpc882 (
      {stage1_12[127]},
      {stage2_12[82]}
   );
   gpc1_1 gpc883 (
      {stage1_12[128]},
      {stage2_12[83]}
   );
   gpc1_1 gpc884 (
      {stage1_12[129]},
      {stage2_12[84]}
   );
   gpc1_1 gpc885 (
      {stage1_12[130]},
      {stage2_12[85]}
   );
   gpc1_1 gpc886 (
      {stage1_12[131]},
      {stage2_12[86]}
   );
   gpc1_1 gpc887 (
      {stage1_12[132]},
      {stage2_12[87]}
   );
   gpc1_1 gpc888 (
      {stage1_12[133]},
      {stage2_12[88]}
   );
   gpc1_1 gpc889 (
      {stage1_12[134]},
      {stage2_12[89]}
   );
   gpc1_1 gpc890 (
      {stage1_12[135]},
      {stage2_12[90]}
   );
   gpc1_1 gpc891 (
      {stage1_12[136]},
      {stage2_12[91]}
   );
   gpc1_1 gpc892 (
      {stage1_12[137]},
      {stage2_12[92]}
   );
   gpc1_1 gpc893 (
      {stage1_12[138]},
      {stage2_12[93]}
   );
   gpc1_1 gpc894 (
      {stage1_12[139]},
      {stage2_12[94]}
   );
   gpc1_1 gpc895 (
      {stage1_12[140]},
      {stage2_12[95]}
   );
   gpc1_1 gpc896 (
      {stage1_12[141]},
      {stage2_12[96]}
   );
   gpc1_1 gpc897 (
      {stage1_12[142]},
      {stage2_12[97]}
   );
   gpc1_1 gpc898 (
      {stage1_12[143]},
      {stage2_12[98]}
   );
   gpc1_1 gpc899 (
      {stage1_12[144]},
      {stage2_12[99]}
   );
   gpc1_1 gpc900 (
      {stage1_12[145]},
      {stage2_12[100]}
   );
   gpc1_1 gpc901 (
      {stage1_12[146]},
      {stage2_12[101]}
   );
   gpc1_1 gpc902 (
      {stage1_12[147]},
      {stage2_12[102]}
   );
   gpc1_1 gpc903 (
      {stage1_12[148]},
      {stage2_12[103]}
   );
   gpc1_1 gpc904 (
      {stage1_12[149]},
      {stage2_12[104]}
   );
   gpc1_1 gpc905 (
      {stage1_12[150]},
      {stage2_12[105]}
   );
   gpc1_1 gpc906 (
      {stage1_12[151]},
      {stage2_12[106]}
   );
   gpc1_1 gpc907 (
      {stage1_12[152]},
      {stage2_12[107]}
   );
   gpc1_1 gpc908 (
      {stage1_12[153]},
      {stage2_12[108]}
   );
   gpc1_1 gpc909 (
      {stage1_12[154]},
      {stage2_12[109]}
   );
   gpc1_1 gpc910 (
      {stage1_12[155]},
      {stage2_12[110]}
   );
   gpc1_1 gpc911 (
      {stage1_12[156]},
      {stage2_12[111]}
   );
   gpc1_1 gpc912 (
      {stage1_13[72]},
      {stage2_13[45]}
   );
   gpc1_1 gpc913 (
      {stage1_13[73]},
      {stage2_13[46]}
   );
   gpc1_1 gpc914 (
      {stage1_13[74]},
      {stage2_13[47]}
   );
   gpc1_1 gpc915 (
      {stage1_13[75]},
      {stage2_13[48]}
   );
   gpc1_1 gpc916 (
      {stage1_13[76]},
      {stage2_13[49]}
   );
   gpc1_1 gpc917 (
      {stage1_13[77]},
      {stage2_13[50]}
   );
   gpc1_1 gpc918 (
      {stage1_13[78]},
      {stage2_13[51]}
   );
   gpc1163_5 gpc919 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc920 (
      {stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc921 (
      {stage2_0[9], stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc606_5 gpc922 (
      {stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20]},
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc923 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage3_5[0],stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc606_5 gpc924 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[1],stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5]}
   );
   gpc606_5 gpc925 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage3_5[2],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc926 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage3_5[3],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc927 (
      {stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35]},
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30]},
      {stage3_5[4],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc928 (
      {stage2_1[36], stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35], stage2_3[36]},
      {stage3_5[5],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc615_5 gpc929 (
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage2_3[37]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[6],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc615_5 gpc930 (
      {stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28]},
      {stage2_3[38]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[7],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc615_5 gpc931 (
      {stage2_2[29], stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33]},
      {stage2_3[39]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[8],stage3_4[12],stage3_3[12],stage3_2[12]}
   );
   gpc615_5 gpc932 (
      {stage2_2[34], stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38]},
      {stage2_3[40]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[9],stage3_4[13],stage3_3[13],stage3_2[13]}
   );
   gpc615_5 gpc933 (
      {stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43]},
      {stage2_3[41]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[10],stage3_4[14],stage3_3[14],stage3_2[14]}
   );
   gpc615_5 gpc934 (
      {stage2_2[44], stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48]},
      {stage2_3[42]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[11],stage3_4[15],stage3_3[15],stage3_2[15]}
   );
   gpc615_5 gpc935 (
      {stage2_2[49], stage2_2[50], stage2_2[51], stage2_2[52], stage2_2[53]},
      {stage2_3[43]},
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage3_6[6],stage3_5[12],stage3_4[16],stage3_3[16],stage3_2[16]}
   );
   gpc615_5 gpc936 (
      {stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48]},
      {stage2_4[42]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[7],stage3_5[13],stage3_4[17],stage3_3[17]}
   );
   gpc615_5 gpc937 (
      {stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53]},
      {stage2_4[43]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[8],stage3_5[14],stage3_4[18],stage3_3[18]}
   );
   gpc615_5 gpc938 (
      {stage2_3[54], stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58]},
      {stage2_4[44]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[9],stage3_5[15],stage3_4[19],stage3_3[19]}
   );
   gpc615_5 gpc939 (
      {stage2_3[59], stage2_3[60], stage2_3[61], stage2_3[62], stage2_3[63]},
      {stage2_4[45]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[10],stage3_5[16],stage3_4[20],stage3_3[20]}
   );
   gpc615_5 gpc940 (
      {stage2_3[64], stage2_3[65], stage2_3[66], stage2_3[67], stage2_3[68]},
      {stage2_4[46]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[11],stage3_5[17],stage3_4[21],stage3_3[21]}
   );
   gpc615_5 gpc941 (
      {stage2_3[69], stage2_3[70], stage2_3[71], stage2_3[72], stage2_3[73]},
      {stage2_4[47]},
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage3_7[5],stage3_6[12],stage3_5[18],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc942 (
      {stage2_3[74], stage2_3[75], stage2_3[76], stage2_3[77], stage2_3[78]},
      {stage2_4[48]},
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage3_7[6],stage3_6[13],stage3_5[19],stage3_4[23],stage3_3[23]}
   );
   gpc615_5 gpc943 (
      {stage2_3[79], stage2_3[80], stage2_3[81], stage2_3[82], stage2_3[83]},
      {stage2_4[49]},
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage3_7[7],stage3_6[14],stage3_5[20],stage3_4[24],stage3_3[24]}
   );
   gpc606_5 gpc944 (
      {stage2_4[50], stage2_4[51], stage2_4[52], stage2_4[53], stage2_4[54], stage2_4[55]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[8],stage3_6[15],stage3_5[21],stage3_4[25]}
   );
   gpc606_5 gpc945 (
      {stage2_4[56], stage2_4[57], stage2_4[58], stage2_4[59], stage2_4[60], stage2_4[61]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[9],stage3_6[16],stage3_5[22],stage3_4[26]}
   );
   gpc606_5 gpc946 (
      {stage2_4[62], stage2_4[63], stage2_4[64], stage2_4[65], stage2_4[66], stage2_4[67]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[10],stage3_6[17],stage3_5[23],stage3_4[27]}
   );
   gpc606_5 gpc947 (
      {stage2_4[68], stage2_4[69], stage2_4[70], stage2_4[71], stage2_4[72], stage2_4[73]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[11],stage3_6[18],stage3_5[24],stage3_4[28]}
   );
   gpc606_5 gpc948 (
      {stage2_4[74], stage2_4[75], stage2_4[76], stage2_4[77], stage2_4[78], stage2_4[79]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[12],stage3_6[19],stage3_5[25],stage3_4[29]}
   );
   gpc606_5 gpc949 (
      {stage2_4[80], stage2_4[81], stage2_4[82], stage2_4[83], stage2_4[84], stage2_4[85]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[13],stage3_6[20],stage3_5[26],stage3_4[30]}
   );
   gpc606_5 gpc950 (
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[6],stage3_7[14],stage3_6[21],stage3_5[27]}
   );
   gpc606_5 gpc951 (
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[7],stage3_7[15],stage3_6[22],stage3_5[28]}
   );
   gpc615_5 gpc952 (
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64]},
      {stage2_6[36]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[8],stage3_7[16],stage3_6[23],stage3_5[29]}
   );
   gpc615_5 gpc953 (
      {stage2_5[65], stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69]},
      {stage2_6[37]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[9],stage3_7[17],stage3_6[24],stage3_5[30]}
   );
   gpc615_5 gpc954 (
      {stage2_5[70], stage2_5[71], stage2_5[72], stage2_5[73], stage2_5[74]},
      {stage2_6[38]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[10],stage3_7[18],stage3_6[25],stage3_5[31]}
   );
   gpc615_5 gpc955 (
      {stage2_6[39], stage2_6[40], stage2_6[41], stage2_6[42], stage2_6[43]},
      {stage2_7[30]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[5],stage3_8[11],stage3_7[19],stage3_6[26]}
   );
   gpc615_5 gpc956 (
      {stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47], stage2_6[48]},
      {stage2_7[31]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[6],stage3_8[12],stage3_7[20],stage3_6[27]}
   );
   gpc615_5 gpc957 (
      {stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52], stage2_6[53]},
      {stage2_7[32]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[7],stage3_8[13],stage3_7[21],stage3_6[28]}
   );
   gpc615_5 gpc958 (
      {stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57], stage2_6[58]},
      {stage2_7[33]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[8],stage3_8[14],stage3_7[22],stage3_6[29]}
   );
   gpc615_5 gpc959 (
      {stage2_6[59], stage2_6[60], stage2_6[61], stage2_6[62], stage2_6[63]},
      {stage2_7[34]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[9],stage3_8[15],stage3_7[23],stage3_6[30]}
   );
   gpc615_5 gpc960 (
      {stage2_6[64], stage2_6[65], stage2_6[66], stage2_6[67], stage2_6[68]},
      {stage2_7[35]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[10],stage3_8[16],stage3_7[24],stage3_6[31]}
   );
   gpc615_5 gpc961 (
      {stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72], stage2_6[73]},
      {stage2_7[36]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[11],stage3_8[17],stage3_7[25],stage3_6[32]}
   );
   gpc615_5 gpc962 (
      {stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77], stage2_6[78]},
      {stage2_7[37]},
      {stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage3_10[7],stage3_9[12],stage3_8[18],stage3_7[26],stage3_6[33]}
   );
   gpc615_5 gpc963 (
      {stage2_6[79], stage2_6[80], stage2_6[81], stage2_6[82], stage2_6[83]},
      {stage2_7[38]},
      {stage2_8[48], stage2_8[49], stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53]},
      {stage3_10[8],stage3_9[13],stage3_8[19],stage3_7[27],stage3_6[34]}
   );
   gpc615_5 gpc964 (
      {stage2_6[84], stage2_6[85], stage2_6[86], stage2_6[87], stage2_6[88]},
      {stage2_7[39]},
      {stage2_8[54], stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59]},
      {stage3_10[9],stage3_9[14],stage3_8[20],stage3_7[28],stage3_6[35]}
   );
   gpc606_5 gpc965 (
      {stage2_7[40], stage2_7[41], stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[10],stage3_9[15],stage3_8[21],stage3_7[29]}
   );
   gpc606_5 gpc966 (
      {stage2_7[46], stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[11],stage3_9[16],stage3_8[22],stage3_7[30]}
   );
   gpc606_5 gpc967 (
      {stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56], stage2_7[57]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[12],stage3_9[17],stage3_8[23],stage3_7[31]}
   );
   gpc606_5 gpc968 (
      {stage2_7[58], stage2_7[59], stage2_7[60], stage2_7[61], stage2_7[62], stage2_7[63]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[13],stage3_9[18],stage3_8[24],stage3_7[32]}
   );
   gpc615_5 gpc969 (
      {stage2_7[64], stage2_7[65], stage2_7[66], stage2_7[67], stage2_7[68]},
      {stage2_8[60]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[14],stage3_9[19],stage3_8[25],stage3_7[33]}
   );
   gpc615_5 gpc970 (
      {stage2_7[69], stage2_7[70], stage2_7[71], stage2_7[72], stage2_7[73]},
      {stage2_8[61]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[15],stage3_9[20],stage3_8[26],stage3_7[34]}
   );
   gpc615_5 gpc971 (
      {stage2_7[74], stage2_7[75], stage2_7[76], stage2_7[77], stage2_7[78]},
      {stage2_8[62]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[16],stage3_9[21],stage3_8[27],stage3_7[35]}
   );
   gpc615_5 gpc972 (
      {stage2_7[79], stage2_7[80], stage2_7[81], stage2_7[82], stage2_7[83]},
      {stage2_8[63]},
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage3_11[7],stage3_10[17],stage3_9[22],stage3_8[28],stage3_7[36]}
   );
   gpc615_5 gpc973 (
      {stage2_7[84], stage2_7[85], stage2_7[86], stage2_7[87], stage2_7[88]},
      {stage2_8[64]},
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage3_11[8],stage3_10[18],stage3_9[23],stage3_8[29],stage3_7[37]}
   );
   gpc606_5 gpc974 (
      {stage2_8[65], stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[9],stage3_10[19],stage3_9[24],stage3_8[30]}
   );
   gpc1163_5 gpc975 (
      {stage2_9[54], stage2_9[55], stage2_9[56]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage2_11[0]},
      {stage2_12[0]},
      {stage3_13[0],stage3_12[1],stage3_11[10],stage3_10[20],stage3_9[25]}
   );
   gpc1163_5 gpc976 (
      {stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage2_11[1]},
      {stage2_12[1]},
      {stage3_13[1],stage3_12[2],stage3_11[11],stage3_10[21],stage3_9[26]}
   );
   gpc1163_5 gpc977 (
      {stage2_9[60], stage2_9[61], stage2_9[62]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage2_11[2]},
      {stage2_12[2]},
      {stage3_13[2],stage3_12[3],stage3_11[12],stage3_10[22],stage3_9[27]}
   );
   gpc1163_5 gpc978 (
      {stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage2_11[3]},
      {stage2_12[3]},
      {stage3_13[3],stage3_12[4],stage3_11[13],stage3_10[23],stage3_9[28]}
   );
   gpc615_5 gpc979 (
      {stage2_9[66], stage2_9[67], stage2_9[68], stage2_9[69], stage2_9[70]},
      {stage2_10[30]},
      {stage2_11[4], stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9]},
      {stage3_13[4],stage3_12[5],stage3_11[14],stage3_10[24],stage3_9[29]}
   );
   gpc615_5 gpc980 (
      {stage2_9[71], stage2_9[72], stage2_9[73], stage2_9[74], stage2_9[75]},
      {stage2_10[31]},
      {stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15]},
      {stage3_13[5],stage3_12[6],stage3_11[15],stage3_10[25],stage3_9[30]}
   );
   gpc615_5 gpc981 (
      {stage2_9[76], stage2_9[77], stage2_9[78], stage2_9[79], stage2_9[80]},
      {stage2_10[32]},
      {stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21]},
      {stage3_13[6],stage3_12[7],stage3_11[16],stage3_10[26],stage3_9[31]}
   );
   gpc606_5 gpc982 (
      {stage2_10[33], stage2_10[34], stage2_10[35], stage2_10[36], stage2_10[37], stage2_10[38]},
      {stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9]},
      {stage3_14[0],stage3_13[7],stage3_12[8],stage3_11[17],stage3_10[27]}
   );
   gpc606_5 gpc983 (
      {stage2_10[39], stage2_10[40], stage2_10[41], stage2_10[42], stage2_10[43], stage2_10[44]},
      {stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15]},
      {stage3_14[1],stage3_13[8],stage3_12[9],stage3_11[18],stage3_10[28]}
   );
   gpc606_5 gpc984 (
      {stage2_10[45], stage2_10[46], stage2_10[47], stage2_10[48], stage2_10[49], stage2_10[50]},
      {stage2_12[16], stage2_12[17], stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21]},
      {stage3_14[2],stage3_13[9],stage3_12[10],stage3_11[19],stage3_10[29]}
   );
   gpc606_5 gpc985 (
      {stage2_10[51], stage2_10[52], stage2_10[53], stage2_10[54], stage2_10[55], stage2_10[56]},
      {stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27]},
      {stage3_14[3],stage3_13[10],stage3_12[11],stage3_11[20],stage3_10[30]}
   );
   gpc606_5 gpc986 (
      {stage2_10[57], stage2_10[58], stage2_10[59], stage2_10[60], stage2_10[61], stage2_10[62]},
      {stage2_12[28], stage2_12[29], stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33]},
      {stage3_14[4],stage3_13[11],stage3_12[12],stage3_11[21],stage3_10[31]}
   );
   gpc606_5 gpc987 (
      {stage2_10[63], stage2_10[64], stage2_10[65], stage2_10[66], stage2_10[67], stage2_10[68]},
      {stage2_12[34], stage2_12[35], stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39]},
      {stage3_14[5],stage3_13[12],stage3_12[13],stage3_11[22],stage3_10[32]}
   );
   gpc606_5 gpc988 (
      {stage2_10[69], stage2_10[70], stage2_10[71], stage2_10[72], stage2_10[73], stage2_10[74]},
      {stage2_12[40], stage2_12[41], stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45]},
      {stage3_14[6],stage3_13[13],stage3_12[14],stage3_11[23],stage3_10[33]}
   );
   gpc606_5 gpc989 (
      {stage2_10[75], stage2_10[76], stage2_10[77], stage2_10[78], stage2_10[79], stage2_10[80]},
      {stage2_12[46], stage2_12[47], stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51]},
      {stage3_14[7],stage3_13[14],stage3_12[15],stage3_11[24],stage3_10[34]}
   );
   gpc606_5 gpc990 (
      {stage2_10[81], stage2_10[82], stage2_10[83], stage2_10[84], stage2_10[85], stage2_10[86]},
      {stage2_12[52], stage2_12[53], stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57]},
      {stage3_14[8],stage3_13[15],stage3_12[16],stage3_11[25],stage3_10[35]}
   );
   gpc606_5 gpc991 (
      {stage2_10[87], stage2_10[88], stage2_10[89], stage2_10[90], stage2_10[91], stage2_10[92]},
      {stage2_12[58], stage2_12[59], stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63]},
      {stage3_14[9],stage3_13[16],stage3_12[17],stage3_11[26],stage3_10[36]}
   );
   gpc606_5 gpc992 (
      {stage2_10[93], stage2_10[94], stage2_10[95], stage2_10[96], stage2_10[97], stage2_10[98]},
      {stage2_12[64], stage2_12[65], stage2_12[66], stage2_12[67], stage2_12[68], stage2_12[69]},
      {stage3_14[10],stage3_13[17],stage3_12[18],stage3_11[27],stage3_10[37]}
   );
   gpc606_5 gpc993 (
      {stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[11],stage3_13[18],stage3_12[19],stage3_11[28]}
   );
   gpc606_5 gpc994 (
      {stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[12],stage3_13[19],stage3_12[20],stage3_11[29]}
   );
   gpc606_5 gpc995 (
      {stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[13],stage3_13[20],stage3_12[21],stage3_11[30]}
   );
   gpc606_5 gpc996 (
      {stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[14],stage3_13[21],stage3_12[22],stage3_11[31]}
   );
   gpc606_5 gpc997 (
      {stage2_11[46], stage2_11[47], stage2_11[48], stage2_11[49], stage2_11[50], stage2_11[51]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[15],stage3_13[22],stage3_12[23],stage3_11[32]}
   );
   gpc606_5 gpc998 (
      {stage2_11[52], stage2_11[53], stage2_11[54], stage2_11[55], stage2_11[56], stage2_11[57]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[16],stage3_13[23],stage3_12[24],stage3_11[33]}
   );
   gpc615_5 gpc999 (
      {stage2_11[58], stage2_11[59], stage2_11[60], stage2_11[61], stage2_11[62]},
      {stage2_12[70]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[17],stage3_13[24],stage3_12[25],stage3_11[34]}
   );
   gpc606_5 gpc1000 (
      {stage2_12[71], stage2_12[72], stage2_12[73], stage2_12[74], stage2_12[75], stage2_12[76]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[7],stage3_14[18],stage3_13[25],stage3_12[26]}
   );
   gpc606_5 gpc1001 (
      {stage2_12[77], stage2_12[78], stage2_12[79], stage2_12[80], stage2_12[81], stage2_12[82]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[8],stage3_14[19],stage3_13[26],stage3_12[27]}
   );
   gpc606_5 gpc1002 (
      {stage2_12[83], stage2_12[84], stage2_12[85], stage2_12[86], stage2_12[87], stage2_12[88]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[9],stage3_14[20],stage3_13[27],stage3_12[28]}
   );
   gpc606_5 gpc1003 (
      {stage2_12[89], stage2_12[90], stage2_12[91], stage2_12[92], stage2_12[93], stage2_12[94]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[10],stage3_14[21],stage3_13[28],stage3_12[29]}
   );
   gpc606_5 gpc1004 (
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[11],stage3_14[22],stage3_13[29]}
   );
   gpc1_1 gpc1005 (
      {stage2_0[21]},
      {stage3_0[4]}
   );
   gpc1_1 gpc1006 (
      {stage2_0[22]},
      {stage3_0[5]}
   );
   gpc1_1 gpc1007 (
      {stage2_0[23]},
      {stage3_0[6]}
   );
   gpc1_1 gpc1008 (
      {stage2_0[24]},
      {stage3_0[7]}
   );
   gpc1_1 gpc1009 (
      {stage2_0[25]},
      {stage3_0[8]}
   );
   gpc1_1 gpc1010 (
      {stage2_0[26]},
      {stage3_0[9]}
   );
   gpc1_1 gpc1011 (
      {stage2_0[27]},
      {stage3_0[10]}
   );
   gpc1_1 gpc1012 (
      {stage2_0[28]},
      {stage3_0[11]}
   );
   gpc1_1 gpc1013 (
      {stage2_0[29]},
      {stage3_0[12]}
   );
   gpc1_1 gpc1014 (
      {stage2_0[30]},
      {stage3_0[13]}
   );
   gpc1_1 gpc1015 (
      {stage2_1[42]},
      {stage3_1[10]}
   );
   gpc1_1 gpc1016 (
      {stage2_1[43]},
      {stage3_1[11]}
   );
   gpc1_1 gpc1017 (
      {stage2_1[44]},
      {stage3_1[12]}
   );
   gpc1_1 gpc1018 (
      {stage2_1[45]},
      {stage3_1[13]}
   );
   gpc1_1 gpc1019 (
      {stage2_1[46]},
      {stage3_1[14]}
   );
   gpc1_1 gpc1020 (
      {stage2_1[47]},
      {stage3_1[15]}
   );
   gpc1_1 gpc1021 (
      {stage2_1[48]},
      {stage3_1[16]}
   );
   gpc1_1 gpc1022 (
      {stage2_1[49]},
      {stage3_1[17]}
   );
   gpc1_1 gpc1023 (
      {stage2_1[50]},
      {stage3_1[18]}
   );
   gpc1_1 gpc1024 (
      {stage2_1[51]},
      {stage3_1[19]}
   );
   gpc1_1 gpc1025 (
      {stage2_1[52]},
      {stage3_1[20]}
   );
   gpc1_1 gpc1026 (
      {stage2_1[53]},
      {stage3_1[21]}
   );
   gpc1_1 gpc1027 (
      {stage2_1[54]},
      {stage3_1[22]}
   );
   gpc1_1 gpc1028 (
      {stage2_1[55]},
      {stage3_1[23]}
   );
   gpc1_1 gpc1029 (
      {stage2_1[56]},
      {stage3_1[24]}
   );
   gpc1_1 gpc1030 (
      {stage2_1[57]},
      {stage3_1[25]}
   );
   gpc1_1 gpc1031 (
      {stage2_4[86]},
      {stage3_4[31]}
   );
   gpc1_1 gpc1032 (
      {stage2_4[87]},
      {stage3_4[32]}
   );
   gpc1_1 gpc1033 (
      {stage2_4[88]},
      {stage3_4[33]}
   );
   gpc1_1 gpc1034 (
      {stage2_6[89]},
      {stage3_6[36]}
   );
   gpc1_1 gpc1035 (
      {stage2_6[90]},
      {stage3_6[37]}
   );
   gpc1_1 gpc1036 (
      {stage2_6[91]},
      {stage3_6[38]}
   );
   gpc1_1 gpc1037 (
      {stage2_6[92]},
      {stage3_6[39]}
   );
   gpc1_1 gpc1038 (
      {stage2_6[93]},
      {stage3_6[40]}
   );
   gpc1_1 gpc1039 (
      {stage2_6[94]},
      {stage3_6[41]}
   );
   gpc1_1 gpc1040 (
      {stage2_6[95]},
      {stage3_6[42]}
   );
   gpc1_1 gpc1041 (
      {stage2_6[96]},
      {stage3_6[43]}
   );
   gpc1_1 gpc1042 (
      {stage2_6[97]},
      {stage3_6[44]}
   );
   gpc1_1 gpc1043 (
      {stage2_9[81]},
      {stage3_9[32]}
   );
   gpc1_1 gpc1044 (
      {stage2_9[82]},
      {stage3_9[33]}
   );
   gpc1_1 gpc1045 (
      {stage2_9[83]},
      {stage3_9[34]}
   );
   gpc1_1 gpc1046 (
      {stage2_9[84]},
      {stage3_9[35]}
   );
   gpc1_1 gpc1047 (
      {stage2_9[85]},
      {stage3_9[36]}
   );
   gpc1_1 gpc1048 (
      {stage2_9[86]},
      {stage3_9[37]}
   );
   gpc1_1 gpc1049 (
      {stage2_9[87]},
      {stage3_9[38]}
   );
   gpc1_1 gpc1050 (
      {stage2_9[88]},
      {stage3_9[39]}
   );
   gpc1_1 gpc1051 (
      {stage2_9[89]},
      {stage3_9[40]}
   );
   gpc1_1 gpc1052 (
      {stage2_9[90]},
      {stage3_9[41]}
   );
   gpc1_1 gpc1053 (
      {stage2_9[91]},
      {stage3_9[42]}
   );
   gpc1_1 gpc1054 (
      {stage2_11[63]},
      {stage3_11[35]}
   );
   gpc1_1 gpc1055 (
      {stage2_11[64]},
      {stage3_11[36]}
   );
   gpc1_1 gpc1056 (
      {stage2_11[65]},
      {stage3_11[37]}
   );
   gpc1_1 gpc1057 (
      {stage2_11[66]},
      {stage3_11[38]}
   );
   gpc1_1 gpc1058 (
      {stage2_11[67]},
      {stage3_11[39]}
   );
   gpc1_1 gpc1059 (
      {stage2_11[68]},
      {stage3_11[40]}
   );
   gpc1_1 gpc1060 (
      {stage2_11[69]},
      {stage3_11[41]}
   );
   gpc1_1 gpc1061 (
      {stage2_11[70]},
      {stage3_11[42]}
   );
   gpc1_1 gpc1062 (
      {stage2_11[71]},
      {stage3_11[43]}
   );
   gpc1_1 gpc1063 (
      {stage2_11[72]},
      {stage3_11[44]}
   );
   gpc1_1 gpc1064 (
      {stage2_11[73]},
      {stage3_11[45]}
   );
   gpc1_1 gpc1065 (
      {stage2_11[74]},
      {stage3_11[46]}
   );
   gpc1_1 gpc1066 (
      {stage2_11[75]},
      {stage3_11[47]}
   );
   gpc1_1 gpc1067 (
      {stage2_11[76]},
      {stage3_11[48]}
   );
   gpc1_1 gpc1068 (
      {stage2_11[77]},
      {stage3_11[49]}
   );
   gpc1_1 gpc1069 (
      {stage2_11[78]},
      {stage3_11[50]}
   );
   gpc1_1 gpc1070 (
      {stage2_11[79]},
      {stage3_11[51]}
   );
   gpc1_1 gpc1071 (
      {stage2_11[80]},
      {stage3_11[52]}
   );
   gpc1_1 gpc1072 (
      {stage2_11[81]},
      {stage3_11[53]}
   );
   gpc1_1 gpc1073 (
      {stage2_12[95]},
      {stage3_12[30]}
   );
   gpc1_1 gpc1074 (
      {stage2_12[96]},
      {stage3_12[31]}
   );
   gpc1_1 gpc1075 (
      {stage2_12[97]},
      {stage3_12[32]}
   );
   gpc1_1 gpc1076 (
      {stage2_12[98]},
      {stage3_12[33]}
   );
   gpc1_1 gpc1077 (
      {stage2_12[99]},
      {stage3_12[34]}
   );
   gpc1_1 gpc1078 (
      {stage2_12[100]},
      {stage3_12[35]}
   );
   gpc1_1 gpc1079 (
      {stage2_12[101]},
      {stage3_12[36]}
   );
   gpc1_1 gpc1080 (
      {stage2_12[102]},
      {stage3_12[37]}
   );
   gpc1_1 gpc1081 (
      {stage2_12[103]},
      {stage3_12[38]}
   );
   gpc1_1 gpc1082 (
      {stage2_12[104]},
      {stage3_12[39]}
   );
   gpc1_1 gpc1083 (
      {stage2_12[105]},
      {stage3_12[40]}
   );
   gpc1_1 gpc1084 (
      {stage2_12[106]},
      {stage3_12[41]}
   );
   gpc1_1 gpc1085 (
      {stage2_12[107]},
      {stage3_12[42]}
   );
   gpc1_1 gpc1086 (
      {stage2_12[108]},
      {stage3_12[43]}
   );
   gpc1_1 gpc1087 (
      {stage2_12[109]},
      {stage3_12[44]}
   );
   gpc1_1 gpc1088 (
      {stage2_12[110]},
      {stage3_12[45]}
   );
   gpc1_1 gpc1089 (
      {stage2_12[111]},
      {stage3_12[46]}
   );
   gpc1_1 gpc1090 (
      {stage2_13[48]},
      {stage3_13[30]}
   );
   gpc1_1 gpc1091 (
      {stage2_13[49]},
      {stage3_13[31]}
   );
   gpc1_1 gpc1092 (
      {stage2_13[50]},
      {stage3_13[32]}
   );
   gpc1_1 gpc1093 (
      {stage2_13[51]},
      {stage3_13[33]}
   );
   gpc1_1 gpc1094 (
      {stage2_14[24]},
      {stage3_14[23]}
   );
   gpc1_1 gpc1095 (
      {stage2_14[25]},
      {stage3_14[24]}
   );
   gpc1_1 gpc1096 (
      {stage2_14[26]},
      {stage3_14[25]}
   );
   gpc1_1 gpc1097 (
      {stage2_15[6]},
      {stage3_15[12]}
   );
   gpc1_1 gpc1098 (
      {stage2_15[7]},
      {stage3_15[13]}
   );
   gpc1_1 gpc1099 (
      {stage2_15[8]},
      {stage3_15[14]}
   );
   gpc1_1 gpc1100 (
      {stage2_15[9]},
      {stage3_15[15]}
   );
   gpc1_1 gpc1101 (
      {stage2_15[10]},
      {stage3_15[16]}
   );
   gpc1_1 gpc1102 (
      {stage2_15[11]},
      {stage3_15[17]}
   );
   gpc606_5 gpc1103 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc1104 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc1105 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc1106 (
      {stage3_1[12], stage3_1[13], stage3_1[14], stage3_1[15], stage3_1[16], stage3_1[17]},
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17]},
      {stage4_5[2],stage4_4[3],stage4_3[3],stage4_2[3],stage4_1[3]}
   );
   gpc615_5 gpc1107 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10]},
      {stage3_3[18]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[3],stage4_4[4],stage4_3[4],stage4_2[4]}
   );
   gpc615_5 gpc1108 (
      {stage3_2[11], stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15]},
      {stage3_3[19]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[4],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc615_5 gpc1109 (
      {stage3_3[20], stage3_3[21], stage3_3[22], stage3_3[23], stage3_3[24]},
      {stage3_4[12]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[2],stage4_5[5],stage4_4[6],stage4_3[6]}
   );
   gpc606_5 gpc1110 (
      {stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17], stage3_4[18]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[1],stage4_6[3],stage4_5[6],stage4_4[7]}
   );
   gpc606_5 gpc1111 (
      {stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23], stage3_4[24]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[2],stage4_6[4],stage4_5[7],stage4_4[8]}
   );
   gpc606_5 gpc1112 (
      {stage3_4[25], stage3_4[26], stage3_4[27], stage3_4[28], stage3_4[29], stage3_4[30]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[2],stage4_7[3],stage4_6[5],stage4_5[8],stage4_4[9]}
   );
   gpc606_5 gpc1113 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[3],stage4_7[4],stage4_6[6],stage4_5[9]}
   );
   gpc606_5 gpc1114 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[4],stage4_7[5],stage4_6[7],stage4_5[10]}
   );
   gpc606_5 gpc1115 (
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[5],stage4_7[6],stage4_6[8],stage4_5[11]}
   );
   gpc606_5 gpc1116 (
      {stage3_5[24], stage3_5[25], stage3_5[26], stage3_5[27], stage3_5[28], stage3_5[29]},
      {stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23]},
      {stage4_9[3],stage4_8[6],stage4_7[7],stage4_6[9],stage4_5[12]}
   );
   gpc606_5 gpc1117 (
      {stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[4],stage4_8[7],stage4_7[8],stage4_6[10]}
   );
   gpc615_5 gpc1118 (
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28]},
      {stage3_7[24]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[5],stage4_8[8],stage4_7[9],stage4_6[11]}
   );
   gpc615_5 gpc1119 (
      {stage3_6[29], stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33]},
      {stage3_7[25]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[6],stage4_8[9],stage4_7[10],stage4_6[12]}
   );
   gpc615_5 gpc1120 (
      {stage3_6[34], stage3_6[35], stage3_6[36], stage3_6[37], stage3_6[38]},
      {stage3_7[26]},
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22], stage3_8[23]},
      {stage4_10[3],stage4_9[7],stage4_8[10],stage4_7[11],stage4_6[13]}
   );
   gpc615_5 gpc1121 (
      {stage3_6[39], stage3_6[40], stage3_6[41], stage3_6[42], stage3_6[43]},
      {stage3_7[27]},
      {stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27], stage3_8[28], stage3_8[29]},
      {stage4_10[4],stage4_9[8],stage4_8[11],stage4_7[12],stage4_6[14]}
   );
   gpc615_5 gpc1122 (
      {stage3_7[28], stage3_7[29], stage3_7[30], stage3_7[31], stage3_7[32]},
      {stage3_8[30]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[5],stage4_9[9],stage4_8[12],stage4_7[13]}
   );
   gpc606_5 gpc1123 (
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[6],stage4_9[10]}
   );
   gpc606_5 gpc1124 (
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[2],stage4_10[7],stage4_9[11]}
   );
   gpc606_5 gpc1125 (
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[2],stage4_11[3],stage4_10[8],stage4_9[12]}
   );
   gpc606_5 gpc1126 (
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage4_13[3],stage4_12[3],stage4_11[4],stage4_10[9],stage4_9[13]}
   );
   gpc606_5 gpc1127 (
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage3_11[24], stage3_11[25], stage3_11[26], stage3_11[27], stage3_11[28], stage3_11[29]},
      {stage4_13[4],stage4_12[4],stage4_11[5],stage4_10[10],stage4_9[14]}
   );
   gpc606_5 gpc1128 (
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage3_11[30], stage3_11[31], stage3_11[32], stage3_11[33], stage3_11[34], stage3_11[35]},
      {stage4_13[5],stage4_12[5],stage4_11[6],stage4_10[11],stage4_9[15]}
   );
   gpc2135_5 gpc1129 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4]},
      {stage3_11[36], stage3_11[37], stage3_11[38]},
      {stage3_12[0]},
      {stage3_13[0], stage3_13[1]},
      {stage4_14[0],stage4_13[6],stage4_12[6],stage4_11[7],stage4_10[12]}
   );
   gpc2135_5 gpc1130 (
      {stage3_10[5], stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9]},
      {stage3_11[39], stage3_11[40], stage3_11[41]},
      {stage3_12[1]},
      {stage3_13[2], stage3_13[3]},
      {stage4_14[1],stage4_13[7],stage4_12[7],stage4_11[8],stage4_10[13]}
   );
   gpc2135_5 gpc1131 (
      {stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13], stage3_10[14]},
      {stage3_11[42], stage3_11[43], stage3_11[44]},
      {stage3_12[2]},
      {stage3_13[4], stage3_13[5]},
      {stage4_14[2],stage4_13[8],stage4_12[8],stage4_11[9],stage4_10[14]}
   );
   gpc2135_5 gpc1132 (
      {stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19]},
      {stage3_11[45], stage3_11[46], stage3_11[47]},
      {stage3_12[3]},
      {stage3_13[6], stage3_13[7]},
      {stage4_14[3],stage4_13[9],stage4_12[9],stage4_11[10],stage4_10[15]}
   );
   gpc606_5 gpc1133 (
      {stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24], stage3_10[25]},
      {stage3_12[4], stage3_12[5], stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9]},
      {stage4_14[4],stage4_13[10],stage4_12[10],stage4_11[11],stage4_10[16]}
   );
   gpc606_5 gpc1134 (
      {stage3_10[26], stage3_10[27], stage3_10[28], stage3_10[29], stage3_10[30], stage3_10[31]},
      {stage3_12[10], stage3_12[11], stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15]},
      {stage4_14[5],stage4_13[11],stage4_12[11],stage4_11[12],stage4_10[17]}
   );
   gpc606_5 gpc1135 (
      {stage3_10[32], stage3_10[33], stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37]},
      {stage3_12[16], stage3_12[17], stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21]},
      {stage4_14[6],stage4_13[12],stage4_12[12],stage4_11[13],stage4_10[18]}
   );
   gpc615_5 gpc1136 (
      {stage3_11[48], stage3_11[49], stage3_11[50], stage3_11[51], stage3_11[52]},
      {stage3_12[22]},
      {stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], stage3_13[13]},
      {stage4_15[0],stage4_14[7],stage4_13[13],stage4_12[13],stage4_11[14]}
   );
   gpc606_5 gpc1137 (
      {stage3_12[23], stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[8],stage4_13[14],stage4_12[14]}
   );
   gpc606_5 gpc1138 (
      {stage3_12[29], stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[2],stage4_14[9],stage4_13[15],stage4_12[15]}
   );
   gpc606_5 gpc1139 (
      {stage3_12[35], stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40]},
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17]},
      {stage4_16[2],stage4_15[3],stage4_14[10],stage4_13[16],stage4_12[16]}
   );
   gpc606_5 gpc1140 (
      {stage3_12[41], stage3_12[42], stage3_12[43], stage3_12[44], stage3_12[45], stage3_12[46]},
      {stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage4_16[3],stage4_15[4],stage4_14[11],stage4_13[17],stage4_12[17]}
   );
   gpc606_5 gpc1141 (
      {stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[4],stage4_15[5],stage4_14[12],stage4_13[18]}
   );
   gpc606_5 gpc1142 (
      {stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24], stage3_13[25]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[5],stage4_15[6],stage4_14[13],stage4_13[19]}
   );
   gpc606_5 gpc1143 (
      {stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30], stage3_13[31]},
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17]},
      {stage4_17[2],stage4_16[6],stage4_15[7],stage4_14[14],stage4_13[20]}
   );
   gpc1_1 gpc1144 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1145 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc1146 (
      {stage3_0[8]},
      {stage4_0[3]}
   );
   gpc1_1 gpc1147 (
      {stage3_0[9]},
      {stage4_0[4]}
   );
   gpc1_1 gpc1148 (
      {stage3_0[10]},
      {stage4_0[5]}
   );
   gpc1_1 gpc1149 (
      {stage3_0[11]},
      {stage4_0[6]}
   );
   gpc1_1 gpc1150 (
      {stage3_0[12]},
      {stage4_0[7]}
   );
   gpc1_1 gpc1151 (
      {stage3_0[13]},
      {stage4_0[8]}
   );
   gpc1_1 gpc1152 (
      {stage3_1[18]},
      {stage4_1[4]}
   );
   gpc1_1 gpc1153 (
      {stage3_1[19]},
      {stage4_1[5]}
   );
   gpc1_1 gpc1154 (
      {stage3_1[20]},
      {stage4_1[6]}
   );
   gpc1_1 gpc1155 (
      {stage3_1[21]},
      {stage4_1[7]}
   );
   gpc1_1 gpc1156 (
      {stage3_1[22]},
      {stage4_1[8]}
   );
   gpc1_1 gpc1157 (
      {stage3_1[23]},
      {stage4_1[9]}
   );
   gpc1_1 gpc1158 (
      {stage3_1[24]},
      {stage4_1[10]}
   );
   gpc1_1 gpc1159 (
      {stage3_1[25]},
      {stage4_1[11]}
   );
   gpc1_1 gpc1160 (
      {stage3_2[16]},
      {stage4_2[6]}
   );
   gpc1_1 gpc1161 (
      {stage3_4[31]},
      {stage4_4[10]}
   );
   gpc1_1 gpc1162 (
      {stage3_4[32]},
      {stage4_4[11]}
   );
   gpc1_1 gpc1163 (
      {stage3_4[33]},
      {stage4_4[12]}
   );
   gpc1_1 gpc1164 (
      {stage3_5[30]},
      {stage4_5[13]}
   );
   gpc1_1 gpc1165 (
      {stage3_5[31]},
      {stage4_5[14]}
   );
   gpc1_1 gpc1166 (
      {stage3_6[44]},
      {stage4_6[15]}
   );
   gpc1_1 gpc1167 (
      {stage3_7[33]},
      {stage4_7[14]}
   );
   gpc1_1 gpc1168 (
      {stage3_7[34]},
      {stage4_7[15]}
   );
   gpc1_1 gpc1169 (
      {stage3_7[35]},
      {stage4_7[16]}
   );
   gpc1_1 gpc1170 (
      {stage3_7[36]},
      {stage4_7[17]}
   );
   gpc1_1 gpc1171 (
      {stage3_7[37]},
      {stage4_7[18]}
   );
   gpc1_1 gpc1172 (
      {stage3_9[42]},
      {stage4_9[16]}
   );
   gpc1_1 gpc1173 (
      {stage3_11[53]},
      {stage4_11[15]}
   );
   gpc1_1 gpc1174 (
      {stage3_13[32]},
      {stage4_13[21]}
   );
   gpc1_1 gpc1175 (
      {stage3_13[33]},
      {stage4_13[22]}
   );
   gpc1_1 gpc1176 (
      {stage3_14[24]},
      {stage4_14[15]}
   );
   gpc1_1 gpc1177 (
      {stage3_14[25]},
      {stage4_14[16]}
   );
   gpc1_1 gpc1178 (
      {stage3_16[0]},
      {stage4_16[7]}
   );
   gpc1_1 gpc1179 (
      {stage3_16[1]},
      {stage4_16[8]}
   );
   gpc1_1 gpc1180 (
      {stage3_16[2]},
      {stage4_16[9]}
   );
   gpc1_1 gpc1181 (
      {stage3_16[3]},
      {stage4_16[10]}
   );
   gpc1_1 gpc1182 (
      {stage3_16[4]},
      {stage4_16[11]}
   );
   gpc1_1 gpc1183 (
      {stage3_17[0]},
      {stage4_17[3]}
   );
   gpc1163_5 gpc1184 (
      {stage4_0[0], stage4_0[1], stage4_0[2]},
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_2[0]},
      {stage4_3[0]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc623_5 gpc1185 (
      {stage4_2[1], stage4_2[2], stage4_2[3]},
      {stage4_3[1], stage4_3[2]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage5_6[0],stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1]}
   );
   gpc606_5 gpc1186 (
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10], stage4_4[11]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[1],stage5_4[2]}
   );
   gpc615_5 gpc1187 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4]},
      {stage4_6[6]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[2],stage5_5[2]}
   );
   gpc615_5 gpc1188 (
      {stage4_5[5], stage4_5[6], stage4_5[7], stage4_5[8], stage4_5[9]},
      {stage4_6[7]},
      {stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage5_9[1],stage5_8[2],stage5_7[2],stage5_6[3],stage5_5[3]}
   );
   gpc615_5 gpc1189 (
      {stage4_5[10], stage4_5[11], stage4_5[12], stage4_5[13], stage4_5[14]},
      {stage4_6[8]},
      {stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16], stage4_7[17]},
      {stage5_9[2],stage5_8[3],stage5_7[3],stage5_6[4],stage5_5[4]}
   );
   gpc606_5 gpc1190 (
      {stage4_6[9], stage4_6[10], stage4_6[11], stage4_6[12], stage4_6[13], stage4_6[14]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[3],stage5_8[4],stage5_7[4],stage5_6[5]}
   );
   gpc2135_5 gpc1191 (
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[4]}
   );
   gpc2135_5 gpc1192 (
      {stage4_9[5], stage4_9[6], stage4_9[7], stage4_9[8], stage4_9[9]},
      {stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage4_11[1]},
      {stage4_12[2], stage4_12[3]},
      {stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[2],stage5_9[5]}
   );
   gpc7_3 gpc1193 (
      {stage4_9[10], stage4_9[11], stage4_9[12], stage4_9[13], stage4_9[14], stage4_9[15], stage4_9[16]},
      {stage5_11[2],stage5_10[3],stage5_9[6]}
   );
   gpc2135_5 gpc1194 (
      {stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9], stage4_10[10]},
      {stage4_11[2], stage4_11[3], stage4_11[4]},
      {stage4_12[4]},
      {stage4_13[0], stage4_13[1]},
      {stage5_14[0],stage5_13[2],stage5_12[2],stage5_11[3],stage5_10[4]}
   );
   gpc606_5 gpc1195 (
      {stage4_10[11], stage4_10[12], stage4_10[13], stage4_10[14], stage4_10[15], stage4_10[16]},
      {stage4_12[5], stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10]},
      {stage5_14[1],stage5_13[3],stage5_12[3],stage5_11[4],stage5_10[5]}
   );
   gpc615_5 gpc1196 (
      {stage4_11[5], stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9]},
      {stage4_12[11]},
      {stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6], stage4_13[7]},
      {stage5_15[0],stage5_14[2],stage5_13[4],stage5_12[4],stage5_11[5]}
   );
   gpc615_5 gpc1197 (
      {stage4_11[10], stage4_11[11], stage4_11[12], stage4_11[13], stage4_11[14]},
      {stage4_12[12]},
      {stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12], stage4_13[13]},
      {stage5_15[1],stage5_14[3],stage5_13[5],stage5_12[5],stage5_11[6]}
   );
   gpc606_5 gpc1198 (
      {stage4_12[13], stage4_12[14], stage4_12[15], stage4_12[16], stage4_12[17], 1'b0},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[2],stage5_14[4],stage5_13[6],stage5_12[6]}
   );
   gpc606_5 gpc1199 (
      {stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18], stage4_13[19]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[1],stage5_15[3],stage5_14[5],stage5_13[7]}
   );
   gpc606_5 gpc1200 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10], stage4_14[11]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[1],stage5_16[2],stage5_15[4],stage5_14[6]}
   );
   gpc615_5 gpc1201 (
      {stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15], stage4_14[16]},
      {stage4_15[6]},
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11]},
      {stage5_18[1],stage5_17[2],stage5_16[3],stage5_15[5],stage5_14[7]}
   );
   gpc1_1 gpc1202 (
      {stage4_0[3]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1203 (
      {stage4_0[4]},
      {stage5_0[2]}
   );
   gpc1_1 gpc1204 (
      {stage4_0[5]},
      {stage5_0[3]}
   );
   gpc1_1 gpc1205 (
      {stage4_0[6]},
      {stage5_0[4]}
   );
   gpc1_1 gpc1206 (
      {stage4_0[7]},
      {stage5_0[5]}
   );
   gpc1_1 gpc1207 (
      {stage4_0[8]},
      {stage5_0[6]}
   );
   gpc1_1 gpc1208 (
      {stage4_1[6]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1209 (
      {stage4_1[7]},
      {stage5_1[2]}
   );
   gpc1_1 gpc1210 (
      {stage4_1[8]},
      {stage5_1[3]}
   );
   gpc1_1 gpc1211 (
      {stage4_1[9]},
      {stage5_1[4]}
   );
   gpc1_1 gpc1212 (
      {stage4_1[10]},
      {stage5_1[5]}
   );
   gpc1_1 gpc1213 (
      {stage4_1[11]},
      {stage5_1[6]}
   );
   gpc1_1 gpc1214 (
      {stage4_2[4]},
      {stage5_2[2]}
   );
   gpc1_1 gpc1215 (
      {stage4_2[5]},
      {stage5_2[3]}
   );
   gpc1_1 gpc1216 (
      {stage4_2[6]},
      {stage5_2[4]}
   );
   gpc1_1 gpc1217 (
      {stage4_3[3]},
      {stage5_3[2]}
   );
   gpc1_1 gpc1218 (
      {stage4_3[4]},
      {stage5_3[3]}
   );
   gpc1_1 gpc1219 (
      {stage4_3[5]},
      {stage5_3[4]}
   );
   gpc1_1 gpc1220 (
      {stage4_3[6]},
      {stage5_3[5]}
   );
   gpc1_1 gpc1221 (
      {stage4_4[12]},
      {stage5_4[3]}
   );
   gpc1_1 gpc1222 (
      {stage4_6[15]},
      {stage5_6[6]}
   );
   gpc1_1 gpc1223 (
      {stage4_7[18]},
      {stage5_7[5]}
   );
   gpc1_1 gpc1224 (
      {stage4_8[6]},
      {stage5_8[5]}
   );
   gpc1_1 gpc1225 (
      {stage4_8[7]},
      {stage5_8[6]}
   );
   gpc1_1 gpc1226 (
      {stage4_8[8]},
      {stage5_8[7]}
   );
   gpc1_1 gpc1227 (
      {stage4_8[9]},
      {stage5_8[8]}
   );
   gpc1_1 gpc1228 (
      {stage4_8[10]},
      {stage5_8[9]}
   );
   gpc1_1 gpc1229 (
      {stage4_8[11]},
      {stage5_8[10]}
   );
   gpc1_1 gpc1230 (
      {stage4_8[12]},
      {stage5_8[11]}
   );
   gpc1_1 gpc1231 (
      {stage4_10[17]},
      {stage5_10[6]}
   );
   gpc1_1 gpc1232 (
      {stage4_10[18]},
      {stage5_10[7]}
   );
   gpc1_1 gpc1233 (
      {stage4_11[15]},
      {stage5_11[7]}
   );
   gpc1_1 gpc1234 (
      {stage4_13[20]},
      {stage5_13[8]}
   );
   gpc1_1 gpc1235 (
      {stage4_13[21]},
      {stage5_13[9]}
   );
   gpc1_1 gpc1236 (
      {stage4_13[22]},
      {stage5_13[10]}
   );
   gpc1_1 gpc1237 (
      {stage4_15[7]},
      {stage5_15[6]}
   );
   gpc1_1 gpc1238 (
      {stage4_17[0]},
      {stage5_17[3]}
   );
   gpc1_1 gpc1239 (
      {stage4_17[1]},
      {stage5_17[4]}
   );
   gpc1_1 gpc1240 (
      {stage4_17[2]},
      {stage5_17[5]}
   );
   gpc1_1 gpc1241 (
      {stage4_17[3]},
      {stage5_17[6]}
   );
   gpc117_4 gpc1242 (
      {stage5_0[0], stage5_0[1], stage5_0[2], stage5_0[3], stage5_0[4], stage5_0[5], stage5_0[6]},
      {stage5_1[0]},
      {stage5_2[0]},
      {stage6_3[0],stage6_2[0],stage6_1[0],stage6_0[0]}
   );
   gpc215_4 gpc1243 (
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4]},
      {stage5_6[0]},
      {stage5_7[0], stage5_7[1]},
      {stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[0]}
   );
   gpc615_5 gpc1244 (
      {stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5]},
      {stage5_7[2]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage6_10[0],stage6_9[0],stage6_8[1],stage6_7[1],stage6_6[1]}
   );
   gpc623_5 gpc1245 (
      {stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage5_8[6], stage5_8[7]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[1],stage6_9[1],stage6_8[2],stage6_7[2]}
   );
   gpc1163_5 gpc1246 (
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[0],stage6_11[1],stage6_10[2]}
   );
   gpc615_5 gpc1247 (
      {stage5_10[3], stage5_10[4], stage5_10[5], stage5_10[6], stage5_10[7]},
      {stage5_11[6]},
      {stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6]},
      {stage6_14[1],stage6_13[1],stage6_12[1],stage6_11[2],stage6_10[3]}
   );
   gpc1163_5 gpc1248 (
      {stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[0]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[2],stage6_13[2]}
   );
   gpc615_5 gpc1249 (
      {stage5_13[4], stage5_13[5], stage5_13[6], stage5_13[7], stage5_13[8]},
      {stage5_14[6]},
      {stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5], stage5_15[6]},
      {stage6_17[1],stage6_16[1],stage6_15[1],stage6_14[3],stage6_13[3]}
   );
   gpc1163_5 gpc1250 (
      {stage5_16[1], stage5_16[2], stage5_16[3]},
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage5_18[0]},
      {1'b0},
      {stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[2],stage6_16[2]}
   );
   gpc1_1 gpc1251 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc1252 (
      {stage5_1[2]},
      {stage6_1[2]}
   );
   gpc1_1 gpc1253 (
      {stage5_1[3]},
      {stage6_1[3]}
   );
   gpc1_1 gpc1254 (
      {stage5_1[4]},
      {stage6_1[4]}
   );
   gpc1_1 gpc1255 (
      {stage5_1[5]},
      {stage6_1[5]}
   );
   gpc1_1 gpc1256 (
      {stage5_1[6]},
      {stage6_1[6]}
   );
   gpc1_1 gpc1257 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc1258 (
      {stage5_2[2]},
      {stage6_2[2]}
   );
   gpc1_1 gpc1259 (
      {stage5_2[3]},
      {stage6_2[3]}
   );
   gpc1_1 gpc1260 (
      {stage5_2[4]},
      {stage6_2[4]}
   );
   gpc1_1 gpc1261 (
      {stage5_3[0]},
      {stage6_3[1]}
   );
   gpc1_1 gpc1262 (
      {stage5_3[1]},
      {stage6_3[2]}
   );
   gpc1_1 gpc1263 (
      {stage5_3[2]},
      {stage6_3[3]}
   );
   gpc1_1 gpc1264 (
      {stage5_3[3]},
      {stage6_3[4]}
   );
   gpc1_1 gpc1265 (
      {stage5_3[4]},
      {stage6_3[5]}
   );
   gpc1_1 gpc1266 (
      {stage5_3[5]},
      {stage6_3[6]}
   );
   gpc1_1 gpc1267 (
      {stage5_4[0]},
      {stage6_4[0]}
   );
   gpc1_1 gpc1268 (
      {stage5_4[1]},
      {stage6_4[1]}
   );
   gpc1_1 gpc1269 (
      {stage5_4[2]},
      {stage6_4[2]}
   );
   gpc1_1 gpc1270 (
      {stage5_4[3]},
      {stage6_4[3]}
   );
   gpc1_1 gpc1271 (
      {stage5_6[6]},
      {stage6_6[2]}
   );
   gpc1_1 gpc1272 (
      {stage5_8[8]},
      {stage6_8[3]}
   );
   gpc1_1 gpc1273 (
      {stage5_8[9]},
      {stage6_8[4]}
   );
   gpc1_1 gpc1274 (
      {stage5_8[10]},
      {stage6_8[5]}
   );
   gpc1_1 gpc1275 (
      {stage5_8[11]},
      {stage6_8[6]}
   );
   gpc1_1 gpc1276 (
      {stage5_9[6]},
      {stage6_9[2]}
   );
   gpc1_1 gpc1277 (
      {stage5_11[7]},
      {stage6_11[3]}
   );
   gpc1_1 gpc1278 (
      {stage5_13[9]},
      {stage6_13[4]}
   );
   gpc1_1 gpc1279 (
      {stage5_13[10]},
      {stage6_13[5]}
   );
   gpc1_1 gpc1280 (
      {stage5_14[7]},
      {stage6_14[4]}
   );
   gpc1_1 gpc1281 (
      {stage5_17[6]},
      {stage6_17[3]}
   );
   gpc1_1 gpc1282 (
      {stage5_18[1]},
      {stage6_18[1]}
   );
   gpc606_5 gpc1283 (
      {stage6_1[0], stage6_1[1], stage6_1[2], stage6_1[3], stage6_1[4], stage6_1[5]},
      {stage6_3[0], stage6_3[1], stage6_3[2], stage6_3[3], stage6_3[4], stage6_3[5]},
      {stage7_5[0],stage7_4[0],stage7_3[0],stage7_2[0],stage7_1[0]}
   );
   gpc1415_5 gpc1284 (
      {stage6_2[0], stage6_2[1], stage6_2[2], stage6_2[3], stage6_2[4]},
      {stage6_3[6]},
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3]},
      {stage6_5[0]},
      {stage7_6[0],stage7_5[1],stage7_4[1],stage7_3[1],stage7_2[1]}
   );
   gpc623_5 gpc1285 (
      {stage6_6[0], stage6_6[1], stage6_6[2]},
      {stage6_7[0], stage6_7[1]},
      {stage6_8[0], stage6_8[1], stage6_8[2], stage6_8[3], stage6_8[4], stage6_8[5]},
      {stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[0],stage7_6[1]}
   );
   gpc1343_5 gpc1286 (
      {stage6_9[0], stage6_9[1], stage6_9[2]},
      {stage6_10[0], stage6_10[1], stage6_10[2], stage6_10[3]},
      {stage6_11[0], stage6_11[1], stage6_11[2]},
      {stage6_12[0]},
      {stage7_13[0],stage7_12[0],stage7_11[0],stage7_10[1],stage7_9[1]}
   );
   gpc207_4 gpc1287 (
      {stage6_13[0], stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5], 1'b0},
      {stage6_15[0], stage6_15[1]},
      {stage7_16[0],stage7_15[0],stage7_14[0],stage7_13[1]}
   );
   gpc1406_5 gpc1288 (
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], 1'b0},
      {stage6_16[0], stage6_16[1], stage6_16[2], 1'b0},
      {stage6_17[0]},
      {stage7_18[0],stage7_17[0],stage7_16[1],stage7_15[1],stage7_14[1]}
   );
   gpc135_4 gpc1289 (
      {stage6_17[1], stage6_17[2], stage6_17[3], 1'b0, 1'b0},
      {stage6_18[0], stage6_18[1], 1'b0},
      {stage6_19[0]},
      {stage7_20[0],stage7_19[0],stage7_18[1],stage7_17[1]}
   );
   gpc1_1 gpc1290 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc1291 (
      {stage6_1[6]},
      {stage7_1[1]}
   );
   gpc1_1 gpc1292 (
      {stage6_7[2]},
      {stage7_7[1]}
   );
   gpc1_1 gpc1293 (
      {stage6_8[6]},
      {stage7_8[1]}
   );
   gpc1_1 gpc1294 (
      {stage6_11[3]},
      {stage7_11[1]}
   );
   gpc1_1 gpc1295 (
      {stage6_12[1]},
      {stage7_12[1]}
   );
   gpc1_1 gpc1296 (
      {stage6_20[0]},
      {stage7_20[1]}
   );
endmodule

module testbench();
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [20:0] srcsum;
    wire [20:0] dstsum;
    wire test;
    compressor_CLA486_12 compressor_CLA486_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hcf671cde836c875406a3b698118e2e6f4b40420c92c06bb277755f3a75f226de016014f508b854f37e26d5d1c6d9c752db1a301976f37c6dddea2bf873056a7f0d26fe5e04b64cd525fa62b8bc2d657adc0c86fd3bb442bf37ed5262f6ec6f650c1beb04e21f861b498ef601109c017b243b328a50dac745a1041e96af7b09cb85fc4c2ddd79a10c5b90b664c59f1f711a775c7d07f731b076fe2668964b82fbf0a3ad85792f6ecc7a727281ef9bcced632ddfd3d8c68610cc58fee749c7839a810b722f110f54770acb2da5acef244ba0d61a0d87d710258b066148b5e97405e37ce10f97e3619f1fe4b76470f118dc58365f3d2198e916a36f87d3441361cd0811aa71fe01d9af29bba85ddfe28eddced93c55cf2c43ce993e67ba6979df971a50eeb1ad795a211dfc9d59d6073a0968ae86dd6ae7174c00c7ebee767a100f3493178177dd3cb409a6fdd15e05e1285a437e16c45f0d741945be7e49f677354cacdfed89ac23a78c34baf026e80199d59d55f6676edaadca1afb63622eb9f26d45ee7bd98b893d543efe7f0a0b11de40dff1c68daa39a7a92390b9c662aae6aa2ab7ed14769b0b0c11ade5f890fdafdeaffca6fc46b9fbad81329b3b5a02eead723da2bf34cdd59f808aaa0d3db9da48cb0de3a1bd0adfaad253fbadfd9bf0524b20b4cbacf5d7e6c3299acf7861ab61d411f49501dec9720357abbaa5f9df08e24d926e2808a3339dbe6977095e4be4be20542abd6f9fd611f5aa4f2e5756baaddb2711e273b81d5a2905a9307a5ad14ba1b1332a34363c1d9ee2871d8e12432d1cb91a4ac84db0cc7c59994dae4d82279d413d3ea8409ecc40c56b3e14b45486b23d373f606d0eb0f323898626214db70ed5d8d68ee7a4a197438209207d3bfa4ce75e614d2a3ab3cf62b69d7e1ec009467fa01603f162d0c9eca5f983b03db2b45cee7de6e15a8d3d40ab72fe951feff7b74cbb97c862ca5c703db6edbc040cde730f382fc4e8e28a61898f080c1cb1490b88b0e6f57e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h19b7df22870762f71ebde9223689117e5c58ff89284ed4718044358983d8a00276d0594d4f987ddb7db5de710fc152fef64cac749139de3ab78c70209277b6f17f6690ba2804ab87071a93946c7c4bf7efc524791226aae91c11ad45d474bd37143dcf4c9d032897db8303948f29202f0f36d6af05cbb28da9abd399e8810196fbe2cd62bfeb349077ef77fc79c44a4753c12f5959eae479a704799f974d5982f96d7faba93a3baeea2be53b3ed81cf517bce019bef709f1ccda746972ba1193129b1fb8e04a366b4ea48006a6848b0bb065de6f4b2dbd799d591dbf33a16278c5dd9685d6aa0a576d446537291d28b9df391c3391da339526cf3782587e7a72594ecf9b47bb93f2da277ba4905a018785b0e825efd6e4b13b61f69e67d9f35889e67c70c53a4feb09914c149f47f763632f016002e691b30105c91841ea65c31ad5dcbe8dffe75db789df98d9ba8aec3c37e6af1c7f51a1fe97f2ac078507cc8783fdb6e79c6581a8e95b3641a52699f5d56f368374516742aee955efbfa001d42bb03fffc0970b16dd99ee9b0e51d904ceefae8cd27231afb46347fabfa12cc703540776ca15da2008c8cd6148922be8c57b482a70eb5873d12f34d5aa072dd59f55dbcea3447b3593a52b548513d78d16f9ae3af76d7feac2cad9a7afaa9686b4c63912ff7c3215dbe0af44022a7db3c53265d6f2acee072713d6fb478426a523790efbfa4a5d8c0db2a93ae7f62068b472a1c22e98bb7af5fb0cbac31dc2ed8f27121682e6dfa6064e5e23e5f43ef0b2d58ff1e4a6e7c562e6e23cd5c46b6baa6d15fbbefb789b0333fbab739d333680c603dbedff6940b31c20727e42e1de727e835a6ac9d08e5708c2ecf01b4c4dc81f6d15ac233a73cc86f97d922c2c7d676d735b2c4ff0d196cb80ff3280b2e9158ecb983c92ec2f5398d2eafd2b06dbaf34edf9719646c7c9b13bcd498c6998dd91ff99b23702ce2a79e1aadcf4659527ee116ec1ab9ef2c33b4b73fba44875b7170b1336fe838f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h9cf2617147e65774558ab85b8489780a515d3d5bc48cbcdbff43ae1950ea5f80eec7b15410e44adad2132d07afc1654b4d39ce3b1696ce76f179144c2fd4028206614c1d98c51b0658861c1d41361a9c1421a57fbb8dfb8860fa40554b0c5f16fa2eb6585d5c3683c8fee343f8568064ff8ef9ab1b7b49e10f6657d0b9baa3238953c6300466b06d340b3850a5271e10663a1c09f41431227b88c56e3e88b3dde5315fbe801cb0771e729a00ff0388365debbfcfe6337a8793c9ea0edd3a2bb85ec8398d75fb06a709f16d31f30a574932cffef672c7d75474c69118cd72c224c8a5e2e7f82ca685c94a71f3f3ed670deae56c49d2a3a93cf32f05dfd0b065ffddac60b0fda4d49d07e86bc2a14bd3e70cbc2939194daddc87be63661a28ed18f96baec54ca78c5e22ce3c612b9de3251c255f79c9301505df5b28ef8f90e42aa31fd9125db96c9040528562b1477ff53ee2e961fdbbc0aae78a459b3295ae2caaab91b8ef63896abcf5e88585ef1187fef4ebbd90f2c073be48b55c339d76dc3058012786d47008e5a783dc80a47c307033d8c50ec757b09ba07fe8b0961b2aa7ad4a6fc4de06247d84093e2f7c1b5b162bd42f9aaf4925e51a6c590f67a654ca9259aaf75c8db8c791c45a9596058c4a62930e09bc682eeb58acf656781fcc5b2c46101e5d2ed7b1a2f41ab46ff168721db915ada906e59eb150ad87e1c7388edb25d883846e275b1f5ad1daad1b0e17825f1583b2a9931b7c7a9f85d59d141261a5ab4309a42c7453b3614ad66f147b3895751eef36f1f99e58850a8823070af5f2922efe4fb8ca1a88ead051bf74a08d6759f8115a33d740ca8563d3c1d79cc1d2627ba2f142287e7fabdf10dee8364512cd4c106a739e23ebe6616820bfcaf68da5b0accf0ca0274cfc61a5e89c257da8ffe80668565dc70dc1122cc54590ea52e41f241c0f8c4b1812ee74e185aabde13f3b055ff3a2d3f357eb0a8e3e6d438c8fad7827e45c417849d84988dbe00accacad0f6fa482;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h55e5705a78225f20e177a67b86f527ad6625a472aed81b902bad4ee3ad70d40a160a23dd6092248bcaa6dcd0cfd5726cf4f146c4550aaddc44f3fe42d7e9db855a025e8bf346340c9698b01efb4cba430c6e88a230670482801f551d6ccd7866fb8684e777462e00b0336eb38dee0d7fd1219fc876e85f83fcd17a848d0d6c8e8f11d5c8268039baeb7d00947f0f3ed80b0fe00d425c71c7b8e1269e02a9b26f21159bd8f4c081fc04b547f65bed728fca9f672bf1eae5b3e09fe650085658e47331e7971033f1026545ea538f7cb1318cdbb8b9cd648347f21acb4c0a18ce518e8f7bf9459d612a55994f29bf070429341d5dd7c0768f11e10830dc03c437be655701105147fe9a00b57b623873d3c81edc22d61d633a14713acf418004d42a4cdc1a4ffd75577ca2611ae704776742bc0220f6b53ec1428d2dcd29ddefa3d078efb6bff528dbe40997665993e882086f21811b6c6a8832d38492fef57a55741cab14d8d86d97ede68de6bfa293f974a86a27cf8294d43b71abbb02d120dc0faad917a40c7b74f6712114e176f4a2ca02692d3db071cc1f6f75dddd262d3b69dcf478128a27c9eb2cc4d8d19f06c98f51e213de6002024ddd33e8949dd9ee2d3e0ad112c22db978682449bd266cc2988989c0f7a938f4169a69ccfb0d22aa6f31765bdade8c615d2c60b746e1963b255868e4dbc4551282ebf636385c5827f58988b8eec920b6b0b5968fba94dc5fc542b6e8768894055d14b7100297deeb8dc609a109e672f3ca5a45f9e00762d951d001d47f23e30c2391952e02f9ff88fec0048b64b089925579fce335305ee90e0283e437e5334d61251be9ee0b299beba6392b2977393dac90a829cd97b1838a44a3f9dd287148220f3b00b2ed18b6ad0b3c7d3614c323dbdf14bd79f05cf9c07c3a930250e52e004376f3098e3f3c5a36622e99e3f96bffef975da981c6a94a4f65b2ab48b2b598a3af3e5b3a9e59a3a7a3a08d2235fc7602b073bd9ad59dc5dc64dc365740805cfe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hde3b4553348c8301f846f884a8ab8a6c20042984f6e83e1d5ee2795701b8e3756137624cbbe3ada61c8ffcf0d872344d64b9621e819b443c69e041154c91e724ef3163277199e5718ef83614dd12993a69aeb44ee28f419677afe36d6f5452bb9779f775941f9087a35603a157b87c3269205d8b19bc7e92a051a4991051b514cbbbe1377ca875fb531e7422a9fcb0989d1127d2539aa3cde0197444a6c5a9a071e7fdec40eb8a25f140c76da5df32b925b7b6556ce3e5bf0e57abe8b863cd80a4baaf875b3ad674061c8b8b7a4c45187efc9c43b6a623f9350338a88713047b055aaa9ecc89f8bec922c6248edcd0ae804bda61f4f1eaf36ff5bd2a0a96dca246388cee75c05f614088389c3c9d5399ef5070960179ff5ba3b2c86addcb01e936d58c64d8130ac4d1f3c0cc9caa6efcd7c1713678daf4f3475b1f65a4c3efb4ff5d70dd843ba663890857a20225c8d72c1df773ba4a6dc62ad9d9e41317aec40422324806b8d496a1bd0c4d3fd321e65fdf7fc95cc565b5d5262a702ff174bd27d521675b69080b409bda9d120ac64949168bdf750fba4398f72e5d4f9c8d7a969a4d34e6d1635de7f5b9a712081104c29037b6d5ba7a7f6edd37d379b4122a7cc78124b8263b441f3b58fa93f0100a76a27b25a0bf49de72901859397c6610e9b23ed8f10e50596eaedb93ec1fe663b5a6ceb2d8993260955e1d45de11d45073f2fc779bb994804bd12cd4b1550ff05fb1b18f59f394c72941e1dadc697644c6c046875706f7807106fa171ceb2e9e92f7d1d6307436a162b517a6825b691232e1a354f2ace25ad3ae122e7bf7567cde9124e0bf0605708318af63efd954c918a585a184b2cb259e7e8a067ea1765e73dba2ea4c70f48c4d58345e2d4fbda8dba697330a026e61af73ecd7cc8460ec501262e3273e7ca10ffc4d818e3af0419828a8cdbcca26b10f3bc45d624129ffb5617608a98279ed0e4111b1b35615219c6d50e24522c928726ad9297dee47e839d29ceb7cf7104086;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h5c6cb8960c43a75e1ba754b4e95bf973f32b6b86598e88d652e60ec27ba8586bc2fcb9e8b1da57116e85ef59471a8f8b3415ee49f6df11fa9873a405a7d4af9cb889cf24b3d21e636ca24218f2fadee29f38d7cd8dd465dcd7b325efaec2a8426bd0f3e4b54e65c18100bf52d6fc603372d35aac0971f917c3436b24492b9850b30e8fd35dba4992d9a5bdfb8c5cd0e5c5285691bef484b76d1446d82bf1f4560b80646b6d68ab07b4dd91460739c983111390fbf675379bfbd56f0ed770f2d93a85c81758ecff86d47ceb0c41f4e253fbdf1f1120ac6dd30134fc22bf3d8d39e11a7ed35cc6c2cacb8f29eb866dbd38ceb265b1b4b7566b4f4f2fa5ed1705f0c1521617c3e2f49ac3b042a95b70166832a170c1e7acfab2d2c2368a63ebbc16954b12184585889c497674e6e3dc95ecc99bfdd0c7e6a8e77f6b22213e9405acaba5a6120d0a21501e8e10bc9e489e547bafac66bfc099d851fbfeb57d9d13fdf9a93cd4e5eb43b6d7e682dbd1702b8bc229a23bf11a64fbeb4b5435b0366dada4eb038ff3dfa77a8e7c58bc255dbe31af17d7baf5306531939ccab54863828e4928b9de74f455d3b52a294b85a5b8b62240e9b2242e2e6e091cd2bd19f8513efae763d1cce93e7055c4e26d7ae38906f83eeb657ca6a6b899614e8fa367abfab78267d6b948fffbc0e1ed20ce9f906368fea949bcd0453279c30d14018bb2bc9e6baaf6a24c7b32ff0a23e863a96ce3a669e2bf8a0dc9794ed2a2287dd5449700ba67304651b1a7408f30f3d2769f737ac3031e058faf8ce1fa94cb93ab56f26a319dc75f4156b15f1c7a47603cec53e77c8f3ff56f3b8a885657a626220012c4caac26c6e5c833a6bed2191dd86d9640000338643874a264bf348ee3f4f3e5cb8d40018dc26e4c29178031ef7f21f97ebdcf1162a76e29532ea86dc1167150ad9cf9401bae2e73619aec0be130efa6437c095e4a004dcefa22264f4ce4c31ec528dd3aaf81635b5538003fe017b4804a6a28aa61b99777b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h1ff8aa5287d6001b39f39827c510e7215ab22cc6bf6a22f6d7ca7006acec1e6bdcbd0217936512164e9311c83d563df37db52fd936f396e2b64be64cd0850e713632962f4ced796dec3ccef29aa1839522704ac4d09cceb52d4a9d297ef09a6709d1d0fbe61c2f413e10babcb0b70d7bc0f8a20040cd19e435c7e22c5be0825bbbce6729d30b43118fb90ad3ba023d8ef1371eab360a79ef510089c90b7b8d204df76e3ee131d9450cc2c00cc932c203a5c43c2f9fe8d340f9d7d919f1c81e45111fe0a1e6fed82a94752960ab584076166f3864def75e71281dad9fd949f90d0f64b44d1fed940fdb983d5545950150f3d133f1f74472dc6b318931bdcc14e23730c87f0c045d704fb2a82cb1f52bf85510e17385aed899860fce6c5e601bb897de771aecfa9036c2c5162136b495b6ecc66b9524a5f7630e8e52f3e79d7678a3ff4dacc8ae21e59ead9267e99d395280635ff112e4c48849589d6a1133ecad03e0156ddae0d09e5475165ab66fb63be559c5e304a6dfac8b951f0e1f71135db90ff3860978240c742cbaae6ed7da8694ebc16296e375c4af4cb801238e0223f49e81b5dcb6bc33eef78d0ac895a7a33657453c988bc54dee048f4a6cb60019c761b2ed4284191176a4efc188f60cfe03b2b40e25ad5fa0ed8676012fd76d17e33afeb5ea09fc331206e97fc91348d62f96c12209e656d886d4bed088fdabe0a51478c6e4f9805ca0b75c27f175df6cca716e8cd33357ead1eea6881d7ebf985ee2d38801474135034e80d843c4f6d5c3d0b4724eaa9d026d1a2ddb4d27bbbd54bd11f611ba5bcf4abd95ff365d118145c21f4560abe25bccf1957a09b2c549882bbcd1c4f4398bafee3ac33e94f73fa5346a4732481c8bdeb08608f6240d6a3c209de5229906f977f97422fba9e2ca3d008f3260e41cca14510dfad02f21011e1d1aab89a070b5ee2f633482d21b4fc4002aefbe9969ef75aea5a83dc11ebfa2379620bdb6a8fd6c0607e769ac108530aace88bbbeba5807;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h29f664ca5046d13eed39af4450b84c24b2a62107d31e8972ab2dff4a87ab249943751689632d8b65e779c9426a1ea994a28103b23622c1378d66fcba6b1474760a6312a0bcf990b061ab08227390b47ace186a356162dc930ff5e64687dd0a9238ef89d4a3fa4a9379f89351fda8152781b25c08adb787a6a0c6890df52caec61091a5d99a7d7915f6cb31980dbd47caaeb5130c2919f9a67b325deaeb86717e6e45a62d94a4fbbc127fcc93ceed35e5f731381d1a6449f324fa6caac5a25a3d3f548e9ab4f3b07b1fedcb1f06cf7659d263522eb04793681335b141eac84bf293a3f9a2e24b34374afdd15f4c2245c99e5f26154de6f5d702da2e49a237506869f56c42e1d7c6ad2a943416425df09da236634b52d1b8d8e162f650e2187f93f8dc265d1bfe83a01f89d5ed5a70e1141f0560c57e1dd5d51fd3c31d01155cbaab47782462cb50ca1fd6b5b18c8418cda53eac57fc46be9d0432032158b974a15303a3e0efc2c29fb0a72afec133751da25023358ebb178ff1bf37a915bf99c0723527f023b12a480b8e18c563eaa07af9f5c07f4b81a6a1b432596acef0ba41264da226a34cb5599e74cdbcb4ec6afbfa380f09fb4deca25507dab6a1c1b18a5c67f32b89dd092a38e0a2dc97fc9c295a757a7cf8f58076ef4191901367039f6b10d7dec65f37e38727e9b16f8aac7a28c7e176d92be35139d98cc28e8879d8e141d083866ba282b932586fb50114d56dad73d01052bb339e570b97f8e4b3569ab42bcb364264960f0e4eddd3beb9beda93ce9a8b57786574f3c72adcce2787f2a9b24e9b7ad14364c1753af7f0b3200c3d063893b8b78f4224622edc3a9000187c731f47f11c822f5f00e8318bdbbbf8fede6c961824ae99f0364644a8302e10c91e474f9eb6dbb33e0bec01a103a5ba42152e4a4e1cd4c59dae5904590c903094dd056d428d1049e61a871783bb4fb75292e7d6e8756cb1b52011d0286ded0c14cdd1cd66adc70d2ffbab8341f497a08308aabc7926dc02;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h727a8914c06403270a75f6e18eb2d0720c845f05908c0b0f3d5188bfd902a9393c43f7dca5f3eb2f3cc96969ebea865791fef15b43d2b67352bf041f280e4046a3df38718c97e85eff35de1eed7714208d0f464de0588dcfb6450a8702541547a758fe009bce6adecb1511cc5503c6a7c5c6a9c2b89e566c7570a19d45b673f01d7222a3e9306a14a94d773ff9b7c2be70971c87862c37bd4f730f38f9f28769b912f054dd2796c68c794022843703093032d4c7f6f0ae022aa5fce74a2bdd9f723ed6b9cc3647e4d9f56ae0f2f50d3f2326f23a7ba7a85822c93fdb6da1224001aece5d812e28ea4672219932b10468adf093ecc4064572c1ec0ed712b1037cf148649baa4949be3eeab8879099934e350507c7db3c411258e89b133a9129cd32eaf4d183ca75a571df53b70525493d0b967639ebbb409de0cfbca05afa2b9959290c884966fdc7cd31ddd8b9ddcfe2f1217ab6465a4f28c84c395e4e94357433eb53b713c36922da51d53a2fe664e7f3a6bce17675029c05237b8ccfc86c878a659021ee79e18ee83a3007f661e401633b05629a5280114e948a500594df0febc028da2b63ca6bdf3914061777d1186c05032e03e5a07c12e9ac0fdc6a361131be30c7d032f2a46fb1757c7741d3dd0555398a2d929d740ec627293fcbab3da2355995b90dc50a780f6117aebe52a0f16389ba0d058ae5a1afc4e3671e4e228cff6b0fb2c2ccacc0eb131967036b3a78f5b50c5ed48382d1f2c6871fd04b7c3ebab3c6e2f47f0442f0a74e83446fbe45507d4e7b3ca883a0700d313adfac2dd6ac9277ecb19dd839054761e4fbff95be88493a404ebfa6575abcfe90aa418de5d5df6b666272de997fff54b634635dc5ea9e7ce4c9f7bf5e1850519366c72a0034e6e9a0a227d46e8e254e4a807d73d5e506c4000062b126f7e7c82d85f799194bb6f237686ed6cb83f7ac54baa9b0e2b286bc61b745116f95a3191473ece2db3f343e87716b65e5161e8b650b6e4df8f0beb4751057742a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha1a1ccb8edfbc33d10bf53d115b9c37f3dc0645a637638b14323ae30d6a1d557efbad310fd7f26e5a2ef0f79ac5cc14f21016bd7608e9a5c28a96502b328388daa9182d815f806a92cf18797530ff11398193ad9fad1fb1bd5852f4d63c9103dccf707ec7079859f3d98f6db5fa0db8933e4466189d28a0ade3ebe3547320530a032cce73a8892f7e7741522ecab76d3681c1cf5f3a371d8e689c744738748e75221580b2ded4287087ec3407db552f188184fa6328ce567081da8539b0c502243f752cc6b6f68e2062552ced53e1680897b16671ac4d8ec34621dd62a5701c6372121028a4859b4455b0ec2596073761ff0fc2ce11540c26e10bd30c5914aff2d517c7109299d2290fb9408acc4ba9c902002e5b2a5ed9b138400228881639ace4b602a681dd83a8cf4a945cd9c1d636d6d5f4440fdbdd770db2a6f8685d8d663f88d07c3652abb9005c39684840600d81fd1ad6e9b927037c870d29216700d27b3613f1bfade20ff0ed122c505f138a512d20923987d3a010149be611ac1c9a182edef363827f199153ce8db808a331c00f3b61e6c27d879c977d1489f0a150e6c4b5560ee0f14e0211a7d51600f17ba511a23f84b78ff8b4273a6da44c1b89c951443564991cb84c22ea9ca3aa5a5344c57aa3d3c48c731cf9594a3b6a66149365c095809d65dce10a81cace45926cf08c26c13c7edbf5dc114ecbf4ffd32e2691c224842c1e3d2895d81c912cdcf7dc3c9050a209d4c7be1eec9290619d098ec373389225e8dcf1cfe0e9869a1b02c79a405ee04dd34531abbc3730e2344b25f247d7a641989267cc613489d2e8b6ec569a905eb5534fe62dc1a672fbb7c1f7577522564510841801b5c1837229817fd775e44cc42648b63eef63b2b408b3c394d9d15dfa0bb0e93dae58937231b4241a384d6ebe1657b78aadfb72fcb1fd6e49f638b3d1cccf16cac6a7e73c6ba81ae4a3cd48252aa480ce4aa7ca3d82367974121d20e154678707dc278861fa43cafe0c56bcaa5ebeb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hf883f581bd0955e8084854555f5543f4d6e589cc47a2b1565933b48ae905167df03fb1add4dff760be280e9fa2176fa88842b83985f4167e49036c43622b58389c0f5090a76f08ab4934629c973ded30afd075b7031830e53ad72e3f47b85e6fe12bc36a36a051d2718ec4a2d4a9c53ed9417baef4ac9763f8c99717d246790522810cbab4a561278bb87190314e549abdb13642b6e18ef267b27b0f0ddeb156dcfdace02d684a03700996559ad90e9eec028db2bb8b1e3e62de36c34bc89e3a7331b8430b4670e63965c46ff55ed4ba057dd7447a0fdd8b28c79e890e030db44d4f9a7cd598f785d5666edb9ec3c785850664aef582b9a2db122f4172d73806d05b3665efdca85850a0562a618ccfec5a46048d4e6350e16adec5b09470165837a9d6fb0e89929aee90f71bd2dffa08ab00655d09acc3da71c6567712d1c969e9e62057063afee87e95043f13e36362ddeddabc33a099db95732d1c10b992d7501e3e011f18c39b09e5cfc6c1835a319ee649befc70065c6b8176b85ebf8f0286fbd5eb66ab3415c4e6ff514b606139b469e526bd17dde2c7c51c751bd9646b6316bce201b0bfb81c69fa9d4a6d55f97b9bba39ec48ec3e0ad810ce01bf1f43aa8417505877976d0adc8f5139238bb47c278dbb17f11562e2cc6f672edca7ce95318081c24b250978c41b6805bfe69ff53710601168039df8a5c8a8b8fd1d3f5b07b7a1f5de110812f41bbdd9021f1b7f6c8965726a4997f858f235187061da603af3698027ddff2deb14a961aa04d3148b0a5b7339755666f46b8585326c6b7498978d6e6e56408783bba01276ac876ea18817b61feec39c917aa6133919ab32274cd315f0e433af8c91f6a2a0ee4ecaaed3959fabef94fbbf7a875d0da612f03fbe19e785a9e51da11b7969b9334e61dfd2e8e8eb039155b4b994b43ce7946c03fca13fc6b8d03fdb2974060c1bab99aa494852fb5f9017761c1522cec47ae7d2eea1fb659eaf9104a275296d7f1132c9d5e2104597b0f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h1308809e9ee355e3a6664147954ab6f4a2e622c170e33ce7ccec5e3669710014e1c391951002dad6dfa3ea79ae08881cf23e13a01d27eb42714fc53fdcecdf9d8f80d0eb68c7b7be05493227d1065d6de8927b2a224369fa9254c9182e226dd4c82dc18c9204824f7d34627d80b826a465782fce8c1d2c413f3d4d88da62d666c46f1f1904091e7eedaf91e7f1a60b05242984231966f5d3fcb183675bd94ccab1abdad47f30f4f968cec06728a713524a3579f9c3874f3189085003cdade449b33635864bec9714887c185d0d99d36e839f1e4aa882e18f349bf7fb1511d68cb1d1cca5ca1d311077d0f6475392c9b367a596ce2925d7d02528175efd33d93ea408d7efbd7e0156a93edcc3c72bb3788b6570e10b9bc31456ccc57d4aaff3ecc66bc8f4dc093deed25a2d8da51e37c7fca964d50122a2f8a906c621cb70e1ce4944e0b319213a624293204b331e351adc7d9a5bfc5f7cd9b314522d16ce707a39e851b8afbd00f99c8d6b42901b90b79127552e075500d8a1f8490531348e81993e8efeb4ec1e556ba98dd38192bc2ccece01b4540e77d8613d63f06aa64a2a9d9f3ccf63ccc6b03db891c356438cb8e6f82223e0ba7d69f10ec59cfb8ccb277a5f0a7ffc9cbedfe577a00eb4e5bbe4a3019def246bec2ca0701fb54be8b1bb99ec904be9fb99ef85b117ebe0b74db6b26490f6bdf77cefef4349db95f400f8d20c5efa3a82e5506802d274d2e0e92a4c071bc01eca58a6327caebc8b14d18f914f040877dcbf2bb69ba2402bcc32cf2d1760a8b867f0c0cd201859d2d6f335dd0b4187dd158f8977b42699320d98a3b2b2f938592e7f5980f4a07acd866b0883f7382971a6fac17c1cfdbfdb3fc46c97f676f47b7850d25a3160b898ef9237cde2758e06ce20c2ca857bb37b95fd9d96b99eab5fbcda30842a517f3e169526297abeeeec30e833eb2eac0f6b1c65bed856a7647230693beadff1017f7bb82a4c7c366f5f731f6841676201fcc705367d2d7fcaf262ce7f61;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h42f24b3631115a76916f238f038a1edefb683331816ed508409426082fc8fd9cf686619a4ae8a7068f39a2d75ed32815f1b3b49865c9f7638fc16fb51d42fb5ac667014323014d069706abf9789d7b433b7968df0ffcaa08e4c25a9f89d1b54f8e3972ac44678146f893dcedf4ddad69492bb1e7cd3a7addc30fb0c87414a998b4eb1992ab72b935966b38e452c6012a2da1464e776e837d1b19bf30e8833a2dc59aad3c3c1317eee31b45605f2244a083477313cbba381ee0b2883bfffcb44b445867ae58e1fdbd81076e1fb8c60992c95f9453a11c9c164d8d2d3282d3ff34f720dbde63fe2198d5ede933612aa84c013f14b2ae61d06b10e28000eaf912b0b350569737e865138fe0522e9a5e007bc11107a3d47fbfb5b43cbf85ca42f7e8477757b3d3ede22e6a09068a32b7fdd3ed2ff716746f43667170106ef1a0f1670665db8bbc6cc502b2a1a86489374e2c36dfa4577a8c50a0ba65632ae98b6d321d0be9db98911ce29fbaad056f2a29a824d0470cf0209de9f448d6c3effb3fccad40b49a27a805cd202f803be32b9d071a9717859440f16be9ba9c2b7bfac4b307f144ac6ae5322ef2b63605aefb4a2884ed3c41769417a49116bb386934d5563d25a272a881abb33ad581f2cbd62e8ffcf1f5e3a9e4de55516548306140c4ae1c04898c64f48e840f4eec0e9824e6faefe433e11c369a82b95950cbf6c8c99b03559d9358382521382e5047db50e5e72a9db58b084d4cc3d24891eb801a26757f17df7f744a29819f5475bdc0efe76085f710307544f18a159383044ce33038fa545e28e4d5966d6a5ce65e21f824e5dcad022cd818e4143f1b04e59dc68387e15db4801552d3b6bedf976d4fc0afa535d55ee0c8674650d0091e5c410251d1ce573be5f76b0e693b558f2d63cd3349ac9d037f77b2c83f48ceb7e0db90401eb68547621093cf0ad2381c08345a109d62db45840a796aec276c78a1b83a9e7a1f8684698fbaa7093ca68f6414ac6cf9b3ae618eaa35dca59c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h2d9da2267cd7179469cbdf2be5889546f5484e83cc02d5813e1af088978f5320b9b9d24ee4ec17ac928d6cb6b6f99be09c25e42a884b5f973a70b4419de0886e11b38b01f2066d6b6b5497fb6b82f9ecc28b4286f5980e70f1d29df4759942a0edd03ab3c86a8661742c430b717981b461b1a3feddedc505fc27cd0e42dc1a8a64477d7c97567d3689252ccce134b3406feefbad696dfc83fbe4c51e99b1479b1543302d679600a18f08f06d0329ce15340c98dd588bf5c54c66555086f3ba30607ab65812f66d5f8ec47012ba6b046177b98d7c9769d32ed590d04db0b34345a028a194a6c15cc65ab6a76939cddad6686de76eb17aa6f80402c240a8c52c9f40c90135715b830dcc3c0e1a3c33d9995e1d33bbdfa283401f09498231d53306f7b723a1c2448f06a75723bbefff53281ca65cc6ffb3f37b9de3cfc0dbb0df18920c977fda8302de45dfc0441d8a5c155acb8b860556ff14d879c99f80bfd690a8d2e672d5401641d403fafe42b36c15205757b8570b1bab855c3453a32e468b20b9c1ff9eac4d1b0617063f3c8a75155f17a835b2d9c3ac609f4294c08ca09bf16781cb214809285a1c44626090a51571af660cac0b13906322dc8e99631a5c60e1c2634b4d7329f047c8bc581d454d9823b40b0c9ff7b9688e007b15d8275b8191a63f8a99ccf5c5bc2a533e83e19aadea82219d109a7e807c3cfb05ebbe2fa495a63845b1db7564ed4678add8c045547ee2f989d48cd482178c18fc24c9c612f02cccf0bbbaef1d5371f1c835b38d7e1875cffab1cdcb726ee21f9e692081fbb580c66d6b31de00c791e82a8fa6d267e9de14936d3609c5927952b6fbfcc8ebea5438100e47f8404d951cabcb4de8c143cb2250c09a4c4ab6367ab5f8058ef0c464fee58527b1b22d80b3beb5b296b8179d27e7b97e6f7370d1d0f860f28dd879f7399e11aad9a11abcd4264b9e273d9a10b59339f62d7cb701c87a57dab290cbacd14d56369e9f6f7d0a9d15f82f84f3fd9e1cf98df7e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h86134ed8623fb27cab62d6d4def6ee4555838a8e21c31d951820414b36a40aee61404cd8982dd006c5e97e188971dd90c9f26c112d263d6cc3a1fc1117d38d4f8956668a886ae8b1c04f8bd4b80e56b7ca2b496f76e3ba55bc3f5df0fab7e9648938879d0eeaa840a38e1bcdad0195b1a32bb82eee5f0e4939cf626c2ea6eaa7bb056fe129c7a33de4f721f462540bc7d129300539705e9e470c6c42c7c6b574eb16c5f50e23a727b99d2dc289236629c2ea6ac9febfad56b1ef9e96ad948bb34d8aeaefe35c3ffbc8db78884aaf25199ddb04e27526a6544e965cdb10ce6dbd3825feaa56b08d6b028d74bb9e24e20aa9783885c14c912216bb745f0efb4d78f95739b9c7d12390122cee4e1ba2ba127396cfb1a874e0e913f0978afc68849f15aea426be04e368a48a6022574e6a5f826d7215facd91e958bc242078f9fde00d80bdfd8336e3a45d5b07e59577e92fee59ad420f373d01db1d6ddbe3a193759529b38d115a6d21e9bab06148e6b3eef993777481f7f9576be4dc946f71c6ea0cd52466d8afa08a25dc57cd1eae84209df5fbd0a1bf59a356468edaab8ace13a466b0d552020845776bb6536b92ce633c317a62e5334f23aba74dac63669b0359d71ab69cfb1578c4e28dc92e05b6269a0890377f122928fd7ccf0d499f46935cc85c873b5e8e9b8df61584802e7505acdf07272672bd7aad6d16cfbe501ce99f26b3b0117fe1239df0b4db03e56fe6e1ac3bc989b5790f24121577f0bfc1afa610cd116bc2f8fd30444976f2992d2ea58f2a21e3441bd09239b8518e7bee070b6cc1764aac0c0c583fdebc051587b7a682cbd7c5de3de8021a80d7696e50f42929e09bc664965be1074cb21b60a5755a256791cb3610baef2aa4569d36e8e9d2215643205f5e7293d958dd0ec39623662ac14f471999804143145309972c9faa4fd2c6a9ea29f958345d948e6e610366e19349474628b51e57fba77d2fd2b99b8f1c8f4ce45058654d27a38a569dc6900e7664be0d42bee0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h20ce3f154a4da86e31648fcf5871b2155d113c0a0b168a702b997dbcd6e12a62fdbed914e19b6a4a7298d8e4951c41d9d979ff4b38539aae74b7044996f2adb3c601b7e2621a333f0294d6d89f73a2388df3976900401a942e0edb4a31cd859399c421f2494804b4ed1370bc9d19fc39608a7f9021922601da8a6c4f161f0ba76f4f9fac5c02812533b8c83332ec337778fb2148e9cf03918655ee0050c65131bfb17c6e44923ce0a469e3bcad62da886186b171a7373451080389c729966375f63ff9755011eadc9896115a650bf48cfa0e6b83ebe8eace90f2e6d3465fa7b279867b01bcc8e128faadf420e4d0c1e8ab54b8646863d8d20afe5611b5959d691e226f57a6e99ee18b695f496ad565d73194c238ca760b00675f524dd90b891bfb470af33bf86786fea277e1b936925fc0da6b09aa2f395aabba38251e2cb04a7fffd04b81f7cfe1e83227d73315cada4a316aa7dcdfd1cec0f441137efd2cc17d66f7e2dab965dae49cb24fb3cad4d268da7d3856fc76cb6dd62d421e94569ebb1f4d907bf4058d3b684d0e0f5d8f6680c712a94a6e5a137b7b931fd1aa247d7fe6741ca8ad683bff3a63105f18b3528bca397dc38e070091fc4cd04f341267064e8379f445b7fec75f2de751aa5cc55de39492b80ac57c1c7c7c46004df8a7c2fdbf6e0494b8d18c1390dcc2ecccd514f4b2af2ed670b8b78154aa09eab1d5ab0add85c4241e24b07332255b7e3a371a9212a10338c362fda565d18a9aad04cb7b4b960cf2008ac734d5a7229173cd99f0a32a4d04e25d72b3a59aab4ff1ae3f7deebc66d342ae494c38d0dd72f1efea42eb7ae0f476e16b78bdca7f59554f09cab00199e90de910db174adb0c01715905680921be13eaa71bf32a436fd2c08663ac1861a9b8b4a2ae1e84d87348e498923770824490fe297967d0029d22ab011bbac06bf8b58073d18611e24a10df9a2b981328b2cf8793886397019fbd1ed81f0403e62c2dbb9c9617d6ffd821d8b0cb1d067ca37f311d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hd215b4a3684f496ad8fe2b667dc31135bac5906d375cca808d50a68081da4f07e6516866096ba54aff3b1f27001f0fe1d930523a737bdc1b2dc9d52a88376fe81b11b861cb9b7309f958ce48830cd0c69b4a5da966c02a19a474d63a2b5e5e0e79b68d36f0036d77b34b26f90d319fec2ac9a5a8cdaeaa4c34a0a8990c90cb88893da0704d101cf925696b9355e8579d04f8fa6898956ed69c20fd2e7ee7ef68869484ff24e014e173960062e3b580516326a19acf2093be7d60cfce9869d814ad3ecc6b4b01d7b9bdc5e8dd784115a7ad551db2dddac74186eb011d037e89ee9b0da135dd45543d2e33a65b1b917dcc80e0c24beafbd104db6bf352a192b37497c2f17b701871d6f219a273d3cc6b355cd997efa344e43551d6ab2a69f221ec19c5975e8ede5a37408630044443bd2b052de5c90820963926eae2690877201e5b4cf3d5fcbeef4006604d51f93367dd43ee04f09a2af2a742550082426c375560abfeec38ffdf9659b5151ef8f8719994040d016436773cb7845063d609f573fae561842099fe9caedcc17a42fcb0da707c132c06d4a39019159fd0331e06c23ef9d2e2cee36bd28672b475cd69e770463c434fb40deb761230dc26efc900f7273bb4b2542c0a7108a51eaf48902e8388b75292ea4ff521536d44b4481c4e9a0bcc15c3e0dcf49e78b4a37cefb5f22aa1d36e06a6e1100a619be19e97466f582c9a67eaccf6c1b1d646a7c0ac192257ce2a1c07dfb24f427e7ed3eca815de0ee6e03125c3b303a413f21e3e1768febbc873f8d3ac1f53e85fac7770638ceea12ab65ba5b6a4fac94dfa3ee45940ca7e8b45698ed13370eea95583dd486ebe19c078f5d0e29e17b629a0b29a252b053ba225181776839a1ae965f90ff1efabc10c56851da35ec3cc2448ba10ac1754b8176b7073a1fd37bed80e25220f8687cfbedc64828bb4ac89c8530760751dce01a885e07a37d96edd1fc346ba083259c56ef66e42ba8875d9fb71494eac9db3aa5b8753ea6598eee3a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h37acd547463df61fbd5591c6c22415164265192b07f4a5865601302f7c50d53cce4635077ce9a7a3efa2c02a2b86f5b356341b61549cb341a8d2fc4d7420990959494a1218228499b0d963542ff82d3a8c0e89e03881072870da57790b1685df1de07fc22a3baed069b7759db6d153be6c4be61d2169c132a2e6737a953b48ffc38b75de99db34a800756f2b512876f9a1c69532d4573a9fd4a891e07233c95f641b4d2011f2f4be1d5fa8c9d1642123b0147a2d5c2ecf6f1073d71fc278bf5123b31d9bb7456088854f30d053cc24cf2c01f4648df74e2202bd0aafc1f58ec9880cbf512550bf93e7b49ddee435d69f61521ac800598607eaeb963e2981d5169ae051ba73aaf8e48359b285a5c17c5d63a290e25981ddee30edfb746a987b0ed12feef5633a7488df62b71c98b0c1d8af863c15ade4c2a68a03074725187a883d76601f26876899590934eb8788dc5f2ae3f4a4256dbe8f5fd54f4aff614f721152d632038805a0e208a32126597566d42edc97aa6b373a3f279296109977f6ac3b8bbcb55e1844f3e590e5707b19ab17c9689ea9f3b0181af004a6945ef8860e33a70ad67942e545ba48948729ef6f38b6e94f21a07f40d6d1848a4a34a2308a394e67e888741c3eb30d0657a5dd79abe9867deb4154a27786bbf746880f2eae82de5dc115c20097e18eb50dd2e42596f8219aef7950b50c07a34ac78845aa30367e55f5b3c0227793adfd6e55886d88a15a313b3c670c8af9e29536e96bdc50b3d9b45b2e56e9023d3fd52aabb9fb6d9d45874d9eb5380ef83ded786cfe09ec49d3ebb8cfa9e15b3d27fe9f4d4f0355dbd5ce3663e534f3bce656bf3cb12a283ee38280e75a7ca71c5908bd7f24c949a304631ae7ce26dd21784c499af8afb6af3cb1eb2d57d03375e35643fe290ee669b50e84aa448c8de00ab0e7f871e534129489b67aadc6ae01b721e1dc015735c1dc5729a744b749b31b9f21acd8b94e0773ce66bef5aec859d645f3c73932c443ce2149b61107db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h6237f713b1a865946de298b42c9183b20d43c8295ee6da819f70df57e718d9d7766cb8e20026c1bb860dc58384d15867b1f1cd9d9bb7e7e9fa6ddfd1786ba93827df39ea4eafdbe0ff1e5f21d50b15bed9b0f77f8d58f5f3578a3bf6b159308ce6b8990a2b9adc7b5f154b363ce60ee95b522e56663b7a93c9d1120ef044602a4363a639700060a18249d9b8f8e8181128c88509b8995828d35a1e02080a453c7b13c4bd14e1886bf03384ce6fcf08b0f8e198223cd7b509cf257ca0d2308a2e4847a7ddff4153aa89cce136ec33f28ce3dbe489d71ca27225bba3ac8063b7b1c26c965f70321b44e0b9ddb73ef3d7d2ad326f17fe6ed6e0a8e233012238e3c3b08e28421506f29177863ec3f5340d3e5c5e324b4148b726186e2e5b01060bc91b4b89665484ae66e428e37132a99617ae2bea44c8c2cc66ca0b95d5c67cd212d181a4297952f090f656814c0d07ca8f371c6ca70a519cdb138a594e328e7889653bf775eb6d1b3d8b4258ae14a8383eee68ce2ec2dbd9db87f0e46ac33b95bec7f9a0d0ba7ad0d3d3d6da7acf35e3f132547699991a7bab08dcc4bcb4a71c21ac69df1e4cfe75b041fb043c05a69b6b23e80ca7d7f062779a41aad0c518085ecdbae9b136d641c24a91c4a86654a4fcc794f343cfbf08d5b2ae1d05f557648aa0f3195e09028f7a539eb08afde9b1d1a96913c334a5b17ccfafcdbb115b56e803a41f477b59b8ffa1b4a3bed23f40fd024507211c1a84d0143669571db01b6de7716b08a867a75f5b88aec0c3968bc68d7ab1f1abfd787bf864a3432d2dc4bbbbcd34f51da75e87d6a28e94e26690bf25fcf99a056c08ab0a66d9d8028d0f0db7bc61a312918598217be4b78b8a5fb18f29c0697ed64f88fb37461a7305a0b2c6f4254bba022532d7530257547f2bf6cb1204196f8fe5ba4c88e642d3215a978f7e675681fedb47976644e5962cb384dd777860787e21ff6480ac4110bb8ff300a001d3d8ff6c2ec8ad373900e1288f75d62d9174897b2f26;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h54b7e64055114bb01d599326c5c4a1d3f96d03e2dd34a17172376e93c3203678ab48619df4cc69a4cf5687643027d328bd202559cba44bba765b63c4f0a2db80f5f1c1d0e963fb05cc3aab4d96bfc5491fd44168f90ab3bc1ba016f7e6ccbf59c6983ee21c9c4221efb35ac0fd89b283bffc8de84ede346d6ffc4f0afb51f45b05459eda70fa6ac3785f392bc237941afc37b9d8e30622cb1077187f3d8aade40ff2c1ad85c06fd0f71a68d3ca998caf70d54eb66af2af63f0b35ae3b9a1ec819d7f990c1acc840ba36c3a0014e977b1af0cb48639b411a2bb2065af9630bd85fb6e5b0f20d4dbea9046d751263657974379de55725483e037dfca63f902639fa37a340fa60b104251b6f22b84c024adc5dadbc9e681ef273ef126e004bc1428b6b5f596a4cdb80c89ee0ff416867d50320e6241cf9c2a7f090482386f428bc170c03bd31d25a9ffdde5006768cfcb7de163b7b78ee78ae32e85600d80b32ab69ad3568101f0f6d85217e65f1e05842c07ecc90eb3fb265ee99e02841ecba8a55bf982853067b2a10cafc9c0bdc5b128a2c614dfbc2894e6df8bdd5a9b60f1f17a539c7256f1957e36ca00901b19c977b9870ea3ebd01da8d396533b71c226cc6b4731a87fedaeaca25059ee956f5edd9d45011709e5e6ad65dfdf0b8db636e6d119e9d322af9faa6e9c6d33afeb4be642f1a7bb2971c4cc0ee7292764bd2bf9aceb1b256b1177f3c41695ccc18e8e3dc9e0918d6456fb66d37cc2af79bbf2c68dc8a7fa1b58d938337eb3e05e71ffe16a5b239247be9b0b456954e369880dda95e624c89d6f306812584646533600ced6404122c389a4bc8e844ddb3e4848183e604ddbeff11221d21099ccf72516a7abeac96973f6dfe8083663e2adab3e4723843fd0b1a4aea06279ab852d2638b7e5994462074cf7ddfff6d6eeedcffb18cffd6127fe70079e5ffcdec89d58e0895410d4c82d48140a2bcb0881c182e7ee7b4b24154c89467d3da81e14a5867b97fb376d41c73ca09d28;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha80bf239b95f4028157d1e8bbddb2ce69a72388b92c6c4355177c5605376b10961e7f62099200ccba9969abc4e1a5cd401dbfa5c6143cdefe36303ab3241602d8c020bf44ce8350c01f0b57acdf0c6c1f082c07bb9b488e5d8e62c3c5f23a172c7c26d7cfe40728dfae31948c809e86239555b7e928b265352bfadcd8fd73f3054914fc52adc2a775cf9a9d25630221c277a2eb3ef07010bdf409c24edb3bfed251771cecb5c87c7534a2f1a97ea41b5e7a5ace4204c91f99fc699ce8c45d69a8459acd8264ea7207ed526c3f3d56073c21014c8f79a7e2d406d58a7f20db180893856f169fecbda3dc91d3f2792a95974eb0dbb605caa813e38223faa422d2060efc9b7e7fb2eb5891572b392dd782424afa8f1e99642e4b69ec1a54d7e2d569f599caf43e885b4d0321fa53030601675b1db4fefdb6cbd6eb2a32979b5e7fccc5f7b82e276a0729552c6d924f34ecf72812dfa52af429bf6bf6a97d499a6f64d0d9d52a618b223fcaa332c7c47d851fffdaa410dbfeaf3db2caa0e4ee377c9bb48c37f2294ff2c878875e15fbd46eb625b0ac129ee5ee6aa4c82f0d11d51960fe18c5da510c44dfbcd2b294555115a0f1b3d9a530e75894880c0c5b3fb4a0b14cc1ccbf9c09e7a32aa8a34bc2bd08e90fe11bfd22fc55f3fc94276f1ef7185a2dc945c6c553dbfb00d98fb7837b770db57a5fcefe049ea838cb48883f5d4be100798b0a59be7ce2d9fd03f164f6a96bff9809f09815a6415baaaba00888ded8da83da751daed1af06ca361ade16023f837d360a054c0581050fbcf3c9136cabbff939829adc59c6055ac09fff15611f780498fb7633f413d30cda53db959ab0d0b1e9ae180f4a0b6ac20adb35700976ddf3753dc8bf08370ef128f5b2845cf39be78ede2362908ec0745a80f5756e841661a370a827b7ff4087b8a47a2d9c1183da3df9fcafcecc64b17fab26308cf0f05e7abcdcf936cb2a7e305fb4ef848e7b9ac19aee329451938389ccd53ec9b33a9367ac4524aee71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h623c30eb3008b56cb1dc9970a8b43a887f453e1ebedc652446ffc793e09ff4995ed9171c498dad489cffbe38f00b9575e517eb7e603a59cbefdb77f4332b65b330d633361f0aefef23a3ffdbcf57a3e4560886c7c2d51c893e9825df3ca7d07cd77530c07fb9cef3c5dfa3c3662a50e4e66f892183b7000fe1fa3e340c7500312fda0a4f37165a11102270655c9640ecb2728173331604d0ff94c49f745a47f4c422d5791e4ce7bf9a652626dd14a1c3f3da6dd3fb3ebd0c58e4b69a4300aa391da2695bfcd04711f84628a36aabf3f4b12611fb244bdcabe039093375edd907650c5749f7501c5db9e1c8e12c1d9e3896b2dcb97b5ee9e39533b78853d43d5b0dc779c75534e6a94c84cca54781a36a94386de592823a5f3ac659e9cd264b4e0d538e0dcf75a76bf2344ba5eb69e61158c697302d8eeeefe2ec8697cc63a4a00eab7050744b4fda1c3d87163bd95a504824117cede2cf0c950c1440a442d5b11c0bb2397fdd04a683afe532a9aba4ebd944b054c936e2c2ba7f54e0a8f9480e5613e1bfbffe7582cdf74580a13b9be010b7bdea0124c7aae01ca223dbc825ad767c52e9e1ef98c45d63ca5fb7a0d3d733df78c5d72486d5f76cb83e611c5714425f1d8a3627db3aaefc5934c07bcaa6963fd01e2fa19f952dc6c7ff0b8edf7d4c3acda55390cef25c7acc504a0a999fdda2adeebd6c5cf215527e7c146b0bbd472bd3f247ba37b0f5a1acf00e7328ece65b8fa5048649c5fa179d73234de4618c6df216cbfc760455fc3e13d89efefa55a3414b4db14c607353bffe466afc55c9f30a0e7d893ff33852b505bca015145bbed2ea653b01df4ba196181b6ed9a7624cc90ad6f7ce1af41147684cb04e666eb50b1c8fee358d044257fa86ab5fea49fa1020fd3813c0890ced1b1374bac3d2f109825a9eb4bc776c8099dfe0cdc94313b82636081c2c5429437fb3f7f74d9be231311ffa073fa399d01cfcc1093d710683ff336d626fbc38852b8647438006f8730ae7e97cb6f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h84c73298fe0001e2c8ff78bc754f132269019ca5a947be44d5e2a7d89e2cac8fb83de5de53b37471136ab9eed598069ec88b0935a7497e3af3ca3e1371d9e4ba29c1eecf86be05dbeadaa9b4e7b6f5d0a639a5a3501a3bd6818f7b55a3d2fd43d6ebb0b50dd97d0732040cea6dce5ca29fd15300c04673db6add7b098da671a391e4d994791c241c35720f5b206e99736be9d7a7955613b6289ec67f14e9925c30cd04996ed3998ebb39799854cf56099b8734e50738db5d4bb0a5709da8e2f6fe2694e086e979d30e926abbad25ef013eaee8acaa3fa68a4bea667ac11e78fd4b8fb805b83bcb96d1bdc5f63fc640bc0e08404379ca954349e42c3828206884b1180d9d41cb9b5ea914cec3d6d52d488cd6920554af875242b219a5f6941422a943392a5f4d510506efe06bd0d7aebb699dc8199535166d474737cfeef03c34b865f190f754d5b4211cf62cb743e286bb419fb75bf6b2dc094b3a63dcc0751b0285e5e6b82bfa20153a234e0aa20bad420be62a6b6bce69a5ac3af262483149d3162dafed69d96cf0e74cfe69ca75528983be71d8feda62643b4255634c681024be86b3d1837a13f833b51497142edc6e575b37e92d01a6d88c13a4fe002fda66d14fe0b60ab4d8e336ce9844274682435d7dcdbc88af8719be4b7c59724d3ee7d3786a225b518026fa9bf9a23253c9b9efb8289eaae2f6e7e9708da6593f8ab72fb288882c15fc9379d9232c074fee981bf180128e0ec4e701deee266c93016e4a6e2249578cdef73a86068192915ba32664b10f3178303964ee528261b318c9b418e15f3432eb7e133c3d55edf76e76a8df362d967591d9320d05a612378c1fd1da604342ce31a420f59bc7c37d635d2e6dc98bd7a4db9781aca5c25a53c9f2411c898389c6ba34bc25e63bd240d846354a6fc859cb3870660d74c78da869cb7dfff3569bcb32c49deb3dd6eb5b4c0905073615c42aa9d4c990e44ceb4a6b2877efb722c2e2894dbdf73a4b55c1d67ed6d8cdc8ebd00041;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb9bda960e4f03b1d9ddf08716a3eafea51938e6aaa50c2a10ddd6ec9b5a6df7cbc4d850ebb882f52589bc67d75b23c62bd6f0d0840f5437b746349727ba9b7d0fb62eabd56b62dcc7eabbf999b5a30ea1a9bb3a8473fe49fa67efccea1c2b64e3542f00f384456f65da64ac0e7176ac21ec91f89e01694d8fde960fca4ad728198bcfe41a6367d5e10b920b6123d6bcf16d6cfc30117e420c2d0fe8237b02254b4cea367754f2fc43b5ec22dc03ab028ebf31e7203a64c53d5d1c0f179920270a729734b4ec92641c9b1c5dff08196a4a6c0f0190af9f507960b9911a86e316739d36c7cbef6e08ec5f3838de2c6b464481f820ac96da4f8caf86b30e0b3f5c0916f87f2a48002f70d9f5af0a5c5efc76549efa169c59c7c3dcccd1ffeb7860a8f57e6952b43a0c43712a9fef38cfe8aa6e82da612116ebd23265c036ed0b1930464b4ab4d442a099f3d0936f7e6540b33f94df96027dac18d7d5e05d5c397e63284ac42131dc302e723b5745a6028fdbd6d439207f61f0c2f9e6abea70b31ebcb999b61986a935d52d32ef6f6a989486ced6551971a647fd72cffcab50bcc3b338ce62a32d47224fa6f34724c0836a7a5bb3df41f4e338b30a876f7451fb1f7da664852a30995e295a9f695a4e34ce4ada1652abb42b6dd5a72fc0991e79fe1c56f29359bacc935bf29dddcbb34623789c6ef6331219802fea7f0a956e6be01490ffe1a0bddd73726d99ab8b39ffed4a67e7c2191d548c69cce8ac4ae791c64ce9064dc860c41280e5c6dee1972d710bbd3ce9c62769ad6d486f2b166d94217f63f32e80d18ec70d1de2329e497b6f04d00252ed269f64860be2aac3309e42da40c99a96d72c3c83bfbecabc635926cabc482c50090028156811d1dd2964662e668c0a1841c69a4d6030805ceb21053ac051f4443603fce3fd473bd20199237fc1c3bee407af89c2c99f04419c474edb0e52cad783a34554e7fa216a2bfe92a8ebb6b7bd05272e3180d081d4d9e275f55fd71a73c5d5ce818;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h916bbd9c179abae47178a4eeada64cfa917224c7e45620f6f2c2c8032e3bea7f9e8962060ae212e2a9f8a1cfd2ba0014efb2560d608715df65352b300869f9a2b3f47ee89e894aed69f00a494a4d7ed83249952c97de302cca1b46a888cef34f0a446320b2df9eb04685c54282f8fe49b049539c3f4ccd7593048a48086df354b1b741e32b547be76c84c0728d0e3dff4c8b2e268533d4e80b90165a4178a2346b9489c733cd94be2c314d9fb54c259eb28c9e5e8bc75a87fc245e0d19a2a69fe90f13b1af9b2da51e5e496824536dc9ddeb5e49ac659fcc139d1115e0c1ab54116798265a78c11668f2f97d07b3472a6cfc9e6907db2ad65fbc2a0d90c587d96def5237e644114a843874f2828305fee7fc9a5c4ad6b4af664d9eb82124a19564d7bc0e8ce96ca94a2996fcaa194f7674792f35a5a62d09255a15e0f2305444c7fb542a588ca7e4868cdc6a3bcbacd109daac2bdf1cb5c2b1ea848708f9fbfe686f08a1d8679ab856c2b7c9e4cf1070203b61aaf8a78c730c7e1216a3b68702460d009ca97227a301fe13ba1ec381d95787772e119f3ebb7caa2b1a2631a6dabb630eed0be68ad6d43f60df95fc105e4c0eccf3505199079d5b50aafcfc3949d7c0d05d5d66b5210e8c9490de426116d1a6721bc37a052c96f10c0dc6d56ef275c63d752b0b3c4ccf91cc5e387d9eb85a5b72de1989bdc1a33615fa756f0ff0ca64575cdbb7ef9f295fd419456b6d54c16ca74958013ec607fd3194fb6b3727f4243f4e89f996a4da4a68fa352ba3ac44a980c97ff61984a05e3b03ca4a028466bbdccadc27e73090ea2699454c7fab1288ae2c460de32137fdb3709f55b0ea8cb669e6059e609259243410bc065d2e98ff72a626dd8174af721ca42a8e5b5ce71d977f76325c2282f922aa5a24879e3ef6dbc0e8b03a8cff0434708931cc8f65fae6dd89d562d81b7e6956e63cc6150b82b736c648d30bec6af177c13504774b689580a921e1339320933f11cf193a80f8ed02a8ab2753e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h90c0e9b8cb7e5fce7c2dd109c921f58fbcf86a4ba0cbc36df70cf3f88f7cbd82eaf640eee79e9e89321373a8e6506349f178d95d835d333a12b3840bb1a658229e1bf00554ca20b5b44db0d476e9226b26796bf29736e97b5c8d96c600ab886e07b978426f420cea0b07133a901ab515c1f9e36402868a2be502ec71055ca4e25451247a53d69100f8aa6d6033dccacd2c7e1e613e971b361f81754f2a2b1240c85691caa293571549da687e8296487b9db342baa6f32ec408cdb30d12ecec8f26349d0b859904f778a5ca75ed1586a420dee48f2d07264c3d03639df04659b32349d5d79481e4eee66882d07b4710eda4ddd8549fa4968ebf59abeace597682d6ef92125ee792f45cbaa23e020d498731451115b144c5a0800ab6e33a088c6bd3109a4e346a36e2dff6a586a1f7e2e4bdbb2887bc50f1baf53da47278e524eb3f255c74ef59633cd51e80c0112f355f32d0817b7af735392cc74902808baac4dbf854113401ce50997a70a0e61c18adbe5fbd628244e773df87aac258881cd6791f5195d42ad6c875fd35e5a332c0e3b94a2495b62bae67ffd45757f58a819b179b0f3afc38e55938d2a01ae42b7fe525b18e11f2dd45fd8e6f49902db5e71578794c7c183b27c3f7a47b6ddcd1996c161a2f2909edc3542aa71c80a7851a055f8c0125de7bbeb21a7234f3f5c2b66b4c0a5e65138c9f0b6d380f00faba1a546dfc34697067483a3b81492f53c331db1c1b35de10a81713b7322cedac159602ada8bb7d041bf9daa677b848b868cb857488e82c5ea52dcb303573c3650903dfa0f898a70a35cfd5dd53a876de2f43af2122a9bc938c4b5dcada85a602e52150013447bc9891d83126cd8415cc7658b04d9ba7b647664d9f9daa2cc9e0d4200f9a9e29bcfa5f6bc2dd67b88b74732bf01517738d14c01491c8d803b89b138c866bd66a7e33581feb1d4d6f6a484b6f46d43ca63e6e3d53b9c2b2a5839f351b71875b92aba1b7d22e789c900d42d97e6f269760c16e2a19a029;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7d683845145cdfff783a93da9615fdb1dee89525bb1e744d3096b038039eab5aa883d89cb13d7d7278d8a12459e1cd17720d173e2ce9fa0a4a54c8a2f5118bea40bcea2a01bed7b734ae62b31ea2569983ea87e78c9f697f21a71d325bee7ab4cf44b48ccfcb5833e053f8a4c722ed0c6cb02de65c35754ca6fb9b34e2b12a847c9a1f2e3890ed656fae348ff410a237005cd9502248c6cd27703d472f906469d7a1fc6c894fec64a5988bac813cb9076d8df49a02de6c56a908f21f2e4a5f36291352abdfd7784e30f43d577888e6f70bcff1c929cf72d4eface2556583f77b1d05f1012006fd6147722260ef116cb58b85f307c5f3c683bd07c5563297101a31b7c2ac60f5ed70234a28c97d4fcbc78373e1025e7d77ab305b7a71bc0b875964c72a5d37b90796828af7dd39f56c150ce4903266586bf8413602071d9298408bc39d70bdb3a7658442fe6c5614fe78ff780246be41ae6df9a0a9c2b82a1441b3b9b0b5377392878b873a236b7435fdddd625abbd141370d9b5c9084ad1ebcef5021906909204a1ec380e73aa44f464b5111c1c072aa9d8f71552582c7cf3a10f207692e306fff609f91f7ad45473a77bbd2b075f6530c14c36133f04163b740941875159aa4d5ab33d278a3fc6090382193bdbb79f7687867bf60649e984c50a32651d3c9516a3334f9075607af1240224b610acc97fedfbf892508bd39d45c7b025524a88b72e6794c696893323f67754e46b884797d8904637da1dd49c9520bef916c5ce0526640cfe974702e60de8632eeb1bc22cb221b5c66ba4aadb1acaddc0a4656426492c55e5098252b215ec404eec141550887991f3f67dc11d0f7e377dffd8c0668af75c197b35ea0b6c59fc677a8819226f511cf46cf88bc0eb1068c3615dc2814c389867a5b78553f19bc3bddf64465c74cf4876540abcc21c7c332d9c6d6ba20b3692077ff35a986545c00d8ce45a3b0d5b393b756ae64792a487aeff7f53749ba8fd0c3458d83c99ef4f3821187568c2fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7e1be6d521d90ac6a3019ef102bba766c913aab8536faba5a4f52189706c6c643e2e8494f2b5731657d324cc6755371c2ab32eef4a806a7020315ffcf4a6a271e9d30a9e9f04f833c9baca76287532c3476b10f60762da4e944a350b87cd4258e545a37ccacf7febe08bed66366a41d6c5b7192524528f26c0e56f19720f41d4f5b4097f2653739a231ca3b84d873090dcb21f3ac90e87e5e07a0bf9d601513c4c48044f82398ec0956645dfece0dc1a83781fdcde434374e19b9a7a58d92624d025164fdd3efe91f541e34062cda39c48808874859a213621b2c4827f18d79e54805fc6461e49764242120dcd26dcc4a05d36c0e1d8f23356b27e7f06c1e817cbc4446493d5e7c2662321fb4efccb0eef661bc39c6902cdda68a9c5895aff1502262e21dd1a6d8ecfb63a0b4cfeac60279bd519201ac4873760fbdeb5ad56ce02ba15a2d58f9ddf4d576a9e41542c940c6cbfe533d08b2ed946cb3ac3088d1f9f6c992b1e4bb6a09e1fa567561e05ebbea95d9fa7d911f2e3a2a65400f322e2b1320d06ed4b8991d586da01df98933bfdf220b12adf618f31f2bccc122220ccfd400dcf97a708a48567eb5172138b1a063add51d7fcd1439ddce88f003a30864afb6b207f8b675ca4cf206fd38c2b79549f6496f1593d90baf12be644c08c7967766a0cc184b28d750ed93afa55549b0d6f3953a33b4634f9ea04cc49eee2cce1245aee3a7bbf1fe67ab4186645db42052b53cf0c2fa83f144500ecb6962956d97e0c3fb7d1bbaa9384bd0991ad54fddad7ea553a6a102b35b0259686120bfcdc6050637cbe5003fe0b13e15c7800433a8c289cc17d970c7164e70661403652807aadc45fc0a80118b12d0be0d63834e269774bfb4142e60a988efbc4a00ea8072bea2ebd54a9a954f610bd54d5f5816b00b49cf69c31d46312f0332eaacae8c908e17bcdabbf3585452edd27dd7037f20850d87e6d05d40b91fd01eedd575e958186187ea0f90f090a15efed73dc44d7aa55513efa4f0262;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hf752f89eaa698eb6f95bfe9633755cc8ea87c23da0d711df3550f4c3b2e9b90148ebdc41c803cea7e5de45bf3b78651c48af20d5f97ba7e5283eb5b87dfcd3e2d63660998988e05e0e9136616bb472825e17ca9860819cb0c70436eec2b4284db7d5c23b9da2d73da2535130618d2886349fa586cfdef5fbbbfa62bb8545d68539c811debe422acf38fc05764b5cab02d2e3f62c92b163b9fb6984901f86d7dee4646275e51bc6797bf126e07958bae8bf61a2f1a9ba387ff8f84f3d0a8bc250bc1bee4dfe6a6f7ec5dc2019638830ad99cf3b77d5eee948715c5af448f088bd06ff0180eb59ff2f7e08a6def388d51619dae525376fec30110466aa845441f1d8bb540e9e755fffddc197966d805db0651feb074ae66cd116abd8a6327b905424e8adb719348790a557dcecec6a900dc5ca60e352c220583500e574b8192b03f357d2478f642c210e8d91e132f53addd97bb325fc0cd93bf662195abc0a8fda93754c600fec7d3907fcb4e3f6062a737ffe5c0967f0f216cc9f3262e6403aa9c5e10c55830f66b9af37300b69c07736882ff23fc65bf041ff4561dd2282581d6abbbc48de4239862fb31a6c45f3ee77a8e3385e5f51fd0f7871ad4f6f9bfcab9825b6a483017be2f246e2e162ea57c65f2e119b38b84b418c53bad0683476e83f59efae57da285d161978e69c6f02c2d3f81e8ad45e87f70299fa3406d4ed5f31b9d33da1dfb15b5f2b31a637b9d5f19007877f6c6f30ccae905ac2eefad55ee5d044e0f47e8309ed818b9a926038fe48969d3b4e396d21d445ab953be357969ca3af59ae99e62871130c363ee7df7edbc4fe69f970560e656e350268bee8a2a084394e6ef924de5853597c28869bf25308249128568cb99996c5000d865bfba952a4e351b67e737e650821a96c9ae3df06de5b359c0be5e5408384db80f2d3bed2ec2e17d64c1c87502ac936a361c0e35502745b0853acf41580fb8819bc3af467a8f5267be92d6cdeebf2985b4f834fad005671550ffa91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h58a0c58a7bea4e9f4759da9507598e728b68d7847744b5bb6c65ba83a82e6059fb39fe6c502ea3e3ca66bcfb2ebeb9f4c3a2134666c23db4dc3800ebb759e716220dd918eaec6501d253cca83dfff5349ba423029641790e5304d621b69df159b1d6c996df3a36bcc415c340ddcf7e7038889adda8eb9781f1b2af700614228432b71b5a85f8e8b67417efc03086169d75a8f4144fc7c8f0f45dce39b9d193b1aacccd9718a7d58835bc850aee57c8a92f7097956a69dd1f1a3a38c68ec1441c1fef2aca313d62403ec554edb66c91f174e921bc5699b06c8abd68a61e337949a7cb0d332532297e5ff525c22b193ca249fe29d8731d99354de2a74d1e69cd82924774f439548fa9859929adef942514f25e7f59123f0cbd18d837ea1d335224058f8d21e2bd9a105805e14f74b272332197be548317b89dae4baf2aeaf07554b00d542d5fe47e66112ee22a0162f2227a079276939bc483fb854c9c1794b360852d65dd83ccd7c8b924498da64378c36b73b2cec2e9f4b1df71db921c16834bc05bd72c6cf2597228c979a4f58f7280767e3e4f11e8ed59a0525c6c20ccc59baedf260e42ac5a1696e543d917b70786c88af65ab096561dbcec31368eefc9b1500b41d7185755efb26a7824287bf475dbae66968aa7336356c8578dbdbdc50d151655a9a3accdd007364a8f0fbe349ba773c243d8388c4ee3d417e6a736cdc2855c42073ca275615bdc954b3e1241e6b0fa55e96b52c4e83636e795df07de89888c5b8e91a32076a7f3ad2d8366fd9f383bea2cac08cd159231e28bf62921eeec4b31d40dfd0f6d2e5c45b598b0eeac5a8af6e8f9b588ae86f421c9a15e0cf40eb59aa6d2888c51726570f8f5cd8bcec928b347958b6304dab10323deeb02fd8c3736ae46d7c780f8a27618d2f0b0d71a58c1c75cae80009479e4b0a35db64e62daaab7b0402c8cdfdd490273575790a3c79720d65794d2dd1477bed14429f2d8905b38a644a66947b6a05061e68251281be680f7454123ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h8d47e56e1eb7a8664197fd2755ad7726507618dab188246a0428e7d1bb64152580a252af87ea48847eae1f8d847d451edc6569240d075090dfce6558e7858c35d5b98e74058bfccb0b171dd688031473b7250a0ffbb7b0c23637f3cfa7290342a90c8265d9f57480639675d7dcdce0dbddfec648ae8e38968307e0c53e4a853a7f487e327e45c63f4338d3c185562fcb327f4e6144e43d13e254f4b296de595a67744c60a93d99c78ac8414a89e728a259bb94c1f1ec1d606020a0f0f1439fa13e04d51ebd1c70df925a44058d12a25fdcd642912424844873c87a4b6a6eaa8d8d5f0c54f862ccae51b879c045b0fb76179ee11d48eb951f45d140c90df9c2920e53dfd52528328debd16439bb64edc7017287c0a73238ca0f3e4a5490769e78343ef4f22bd3f2c932c49654e1a28bc64c1da070f2cc67e82b071b5321b624cdba973ca1f23e9116d2d14526a0a9075f934041e246f1d334b0dfb16814c6e5c56fa1d65eaadfc4c1b4516c03d94630cccded5fe999bda92cf844eae1e822778c663a5986bfe104063779b8ec55584690d9507cd11fdd9974a255598e109ac7588b4651a02d4a74b5695c7116a0e785585407c47295b051e101f26bcd9d06361abf13d24e14ce5effdaa90a09caeea66ebb7f2e9708f9c731d26c142950686b911d28a2f9cdc999ffa6af034549a90cac267102b7822d85f9e8c0a0c9097d2222b495cefc02537c543187b52a9c64901238e44fc3029ea669b61bdee36c564a09463d62cbb48530c31ae3f78edd5221cfd7806300503b89d2f82aa8fff46e7bbcfb36c0b6d5a01acc4a69250b645b475d378800073891deb3260751b8e3cc38d5e76ea9548a31a74f8fc22e443943dfceefa332eb25dafa919457322bb0fb9b2b8f188465d176d91a533f7d703bf9a3efa261190de8343b69dc5c723e1ef7779b08b55fcdb90ba0cda00f9e990d4a1cd0554412594585704cde8b43c584512ae5575e2a54516b90e30028dd16105390c661062947cb2a9b28e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h9f858303704bd2ef2abad8ce0ad42f68856108688327411fc23e69097be8af5c1d0ef753a216c4316826b27c19d363dbd6b954c0f3cdaab0d9e5c8bc8768561079977ab0ca68351b97af5af1f3fa926eebab968122427a4e1543c85bf0b1b9b2efbf3ef9db2b399f0c48e88aec7926309bd0323327cc7e78663cdba0e3919f099902d557ae67c946e03ab36b43901efd3e1af36a03318bff2e34453097b433808832fcb204edad2803253366a39cb8d4fe345ded4210981d3b6638db1a030b8d4df7a3afc7bbce25286b29a4b142ec6cd111bf4c338420aafbb76bd602c07fd907ab35f039fd60ca2ee7bec9e6d52778425df8e9bb4a95c43097d5823229ca04e8d697a7b9d63c9a395c98a45c35e3c04dc724580890d8da56b3cb13d1b7df7fe1668d955e14263575ac17d1fa31534722d904c55fa68be66fa29a7cd6342d0a6fb056db61825d66a41b1d0b7fe3958acd32912a0b2a215ff0367cd45ba11d146b7e363460d6eaced0b2cc11a01096e04206ef13ea7f81e4f7372d4af441089a97a65eff081cc8d6bc017a7404d757a889fc02c311cd3518c5d8fa607548c6a59cb91a7426deec0f24aedfc058c279551ec8d8af1344d04f3e28331e8e8e26292a16e4bf09f53e1d309e9b02340a2fc1feba26cee209ed3ef761894f8ad972b2412551e1890e3c46dd630cc015ca9fb1aaf984c2efa6928682771856deff0020962c690c9e4b3dcca58661301429e5e22805343a0c66ab3e1f301a04b772c0a85a42b150ceac65b5afb86cbdda4eea09a409cf2575d1c7171238f8b069833d187fab099c0b74741d7c021444cf7446d994f6054fef1e5b5e5f68b19bba1d14b7d93d6eb7528c9b33bdb0c2b23304f3197f145a32d1b97c40943d605b9bfb916cbef29d687302e303a801c9feabb46f3dd81478966e104886d772769392430191aaa2014596c622bababd0421072207c707c8a730b682a5af23440833bd2dba7816209fd1c682a232a63e495058e15cee2492989cb1d1cac55f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'habb06df3c0b41845e03ca263a42a0aff66afa4184c141a2514d962ace4266142164a1bd0702a216a3dde8fae44cf54ce880ef0b69c4685d99b2514329717348781b74cc941a051a2dd2d57af5edf9d7490ebbf3b9729104870681de67a5baddd6334eb155935835060c68a10d9aacca952f15444500a9ff5c6dafa54a1011747191954f14255dc9d39d232717bc6da7c99df67bfc98f587bfc15b4b9990ef5d80cd3bd75a9818aa2a73ef08edde2bfa52b8f56c850e44a82ff3b1c423b3ddea0ae62268c02165d795d398ebcce2831927c8001e106b13026a3deae7d5da91c249cd3f20262e26bfd1cb30e1399e5c50fc57e543552bfbd8c410e0c4eaddae3a3d8864d5020a5b7e193f2f5851e52b8424f025feaa86497c734b9a5b7609891e816bd814e718902ad7c6a507993d5db23c1b11e6e4dbffa95572b71c7e31a75f06c4959ffe82f7f05a9cc2a3763b34f461a34fddff6bcc378077eb010bb593799a0e6bcceeb4f6652cda79daf785a20d9082492ea0d37d076a9a3b66b6e8e1c9943ad609b696d66438e96273fbd8a9a47f5f8d1266fec6a1be8a41a37f6f1ab337d0fb891396348fdedd258f93edcd8c89a2e1e3b315f2499b2f07f7a78a764ab8b65ebd2dc68778778ee01df74a64e7c3ce54810ba6b0393c8abac67964583f7ff086e22415764df3c64e7fff5c30e222adeeb700516a714af13c619b633e086b9bb5f1eb2d9c7296a38707a6f263161d75b2393f347e0b2fd5348b00857e3f4b6e9a24a9e0c683a946c0b629061f84831a427d8caab02d454363005a56ab00d01b2d458dff8553b4d57ad87979d7d85ec3d435da798a4a9496191578ad377195c2049c08ff4700d8e24a1f8b2a3cb0caf19dc004ab91bd05e4bf03c80156ed82d9d934d8e30358180760a9ff01ea1c41e5d815c5eaa809e4c26078b79e04d4d408f813b1a24d3095d2a9443c75c7bb71e1d2d8c69ea08549f248227ca19fb331a4df5240c48c989b27df1ff55b4ceacc9f7aa2eaa5b7a0d38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h58de7c53c64f2ccf9b6e289c61f85bf7e025b703b9d987888ea4f97326c68709384a46d1620defdccb69b4d5f939e33547c54f99be2513329d2b82bc78222e1860d971a541a2f9b1f7eed787d0e1a0200729b610f0cac9d96c6ca3b554e03b5dd69322824a26f0787b10d0ce3f87df9443a154db22f37568607088e5ebe27369234743103cf60eb0515065c45afdc8c421c79765b14fd9c5d0b63a6fc87fc68006066c1079e2c7aa484413bd72a78d0588e375062d461408f0c54e359efa2beda80c8b8680713377e1af0172ff6c4e51a04690e45aff13c04194f5f89b8383ecf0138ad83d998472b9392c9bca38b63d4ae98ed5d461277d1859a36f7739365df402cf353045d255bce4679fe9fd7794b3e01e70fe90ffb354f9cffd43801ab9f43c58058f23b2d8df06335d91faee9d7f6c6303c7aa94080e635ee563e52364b03740e90cb7d757dae23ce8b3cf6160dc915cd3717f01f5870f3f5df51a538b573fdcd531293290c29e94b54961c0aed1345e59a958b89e9dfb5f6550c67ed49a1aaf2c4a578eb36beedb7d03780fd4dfe900357b880f15db9efb236e7f348fb8fc7b303d7a04e886c0df457e38dc21530fa65df8a21b149e76894e68f00e85ca38c8ed46ebdb50ddfbe133cdb8f9b08d30368db303bfed3850e94be737c6908bce30dc2a8bbeecc59ba0a00a8fb46d5eeedb29d09807327a13586fa3e331fa5042e6b5b29e3915aaac6dba015a6e130d0b46c5f9d4bc37b55145f3433cdb56faffc53c1693a3accd5070209f4186ee42265b72b660ffb9bb6e44cae3a565ad5ce27c84d2dc9bc6eb72173cb9e64a8ce65f6f7969e284651ebd8ebb71f4e93c241ace87da42241bdd29a6bbe9a4a0aae22dc154138d79025a9d784b7d3655aaec366f4fb1b2d46e536242bfbc66b2f935812b238723bb1888c1c05c2ee0c7afdf2773aca80bc447efbe4fc2ffb41d444ca965d302f317b4a09ac27e6da1d980f0122c4098ca78c35d84966821780dfd5af8597337c26059a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hbc0e536e48de440f392bb7e74536f9d76ddc0b4500e85452c3288a150f1a6cd9fffdfcf79ef71aedb12ef92dd7b3f71c36515d16e94e5c0acbae10f987556a9d426ea96ec8da82c8a3f84dfaf0c73a7e6ad99f0d454d65345edb4f217765e59b3c768e3a89b2240edf62b5a7ee102241c116ad62f9726b14b3421fa17e7bcbd53aafbcd42b43569995b180a987785475b4e8e78b86ba7c273dacf54dd828c45e79666e37a0b8530e25f581fb4a8a231e607b0f78aac0b4c0f5d0ff80227efa08b1f4b2b18c3b18448a85a842904e9d17e23f41eed03f63c30ead5b6b676f0cd4962172852deaf7a828e84490c71a2034ea5f142cfdab9f0964a0e1ffc85611853dce5f80c25bb71964d6345738780836e21f27c38b6a1eef97dc99de5fc093cf245d2e22b5db3c89b23aeb501ef4962a20f99660d270286544398281d3c64a32f2b88cc9febfd1517270e18f71eb2806b171eeda3fedd47ae609602e5c0e5c30de5809d7a65f2993c3a57dffda889c8873ff8ca95cb8710358591c83b357755df604209152ad2fe86253f4659d12c5813f5fe34510f90ae6801ec2249707d887c9be4085eb71edcf93cb5684bf89e06e857e43a997a54c992ab6c191c3325a981ae0dab1eee38a49745fb96f44a2e43ad7afa378cca78b62b63b6f14ed0da9a389fd31e226a274ff22cd6b62d0863bdf0920c0fd624d26009ea66511d1ba4eb51d0371f0b5ec446fc81e57735284f04ac4d8f0f7ebb540bd2b175a771b82037aedfaa0bf70ce5692a695325c203427095ae18fb5c4a7ebcd242a40fc3d4db67adbc80917513a34fbe165bbe39175b2848d1351eeff1576aeadd020e4e3baa5e7c05e0ba199dd30500d5530e98d4c94607ad707c17b1514a57349c8e111f1822acf8d40982695cf5a36c432c31933138311c7d7cdf392fadedba2de8b027987236cec0514e5901ce96f6778dc3471a8e94073f511c36e0b632fb9709086b86255903b369881f8de424d0db0c7710ba13c3123d8d2539beb0725;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h8a7380113da8c45704d7cf318d9483917d86680622c67112fcf2d5998a9cb7b0783d9a1d93956ec0103ec8f64d9eb9d77d3cee13207e34ffe89608e439025c3be8339838ff3273a9ab5ac59981f264fa594411e23d129775e6c53fd0c90058333706753069bccac60310d4636c35ea5de0f7d0612c6449ee428ab041b0d16f37c6ba26e27a7de781926f6c98dd33ae6e75569dacd1457e70a4cda74a18359c06b6ea8fe9f4dfde85fc80a89efb68604f0fc9b576e87d0f0ee629837138c70d9cfbfc086c6b9f0342a70ffcbbb2d9f6fac4d67824a19c64bfbe269217e05f4bf6ca2b94904815f5edc52c5f802925dd83dcafd8a8d49ef460cd934465033ea4fcd08786b8ef4f75f0b434eb85498ce4905440e53b21b03767a98ec0f089dec87d9456d82503a1f264a77347916956c1290a881bd57ad7c458c1412ac9ee9298465ab7cb735680244f27789557342797c4ee0b777f675831a806b17dd89eea27b4c99b80b92060a7cc724a38e92a1b876d2275840410ef68a80892b47268494a0d3b19d33e0e741a04d67a7a53716eec1acfb9cd1808deab89a39998dae155ea32946a0bd44fcee7d1657e0dc42e515450f8ee6fc8990407be6b02861f6af5ce7cb5575bdc47472c4a49e52dbc2b9220b7cc467705f0a2c5c03a48c66d23dd72698c5bc7dd05524b5f9b13e2a7c9c6f9c660707675943cbd2cf5c3ceb96bdf5e916e39a62f832418e8ff9c115ceead4a9d3a9c62bc13a7bb87f40b0f9652aeaf9374c8f53b591f117ea0c8ed8527c6a3e8513af88a25ba95b9b7afc090c930d30f88366f3f9f00b12c8d197703cee40ae55ca23cdf5be1e4f25ed5e2cac9b6c02aa1d5a5cf9dc1da7cf8cf691c8370e476a550429ce270de42354e7a3ff5fd908fc1a9e101a78f05c6cb2120470eb0af73f43638886a47c53728eb354e97f1319983f684ed9cd98ec9d3e8303ec02cdba5c7f82a85ae766540b070ab595516d88552cf127dd6d8f5fd70f779d46c34846c442c6716ce20130fe9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h11359fc96eeb929db6b2ab35f5ebf40aba6c4faf978c48bf811f2868a0597edf4d729e0f55a5c89ed0955401f611e24d65ce16610298c9c7ee050a399175538df8cb12c38db043bc4b5eab541e3278aa5b0f68111404190347cf4f89b021372296ef091890eccf222b7ec175325885ea0489f5cd27d8269dc7b1b22857f81dc200d1e0884f09d9f0d71b73b2ff521d53c7338e06c059386351d172ea1b94f227912b092a629691fddaa431da86f71c1fd20645d60efa719284109d3f405090006fefa981f8e8f3b833deb9e3d7d713af1069c260af5ff8b3e1e55f6ee9f6dc78fdcee36c0fac10b432824a137d96ec487d2bab3519bbb52a660778d0fd2331e89026311d342195d4d7f8d70409b35c17c003e9599568fb356baef0e776303f8fb7c8d91c0cb51795faac65a0bc71bae6fb3a345ea2c4bbd93584d2cb9ffca63c5b6186795499fba09395cb63b1a2c867ec8d6dbafcfb19e912131035b2f6a8a3b9aa00efe29fcc16aa58b0448cd0d35cc34dc65659f42847d6058bbe00264a932b8682fa1735f1ccd88e04b7ae004e2f05b96e7a9d1181987b95acfde6fd8813438fee64cd3b628508a0d8bf963ef622852c0e519254db689c922bcc4de40a63436e2936eac44a657f130e6c854cf4138df34842c414ba3b9b027f58a4d7fbc4de7128693baeb41def78b5d1de4fcf4221c8a468ce5472588e899c8793c971fa17f51f64ce5a0dd6dbef3aeef50a4fee10e172d5a8c0561bfc176525c4f3f3d9220c7b13718ed371a9dddd6d04d704d0122e6947b46e41c42e37d04948237d61c4f2e2001962677ba4f86d9b8259790a23b0f0c2c45b0e91fd6add4a438a3f800661b306cc1b0296ec599f05a347f1e274fbcc4a04eacca5aba2310199d1920ab1cc4af242b2b31b47a8f95cc76ce8568081360bff8a65913abde246d4837b6870cb5f8246a65eccc18870c7654e9c7ad937e1b27ef516dd3f713aabce7327f4e27e791860ed0c6e2dcec9ca9d91d81f52662aafe84133dd47;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h666ed041577f19c1217893be89a7fa8388869bdcad6d1751620688da2ad10c55fbf7305365904dc5a40f4c6854052af7cc3a157b51530d4c990fe6cba4adc1a8e6a92fbdfb6940d79e8dcb73f131865b22f35cee5a97ae76a3f28d007fd779f857b38f426ff22f35e9bb51c7c33ae406c454f35008abdf1e615164f5732db187ceecf3aadcc8da3dfd0cfbd2a2fe26ecc844d10b545ede7506f9847a485e1d434ce9ba2136508fd2905f53a07f532fca500e5102b9914307032c8c7cc8a4550f64a000fd3888214b183141f7253639604c66157f42df14d6ced821615db2bc51989dffd23fba37dd1077e38d99803df4b887ac90cf75a0b5a648b707c2b00d4017542c52655ec9bd8928c9e5a9ecfea20fffeb3c143eda71f7ce1b405b7bd7958bd50d6c9f3480acff41373d0b87c3eb499ed11363c931642c1796a2737cb455dd6b97daef9dc0ec019d69c6c07debd52c209b6b9ea2b5dc843516a11055181fc92171a473d3ad66e0aef2b62f0999d79304db9e7c6f96e4bf5f89f6e16d87be920f25a161e05a31f961ba6ed0f6ae8284195ce444278ae5aedbe3f3405635654b3212d6b162bc6ba8e3f3ab80019e2ece93ba931ea4d45a01297476ce2d2a308d6d930fc21e31ec0423c72a224f9259d5a853855d9c9b2003241bafc1e0ff4bc44ddc34424cdc028b68f9a94e5b4cfff4017ac73d746dadc13df1b80a1aa2c07b8dd3580d2693676bf74b367e21b29bab38b942024f0c62479dcfc488a54a38315634845a9e214aa5b24931a3fa5da318f8f9cb02cae0fb27dba8ac2a08efdecc286e608176160365dc3ae4284c6a2efb0d43237f58cc6aae2203816712cb3d95e876c6d0eebfad58d6b013f5a7b1f58013ff5daef36d0fbc2b59a156676341cdd4574675cac892376b46f5e570be3d70a148354b4ca08cebd805f67ad25019b5f9620d96961d85a489cf4da1cb0193f3afbf583449240f9d06ef4d57e8b8d685d4772b564e709e75ab5e3d560ccbbdfb0753e81a12377643;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h8c2bc8ecc65ca8a7a49a5434d12ed2b725d491252c5af184ee137f3b39e31b2873b20eb3d60cc1ce813657ee706c6e65fbc9c1a85df04184f228c36a29a73b1397cc403bbe5b838731feb86b039b79ba060c23cab46cf79834918ef704d7df4a1debd906ab4f02f99c80938a67db8dea200b6ffedd2a062ad21ccca72412ed91b69624418c991551e2c230006ae73af1744c66cb5ea5bf17145a5b283d265bf27fd10294e68d2a97580d4e8d1c168211fff964d1f170b7e98cad5323ad4f46f5a9a42da6b7d7653b8bde46e546fd38245771d143563f02fc9a5a9e90b444e12cf9009acf37fa24597b4516bc4b3376620082fbce643744497d040036965ca6aa09d2165f5c19ed491da1d4d91254d0841e7863134d3d2de368140c1e187e3a7135e6f4dd31033f5ad025e4ca989ab7b3d5d2ee8ec3c3ca5586267cd22a1112ace6c87726ad32bd7db5cf291e6b4dcef70b4f11de90f82afee5765ebeba23feb9cad6f07d2be6e14f66fdad2d7451e1938392f710ebb3d1917a71dd38c5b1a3a08791e2337c86e04e9732b26fae0b7f76ef9b42d5685d0c4ac6f33cbddda7cfd2446d92b9453e88c618e377ba83c8b7565bc427bbeb3261d78bb2b3c782bd5cc35ee5405708873a0be4071d0cf90bf664c8bb5b90218d7473af96b54c081f073702e9135fb44dccf3f98f72da15dea9edf8a39fea8244da2775dfde6bc8d91480e18ef20ddfbcdbb335d7b5bf641b9f6f755ca893571ad04470bae5ed0748797f27214566e93708baed714832fcc500e4948959b15c3d2e11c5514e75df9a0d2299966384d43874cc82e32e4843ed54e30f898c765f609c57fe2f3af1b377183d8de77d5f55a8adfe1fd9f8f801d1db758acc466004bc4b391623c47cf3a8819c6c0b40ff345ad738b2059e6b2ceee019e227a1c3fbbed401baac10ca136c09d83ef5ba1d04c44a1f6b77477f7bf9b6e11971211d841d16df8b2859d2e20ba2761d1de9e83474f58415c4f176b473823849e0925a59b80dea32;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h402d781146e75a0b8543f625aa156f2f7f8660ac34be7a8cddef8d2c509cae3874b302b020010f353f8532eec619cd0a64ba88f09c88da04746bac49c0a2bc953a21f0837726c05e08587afd2c50a52a5944f739953c45fb8863bfb12188c004e7ea7aeae7cf0997440a0e7f5111a8a68b08ccd11a0906cab53601523927f9294131e2c6ab596fa157d1f8c990c7e7053f057e0d6b05e950165b4f3f124ed3fa2d150c2fece0cbcd3c1c87422ec4771264e18ec45bf4aa81b37b99870ede1267a077ae097ca1858781d0ef58ef176aa9bdf596b0c134d654fd3338336cc34a967832d4811c62d5dfa6227af161bd6cb2d6fffc7f9ba7b30fb44b2b65fe03b8e64a354695d7f4d560052aa23a53d50ec8de60753caac4db3144f576ce334b19f923e99c69b6666b48f829b102f7635b7328b7429f4e37db502694df228d92bf1902ff8c338a71bade08463214d8c95297545b8b378a76f468ec14d45877e201dfd4e3fbe1f066ff576535e2298d61554f93639946e9e3a557339eea5a35c3b2c71516d834c3982c8700fff06eab79de68a8c715e17eed668aa50e81781c5be29b0a497a6420bb2556145910e0280c93e03b9a220d9206bfe02a93b8c96bf21ba46c085419bb07ec89ba038cf8320fcfb87bb77559acd1e2f0224c721105d7356394536a5143bc641bb5e45fb5e45eca50a9410f94625fd64b1d853381c8953c87f3a8bda5cbca3e570e5f16b695a1dbf7ed404f59d9629117ca6bbb541ebfda4f5d5e6099d2c876ccff9886b13de6532a38950480e149f612f6f5af827fb0dc93165119d6a9a26f4eb149e20121756ebc77ff8f866298c846ac51b5ed76ef08093601f1094e80f935d0fcd501407e98b0f429358ab8d711d076c1093f3ef314c285f774e3de1dfe6c87e35155f6851dbbfd987c6922aa597bc715e00fdb3c5ef4b406c76ba1b370b808afb14fe58307b2ab313864e1dc75256ddaaf7ce2516af2f4ff0d177a50043a9a6efd4dab1989d6c045eb4de507282e99;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb74c0cc32661108a99109e986f0805c14a1185f13417300d8b392aa3972d55d053188579c49cbf4addf6dcdce4ecccc32d09abd4edda63f5815d79552f6581450183f01d49eb466a71a5cce38c9950818e2a56f9356e62dd987177f2c8a438416ccc6ab76208d84f02c9fd97381e9c1cc1d7fe889104c0e730aba7a29dd4fdcdf42f563a924d2635fbd128eda48f67d0c669b93b5c33acba2f40bdcf7f3356ad1d9be658c0608a326ca05983a5a70781133e26223b625a5ff0d8bee0a0271cfd2f26aaad13d9ef9cdcd048506b0eedc192d065e9fc73e93ff22e37a2132d6f0bbf6c24702e6328a35f2a054dbfbdab4ca65f879ec29af9b8cf119bb0b2ce9d7dd6cc7f589ceb94eeb785f0d504c8619f776ecd9cde001e6b67deda8b383a5ad42af313c69dda2759426534d3e3eb7aab6bb0b1c86c4e6c06d2ef80aee52a4102488b45fad325189fb23b068eb1d1ff20c781de89ad099b953b2752583c0b0f9ac30d684bbe8e005b47d70371f14fde9944284ebfded179d6d3fb297d44ce8065abc4d08b630933c8f153aa62e3b8e1ceb52d34c0da48784ab23513749e3a5385ed310ca6a674612c89c0f992d811db7ba586590b3179805855243985c6e59c8fecf4d0dbde0c8cb66dd43ec22da4eec1b634153631c3782d65a2e8fe6addfb1aa7aefe7a2ad1572048afec582ce1550e4395f16f9827e43d6060acecdd7fa4427ec006170b63195df068f989fb2976eaf58986b6ec3731ee574991fd31e81a2b5dd6f7a14e02d70895ac12181e095a8b6d46a58fc488ba17de4d03071272b294e3135e81baffca9f1902c9f6f4c59c2ab8e17ae67c3d328a894cbad56930dd24177b3ebc44d7da89720f2aa35f186b558be84f223bca06e0b69b1e40eb8928c8da02d39b2f96cacdf02deff7a1ba4782199ae0b6c95e08327ae838b030beef8d5899a6c8b7540417628f8428abf27b7389b72b0698316f9aefc3154e9b725666d53348d9907aa2184cf2e69be5337d6c7c13413ac1c871afb7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h8c20748f71b8f5cb30ac2a8f03dc8f43b4a315968518cbc1be29c62aa2ac1b02a9df1ad33d17fd09e627279b6371943cacc1c2601e41d2438bb0bc4fbe9a51f013b445d81d132705ef0140616d829bb16fff92b7a29d9f998fa81af2250985c457d78c558149395a23f0c57d06e7ce4dd9e740d1aa497a9de3ac337e80d48ee808d08a5348957761a76c80cf3828799fb97151f0c46cf73b220c0395ef6ac883af8992a9ddd79c88e3be4d969d2950f41b8c5439903093220b195db9119ddbf9250af7b5f1bd0a334648165b7c656a4a3644f874f63277b633be7c60236469f9c651bd6792e4bf83354496de41fc787f68f7f1242c8e3ee75b7abd8a9dbb5db866eb73f84ab108c276f34789cbf104c83da3f9fa6544f42c431e303edc39eb6b6e9707c843ff9de9a1b3299d548f22a2aff4af60a0c79e6309e5a9c588a50e7f5471b2c118751c32de933138086f7373a301224f9f63ec2d0efb632a02eb077b1d37c5e4324e10b7e983756cf1732c87fdb65afbbe62a04bba5efab69d8f7c06cb6e2f4d8c1d1d431637be452f913f67a658b096b0ebef9935cf6ac2ec867ef02ef8e9e828921b215bcb842e6561f5ece429608f9f2942b7206b00db7b0d7b2cf72a05e88a34e72e0d49d5beb58fbcf94e3f3267de172eaf4da9160e6a862fb6b00e24270544401f66bd5a173250a3fedccad74994ec8e94fdec9a0500e1e6f864e1617f213f91b9445deceedfbe7818315d2c20a63c66032b94f3c68b6c6a8f38c4a36ebc135526500fcf0daba01e615511f7b92839a917cdbdfe3f4d74a8114f8a640a999ab57ba05fc392d4bb2d5cc875196b7f1cfc6e8e7e74fff53eba94506121d9aafd76ed28367b86e7d7c019f937fc5e8b56b3b1f18ef801281e99c4d1877341b1b7f431ddef839b757bbe30a88b73761e746c6f99d4fe8674e289dfd52a6d607e467c5f1126deb1d9728a448a09def9cc0ade81954655bbe8101ddcb4c63f57058cb75d68e52b38975a57f430124b2a021fa61f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h1cba47474ba804373c607755604d964d001a9c522e17fc5a8a99b28e25b1871c0658dfd9b2c30a0be2b66b56f2d3dc105a86c15424b95ed0676f597b77f128e56a034d951623285d994faacbea0cd8bbb093a460e64fa156653b9e9b5666e1fd3257da4c41da951ba5128c91ff9992759ac6de00ac66cbac50c93874eeac59726f743b0b546e88e68d2a5336aaded8fca5137646da6c0f9424bb975462591d2294e65d6495bba2db0df13286f061c03aa6194d9b00bd496faf40e6880fee77f7bcab653f70fb1eb5a8a151f79283304e2987e89e08c4cda42bef5728f4d215727bcac050cc0853d7fba8cfb6c75277ae3f9ef8c28d739beed3b7777770550767877fa2bb50a3a999d50c774035a724ebd3ab06c94d5f758ee0443c8db147f1f72ec27d471cfc5a81c249b5bc4bd7f0d7ff68bafe4ad486e1cf522a5cd3abc09a90d8786f793e643bbcd58c192d1c922e2de140938cda69d6fd0d63efb74b9a2eab4b5f38f90a7c160a5e5cd57874e38ece1114624aa39c5c4098e980ea10600e5093017ea735d4f796a640b1742c87ca103d70d31e92abaf4df1642cc88aff76c17009129be5f77c2825eef12acdcc75ef4f189988806e1b592b8d9f0eba15d84c60c83e0879b9e6244b6fb49f889da799a48ed18ea0b79939b96b0677ba9f0387b01ada292c978bbee40da73983a542ac5a74c3c859f78c0c0905808750ad897b84ceb713092a3c84f690240f55bd20009b6ca64a7a2b303a540ebc84566f58acf4c40506df51beda5a331e2f63158495c5f42d45f0027649d7ee814a2e1a3680a3f5fdcffa5f26e61ba93da347c9c8de1c8ff5840cc84b226ca9833103e84c93e12e0a78ec13af1a55428a4883d4c01febfefb78471b10f264f90be978171b4ad62a3521f8ce98affde348d1d216c15b6b1f82d54c3488765338002d1c2b60f0798b03179f75105c57d69504dac35d8847fd83136fb785192eacbc471c8050c6493c5cf0539da37583126e6ef6a2a0d752a7f2ef7c15ede6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h4a17977a0e67601d68d420b1d72333d7437c35491eca355cbdb880f011fc8442cfdea61a86847faf46b6124c1bd149afae4f6937ebe943122f8902c133464cc96d0782279ed3827eaa2a0ab7830b77410adbebdef11bc2b3218f1ec769f9aee08bae10aeed9820b8134eff2df9fd05a9431ca7b51deeffba65ca885e522e59c3baf51ca805a08ea40547fce0995dece5f18ce238d9462ec48f9ae63bbfaeb31b3ae530479c6548f519501f095b012c921cf03b6789759bc134506273174277a68873cea2f9e0f47e3d28027502302e695dedf771ab33e26b34d30f170a12adbd2a58b627fde6bfdfe473bfe39e42987eb4b2deedd52dad0b4664d5e9b6997e1fdc60e18f7f5dea0d4eeaaeb4588af732c38a5ec07ec47654b63fa1c547c8d2a33f00e1da6564dba0b3fd8db18c60ff29c7b4d2c6c80a73136079e88167446550091601fb5e9b03763bc256e46d00abf95ee9105619cb542ff0a805b9792149e994c71c72eee162c0226713bfc496364ff12f870b0a733d93734b80c08aa3b57187eea78b5f8a2dcfeb727f77badd34c67ac2cef270a83831f8792e7233347f619429d995e7f865582ac447dc2b52cf79dcab6c6113771f116e19ba261861d0f8187b5423171cb291cf59aec805df4720aa995eb4c9142d5c76edc58d5be6556cbc03fd59a30c1efef727e861d9a3c41ae743584efe8e7be78980552949a31c5a9c288a5a8de26bed106abde7613faaf013518aecc94889db477d47a21371248fca595bef4b3d1c154fc4e6a48f93a0859ee571f3412c9e18e187f4e47fdde01b118dce2162fb8dcec79968877d43614b23c758147e5f43ea25f0f94632aa3750d1e42f23c9368e669f98438b88c21df6f1cdc5e3902bfded0c2520932e52043e4ca1f0bfa3d21e7b188305c85757ffb4f51307418796e63aba0ab0358bc7025469fcd16b15deb579cabc1c7c512599401430307f56690f4960d910b6e66977c8fbf9512459ff3af99d32501325190399c8a9467d951eaeaa7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h8420155858d203b913b48e211e5a6226334655bff39fabf49311e2fb40f2056a857aed868391393746fb2fe8a57ff86f8cccd4ed5283e9e9d7cbdb51103e1cbbd67f3673513d01bb16ca8105ad47c91be2ec894b0d0dd80c66ba653499844754de6afa586c9d0e1b79ea6b8e94c6dbe9c7c7e032e4d3e6ef8aaf30f366bd89c970da1c405a78b8099cea902457b4982117bdc6421984119adb97e13bd4d692f53c2199735007d866c54f4620f61cb77b6139a5255fea38c92d1e60260616b1ab5d66700fa39d71fdcbcb97ff65af6f568089ebb726f6ca9f339d27da350d52dc84f3736f431e202a404f03eef9d2dce364838a7f394f0a6be39eed2e130d04eb292f0019d0f0243fc1e84e18798153d55c27b0b77f98eb3a9391b78953006972503490725e55f2e997ac5b6dafa52f5c6a37dfbc66fb770810643491be1020f9915d5742f119d98a94f8ecc32d221cb7466e0402cccc2ec0af5448e049cf58ba61ac54f563ffd82cb5b4b98dac3848acec2ea7e005ae7a2ba215b4632109a5add63d894c0e6d61f102ae131e70b0a4f23ad216c12b63336fd204165ff4eb6c0b20043b2b734eeddd318853babbd165afb4f7b04033477f2c0c13f436b1ad09a7c61ca07119b9377c6a908a610ac133e8f59cc47ba7e846dc129b1dd5a5059e1b0f6492b48cffa9eb1016f277c5cf96d7cdd9683fc481b60c6683425e2fffac5ddf5bc71f269111d8ced2915e21c651fcc2db14dac6ab9704ab3d11a1059185e6b9ed6dc200acfc244c31dae60218958c60de3146418f298ac1bab0865b723765ae2141dc477ca6a74fd01834a4e65f7d427560721bacbd0d9b8b2bf247db77ce3d8fc42923b104d33d29c76a4e58280c7f323713e8e5b0a27122bc8199d4b79331049be3db455ab7194a6e805d3362337de2ccaf143701738a40d05c4d9d829967a68aa817e2266e35bbbc5a2e6de8234d88743db37a1ed279ebc2f97bceaf78c8656d32645f87e0ab679dc4507004d17d0c44abda8a8c353e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7e68cc74e2027e902a032f61ae2dc1980a92f32ffdd2ceaa6660f53b137f1e9bf99beb7928f1c641e978afd5a46b510963f585fc8e98bbeca871ffa841ce46b84757e05b73f3c37140ea11a673f40cf1d192b9c429c18a8d5c020c94b9735a93772cea043632cea1f1c8c83fd5567ae64397429530f89eeaea8b472695110c9da93f253b0fd80f85f8caba6f185ff79e6f9a520a62b3e60151d9ad416833de5b3d559c52b0007027251130da0acaae5d2619f427aa348b2b7a55238044a5ef1a30589389965ff5ca00b3303b0bd42f59303ff051c93aaa79ba2613a6f08b9a272e7166a06534ef849a6d1defd5e85959175098358aa9e7abb4f4d85b071bf3c7b2ecf0c29a02320400f5593a95ed7164122ca85fca57470559f5eb0db20b6662581a35734e90d3c49b73ba8843892bc50a00d5014d6772fb5aa095227f8f651a553f86d0fd5892b989b43e0dce61e6fb055cebdba00e0f9fd77208ad8a27a4b95ff65a61f47b25f1fdc7aafb2b4cf2c314e38d8c4f5f71bd8a121554f633c45806cc81d50ea97817557b23ad0b7b46689677646e1ba4b44c7350227207da25592fd3d46b5289ad19fad89100b7e13b472bd6212e562556e30d5eda14577f0b0b00887f2b08acc69a283bd2007118d4c44da31ebe809ba62624baf63ca20ac5d8a0f99c679fc844939150c12b518881f17e13b37480b41635526af3e55de110b93ab9d499515d1a0d36292b2a4722ec45404f55ea2fc595a7349842f86e9367f60bd5f71c80933f4f1fb487be6b4db4b29fa7d528f0e5f9220cea1cf25f33dbc97abaa8949a30fad2cc2e70d821f70179257b9d1e17e56eb6c5ac09934c296f5e345fd61b618145ac02794aaedb751e7aa29c8c7670e50f939fdb0b49624a9fb18627fe4755532b06549373a1f9e8235eb1c7d0e459d015f334fe62cfe47ec88bb53589ac20ab98584f31a6c5567f1c2e93337bdd521b265cba9bdab46ad2de138b87c8917b997bfed748a9562b9279399154fc3e9df2c60fa5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h9032ee1a6beaaa3a663a03f2b72e16662f07c4be70635fc7e85060cfd9f9f4659c6778a8f8eecdd4807043467ffe1ecd702f626c2fcf066bbb4be4103b42f4a808f9065f7e7a8abcfd04a6d6fcce272fd406cf001053151104f653bee7da2b53a26d55adf57eebfb1bdef2f234fb8551e1e416c4c62db72f373af8707bfc2fbfccbc3205d30e9e3d25055fabd0e1c6dda5a736a96562b9e77ef03ec833fcebe7a7102797e2a25a9ca384264b3911d03c87e1cca8faa0cdfa857fe8cd6dbaa51dd19682c9db304a35669e49dea1a8aa8d5bd07ae579299a9aff21bba3a4c7020fec186a900bb1da847d90e903890fb9193c452278ed9e244adb946ff14c6f2a2ddb4b1d02b41dd9e3149912d2912728cbecd24fc608ae8aa26b40109135e40397d482f162c2ae8a8cb24ae8d8f8ac525b424fdbf2618c442838586c3f8bfd7a4079aae54d5d90af61f4d45eb57c7b36f680f80bb3d584a194239ab723299cc0903235401fd5e945432563000fdb6f5114ba740cdec603c47c1c5ff61c945a70ab785d6aebc84a04fcefcebb953bb6e02f2a08a1dc265bf4df5dcb35833874f2c8cc3e711ccce1c9d199930e67f6e37b7395535883e416fc5675baee180fc0346251036266fb553314771767eb61b2613fc65b41817cdf0eb37696196610ab383578320b777f262835d21a8968cf3fc8a49cbeae037173e62e27b923b09c4611908eb84d5c97218683d36ffedb00642f1fdc8a64125b14c852285c355524cb79f547b51ba0899260c228ca3c0d13346a3162f82d932e696d0f7dd46bd07876b8d87d1ed9234106a3ddde82b2401fac89b4278d9b0553909dac8914ca4f95327c9fb15d5efa4a0e77de855213f98bfca51c2d3d69845996ce3e0e9d80bcd5013b935ac32c64aa875737edb09b9204382a82bd97315e4710bca2dd274157128c1cc979b3a22691f4953c005a6cdf5fd3950c7e6e5e5e27128e3b6562df246bee14a0c05a4c09e1782d7779a828b34afb338c648b0ee72ef3600f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h5a0d2acabfad272c0e564b537f08464bd1c70f33660bed4106dcf7b4f0749b55b74d9d363a265fe409389f71eade7a1cef6d72c7bf95f0d84314cecb0c36bbcf730a564c126b4b505b71eb9bddec615b8c34673f8d665d12b3909e918d2f86c9abd5e09b7953b9c4e4968fc436fc3e16b1fb61560aba7446d82b1f3739bbcd136754dcd34961227e80c9cef95f0d4d1d66f6b98ad0e012aabe45aa8a91495aba3506fa4fed7d948d842a4562881090a3d00cecdb62e23ec77f301c77c2ce3b079be558420eba2a31a00d5699e44e34c0c6efc00a87bb43f07a91d8eed168a74b0ce79aaceecbdd806b9423530e03ce7086dc210a4861622d5ee4dba9ecc9cb8ef306d4c2018ce5a3ee11df92c8ada48a4c7b806c58fe9311740790ce605824cc81b82ea87ea732a0e70767f0d876cb4e3d5e149c70311cf4933cabe374b550a1ebb5b2d1f713b8be966594e8d36c36d4ab629ce37c3d9a5d6745148ffd37e658174fe605af5a6503720fb9ebb0f14b0d67bf1ca18da749512381305a1dff40ea61a39989ed606d81e40d3874b429d57d09ef6a5bab452730ab8781255127697349bf8946666d3b43f1b77af107dad2b67c429c7169ea5e7ce2ff7f9d21c57daa07be260d36d7eacd086975c36ca5a52ae423a97da1e2034b3616622ae3a52b738810cd0b5ad78b21b396b19771080918be0ad05bdcaa76bc5976826ef80b0b86c88c2e3027601f6e7b17df05dd2a8442671c757492058e52ccd62d057307f47ffc42bcfe8d61ca13b11a487a49bffc497fc8532c1851cb10763335044f1fdda448046af84b58e05c3f43eb03e34aac1028aeb94f8d773d8456b5966b20c34d69f155f02c0345ff34759b3f2ad6a83e5587bb2999c0c74b7449aee2e779eabd7e2ffa380c66d56f0c187d253884e9df5c61266dafdbb4e093f58c9a62d3e6a47b4c3101bd04db025aea5eb53865fd71006d69713663aeb8d752fda07dc704accdc55719ea4fe7bee65fe7f33f2c1a20f2a625a8126920f1d7f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h2ce6abd7270578ce6d6037b4b7fb75f1a22b5efb9c4fc90b570bb464225cc2bde2f1634d53169359f48dfc02549bbc8bdffdafe4a2c7dbfb4f13275a853889d96980e36617ae40247de0d3924566b02cdc6c13450b191b32feb1547ec4b68288c9d6b9cd9831e0702561f8d9eb784928b9e2ebf379de2aa482d256ef580fec57120d9884e6bfecedbb1fd183918852f9eb5cd93645b4f913dfacaa7e4cb51dd420f55bb07de4fff625745306051fcf76bc8e6410401fe1e312f74dabe7eb4868fefe5a3780385358a575eed41458fe3d3036b44ee9a69528d2419ccaa21fc2fd7c108cc136b8d9e739c2ca6c087f4fd715150294d9db8af8532b88f3370441ec6c633981e13295dd4d910417b3f3461a5b8a13c510df5c88b791029216387ce5b4e3983df3319aa221eb9d47a7ff05d841967b921c1e06fcaa3cf70660cd897a47bff44fe512e9894dd4c334ca4dda8fba9c152230c4df7d0e449fb09d306b2e6097bcab292820dd277ece4e2fda2b45391f8893e2cec99f1b33a41bc052148eff88bf4b96b075315c11d0e603afa94dc2da8c7ad0ccc1fe802f9e40ecbf448550adeed68e151ab7b90787fd3def726f2676904374fc2240756a2ab4ce60018f3d7e18b8e71114cdd9c012905e8fc9bf45af2c90c017cd38492fb5689c78500f9e80fc4fc44aa2de7fa7f1a1c2162d2f08ba80f085f74b685867db0b8c412de0fa13025fd4eb823d14cf9eb562bbe5b445b5092b7e69a3f80a5b8da3315182d38a09c59f8e7b2ff49584dd886360f382e58ca74af9479fb0ef9ee3991dd7935e0208b5e4915d79d7d3c2fc6969c9a84cd51300a04517a619869e6b4a8c422fef9f0b32240abb808a08372a06b669f432434ddcdb58c39ee068ba2a65dc4a0a196402e1c45a7d32362b6c9e8c14f0edace7f1ea999b360b84881523cf9e7715a9630a03e3b24662014f0362e5e3926e73789417906c054548dd067de8f1f607417bdf525c39e485f9a13659f2534cde1e84a98fc273cc9c80b4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha81ede83b1fc22f61ad184312aff30bbae62991eb3fd07321734094130c69573b24e25129f2aca6ed586d56329995da976978a936af9eb8f148ffd217a694ecf8569d85791fbdc0217d509dd338f091459d1ab50af3e9af44160fd113bf60bc5adcafa13f19a5aab753eb9073be6a831ee765d385041b101d899febdcb0522e5af28096f3d7e22744ab6562d5d0cacc945a1268ffd9cde640a5334675b660dac2619b0583f237430eefcd5533eb418bacbfc5cbc02475ac290613e7fe34552bc456432a7cfddf0ad8ddf43e519fa202861b94ef38d187b0dc2646ad7fb04049e97804840271ebd0f5d5ad2e69b27a8a184a823d81ef08282a455d45932bfd78446ee6eced933c9db406c795575bc3006f6af2b3ff7dda7def37c279e45a5e4b8ead4f70d0f431b3c7730032df88a9c1890705cfefb22cce08fb993c88d161de0e787cd559268f2b83d92e282678a839cb31b795b68f3a6a14044530cd540cba142989b9843b8c559dd9ed9b5d23e672c38b349b3f40735d710c17802608bf781fec3b29f38b922c134111ebad7f44850e4203b6231633c221bfbfa95cd452be29acbac698f73fcb7070ce6dfef2f68b2de1ca4ecaf681d521c36ff21e9a5ff6e3e0bc24b7635b855f37b767c7cf66f73924385a14285763a9dfce1ee0db78686d213d61da55968e9e18f232f08000a2b329cc3322c57b223b8207d4820f0cd348a7c023f2312c3f176455834aa7a0f856590613e50add049fdcef524fdea0c82bae86fab54d8ddd0043b69cf4fd13dccf710be500df1a99f7c66803fca3b4d77ce37f2f9ce106fcf9381735ca0fe66033f2b5c43272918f1bd2f191f86951b487c25eadb219e948f585b9660c9c1565bdcf659736bdaa7b36ed6f117406544849e23530a4e030bb6289e226019c9d8493911b6e9f17a73ea8e14ab6ac289708f3b0c5657926606e6d7ea73f293a508df832e9a55d6da694e6d15a212e51acae2e531ad361b0953a6f7280ac6f9a7bcc452b299eb509c928cf5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h642d532e86d51c8e97cfe0c38221fd757c8e5625b3cc025f3a6f1d4ec8fda98b6573d6b997df4f4aed841f7a72b631d0d4467d5ef4af79fb0b1ac43c61be2ddba035617403a35eeb957163be03202d1446cffd19d938ea887e2cec3f6df0080881105069c029fa3474e5203169378c1e4f2fcea372eba1d671c8421ff73ada9addef5fc4b4064b55890d7e5cf73abc229bc08167bbd0103e255f9265d1785903d76412f9c0e3cf454328bdf7c2f142ab431fb741adfdff24f183ba829e245c69abf34bd0c86aaf53026f2008955d31f19674f5b71f76bec517b5e0cf22ce4acab50d540269fea5091d3374cc97c4e001decca143bf9ff3d78e718f0da1a5f9def737f7fcb71d941e2dfab035ddd8f8cddee983f89f2197c29a555229ceecf40dd703a88563d44a8e3e4a90b6d6a41cefc9f8d3aaea6a785fcee3971b6c1a70c5332e4a21d57f641028314e27facb9e9e264d186bb2adec48b0e26113874ad9eec187498414764f0324121ab51a98acb2009eadf0b08c7eadb06410635d4768621f8e86dd928bf00b53e2bae600b37fd59899a69438a29d985c32fb60316997523f60121f7d5c775ffbc2c30e104e45c3c25bb93e52df6a77c98e5103e479b9e429ddf0862c5696d24fb19e63f139d3f54d3168a64020040984e78b181a9f84ffa4daf032a6f5a4315b7dcafc03c1c45b7fa8578db132cf55b3af4c96fe9b0d0fcaf2e1941989182b18d0358ca18b9c28036489fddb0b2b7490ae5571580159f026b668d77902867ffe89f475829f0f047b90e6f3bcfc007b63c14184df442ee2dfe58f7e65e65955f4d377e4d090d4df0bf3b0f7f8e0d45e1a351a9d6835cd7aa39be327b71656ad0cf91d8aadace72c33e7d769c982adec3c4d639af72d1bd5f24681e0442e719c4da640600a3bbf1777072a643240455d6e9b3e56e9eadb93f4305d0fdb096c32b602806cc801f6d4f16d43589261714fb97d8442ee85f2b3b8ae8b87779c3a767b33ac46361b8b3778832e7e5d615361cf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h5ca0fc559655e2487f605f012652bd61466c38d3b3b968aa210451f30cff0a4223f3606a8766576b026068c0d3513cb27d6b5872fecbc35cb0a2f99e171b06e13941632d019a1223ef7a63455ace971a38b0aa6bfd056f9ce7ebce1c57804ff05a610e96472f537a3f625a3ef5850d483867a5d92547eaffd6e8f8bdf6bb5caca6fe97601582257324d5f10d9dd6e6b4e8a66390b496c659d7d0e5e1296013b50beefd07e62b47aa815885007b96defed49f009ab769176cb7a51af3e748bd20e6d93228c8e79df780e87b06158d2d9acb1e38b949e67ae429e0335b61049c53d3ede8cb2946ef94576b72f84d8bbe830484175d5ce5e1bfa2e96697c61cbae29be9f89368679580da2aacea3370de76f49b024182debc3c36475e55563ee1c0ced4e61301f638dbdd320a7e789d8cc8d1bc1ad817509b77d7963d3154358bd951e3d212a79b7a6641f25619263a134e0aecbc36ec51ee6156cf05519c96d64222cdad2582b948a56648b79719c22191b4b73e07c71eca5e77f009d7e4ca4cd9c978b3d7f4f450df0f1165c76b4d30f017c7c2dbc15ab4f8324e6daf205909f875598773d7e455152307f4b49228cf60ea9779c1cee29b4c1ce8dfbbcd4743aaaa7836d29bbed50927b7b98d9118cfb39c6838c097ce5d39e6c03e11b1b0735fe9f74c73dad2c6401158980af49bc2695ecc682a7539719a4992d66722179e1f9e621c7e5c6c9ab768ff142891853d9e0318e5e12a7eb8b03511a906bdc1435b01f8d340f1a921f468fc1866159fca5c6bf6fa3387c3446cc5b971a34f5680d5aa5d40bd38813502b65e3e7364d843fd9490ceb35d3b1e116dc0cb56caae3af0be7b6b06fda53ff4e5745e0cbfa39170aeb81774af31be9bc135465fd717576555cb358af03474b8d5d1e645978c33486dc161e967ddbc33b9c404516bf1d4efac637a4cb1c532d695a3e6498cefed9a83679768830b460523d80332d3ada3871b077d180018094015faa3c4582bcbeb17225724e6eaaea08d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hafc5013a3e454816f551e3a7c752640f323e2713bb58720f53017be681fddc4771b75a4db27ffb05227a0ca5c6eadf21e6462a9bcc699c6ecd8cb15e390b5a291e20b5dcf02f1b97831a7174496dadfccb5076400b81fbdc9b0364e5450b771d0c7821234fd3da6c8cdb88a9a9e0bc17fe7ead94aa1a20f32a986c29060ad3a712c8e7aef8d35f09b08e47799ae63e1a110a01c78f929883cdbab85f2c41292c781ac5383a8c9eb7cfe7b00741d9d2d65cd1445cfd5f96cc5b5139aac3ac8d9a872612dd800a7955ac7d78bc9d00b39da4ac8a6dd1da0f35ed2c80b66a20986f8aa1b8680f96aebb1ef44387020bd24d2a0985ab9218e76abff07ea0d309f401adfa3a6ccdbc19340f84cba7f41ec8cf03b8a067cacb94b3d0ecf4ec9a632084ae0c76c6867a4717b955c6ec0f8dab78cc5600f77d15ec4279f51eb25ce7da2ffd31aef673fd1dc9755e1336dc8ab3a7ce3162a500700fa9fe632ae83cd4350116d3dc284d93668763918430a927a35a973774c4ad62868cadc630bff409b33a260c5e039fb41cab6fa30cd04fc616dc3b4e773392e9eb48dc373e5f72662c5b809ac9e84173b5f24c0601fb26097ba1ec6d6ce199d83e63731c3cc69529a152dac805ec9b8664b4fbe8f7318bf0fc6e12e7d82bce8073b0d0cffbf950226d043bccb251af80a469fe7c31adfa3c441683d2f4aff97cd74dc162788425bdd4a440d0c173a03180b19922b8f0e0072ea4e8b6bb978896cf816272aad89091d27a8940ee9aba41fdde0bf808a5eafb8c580ea377236558bf4c9d457e4434facda37dfe72b5b24899c3fbd34b636281c68555e3859a7267f596a5011d931d7a50a8d58e69a5f1155a5d21a7edcced8ed05ba5caa75f877bd65a1e3941d81f439cb3d1095a1e84a3579d5be8b7edfc2a7ace240d4a3399b4bd1b5d301aea9928dbfcb27978cdf61a694bf0dd53ba361f8bd415684ad263bf1e79604dc7778b344dfdce74231032ad749dc1cf7d49ebaf95119cbac7f2c25fb203f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hfd104c63e72d01939198d7f1c77f7c60c0246bc54095b78e47091e6e83bb3ac0bc9eab9d41ac7861775777f2f49fc4ad0af1c8cf5d25349a150d2c5e5237255b118b4a44ffe472ef6eb1ea1aca2eb044a50a1e7c591dafe9a38e816c8d3507fd706df6a784155476b63f6e453d0f95d6b266edc086ce807bede5bbec31992d543ca043a4a9b9dc3fce64b5543c7fc6bd1c43513994f2ca1d2ecb23afcea93238db80b4e3f74ff316a44c4d8e505d951bc2a13aafa381f77b84f65eaa2f07efac0ae94fda0aecc3ccce014143209a8f0f5fb7f4da3b6aa385fc422d92a7b8aff837fc3698dab315ec29c928a631ba9c0f64541340e6a5abaefe2a770dee8298608b0e5b6d1269e125ef3a0570ea320bcf5650d5a0c1a3fd1cbf050ea287ed8cdb961c09352e2b34e5dcd682238d1ecbac654608304f70c01aa1d8a69eed7d9fc0d6a50ea437260c6fc91d8031d0ba53a6e48116d16caaa40b99cdc0e56dfec9337e2ba4625d51546307583cf468b935dd080c981ba8f240be275c5f81fc1d1f2591460fd0bc67299a4bfaedea6477598d4ddd52e96ff75141caa6f0805428a3db86f30540c4e418ce977349e669827644403c640fbbbae89d7d874668ed5e77efc5ef29efe8b9852f958ab4319e777965c3a77a9f5fe4185253389a0730cc638c27fab66bd79a6d19575ab9af6e18f1b80b31c01bfdc624f01d7f09e63d5fb31aa929f02a089c57f4ba81005812b4d94118afeb1aced9e60c8d981a9ed1ccde1051a7af4bc478e48b02ce51dfcd8e2675aac095d64b2178707dd83d4d7be3eed001c7184693014b0b3b0df80ac71632a7ae61aadbf44d58f85c4d6aa95828120e2aa88da5d0aa68c9152d726dcbff22fbe2ec4abd36159bd06f0631f6b86a3968c3ae6c65e144415014f21944839752547004a73f85cc87b940b9f9bcb28439076d6eea5558fecded553d28195fd4dddc06532b8843360366fd0ead6be3164339392fa362c92963b5202d6746e71602a96371478ed409248b8e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7a75c958ee46aa0cd43be0a93ef5781e1612bb411954727313e9abe3880b62d9f6765fbff6e1329fce95426f86fff323c0b9811d54bb7dfda806d5d4264e4f7c7036aa720e142be5916abb0e9153dd8da8ad11211bda5b0ee8202cfc1bc92fe1f8d5a984ac7b742febb6deb1abb646318cc830184f102a46beb55b31f438754c342f48c2ec81eeab6e828ca48bd742b03309e75fba2e192c87e5508537f4ee1a5b82ac1bca75dae2676889caa43c16a843885e4358effe1f74ce6d2a26c4bf9bd5711087e1b7466cbbb96f19e5234dd5f1fd3fb42c094eb1931783e1b63c85a8a2e3929c4ad3da57e7988892322cee20b6113fac369a16a37cc738abef865b037b75f37f3315989209dc061577c84fe5d86c5315c51e739e1ed7bad4e54ead87359c52c13c81d0c093ba696dc4ec913e4bdc91daa4ccc3c4c28f9ed4ad45f484bbf79a9ebfb2e810df5b65712d2746c9571a1d77af1aae04f711cb576665b1f4e484b707e426533c464d3f0852ff7bfcc3fdb175ff16d0c899892c839ec448356471f94fee06582c2d78443b865bc4c209bb855092408788d82e65ed31e6efa41268147c3e0705b2faf784f9092cf434a7647576a1125ecd26db1c9ebeabe23e35028d74570ea86a3aa1dddac6cd001f8d4c80453c3468049d51260da3fb4b600089b10b12dcc68ccc28f721a0d33d9edaa4838887b053b3b98cd2d035142f8063dfd8de1e4beccbc7eca9cfeb9e14a3025038289f242db074a9c84b6c659094d8a06036e772174fc809b8ce077a8ec4265d1b0a3a14a64e746a3c2cb29d31b9c638b7b912b2d78d1083c3083998d201537eb954e6cf1e40539a4ec8069290e5b7df27e4591f59944329afbcae5acc062364f5350b804d0b4abf8003d9b25282540d1c1f63389422ff61a29fc2593a1514b8a1433fdb177ee9b2671eb20cf046d8336e1ae13e8ae672c8404f034bd6d0e336149762efc5f7723a3212b9d9c9914d137e6bc64219ac4f19b5557a2c0d32e45284a5d374aa1e05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h2758198056455cb5f79e407f8bc06c48a049d0ecb313883359bfd0d6b9261bf701d75c5ca509c169881537248680d3db2f805fcaf7dc12363a81758d175b8f870e12d73176cb32ea9e1107b3a705a9ba55ab8b4e51f47ddbd2b77357bc49db443d71ef384c180c8645016277c7f952114597a73a7c0adfb64e59e0ca64308936c5796b024725da0ce3d2d4eb2e8256683951aedeac9865f2503e898ac73826e63c028cc19b91826a3b3061d145e2ba95cc03a2b263040253c4ceb05e8ca9e9d2c861f7fe0efb40d46f48722c067ec0cb45d0bd13c94012ca5d422eed6fdba1974e10c487a256b032c27b8af899723474178d49d98bea3414ccc60db8f5a6f2307bbbec56627a1201ade92778874e8bc6f760135903d20ec0a7cecb5aa08ba8269a6852049431995c70bea1e744b395473232e678460b06b2ab7c607af507cf4ea8925866f31c3af23694c94968d1d5ee9062fd47cdd566b14af4c9f24ee6ba89e23437acde932dcc667620cac0c9694296358debfa4ecc3e465db811bf5ea11ddebb05c8beea793c5269b4371d36b75bd91664c3cb31543be4ef90cffdfacd9a6827725c82ed42d33c1bf3f52294de244ed196671044f777f7700f872e0d6666c344b678c24a3762fdc8f45efe37b0f4c0611767f0582c1d8a13671087619ec4a12ad36aac39e8de2adb1ca9a9e8906524ba569f9ef823c48f79f9e9cd73998590aa2e5e56096705ca2313c2af67f314e53ef46a25b984bfe8c6d49b040f0f38abf9811399cec0e4a435e7c12f36725972fb5fa9f805a495bf35f118b08d8fcc0526aeaaae250f21304732cb79b88f03ce30b22ac1ecc3b54a0886e706f4cc531ffc2e5315cbde3615fc98d61dc373401003240e1f95acfe0badce2d649734349fa8df41364a34806204ac2648d619c7f5328578ff22585a0755bcb39d669287eddb985aaaf086ab1cfe8c311b7d38caf9b3f373818caea173da8347b2889f3a1a3acb36f5d0d95aed573b2f0581179a2d9ee601cb7a4ed2a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h814c03682879b61dce5d14cd3ba4d364bf59aa1d38d47916b068536a6b76f5228314ced9351aa436de01cd91391b7db8c4547e3ff0fdd2a312774a37aa7b0540a2ed33fc5991ed67a445b54108edf4ffc4dd8741a9e2c3152d81c16607f73471a797b307aaa09401d45810120f6037cd3ca4485c70872b041e0be7477a2a38909b2201fe8f3842ddbfd3e69a50b0d1ba39e25671c9e417de25bd464c8c9f1220e2ea504f2c2cb32ea9f2f8c6355ea968d645975bb66cf7a2bd41cd986b820377c1baac3f8066d80bdba1434904bf9ef99ecc5390ae0949d16fdf81dfb26a14f2daa7d175e651b1a804461104275f217f7d84493b5aa0de4a30ec2271f92862de188b3a514fb39edfb4351cefeac10887192ade687057add3e3fa5913cb1d6d5db09d60768d578cfd839fd4e84621bfe84be599668fb06ebfdd9f82c43f44349c4bf7efd1b016f8a49d12e3336ba6defffd837f023aec6a018469c47e5cf6e8c9bcbcede87124f570f7b16171a0b85b259b9b35fb48aad1e9ea75c062f97cad10795617d64933c6d0e9cafb01d9b5574cab4d09cb686e98b8bbc51c19220523e20ee24e8a981b399c46573f0e2f7851fb16bf87e4b294f96068f8f1bf1ccedd585c404a0138e4c1895a6fad7c08b2454ae2b138f58172adf6575556895e18eb643005cb58facc16111ec3c96156b80ee9f6df3e749c281a5e13c3c134b46bdd8a613b37dd25ab3a74b676009f2ff97c1c9ee9423aac8e13ada855376a1613fea81ec97eb960b2940849d752f4d35d95df9c9a5b40ee4f28da799e94bc15ad6dc1b8c0c7d9ca826b314ba38da1ca9ea6b090e10d9f7b1aae795ef2eafb9503ed5cd963c5afeaa63f3c18cbc4e3e322e7234ae8677803724bcf58cf14086e5cd829b9e231efc10e2b8c038983a0a735eb4a385a33417481b67eceab6d939825a506045ea2da180600710a4e964bd8ffd3b517c16f2ff906f75335ad379ef419973b9f9f55e2fa0493ca61095733a406edf81683ae1e34bd245923;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h90368def18b86fe1cfafa8c29bd814ca252f8ac324b491dfc4344353e9ba5713dfeeec2adb09937fdead19bf6f6227035b4f248e9ff2048438ae4f75572711fe86f1158fbd349ceb4048295736fc6ef89d1ae4c85cdf2b5de77413cde03dc57bc9e973d0d666275658656375190874420c59a9a7324f6b81d5250cf4c4721c5f93685535e6758ad91da2b919691fea0a2ecdce36c434e3a320a9d5db41e5f45d5467fd46dabcbdaf2f56cb9453fc45776456dd9425c352ab9f6a094479049633d987b2f53eec9ccf2dc4e30e54c713d038fffc39be678308eeb732b49e345f03ad38cda1a0a4aaf935cae57584b2148b27ba46cf0d39b1cbce2feb7d41377ee84b5c5aa133e6bd34ef302765326a90aaf2d84a006811afb5f08d5626e4dc459df2e445b09ac616a8f0ddbd63044eac83c7d358f34e3daba4176e012d3419de1210fe164ec12f080229b238bb44b54ec697524e47cf67c886227222aae16d7409d6f0c047a038e7f2d9f2680e3cb915d018a0db3a266dba1f2cf11d4ce45233c926b0c26f17398277a814d6e865504dbd0894714831cbfd0117592c784626ce2fec0380783c8eda2bf6a5d55b65103443f0b5f33b41d7ab5e02efba535e21712da87b0e543164ed3d4fb26ac0d5157a1bd09a08f4c52e8844a2a7deec9e7262642f56b651d7a2b0cabe27f74bde17977cc73796db155cda5617ef86843c85ea6b67bfba53d498c5dfa414cf81a833cb221d3085a33a21d48ea3b83f63de4044b8c5541b2fac0939a665e9f2d658b8fe06b0b2961eeeb053a316e0b16d81defc7af637919def312e05829c93441c93716236cab960b4f8aed0ae9773685c0d8c5d93279b3e1be7eb14d78c9be50b263af6f40b256518f474f8528969a0c6db5373d99e3b1eed8b7d6fba6ccb4bd5ec1d035eb28ba4cac7c97ed99486d0ca01778e6a55a26320814f53e2157b0f84c7c6f965465d2d7775091e1fca4f630e010b15897c45de8492dfaf51a75f2523bf72c1a83402fb2ac23529e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hcac7a0036dd223bed80faa7258f727753a0b19d52541388e8f04a9870877f0ee79ef872f37bf0aea72aacbf4f86fb1203e2b8238a9b360587cc98c4e75ca622a3da2cc491c5ea5505b3da0759dd9f0cb6532dffb2649045b36e63e6a6f20fdb274d91c3ab7ab344038eb0b490a025973f2a3c7997bd2e247ce475f1a1f9002e3a890deb880222cfae4b0cdd200e189716991f472c29e8e9bc9bc581b2e9a114768d73b2b245d67b53fa8fce4329b121b7381802d1e97fd75261087e5744c81d168be19b243f9a2fc35e6950d4f2553069b2e60778e5bdcfb0cbc471a8393ab104b5fcd3414f75c060faff6786bab6c7bbae4d7d1f87480c4f1ec8c4816746ce6aa5b0bd99583930ed5b71f7a6cb34b641824e4203e548eaab5784e9989835e9ac2214014ba00cbcca3ff2579f3d0a95f662e7e29743a1ef409810f96942c44bdb46701eb76e383c4491f74c65f222d8edb10018132eee6e3f329988cf7a724528ae1417923c3df7c35400698bc577762a3fcf7de645cda38b0fbbfe7dbd9f89dac00a92e96f717218301a6c4e20eebf5dd2002225632677f223b10c017de0ab701399855ed804518fc28eeb86eebb6be2f8484b69283e72d0947a09ed4295050d829be8bbb8bf863d10a247842e8b7fadf5e06fcfd45e1339e9c5b87432e047eb45adcb05bec1578997384beb96c5c9c1c306aeda3ffec1fc95b6f3d67c282bc0f5e2c903ee3fd658fd589b77149a69959a61a03ef1dc70c3479a48f6cecbd22d7c92297f3c8de9c2a1f24854cb1fcb4d067cb5f981b0545eb23f1a95b96f6ac0414facce5adc390cbf4e7101fb4128941936fa4d573f3a4dd6c73ed1ca48fba7b28075cd8c8fbcbed0f3a321537f2201d4328b7602ce946e86637efe95ab5061ce236ddae306e06c5ce011293f52c7619477f2f80dec8c8caa55ed3953159f72a091b5f3a78dcc9a94e6f9f0a77abdbae0a1d04d43e768ac5bdd9ab5efa3bfb3b5a8dda27fa1cc92a385858db0448003ad2a084547ce18345;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hdc988f4d9ef737237fc41b89504fad339d7987d1def4dac0bcef1e9b1ad01c1709b2b40b73b1c9508f93a3e004f59490c80135914538da45ab5548bb103edf8400712c4bda2105a8894fd555345c8a845270c2efa63184531e3910010eee4c16ce76c45420d8b2e2a130294dc67f93c621ed83b53e92c874a5a8bbdec31f63cda6a640190fdd42fd1f4c5fa457f8a845228128c00f05ae1c8cb22b0c28b1a8d078ec1c2cc65c0c23561ab4b7635ec336e65a51ed0af63c2dc2851af4cb40b273f19372d3fc3177543a15cffb0b9dfc289755b7af1a623bbb94e681ccdcdb9544c4bd680ca0fd66b0ac6d21932268542690309a9cd3a53b7e9d21929b2f6f7287d9770840b22a93312baa1dcc486daf6035dbc404370300ec5581bbd1e21ff3e3b35261e51571db6816911b0fd6327511f1971e3f93fcf35c23ea7e788df19bc5c0458e1ebc86a1e9b47b592d56fa8be83febf37bbca99c83a4828cc2a3bbde2cfde98aa88b2fae32780ad63cd577a9d909977bd78af93544cad06ff8727d273a89b094d015b7570dad6638f8c366a78db7eeb6ab520db426bfac55c4abe2264e455ef774c449b2aa14c3ff05d83e73bb47b7e7323dce2d4caa77874ee76561b6ec06e36cdc6cb62fbab1789314e154e41c351436ff3aab09d1616ef8186e367014e33451024974cb1d74731f1fd5f7c4210dbef9e101621669749f9208b50fbd54ef380718ed09ae50cf6d3e5d0c5ea49329e43723a07f8e946d500d2d74bc6d86a724825a9a3fd1d6d895028f3ea8e1bb03a55010bd70e6b4125f012028a1c2ee949815e3162a40f0ccb1f3f97b4f6fafcb55fdc1c3cb61f6321b45b0dc0eba8589080a1dec5acb511e08608deab80a8e02b815bd616ed9d3313349907823ef3a1875a9274a4f04f36c411d709531ccdcc723e05e7cdb7ab74ed18260e08568b6c3cdf87bab739f3be7aff773f43db6ca9f4ebecc20f503b74d5c5d3a6314a156ff7da1ef8c958e215d7c9e647892be098968603e0a9f5f76;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h1e31975866d2e4151b2c520265d07e0b0540382985d4cbea0e9695da4fda381a3bef4581e77e016bb20eed78dee71437417da87b981cbec5bb35cd59606dce645ebf81234256ca7117bd4538f654732a1300f7299e99a6e9c6b476718ce678082adbc766b206942fc32ce22f5682a3e4b3ba2879e74c1e27e6173a9612b77cb585d0d4420baa67ee2e5f7852d5a641ff877ceecf33bebd3ebce884e9029a36b947d30c8d6fee949bd6e2af275c5f57bd2cf3124b477d3ea44fa3a17cfe5d11c220689dad5f3d6b56988d5906ea6702f5d0cc0be2a57a4aa434ba23c15f3f4769773e99afd93356f5d6fbc2fc3a6ec94cd53f83901246d25930deaa1c90393c1d93e974659b55982fd0332d3131deb3710d83cd01cd06433d9b43d39f931d734a08b5a4c9c01e8cb6f304aff5a6b4e267b8652a5eccf59f798b68c4a71e065c58e239cfb8d0bd3177cdd2cc5580a082bf17cd92ed80137f15d5fb01fc5ee7017be25e270bd31c2805e1e7af50347fe64cecdbd605ce66ac4e4cde1825db3083ec7ea01cbaf6d81c0dcde49a5e3133a907c9a5cb06ea4da2f98867fc1e68ec5078fe30df2c4c0a78ce47f2c1c5b106d6aa04bdf42e6c7d481288002720a50e4a3b4a0c1fb54dbd68bb31d1e4659c7cb45d23b6944cba7cae8cb24666c5a4fa1ae00b8ace0a4c49b1b98f564a011311961fd9a6354a241b72c38e161f54a5a73c4d9412b89ff2b394595dfa4aeca9ef0386687bbb1682de719a143a4ea149f136cf498e5665b9016fd1261e5e42f1c5d4d1a9f5129f764586a38563e5ec5c7a24e6f13231c760a348e694d47e210a1defb18a713dd3038bbe0ea5f612129958925874c20bf2e5bb1994dfaacfadfd209cad6c41a598fa3c2ae856b753e5b8c4da63382f7ee82f1e684bc4d0570fb3e5173f5c02f22419d915105484659c31801eaa9b700e28fd433b1f4b7609ddd6b26ab57af71c40df7af3d80a6be992ec0b99f02ab89b782723e6ad971d41bb9891e85816805871a58b62126a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h8019ea4ff8591802a0aa56e76c1a3cc09a2dcd71040415beb945cc38c89aadc3bcc0e35cbb1854d7c3c4f4659df07fe994b2b18be1649aec2a79b9f4914449231e606ceb386e944d0bcc3cbb0d559c02ad6575c8ff0f0cd6e9bcb7441ffb51663b84e0741ba5e1386641ab5fdbcd9cfb5bb0fd3cc58baa2f0d94d8cf3176b90f9f01e9f133e49be04600b261fbcbca29ca9115271764f7df1a4aa6cf32f6e5511274f570904837d9562dc5eba7018c258290880b7f2bcc7ecbee5ed6af0eb5040293d7a9d185317377a55e836a2e6f6cf154c4b09d753c38f814cda46ab978313f0a76927d3ffaed06f8cf332419c650a43602867c5bfc7dd0c21599f46aacf6d0e351ee6a5c1a295d3f8b934d6eff90d37e637de8e7b43b1a240855b27187fc54d8ca309a185767f7e298babe0cbca40377b2ef835588f6550f1310e7bdb69d919f5ee7f548ffe47a4f9aee213687d7b3f113e3fa7e05de1ced28eac86508d152c7cf08d9b58e5cb17c215338c7cb9c255334a5c6125587ce131c097277b7ef9fec429d15349537ddbc379923e39411c9a65c51500e4a52d613ddb29c67ee6123952fd5de0f56123377ea550c9c6169dff217dbb882e082a336ef8e94f53219178c5fc67453fe4092f05a7e1346e6882690082a39cec9154e93c9c4c57c88e69e8454ecd971dbc64a41fcbe050010645ad49404c990b387f78ea0e9ccd11a58d5c95580c8629fb4d0b724fca4edb94d1b07086f6f915ebb41b67b6c257b527e151df26334f059b4e11f2164ba6a0d51936621d9a74cbbe8e3f24d895b1318cde9b254155a0f0650cae22e88798f03c74b657f791d26cc7aaa3259bcc1ecf7393ab023e1c7c75811e25182f6b2f05d3b251a7d5773174d09f98161320fad6faf718bceababe77f0d1eb4fc2a5f0513b69c0fcf456ec0396cb8599473054f95d1f0287e0af8cb4b2319b6aa0a35939c95eb9b6add0d583d332474ffdd6f785f1d47fc766356a695a90d2538cf17b4e71db5798b87347cf94d4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h8362106500f0c80c8f2acb8941aa6a85fa29d4629edc061ee40077e701961f06eb21185fe88f1e9fbef23c252a7668f7f443173e8390401de84f969f7045b3520dfe80085587ae0082fa4569b13fe34b04a12bb22c1ccb2a422ab5203d24c6da09dd2710d9fb813041347a7f771b4bc580efc9486fb9b86805d3e11ed3ee56152ae44be219d3cafc3baa120055d9baa7a680a5d95e1a3e44ad7e6b3c37185c6c9211fd014f95b5318f52c44987fabb4bc709e935f04341e23a1a0d9d819b8091a4bfd8f90e49e0885ca90b8b3050c4d7ae5fa66a741130d94cfb791b5276b650b08800942dc60c0a3824119d4cdfcd1df2a190d797921e45c1f2098e082eb09b3ba3d0f48e465b64940a86b5fcc8a056407ff32001540956e0a42cc54041a06a72d1535960cd7ca9ddb51ee719db00313f79c523dbb8e8b6b291cc42a6a9ef6d14a7a5320968ec09e07236885369a1786f610f443b85b81637838f1a0988e1a9557d9f8d7300e5ba6a73a0486eb9840b03a8251fa5f1e3b8f122292878c75bb93e3313e0aa955882ad8d7812ea5470b7b4e7e009da99da166639458632155c40d5bbdcc7a1070a40cf2b23c74004acdf292ccfe3b9c57387766aa8ef4c8ad33b4f1865b7364dd6516902073ec61c4a7d52b1a2c0d97e3733e162417678f7c2fe1d2230206b6dc65d67789cbfbc6d0d3eee09e523885626f84515b530a14c730fbc45f7ee2573782f2d22ef7f5923beeee361f59f0c0c7c5b6da37f9e8c04b4845d955220194c147d3307dd650185c6223663276dc6dd68d4eaf6da83076cf78cc266592705d27eb61c37356b7d8bce89bcbb536129b2d718946b6931ded8f3a89cf3c2bc578678f0d2739f9813c8bdfb3c5075b3324cde654eaa291c4f91b3e0fd825e0a17f47064e13398d37e124fdc4c2f52c5b2a25035465f05f06f226e56ca8bed86e63d71d9e2e46b075f3df01f93e4da972c0e242e0b364aace68deaeb591a37d4d590e2e688b85e2c0e3c8019b9d1880498f035dd2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hda6b47ca315a6026640056faa6dc9552e677c555a3aa9efec7006395f381af31ab19ceaa2f1829e3fb204cff12b8bc232078fd8f4b63987f029bb775b280b584f4687f3b2a02e401d081ff21e6f1c08a33ffbad8d0e691d0383426276126442860811578f6e8b5aabf51b542dadcf0554c9f0112ee26590b7de7f86a0daa44e45f562f569476ae028c5cbb0562f2e956d37d6636c019232455c4d51d76232c81cdc943b9c752d6ccf5bad70abe9b9bf92e41c81d46dcf6fe1b94e710cb23250c61d8889b2ec2d8dced0f7e366f088a970499ff45d4d9155f919ca34d9e6e954612c7f67208e2a5fa67a74e54475fc2bdc6e95e64d7a083cefed15ea2d8677f89606a991719b77394ca81cc8191f833263d54a8cea5c1a55672bed5eed53d333172d58d162abf9298150170ec7f70e3fec5161c7b39520bd669e1b7a3145a474049cdb5361d3a6a9a68cff86dabd4580b27da34d4031eaba047c5b966b3f2f0c0d6355f6b42ac09dfca57b14e5cf12c1b0952d900c82e101b1417f4f0bcac61792b1bf4603f70a11ff36ce5050137923202c6fa4986ebe140b5543cb0ef6268c5608850f6d926ab23886a2901aeb6167faaa27f4e5c33c6df72997a32f78fdd6998320737b801013bb01dca449e8f13f75ecb345e0193f7e98d965fe24556659cc90a145587f951663bc89d068e430c8c1adc6f6e85239a69154bc98fb1c1531595d83de636649e205a40242beb4f3ca0f5686cecb551d7adc1735091963121d9dd980abe4560e69e47945e98738fd9b9528e94bc7534492263455900cc030c3d8fffdb025685d53657b81246d66ef201327f8bd1033d4d0cd6b3764287e2946e5875c48f0060799287eacc7293585d2861c53d16d7c5ebfdef7c91c4c018558146463e9633e91abdef65814b50fd24728d750ad671af8f3e15cf0fe11e2255a382891682c171105f564e887a96ec148df7ef36fe41561a72610dc174307d2734589c0c4132de3f7030b2616fa979fe14c86554ac1be4d49b88;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7b82f86d94c13841dffe02916c5dc8cd23fc4519e3aee3897a496e965ec07264346a6d8a48f130f9a4f251e0a71c2fb6295c3c370a27983efde2c8615f159aac0ac78ab145f01bb2f43eaa0eaa491aed6576e61d426db999d74218614eb44f894be2981dfe08d276cabf22e4451cde30c2dc20181465ce4277ce1d2307e7069eea30fd0b93ab0768f9685bf549b8176e4e03feb4555ed51b43fb3e0ee0eb1ccda99ec6a16d51cbf8a6e61e31470ffba2ae8ca061a96ee3c8cab5da99dba8dfa2312d304c760b7d32b88bdce9fe2f16d6999887e0fedbd4bad2fa0be7c10ddaba1246db252a48f21689dfa3d662c08e6414e1b28a289d516efd9115e8636dcb04a36fce4870cfca0df68bf0088df65606e80ec481a2728714c2180d0051b7b468c23152e18df740b83b34911be969e1ea744ab92aa6e2d71fd892a8a39979655d344a2628533aaed5019822174e3b01a511d005d5b6adbc5c3b12ef7a0cb33f04817aef889872f61d02f02f831f3e0464da756fe8c05c0492f4995584f822c7cf097a5c1121d4fecdc6bd258e33c644414e8ccdf60b855a0afadbdbe91b2077b57b330c761b6212101705983f8a5f6c7911e90336d8a2418d32ae0345bbe956a463cd4db1c70bd804a1af6f71ac3ca5531c4de61f6dc182d6a29e1f7206af549c2974c4d7c02eddc562c7ab7e508616b86a2d3bf060c2fe2c8702ccea8b7c6417c98d4cd0a6ad4be8483350f9907b1d13a563a8f5b5d588d3927bc32c53a35d5ac317503439c9e56ab29e4ad8bcf01ef0616a8b33977054c1ae67288003baced51e4dfc8b5783bde97ebace9a6ec646ab541d94c046d6f2e7656bf3df52d86fde2a04fd917b310d7e87911c92aa392bf805b5dd75713650b8473e8833367704770073b0a5312154eecb65a4a1e7bb054725110abd2ecebb8ee88471d527da07233d8955c2b4eba905af8fcee7dc19b0f3ad78b0d77399fa7272784c4ae15b6e00b84b7d7c14a32ea207116586001f7461f7375648207b50fdf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h1ee16483c90190376ce87871a04de022c2e3fa94dbc56944b900d58d719be682c3aa479a37d3e5a0192d9018645ebae8424fe5e34d0a6194aaf4e7aba178b03c51cead7daae80a59931178313f77a1c62b48b0e53f1fb1adc9f16410b61326d33bb8825607a697b6954b2b5816f1c9dd186ebf463e37e46b9e98249dccc75fe586b8b2ad48ac9bdcc2238c3ea56e25bd78f6d25880ee45115484fa12614b2828724b7d723ccdcbd89dedb61ac9b5a8484be0be6a06a284e8dd68926a694269b2da39ecd61c84453047a3bd214e67723baf38eca3c5e3f464c1df7c1fed31d8133359cfabaf5f8bc292ddb93d539edc494a941b14141613902b7e1efddc54bd47f4dd955ecec447a7dc3ecfdd6c4e483be287896f275f3a9bd4cb876407a56c3ec44328fcae8982237463c7edceaa018aa6aa02e4567419ac4af8d70128cabbc946c1ef2837da25498c65de563e1e4721183a6376fb513c65f438d518765f95bce0bc21450a64ee6c9c14d4efed585f409ee54cc1b5d02129a42908f29a6f5dc3a2b51668b07b637d543cc3740dda806e85359d9006515617d64cdce849633ea59592a0a3a5527f1afd956e82b23359b373c5c1cdfd2d3bafa076c70a8866a4c6bdbbc2e0c050f537d591df2345376930b1a8bde9049b6ffbac306309ec8a1af8c32a57d9b4333cdcf118ce8cc5b273d784be53492387d7e4bb612475b66336114895df829c987e8ea55e6f106cdad2629a8aff2486e582e34de56327249c426006acbb3311f5fb1a8b164c6d09627aa0e260a4324a680eb8bcafe23a1fcff5afce8144199cf256280599601e0935c5acf28e3cf27c6529f59ad1815ed7b7c8df9d17da75af363ba594705579397b8c679ee905318ac3176620441be3570dd36873c63929548cdda7986771c3e45790be91a461fa44a213d92cf807d8254221ff82693a78aceef99e3d5092bbc908e46daa75bb4fc243257038838365c1e60febbdea6b32b3998bc89fdfd7b2cb4c37de7fd0c700b53fe1d069;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb195f3fccd31fff574aafb482c66bc425aa681403b31c2824a2863dd01f29b682c6a80787dee5981bb00b0ad900f0c96305026577b2289bb670a939ed3f34f4d0318e5f6f389c5f4ff74a0bd85691eb19db5474e1a903b371a225dd9a90d7cfe0266fdd4667108f62ba06c4ee1280844b222b91b737a67d8b9c6616ac84a09fa7c028adfaf05446583808f69d65e1f10277465d2082e1f3d3c5343aa456df1dc0d092722dc2dee6144986c373ebad83f0b0ac2ffdbf5fad87126868878562303bf5b227c3a103e96c68a4fc64d586ca25717172b18c5f54518ba6e44b389581b8d25fdf16fdaa4203766a3b0019fd5fe3cd26aa5b66afabb56d098ee2c21583c053945f56e975bb023499b3eb77509fce7fa1a1cfb0eefbabcbf1f0b6c3e5424a67352df16d47a11e73ca320a5890aedccf43acd82884bc4123d18f0c886411b844f27596efbbe791a01194f3cd054de9a429c23be2b281519b17ad03e9fd7784fae2b88abb333a10328001d250cef661f05a1e57964315bfbf5c9f1e32caed65e8260a62837cf1dfc0267c7f18001d6009f2320ec265becceb2f5defd3c2f4097770001eb5f31f3876bddae2ef33047f419891f4353781bb74a64310ae978659e7eb2030e58dbc0ccc4e559347c7d6ad07db6dc90f5617b8116b44fc62a6040c5bb5073f3f40713dfa4763aee12b1296d9ec589dcb6fb25ffc66b83d91c5214a399a421967dd74c80aa6b7f5877d0a970cc7caabb2cb3c1221eb7deea135dbb90cfdd0c8084b01b195c6ab241915a0212530deae0ce604c6d58425ef942806ee992f601e3166cb59dd27550bc5daa55acf9daa88f0a036e5f8efc617406fecf0ae710538b18975054e501d2584e446e054e2882e3d3d8c910ba63db5c27c6dc8cd41928d60276185f13577eac11c6d4533cbe148bcadde20c7a675f1284ff1a1130cf399b64eb819d482ef008f657e9698dfad7892e2823047e40b4ac4e9ee14c825239a451a3175e839e94f139abab18d44ca57eac652b92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha165128468a877ec48d4e76589fd49badc41351bc020975a81afb42390e25960b15b5401e900523ba4a84acf2f0575a96c2f0367c12b33df25195397761995cbe77f8d4b4c3582ff6b97df031360f42df44abef1cb0bb5ca4615d3e9047d54bd4d3635fb0b412a586a1538471db712caa34689255e03385bf5b7fb3f78a782ea1cd29486f7a440d62178fdf4b882c8d05b355bdb8b849f259b532bfaa639347348a1c56b42aab811b03a3d07c547af941eed0e36a80c73b33ad524079682b7b2135aa27a64f95fcf02746b558d695e0eb92ec96a719f3b6e59fd1c01ec5fb34fc221204fd351d92ebcf8501d766ff3b935039137b6094c19442867dc2f49fc65a8271c51fbb3ee665f746bc77e86bc4ce01e196b51de0a990b4af29e81f4b1be8ed62de777721ad3fb0ec611e24e81186b5e1214ed146e1a237f77e7c995fe7b9b343a978f9b391518c534b210603008cc5a2b4d64db99dca3ce68f6e5d010842cf9c15e530cde024f60f0d449b519c003bb05b10c267b5113e4c06cb605e2769c9c74ecb6bd4dbd16bf0105467a3e3e7c5f2d2eeb4ea1e6ee384890b0303b9cac4f63f1ffb73dca489e0c4afff5af98b2c9492730b48a2ccb04fca7d0b13821811a530e226c45d4309c8bd3b4a0bf2997e11581df3e6c23b95ffa96acc0e0d203b37c0fb119bc0e151ddb778f7611d5a691da202b416fadf74ca724ac93ee1d676286ce6e080d13230f32312d9021f28ec3a371edc04d9618078b975604166800bf68334eacc0376ba773fdd07b2ffe776ea97d893578f5546c42f2c02e0408c2881d7cd1c0e9b82675cca0a6e0eab61e87430b2efe98b43d638c94ca5670e4eb26331fa70cf4c130380360a72a81b2513f08c3ad88dcccac3c6768e2b3b967f91d9771fbfc3e4c998b307aff34df31cd359a2f2ffae8d1764df957b920fd5a85ea1f8606b66061aa44ed66ea43263aa576ce6f5a383e9e887b1de49764689c11c28eedf06af60b4f216bf401b80d74e70295f95bff03f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb161a5218fab10d4e2f0047183c3bbc7bd12dbb40c0ab7c1fdd32bccca5c666e1c3858c630d485e40e3aa22a7a385b5f21b05d600a68667d3b90009970786b4fc8ddbf78b65c7a5643290d07c777dadfcab9b22d183fc45dd6695b2f33ff7d840e7649f45ce3a831132f3d86f01b672cb38bb3f6581121b324f4fd17396e80f05fa1c774fae2dad75663cda316cb81cd7d939a05806c19a56a0d23b7c6581bf56c835a48461d75b8ebc8664f08d9ec2c742bac341e64276f11a6c5da0e6f9af045ff10da8989b727d243ea6c5d992e4fccc9ff8899cfa61168e578cb8cd73b08c3f2d6b99f6826023471f8576562e064303b9022be9aebc07f97e5209ce7efc99374c7938098294783d2c1dcffefebd9870dd41f3f509a587a032193d18e9e5a138496458d18f2fca6236631b4ad472024cbd6e04d019c8824d5712d26401b47b1233e861e6def8dfb3c043863f49d346d45a836892f8a5d3c8692d7aecd1b53ea48c5fcdd22d4f38ac3feaba80467064a90d7dceb111bd8e06bab8c9b4dc0d81e2cacf02673e793558ae04331208f5b8305b5282bf13a2ec9b808ef3ae58b6249eb0d28ad6064617e75a38e5dce452a05f9a6d137a4759df85de148451cc686a625a661ca9a2360b8f68300aaef620ded09f0411aeee96a9f9bf0048a7c9c829314f04be1c4d8222cbbcba84aa5888a26183011ac62758ca36f79709bac53536cb66fa10890073e1d665da3c60347a93cbb672376b99c800025e2244e7447b18ba541d1c2bcdbddb02aa422db818452a12ef2bcf16256a85fe17535c1de955896aba833d60f15cdb2b9b34369257c51bfdd005a73c07dc6052d375bddd22a4c434b3f70b632eafddc8083304731dabd2d7ae133487649954e8542e29ba33986604d6f0dd4c02e712e9996c7e9e399a11e438b5055ec12b5ba54811d1d4bf7538d920ad87906293ae22f97396f88074e63215787c469c729e98c606bf18c667bf076f415976b5bd07856f8b50e119cc4231c508ff4d1cc2642;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h76aa21c11b8126cbcd86b055942758e36db3d29b8080e2c1fad2d629edbb86a13d9d3d2e0c518a8412323b67c7bcc1b450a1ffd6c21acd5806e76003578860f73b9783392666de2ea12820e6ca6696e3b7002b062d088c0e5c4ec072101d3e83eb7864f42f58d5a1ff3e5e8ed406fea22764a49dfab4bb3ab9975e3a488333ba62d8bb66c58fb657365fc5799569fd73f4f9932b9bc779b1112e10c1153c2db569f7e871661b6b3c3ba1a40797948a78fc3f93345aec91d8bcf967ccf8c703d936a1f3196839f956399f95e449f414540f9b0017b2fab29164030c6f68694ccc12a9ad9a4f6e04372e738c5b2b606a2b2e70477cce46291376c28558be6cb2e7308249df2c44fced6d53bf47545a35c7168ac18e81dbb1bf63f2a7ecdd86ba7234b1ec56747c6d2898d10c0a689ec78db180d2ce29b28526090934d61227403033b97fcd4721311c109c0fddd4b2747b9e2c23297c3b33d08a22ab81c52eda96f07ea789ea2680fb7f68e6967f961c682517f19122d39242ffdfe487ff77be550dada194b9f10c4cbb0a971dec7395c7065777d1dff5e3700d18839d6be461b34f76dd812096221bf9659debb04bdca9f382491517ebccc1b524ccc2029d7742aa2b1ec860093b82e3cac8a6c67398ef332deb550d2521b155041631d8270eb1cdb5f42014725f3f9b6a43047f3ee3d6cdeb68054e4d650f194f944fa824f11713625834e40bba95f708f1a1e59ef2a25310840755e39baedaa5184d09b6193b4335856d58a1cfed4bfaded4e1c11ef8f89cae93c482b11e1dce03841ddb64f3c340ee36368a4629e1e9c835c8a244a35bb3e1bd6d98524f22c3c44f7787a536de189c50645cb431129a69e64269a61508d7ae1983a700aa08090a214f034b00fe6dfc7d8e180047df3bec6930d3715fe3a2a981421b3133afdf4d45d7b0bb239550c994f5321fe52ef435df6ef6acd1555ece4312a7da63edf04872e7f8795d12c3ab51603bc3e59763d0ce1a7f822a69d26c3dd7b6e47bf8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hee46557c5988f2520994698657baf3095f3b41140d42c9610a7c1a360b70ae81e639a3826ac4cb2cc975fe1a17db06da0bc16424cab1db6803ef92fe972c40113ddae89ed81c7ab3a4152268d3803c7af19178c5f4a190169a731949a39412731f836db5f19b68cf33e651a73ddd99808b94da4782068a0b3692d168c1b482978a49001ceffede5e9539162a478464bd0d3dc978fa520688c0640536a9bf42e18b8b69044c92f318ff06b11118c207410f8c4136eefd2947dc9ca0b52f76e9410debb1989d1b74bd2cafac47cebe3b5d5ad03c93fe2aa6181c61e391dcd5ba1d344221aaf3107b0a81d5181f4d6460c44b48bdbaf3ca739984cd066393f28d417c1a5053d7dd02097cc9177de52bd4c28cc6986d855ffea965b90d1120f8e0a1da07892b8cb48eb6ede9ba79d26d2b4310092923a57b48ceae8455b2d895e8ff2558b00f5f43f5a56b24cfe235234cc007e91b480fdcf4ba1d87420fd26bbaef01f5f25f0962eb86a177ecca8f38699465780b19f15b4a26ba2ba3dce0858d7a9f7aee8a5925fbafb60d37effb471c0f7598f406adfb53c0e53dfe3c0ac9373f8a6ee9bdcefbf37fd3a96faab670e5374565e32b7ca653a329fbe289abadb69935fa3278798a49390d9ad6a15a63cd99ef6dc31a2dc6ca05a2234890d024fe6f438c8d5b9748083e29ed940a5275d7b8be7f3a8b149253fdea673431b40e159627083096c288f078d999a073be4c9e0e1ebae6f0edd4a0e2456dd840dc813adff52e762c637d8665962bc19b080ea5dc3c37ad7cb5b0a08ff4c2236752493734c23849447b4835af536be5460dbb8abc3da23f092538354be336bbeac8ad15cd034451f7b0cd51ec315bc858f11295cd1d57e3ae93608761dc7f66c301205321c2dfa9fda508a44d094549492f94fdcd26df9f149be4ab22b5ff4a96c967f4b96cfd2e62e8e4da7c93bf8b738ddc469a6795ef486e65eab9cbf029c91902da4c5c286916df4cf7f3e3005497ad48bc6974325cc6318ff6c0c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha6f50cb1113b73661d57fa77a359a6b9060012620d596562a2238008b485d8f7722281b00b8f366e78805282110cfa6b217eddbe7133f560594d9ac1ac87972e7e2d47a19d5ffd3f059ab3542e38d3370f806443272c134161866be2ce1c780c96bdf9a0e8f2429c2e054625a195c970262a2a61702719d94d49af1bbbf8ac51eb14b6c833c2f5f97973827b29655964c447ea3d0b7c93d04555bb6a35d2ad4c380a00f0515ee69f215b518a377d3067a072950b507d81f03fd19769e91ed5971eb9e3366fc53f26fa389187abe99c6b2f38c00c84a45282aed264ea728d9602a3f9a818d2099345702692057f901b6959fc05b45d68e7b4d735470a1b5823aec361ac2cf58e3f53abca5d87ae00612363173ca78a44630afca2b006bfcdea5c6e4b16b53f6af2169194ead5fcfe897b86d2d6248831c1e1e8165bc4fa2ddfd94a2de4da78d678830edbce40d5997198b80db025ee9e2a63b568f5a43174fab26fd912080b300ddda76ebc835af13bec0f5f2edd100860b14f389937a95848bb6bfc1ce3643ea47577037899a8ece64da30b43a4ed9b9e42fa4c91386e1b72c976bcaa26a626cb54337d1f6b29830f4768f1058a055748ef3b7446c011f60923178c74f95217588e6fc1d0cbf3d8d748d9ef147e712e7590c64c53bd795f2ee104a0aa54338324c41e888ad29158db17b9924f833371f46f609c098e7634ce708835c65757d2c1212121b06a689c54bd39897ad347f4ed59c5786f5623f1766456e1cd7ad741f2dc721a9cb857a660d0d7657a941d93702914c48bcc7828a494467589031d9516457bfa16b0375e74b5115d3ea3819762e7b145749a85334e97c1b6e19043d0fc263f42c7b5900d48ca66b8fa72dc2514b271300299e1ab7efce6796b80eeefaa5f35ee617c83e39de024dc662136974d6426ee1dad3472f7ea0d974fe44a33c0976111f189bdbde3da25310e581c43fbffe4a7404540ae5d4cb1e65669aafda50e64b507057dd55a6b453d1b62dff4c5e298;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h35df7ab9bc2f55896e24629da3d0d304e8af5f7e2fbb3bb4dd7f97e6132533e74f405ca6a0176c2a4289f6a0bb11c62b2727cb38cb5b9772c658e61698cd0f4098d4515dbb16338ed473aec4989c994a90e3c5e76b21dea8ad7cf2d8f45104d45edd684ec4379335d9e5f62326c5725859247cca1f081d0c40cb24d97c64b1945f3477115fbcbc0a09c0b4bc0afe7925bda0e9d652400febbfea627284fe3249679485ccdd25761da525814282778c79f319d474bb1a782c4da0dd21981d6de9cf782e74c2a8dcce0c62478abafb9e22a10a98f6b9f269315ca2a61f7135ad4fc3916108479c4f21d21d5d5637f69c35b242b3893cb01797d04ad108a545a483304ff911460e9a868c5dcd275ca7dbc6c4fe1eefecef2222f66f61a862273d2945ba562d12e875fde9db2bb5bbd3c2cc018b06f4eb84d72741b4ab07cbe9cf7847067674b599b0ddad799dc72f99ad6f27296cdf581f8026531407b3e2908304d59d46927f492a73b1f525b9cf0f5346995801b1a047935cabbc6e22b39e2b601e647c03ab49bc149cdc6cccc26a4a0dac0d6e5624f2069703e30929526ac27dd3bb00bdd2847aaa1af2862ee39c50a0590971173f902552492adfbb541504fa697100393ff0cf54f480bbb5ae7f9b93731f3fab958f6eb3650e0810a1c80a2f25bb2cad541e25b462334438780f24e9fe771fde0f23f22c8ee3cc3e7028b9b992e42cc1943da09fe8a8597d79731d233187c7cfd54de85aec3f3d8c96f58d531116f85deb19db8f7644972224feb6d0e3f8c88fc0486a75f4bf7a292572be805190088ded1b0e3bb85f368ab701ff50fe67de1ad6a6133d16391a688afb35954c256a10b5fdd8fe1d0329580a329e6d0011d291febcd66b8256ebe71c8ef20951a8568952cda6243642e884b8162c5639ab08dba17afce0a4c26a6d25c5c0b12f82a6ffe10634a2608573800b95dfe4c4d2bb7616b6120e399844809ce7f3d2055982dfb9e0b815e11dcd30f124e985056ffe3881fc5675e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hdc1a7eaf853b15e3f21b5ef0766c71e197e4047a0110f243d7a072bffd4826dad5318d5242edb92a4743af6073d2cd23c09c7ad9e93d2367394f29643a20acc04982338e9dfea38dfabba2ad276802cb2fba6eb57bcfa52b80b2937705eb3c479ae7d0e4ce0a0f3bbb124ac76889e3758d07e73a099a881902b15ed9cfdf43b769c2f97a3c7ded014f95dc97feac991720e8e1fbc7169621bed8d0983023890e65f111033a82204a7feda89fef2ba3a5daf76f5dd3e92c0e63775a2038629dfa4abb648fd55194cd4aabc805a508b81237d40b687e33045b3bce8d57f42a0d740f820c0a04095514e4dedf641eace1d4ca0048e7f1c86886a45a8eeef2e518cb87c4be16404833e637528f30111722c7941355c4eb7e528ebeb5179bcd64d1b64e6dfc33ce969ed662a44392fe7dcba2bc6065e3db07b54c1f158986ceb41deb9e1d176ca569b301f78bcae48327d599ea13a5ff9ec83b64a9cf11ddee7625f0f4fe9c9701dc278eadd0d542db244c65f33d78e0580d63d91a3a7fde3d6337175cb6c9f652252904d6170706b7f56bdbe05b9664ab7e3ca4fe22b444a194b1b51a1ab310928ee2422a00e1b725f29d08d9b17ddf5816b69eef3c440303ba04e46dc628b9789d5246bd65707ab2c3bece57f0eccfbf79b4ea9d992c66fd69dbfc3c940825037dde265710eb0a6e3a50f2c032ff682659189ee2a596623748e17d047a727ff8faecc479035e5d85337f4587ceaf9884b09a3781dd29ed9d5ed395acd0e8ab5b376fe1cb56140bc4998124e2fab7d9c2085d20644b6287c4139aacc30a44587bf7ba45cdaa34b7729a49e204d00fcd87b8b5640ceca0121cbc48191dbe705133a956e16b30a12493c083312ed3e65c0b6a6e9358a863c3913f22cf384b7705ae58e6f025eb735ce88d85fa169bc243cca1b2ffadad46242d0184547249af6659f54ffcf58ea9cb83c8baf087348263fee1132a30dd6c4bcd49c40b4267cc755a8384976e99a712ce7b451638007ce170d4b98c8e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h209c1cfac045aa4dcbebaa0c47534ef0600e5b6481081c08fbc774ebf0c033e65111817c02f7c5f9b4f30146241ce80719d09a0a1f5243bc39cc85f0596234191f6dee8aa8f33bf27d9010116674fa4fc880fa1022307b314a978e3ff922b627964a1d0b1833545825bfb0c882929109b8b4ea13731c2f3272ca8a0afa4192833b8ac441d42cbf77223418415f79672ce3a5796a5135f2bfb3d34ab2e5343e0950a3a059979c1d7c2bdd13d51391550e25e038dac1b7d83edecf3da0bc7d878614b0239968877e03e0e65799fed68675e3b406a85de713f5ebbd193b9b17f503f123dda29bf4764c86677f01229441a01c3ec6bacedabb89fb3202bb9c0a3e9207385235cb491709707a7d60ae57c21f659a785590bdf753e59574f42e233b9ad8956b4ba6a894faa35b4d2047097b39b5ae6eba88116901d970234ae8ae312674ad85827fc482fd5a89ed1113f5974a204f2dcf31fb48172d65796257c1aae5b514d2fa35dafce60ac88f287211a4fe7caaf9e893334c10813dff4c0d6156ca7c00751d75b5b214b27df34548405907d5955d7eb5e3f1143acf2425a2997e9f628d57ee615c002e3ca8982490e4a1b7c50269656d3092d2accf686ab1179a39911c3d8296abc7d7c896455658d7a64f20f7b49f69e31c3142e069e55b01d0db4333742867a29d05def4cacc9e532921897b300fe1c449ba731480eb4d6d073ab1080e678b2e5079f3285b51c39b700552ba7c427a136d4e8293f2299474fb9da6b6ab879e5de722caae6aeca650f13757fe5a09b7b02fd8b7e01a97682dd092a0d0d292813ab696ba59a45911b2a489cb1566336d6c82c1b6af63910b19c5b0368ca38a8bb28a8f5427bdca8efda244adcb64a83bf1f27a2130586570247b87990134bed88fb8e0aca170a3074229c63d2a15460f35a8f62a99002eb18047b7c6a0c794824927ade0b4204849a86001739d4918a386a61af0d488962c35548a685a309581d05c419d6d382deaff210000cafb3f16aac52537;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h9211c8964509cec50780a03f6ecf442c535e39f7153bbb1a393981a51e36b936c3cf658730cf51e37380103d36ea6cda11009246784a2f574f42bfac349c2ca050f6b394d0c8b4f7c55d62c670211bccdcdd6617dd88175c628088fb5db4608ecbfa04b2e080c804434e37cae8cbac412cfec05bdc981a3b27faef8495ffa8cfc527ddcf8034b852c864a0553534aa0a5ef9c349f3ff90c3a83846c2787aa08d9822af76f4c89c8aafa90b3034a6851fb8be58a662d3fe39e9f3e80e5a2fa16abbbddacdddbd789d8c7970f1d5c3183bfb694c3239c387ec64bbb7c7ca7650acc20980e7e442c5b59a05ea766e6390d99bbc16b590c707fcc6780709e6008dc5f011ae9276d18623ee7864ebbd23dd4d8ecad2ed7e9b5549fd1e675233d2f490e136901ee976f111fa766a05cfc9a9bf5ced73864637b5f101dc0f9536384128dc7f8fe96f9b4c48b2e0ca8aa33c95246cd39cae40897212db80e6898c2f10ce4288b244df4b33d39a4a95eb54b1b53adaeecf982b04fd2b2d4f3b090cdc2fd467f9fe545f0f83320ca984f4d9acfe8c072438da881077d9f6ecd2252d7a8cdd91ee9fef3b5dfceeda8b19739f638727a7e8db06ad094c6083f14031ddc9913a34b568176bc0e6e8282308bb91b2180ba7818edd359a72d4039cbec85a746b4a04fd758329e1d5b7b32e2388025c1fd5ed3fb9dbde316cea918cba3d90c4f0f2838629a6ddfd842c8cbf9df8391ad4fbe37673bfb599c726ed5a6b74566994ae2a9189c0eb3f38920c2f9dab834fbf69f399f46dfcc8af4a42d08f53ba731d0c4a1761dcd90a59dfc9c147459577bc15a47627954c2460ac50db418d276dae54e4c07b85059127c84d7c9b12b88bfe097326c1832568c329c0efe01db0fb1f12f6761a9420285eebfb2eea9cd2583412516d54102ff8978814ac9d89da00749ea506c4389e6507e34b0f4d1882d43b9b3305e57484850c3f5b2fb28186019151eee7193692728a7a256ecc2a7aac0b8a9f6b1229fd520c9146;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h13c423e26fc63c8891d94a7561619f655252c1a8120c389fecf99677135298588e326948a3ba41f8c35f5fc15e80cd8f6405a504951d5cd1447b51fed04b31ad171f2bee8b2584c5d47d4a35b926894be07bd54ceb941d86031906c332d39d539f01a9bf8db57fa8bcc34cf5a040257a107ea2cf712839abe592cb79f65fcfa7cc67390f6dd751d52c2fb9dc85b56646f5eca2833c7e9b4b4901102178574e53e5bb9a36c6560b7953b4028be99c0d18b494e48dd7ebadaafcb94d9e2aa70a7559613ff1b3b40f35d96652110c1854d5ad1dab3736e46db5e83152510bfc1053950eb748df53d810cc2ce9a38bcf71da904085cf4e7b989d1983538353167089424aece8489e8975c03f517ba036017b015a468cc0905f35c8974a167feb8eea20bb0c62ee8ebcbc8bba747874e8cebd1dbff9f3b4353287350848468e4e3e1b98fc020a25d115cf991d11e58e77e0c062d9fb61a1c7723cd5c561f3b900fedf0e89173442ab3b98d192261eaa4536a0b591095f5a5c1648a78c83a02b7eb379847f329fb925b44f0a387c5c7660f5fbefd7af899dc0455f87189e92dc3537a8cf6f8f42705fdb47964703a3458af4ab6c611c5837aa6abacbda72b05a8655cce70b91960ff4817015488c992728c107f4eeb47db04f6f251fdcffa012250a34d7a49c69ead312febdacc0782904d99ead5685a6ae56555a70f1c30e7fe5519f19a2edc641eb2e6bdf3089d17d52ebe506562d713263b46e96445ecbeaa4d42d35ca98c2e90526ab37dd13d2b8c8947d77ba6d00c9e2cb6f06049881e2dc33c5fb8dfc8275cc745824951683c6f43de73de7040bc05c129a00ede6ea2c826177665283d85cb1faf042ca5f2111c2cef9ffdcc8432061db4beefc79c75bbcbde75efe8c7165702ed0dad5025944bfad3ca4a5a45a570af217efb7fcf77c44d0e46619844d8f9779b88ff14a66975771cd259fa0c5031866022b72befb0176642c0b13def8b1e6bc5888c362eced43797af81fec73f88b8667a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hfccad176795689dbe7b31206b039db959bbe12ef6ba91690f9af8b2c75af6f225a5dddaf6a9b3d4fd8f048f09748dfb26c26435b785e8ec59328448d19541549623d46a5cf302f096fdca821614c400e47708b5b30c02fcadf8f346aa97ee65d878982fb6d4213cb8edb80d847da6f506d2364baf10086b21c312940a43c23bdb4ffe6ea16d8ada73872c3c2a11fbc0a90a4815b83004cbeaee0243ed229a24af394948ada0cf1a0ac89ce1ef06a8d6c5431e710848c4caa4abebbd6b7a318fa14495f1d434446420fc76b54c9f44d18dea99088ce4806ad302d8a3a29a61e9ae39cb3d07c2d504fe93c1f62a87f691f169113fdb1d3f7da33c4df71b6ec3a8cbe73fb95bce8bdc739a6bacae8718075660f6260bf9926e27a5e89c52f7d155ca77dbe9290bfe32dd9c5f0a63a3c8de55bea7bfa68fca9461db701c0946a66a749d83f664f4686ffcbe1a4ca6c778c5e567e8a2735183fed43be57df99724de4d94467b35d41a3713d4fb2902c29b42c7c4ed32fc53c9d134c19b5438f9b724142f94a3ca14669bc70cec08183e324147b6e58326015437365f10a9d22c389d8538edd8c5b7792056e49646399146e4147d7f64fc8f5fa3381e88ac5a4129651496495fcef80575586272330d39dc065ae4556006c8f010b818766496744b338f01d8b8db1b5302db17465eb6ecef76a655fd2bedf79612b730b302a4bc64babbf08e4dc9308bb55cb28efb62e60a1424f818ade459daa31543ccac708ad099e026a4c17ea9d9f2e9b0657a6d18fe288694a7fd795da3892e88ed3611a25dca89f724f0a42b0c30e8253cced316998da8fb46e6adca733c0fbf3201cdc6be982ffc1c082856341a1aa7faef6f156de518e69729cbcd265734787861229664f2544e6c233136f659107c8ddd1da1871a1de2873eeccc33d3abfebefc4d6e9b9d70853a882273720ed2732206cc4f9c6ce5b11dbeae03a8b03255f682b010216794ca10eb598909c4bee52453e3143b498c9bfa77804084ecdb1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb89e3c71a8679d4a14cc8fa594b5baa46e950afbbf16fc3f4d328125b7c807d01c3c1d732e7cdc9eaeb49a705fc141654a695491426b14d0caa41493a5025c87d1f521e3b0637dac8b6db933134a166665c8529f68511cb038c6b134fe710c202fc7437dae4e5b461c57dce2792a7da5b4db3e4bd5d750ca3bb691788dc25803f1d11b2c05f811ad78e3702cbba204997905619722a0995d58673b275e978e940a5e3ec3a3deba075e6e3f7a278b2a04c211e1ec0c3e373046728a5abe837fa9287928ccb8ecfb07fa023baf0bc7f783f55ceecc9514a980e80b4143dbb2e26222885c088eed8e04274cf93fc933fe739759c972236e3f4ebb4493b7d0086c099dc836040c2a27aeefd5eaec857a9e08ce8ee94fb69ebdf66fdd145a493fd2549f067a4d612729ce353b9f45f6f431cb5b729e0f663b59aa8ec7234cb529e9427fd2e2e29ca2d56e65e94734c2b1942677835a7b415f169a8d9565a618499af3d692461c18beaa69eee51a153b0551f48fe3d9460081824406013887cd4f80af3a35808e8ccb8d79bb58545cb20311cc0c0373803711fbec7099aba95a5c211af6441131c163c59e54a18c5333dc8eb3cf0778bd06fbd8e3576e631971c35aff85d2350865302dbf58c0be9c4c247f68bedb85d8b4f640a03301bbd75901a830f8c70d85d618e13a665fc6ef77edbfd9cd0b5d763e5249a88a42e5bf48c85837e1ba0dd39159892aa7cfa889c2ba3d473923ed4540e3ac2952843d25d79c043ad7bb08110c4ea022756646c46466bf1e5f1c1e3a8705c19cb810a82f6c3296b349f8e8fc620118677841fce6389f7fe8db253dda8459cf4a15b991fd77e6787990bc9d9331b5fd21c81601f950aceff32a3e8fd23644e0970f3e612033ff775a47d78efe3978ead7fc0e5a5ea5a2990a1244a54ca8551a16be1b37d681285d710dda035f5d26d8c9b108a73555e2d3fc243a4b58431f446bbd6f443a7ae99191a245799b4d6424f21935feb4dd4049ca6713cbfa447acc15f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h45ec866e145af0e24ed295f405f76d4027869d647e0e9a136c0f135169d4bfcdbb03d4b6d5f0e7f99dbeceb7620420d1a54a55255e79578f207584392629ebc593de7f83cd7b61ad352156989ab47982f16fc6f2a6ed0716cf6bc553417b6b6c6f4de3fe6235056070ac7bfe0355f06e1250e3a15c32fa889c5f5c57561da6c9f5cbc9d3ed9a812ee625ebef9185efba78120d866a07e80efb70d70f288859c16dc0c22d44c87cc24deabaf2b9b2b1461b0eab60cc3a5ad3ef0126746ea614570409f396c8d269f3826a637206694a80569f6ce6b3ff666332b38ffc8c3b12984a67be3aaa7a4d911793ceebc4a4ef6cba252f240e83844ab44f807587d5d40b2c30dde30a5a1efde726e74ef40a32d3535a3e5c0060b0c026da857efcb00cf067e629695cd154cb65b2442b965b319107b75fa12865bcb458f58cb05e47d42415208520679c66f0b520c67fdb74332c6b9d6b7e1b453a90ffc77da248aada2417d2a750cef3b03f7596143aef46ab1caec7319a9e79991cab60ca8a28207df80b20a5eeb35c29564b421de6a82527f346fb2bda1f6e7af23cdb6f673ade4f022dd1a963438242b7eb9d3129543693ae8bf7cd00f7e3e7edaf83672bda41ac88730264cd8bf079c16a2a19273dfda13666bf2deba1848f61b0da201a3144ffb7a5619a376b2a354742f2652a70025d66a1f7f0a2a772ca99a820d20726f249ca4d0be26c88b62b6db295a2b4070628323764037ce28f56225a03e6ec8a7b69335c6f5536fce58e4d9439257015feca9637d08f920fe9732f7a0b1e47bb432188098d739031b3e889aebcb37e86919805d1ea3140c7544a99329165062260d5d816e7eaf4a7d7aa37f4ce608c5cfdbb05ea089149b47ea1be2bcbe7fef4475a49af6f3aba6d8be9aa86c974d488c9baf03645faa3b592c6ff4faa425e6f864c8491d4db6f7fabb0e9b2c4d91e6e82e47db0c7e904201258714833100c8d264bed9bf1a1f216ac39b9bf4fdbaa7944a540daa2ad60faa6ba4750;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h9c63e2ba56aeb8ed7501c92df5500b79e61ced5071ff01a8d3fd3ce08a630415ada92968ab5b7d9ef405ddb91343ac4588143c97aa0e9b45b39147f762a12b5fe9913d2274caef238a519c25b243cc0519c609ddbe2d808aed79a9b4982875ff27e0675e056d3215226e635e39b602046377c513f6833324834065963c174d9d432b103ada69fd19770eb131b409221138a28b4c99eaba2b225ce6c6a7f1ce7534b9ce19c31022a86078904fd9f4b8359e980811771387eef8803815675e9c910ccc8e10fb7811105189c3c717577f3fc765d97454a8f7e10e9ffabe91e65f99f3ec425f98190336b9bdef94875bbd67cdf5140949b437c11d74c67d4e24e6e7b8be712122919bdb81b1da59b557c9e64713e45881d8a1edaaa5c6a4af8270578d9ab2a825ad8bcd73a4e6bca5a6cb389bf3a14be5a0c791305cdb0f1d1acceb1efdfe6a4c188c9e38a79d5836c44ca9177ab8afcb737c8aaa97a3a5eabb01dd573c77fdef7ab876327d11c8fe14cf8000b87ffa109afeab454c0459baebcfd2b576597d044a9ec1c9361022998f909413aa2e14ba367b0ca971ee7951632bddbce48ba27107de88e43fd02a1d67f08dfce8c1732e956441287e077627df2ad03d3affd199ae79f3aac4fb8d6d207a966c5e2772aa84a78552bca518b7e28d9df9f5616b7ed84f7c99d4b924c9d8d145fba292e51e045367cc3547f9bb9f7f947a6609827a1ac994651188cc41a15564a7b0981b8ede53a8e3e6bff86c5ca1ed01dc7ff1b591bfcecc60a14cecbe83be5ebb35ef4f98b178eba0eda1b06a79d123ebba5c9e7404a58e435b782e07cfd95c36ad73e0a34c9dc8f33a7411466609f8c3f37f92e668f9d9d68686ea7dfbd63221f0245d5cb65f96faeccb2a1a6992de6c7e1282295ed707c32fdac0d155f4012d255f523656d9c36602bfbe1b9236f8ce78220f4db801cce974badd84de9fbd60334e6deeaeeecf92d67e9a56ae914fba8d620010b790785d3b4d16d5fd572577a7be32b122b278;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hdfbe2c8305aae2af006097059a3d2e63f42cbeeb596ba4fa4de7ee50e205bd7b0760c04c536bdc1b6ebae156b3b336962f795237a459bb6c0ad4e9332f6323f44edde9571d11df171c0c60c2be34ad6ddf34fce0b2447b8c74f2428c25d6e620e9c2c2d99ec92973dbb2bd9ceaa57567d09a7b7d0f5548a45629ecada9af53232a16150778bfc00c76f3f48c5e12a54c32951a9f5f95f244014e2ffa0c908eb703c58d58ea5cf59a1a88d8b7b2dafdfd2a632418d59e9c96b63e24bd5bd5fad7cc842490078a733f939c1ac5f06797a72244716e3ee335ad90fd67a6424e8e957db2667761f2c2ada7eaa29dc77e1fb215984723e6c42c6225c69160ddb01f837099fdd502144e0748ecd2a750b09635a8190a84146036fea8b87b8fc93b30b920e96927dc1af310a38480970b8819febe4aa0d00a7d1ef6c2e72e1d95ff927e27f41410559a405b0c96167eaeb305ab34e0c8ab65ab9c310849e7eaf144619aebf6af101482a87a6c965429644e69aeb119373d7c1f2df1f7a176a4c552f4623adbef61d6af2dcc0760c01f1f91351d087d141b17f0d5be286f962bb8e9eff20b428e48b4ce4e3c6d0806b3f5becf1f1ad3e54de822f037cc340fad8c25b41e645b7e91c54293524c9e6e1d182505379b729eccded7dfdf118c5b2a68a374dcbdfbd64b4228fe755e55d4d45a0bf8bd9690e18010050f5a2346f3eaba657baa2ab3f9f35097edf81628a809a39b2e5cfb3d200b14d44973b59de92bbc2b727518324a6a8843427ed98ad4eecf2765f156b62bbe0ff247f17e179a5b336c2348e97f24abac9078b878394938431739a0bc19981ea98ab11faf2a0b50d04e33388a933733b1da7c9d432fe84c93a84e030c1a1348261386e029a37e32404ecf5ec0bdd817cfd8a3e98f098b3b0e96d2cd61cb5bbc992763f5f29125c742e488e6b3e14ad671d4cd07abcdeb2f55c6d5da9d2a0dc1861621fd671735fb1dfdaecbf041ca9033aa5327ab66968316055aebb156f3824e26f7a6e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h5491c20ba2ba697f5f426aadc7c5bcba54c604f1137a0e3c1a832984652cafdd21b08bbfa81538dd1158957b85ee0dcb27bd5fb42ec71f1cdb63557a430b6cbe07bb147926b9bfd3181a4f9c2da8296a49041e0eaea352cf2c4f921b492f202272a81dda9f95bbc5f061f28af3d2d06e0303d1b22e5593bc405d33180e019f29dfccf76e62e2514e583511c815342442b265fce97c97007667a992d75ca10e4eac6bd4b602a64761c723a3ff78f8518e536e171d3c978af909122a7fa10b33ef6bc902d8423eabc4f850f192f94371e137918cb1bbb18c8e74ebda8c2568832a8720b240afc686fc0c727d8a5f07a6aeab1e09efb4bc34f5a736f1779d80553864570322fa78fb4178324af9159c085be16c42180f05b0eb1a79270bf23adbb8a2ff02b28c03eb0f8bc647b70a88aee806f023ad59edc0a5285ef628a5f2acd32263c540f51549eb9477860dfe704152b04f0c27acbc6ffc9d3f304dcbe13f78d74355c14cc9415494a5a87e288333f5ea4ca62bac870652c6f55368efe95e3640c789c227476576bac594298960cd78600d1b66bd58292457dae27b712c4884431304706b1e844a466314c7baaf9396b31d09c1ffa125110614dc04a7b8931a222a1d52923cf41d590354f7e688ffcf5add08d6b13af65743c6798320c73b81334852fd4d9eb6c5ebd23b627f2184215acd2562ded2811dd82fcd422326206e4e1072412e3dba23a3dc453e8686f5c8b71e55e687e25487a7801a606db4ca481b9850d5d144b8e88bb2131395ac8e6c490a22bafac25b198f297c914e2793ac758868f999cbdee8712217394b678296543e5581069d65a619b0fc1fecf86308b7faea447386d68ccb010b7817a475f2288c39d9488e226903d164954a4813f87d774aae5f78ac3b0da583f2d30e3966f114978b7e3dace03dca3d93273ed1be941b66e6473c87fefa4d836f19efe6032796af489cb2a9c7b4a84b2f7b3ad4e46958446713c809c731c117547266bcb5ba30a7c5b90813f3db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hbdda8d868dcbe7958b363fc3c4a27b426a922e7497a72e3fb83d34d3017eba10a3786762a466a08a0490929733d092c7f848670c85e1b92e9e9f579427bafaff36d4d3c1c5af2c812e21dfe5d52fb26390350474252ef0d510b74a020acdf04b0c0083ef8179100ffa154a8647e6c816b40427f1975c7de3913695e0f8af50dfa28a3f5573e2c83dd74dedd97094e1098134a5219a0d3db7859082ba1a7e3538af61af18ff9c78b7dc15903dae7e48ebdbee2dcdfda6de1bd7ba0b74401c4b02e8cd1790990f6c0712d914f5f5dea4d1ccc223ff0ebdec05f570185be661d7879e4268afe509fbea7bdf52e013ee5b4fb53f2fd714ef29027ec2195b8bf96b00e0d7c25c20acd8c13d052ad96e11d4bd8147688498cc6a606765fa22ad74578f3820e5081244d3cd3e8bec850cd044785c43573c86249ddb03486e9ac3dc2041f7235d675878c9652b7318f61db36ad1bc0ddbffd288e56ecfffe2f7d1d79c4e613d064cbcfff59ed0b4bf5840469dd954eae091526d3e62c6fc18687ff21bcd6cf554216ca0239608b431a52c301cae9eb59eba8b2211fcd89f0953d6a97b30b3ee714e25a54d008dc9337a5c72d15e55a2fead2697a4c69eb731b1c225737ea0f7b529f7285fa58ffbe073c3e72ef3deda6930c0b9c92f6cdf545dbb687073592b8d4831f29ed209ee3da2b0e2bd09a8a6c0c352b16a2a6f6b4c7f87654823743c596d004109a87166b472f73b1a8bce15e19c4bae17b0f2bce136748c20b4eafe45574b84cf981fbe5991be6588449c3af134a96db82f6e8f60e839022db081642eaaa1d3157f4d6dea803a3832aa90f84ef410db2352b1d6cc1cb3bfde176e5adf091e8886260b516a11be44c3f3e5b7112a9071a12d7e34de8166aa2336e9fc4d58f7eb82dbea6a1fd75eb3fbf67dd344d8e08d09c9665c3dfb9d1fbbc93ec9f333e32e10aec7395900b7ea00ae160db9c22b54bc6c44f92bbb82374d3d5c0a65a6bb02e842fa1959b402f84ab2cf168f72ddbb2a2343;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7bc70e002eeffea739bb6a3c937655b45923bd2bfebe1e2cc106d54f0641738c5b0298d77d49c6b20e7e2259e4f89880e1412e3c8b6f266f4f5ff1fdd80bd36db961c27b3a7ef28ff8f0c792d65e86901e3f8d7dfa353becea0096c81d637929c0b0636a88fb84a3c8501d1b54f61cc231ca2d6d25f41aae5da8b927e4c8158226a1190ec3ae2c16d25a3952190c508236f06ea86868f36abe52fddcf7bad27861c13645a0520a6974000288103e60eadc01871b4be0b2f867642a101409f89966581a1930ddfebdc3ff78a0a0501604c1faea6693cd386af4cb70b0946e2dfebf8bb6aeb65b278a471806eebe854a6d854f1661d80a96c6d4a3f6f09969ed79b91e00ad81c10d9013b6dd61a55545bbfc33ccb8509df0ead99215f6301b68098004c8a89223616c5045b022524ed0fc9197e5322404c585718dd7cb1d8a5ba0c20506508fac9b327efed41e57b0919b0a06dafa26fa128848245a7dff85547f46178de870593c4db07e1750bc151136af167b045cffd94d003c3ff4ed75377e901a22e682e0b81e666f0a8ea99b149c154b0d3190625ef8ae7946798f888127a1dd9eca141160bb7fabe62607d2345fb0a851b4771906b44bcef01ab3edd62707f2b912a72b78aa4811759d0032f6cb4bbee2a3d9fc80a226beecbb8d319b083515dced5dd087bab0eca2d17d757c4744f5c582c95eeac1c8d561b8c2dc679619bd7aabb39d86c4d719068c7538b0e6fca583f51fe67572d8a0d69ae771ed0d6868904dc17f96ff8111dcc67982bbeced01fee8263d7f5d85e9bac04fa9bd6e916694d771a252c5b223fe2a5a7a5a1a62ee30cb51eb87c1715c5d1c7c65f24b07796e64fa83321621b8f6244fd69d632e3ab986086e18a0ca81689f80f74f241a8cce099ea221ca6bbe47369333cc80707da097a19d5d6f33e7cbd66a75416db8736cb1c14df1a2531acf708ea7a803d7b2b8662f6c08ea17fa41e4878e57e64d3ac7b69292827b901d2cf1f4d5da657327fea09b25925641;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hf691b03d32f38a9da98e646dd94e5bf612dc17e955c1c82adb83c7126f92862975b4337c3a4a077dafd6718a93646bcf3d4d18527bfc1f16772c9e42d13d290a507f5142114e838fb6cc8219197cf457e5658c296e4bf65fa112e924c20258cb37b61b1ae2b3f3ef49a7ac70ccfe7edb3a313e068a10f8a9f9b6fded0931e03447c0a228664789756d746bdc28f8b45b5c3413c59be8b272f548ca880a4ad71ce190b9174792e711c4cf2e3c815c88eaca47bf817b15888be1e8d5b316e3b0ee2e093891d6ed59cddeebb6168bb734acfe11dfbc9de48a4ed8a6910615d2728a21f94216def0a8f0ac1ec038a57648622ddff7402d3e3a1782b7f4f4157435dbb2bf2ef68626e481e92fe24f18467e51c04ba2c7e6af8df30a830381b17b5a3ff0bc888bb922cb9fbdae08d6487543853c8fae47e6138e7caf82273fd46847a9fec604281bc01ca03116765c4578d90c012f4dddd5af66afdc8c740c7f4542cb409ab7775441f430cf5c608cbd49560d4ac662fe9914ed3d48ea55bd6e2c6f228cce0501381b6cd043d7eae3ba6b96b506156d05d7169a6bba19cad4d831b4870cda2449e542e2c6579540e093c38d33fa663b9c908582b195e7469c77cb862c5cdfb97daec300423c60b9354bbac9c46642e45ddf602be0388865b9b405dd48231cec0bbadcb504b74c5ac9858b6c95a7da1381f22a8a33aa2f3ade7fa5a60730f4ecc6d16d1a3ec617e92e26eed743edabc4fc2cc0552ec40c3baa5d837bf6177135ba61068039f08d562700f5104a5ea112803fb0d7826ec2e262ac1508601e08f34b297239237450852c4264637bf5e8cbceab33d48595012a931718e7949cfbdc36af7d5f1c8603fa066803031db6b40384e1ad8bb104813d702f84256f7ebc3dc9384e9db54282636d55f8a5c764b941cb76036d7aca28ab0b260a66c0a5cacb709ca79b428d37d311e587ed4dcac7fd76d41fc86a7da10fe1bf86c12afe5e518b9ff29f8c44caad8e5c59264879a82d54ad02071245;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha0ce22f70327544ccdb595afa1c26de1308c615cb48e46d47a7d43bf18f568b18c8dc5f3ea91abc18760e5fb09467d100d4240cf6388db3030c7c769a44936c884557aa95245d2c84d92310d055fb455a907fb5dc23ec2634e3f033ba5f52a7e31694828607219ad07f94eaf0240d16d4e32c6ee4592a37127f429c2b9ba1755f32d3581f6479b3174f5ea009fea24d0e363b8a17aa831a8836138f6d221306fb06057a2b48fd0b98af220b8d3a6f629e7aa3be9a5af7a68cc5ffcf0cfcd043a1fe39cb78cd382d017c13ed1213571863bb8746ba036689ecbfe4967adb2074a70e3dea5284dc43d05d1e4352cd012bece4f9b0163094038f6c931853d2bff60d45233245c5b3550d9988016a30fdd80a774ce0223672c21819dfc58708013f5c32025883453b3d3a4fa68c8195c98c7baf50f19fe21882e05ae57c416df5c829d1aaea86445fc8373673521af081ef5b1ac992ee83f1ff6e3582d21c1799f8f8e86253b559bf17eacd0761c2305ce6a8840c1f0992d00b364cd8e253b2a99ccebe0f8061bad1cbd42e2139ad963beb530ce2b671d8b9e8bf1ab83331b6423cd34ee08b9845db0974ea276b672fba5ea9ea37247425e70c5da6d7247ba83feea6ccc06c7d33201bbe8e1e98aaa3b13eadce1f3b88da9193fbd7ab5a6ff268619ee4e122f05187e03097edc7c8a66197ec3a23e626521f150668ed1a6de555f327ebe2494d54fc6ce85dce36ddbc34d8d383bbfb2dc67dbc3ccbfc72310273e7335600230a5b24636d3b9ba303aac3cb6eb101058bb1f09ba23151db32ad83a1efeffe6ef7f797d83453683c52c89933b2159a251af208ff58733f24855ab5b4998b7cf7ee620f8da674f3b700673070cce0b3ffe2f5c0a58fae42853a66e86f2ac75c66e9b67414a1bdbc14e01495faf5ccde92e28d45367e43ecaaee3132b9883d0df3d73b805c3a8959a87600cfbe79f54ea209e76127808059753ebf7265aff46245b5340da1a9d46274de3be687783cf1d294e73afff95;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h7ed982064877ab681996b098e315b5505a42e1fe855b53f00b31aaa51eb308fad7198a65d355bf7799282ea00ba0ce67b0da4f570998cae9cd8960267e723ead138d5fe2bd9831871aab6ac9f25f0dcdd082ca641e06f8ea73cb0770456f00bb04f8c17a1bdb49e863a867ab9e63477d7a85bbc98b77eaeb7d0fd47d3da6affab7d33e0d674d3b70378d0edbb281aaed3a5be7e86316533baa4491fd102dc2a32c620a7e61d52f7435741201f283ebe696cc6b9bc0e233d427d0adeb860c7a762d3eeb9a30b551a68156a63711083788ced210802a219960e1b94fb789cdb50e0bc394db5b9fc331852efb57fe0beb86c46b8b166d80b00b39e3c1f32453e4b00f78617da08967c3843b7aeb91efef3663d61eb42ddd74fe397b87a320d3a0c532605b9afe0d1f590177ba4a9310a22fe08adc7aa848e8e38b7dbcfd76ba07a246bdbae77ef595a2649fc883cb00df9c581821ec59d45cbc245189432f13be1d18c9c460b0f9b33dd9870a7397f8a20a098ea1e53deac273569f754010672da7fa9f5a3bea494c9e3d3c2ec8ea279ea192708cdfc7377494315d163843d5da5a59c585163a9eea085ec1c9544b0c4d4883c99203296b30a6e96e9f5cf04b2bfd16340ef5fa4e8cd4b1fbfc376dbdf0a983289fe1dbddb0e07b11d93854c9e0a58784be9b77110069961b41e54b2432f827690233ed5a686fb6056a90d47843b0fcf95ece2afca4ced6e30b607f8e17d192f1b58b86bff4398df6a831d048f5c3ca2e26faa9ce11fd93ca14754403df07768883a7e855af6df238fa585543ac726b78770fba01600898d529359b0ca7d5db7e46bec2f6653a655ec741e579081befcb960532ecffa1f11180ce3f633a5752c5e6e43df5702f428e6e8a7c9e77f711e4f0a9cc1ed27686c051e884d5596a2758d6971ae21084b976abbd667dbd61da5b31b5798709855b8cd8d9ff8ecbc4dd1c3f0e233f65ced0b5539928f40310c7e894a52964da538c783e84bbe6179e0cefd9047901af0438;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hb8e7240eb49c7b9caf800fea511601de20a6728c5ab3f049dc216bfc3eac023e6c17bda0636a6eb113449577dcf71ff29d8ce160eebc2169a602184c7d79795486817c0ab8f9b7547c1d8e8ce4814735cc3949bbfa173e8099fd2f1165683b239b1a44f8fb731505893e637658e1f1cbd5ea8f8f550060361052057af2619e510c1784ba461eacddcee38d540f32ba4517ff171eade8dec943267b5a4074ed9fe13fb1f93a36a355980a8d7c17feee7cf6127d48101fe1aa93cf268ec07035366469d7ea84327e41943a95a9945fd0812eb1b84b6d0bab1f0dd2fea2436e9f65565615fc2be9a7233df79616ad3c3ffe118f9e412ade47c4845f0a965b493c230b6d49dadfef199cbecbff7648c63120f1f3895bafe5cd964c11e3b2528b2c6a8e2dba9a11b5f8b92917464a95365f7874bdd70a83302916e25f4c8a0cd9d4830b734b0ded492f9a2ffe1e0044765c110e890e79196cd4a21a169bf0606965bcf5e97fb54a5155eea8df94f9016c4b2f803c6c7643f257054b3bfdca41fa437189ca22af47bdc13c5714b72d78b6775ced6ad7fab715b5686f6e69c1ecabf3dfb7ce3a26f79c4de2df5a59e7ea5f282087cfb15aed0e36fbc69ea95e305a7e7c28ec179b1d35f41cfc83027f5bcfe9f61b69842c33f6f3754a2915796332883b02da9c53c1bc66a01d9c90da22284e38854aaf19733117f7daf60012dcc566d7fb2efc32b1780f7c14404a7ad8518c4f9f935233ecf6adb7c1f93a3c7a2104932069efc7c989496a7bbdd470110c4517d95c7c3ae794ab1b807c43986d09f823af7d8a4af9a72d4720fe29d931b87a54e99b1aa5313d2d43d654d02f6c4d953daf082806f3255b260359cb11c7f86af50578207a21ec6936ed00bfdf1ea314f7cfd7fce85e491822a6da56696623a4577147aec3886cbdc846dba61a6557d3c64a6497b34f550c51627a468f53c89af7806d094e6e716ba97e26d335fc968973c8be1facee731f54f061bf7eb900363936d3f22516961e5a73;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h172977e93755fae1da7d9d25689f4ced9fb14b3e98e724681f4891764c2d92ffa5857198957d7bba041e41946983fa5936179372004aa562dc138decffa5ae2c7ea2782c68f2f79519af6a4ea032baee558264dabb401c37d84376dd034881eb7daf76c3ce7319d4defa2f06664e1b83e39adde4c4cb6f09d4157ddbcd019e0db9585ba6ae9c5c94947847142a6a8ced0a232a5479cfc179ad178c642a111d6819fda49eb2b59bfc6270a1f6f0b35230aad17bfc64b9808e10027dcd5a8193e3591e697d6beabb762c06f97357a1a9823de2482439d630d4eba4ca8eeddfb1c0efe292dfba76ba7be81278bbd43af543ea17da9cf8a4759d74a9c097726186946dd49b6999c8750ce9c2ed62beb983adc5ee9aed672252b2e832e751de51a9ffb013d33513d235e1a6439e1d1b212c0b9249ee74275997f63f3ffb2977ac1de439375a36ba3f91250578176804f2dfd26c93963a28fef24cb39e1c84c66ba48c5a671c58417d3e225419f538cc7538598676b227abb83df34797a4b01466e5efb688729942326ac0a14d055a90272b8faa6b786b45253b6a9474120a42870e01d50a98a68c2f8c242cd611dca1a0d4890828ce437289db7c8e304fee8922d57318e286d77eadb98a385b145c368758b416e5517b2f3b7b0c49e18cd725c97cd16e92fd93c07d4f0ad3401a4cdbf74bae4aa437ffa53f7c24f53a829edd4f7327f77d83ae9441dcbde871b9ecd6f4586abb609cc2558d70fef2bc234c06802ebba971d2ca90915e2bf1c2f65cabed3097d58d32e67c340542eee24a87f556120c0e92e5254c1b712cfaba71a53841dddb11df87d8b3195d9a02fe5e7cbeeb6212e41639cc63f3b81bf6a6af13e900f4dae6615c9288fd63463ff2b39ef30117d716a50c3a9dec443b5275ddb2779b52001cbec83c9130960c04a3fbbe1fd8c61527b50b821a0d533a326ee51741bc3ac663ddc17a14a1f93eeb84b2bab4ab6ab315cce1bb24813e32412feecdbffe02f8aa38bc73e95386bb97;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h2f29b441e0016bc5cefac32ff3676c3b37c60ccb7715e44b11730ddb6b79511bc3b6984f51f333ff15bffc49483976044e09c8eac37d15fd71d73566ee36818c6d74454d3c6a2b49fa288d512b55931152958f4e33b3d5e159d9c7676a8046fc039915cb34b32affcc5937869199972d002f0cb96eae8c75967d9720bdb17d943da20ed083d100c09bc63caba914bebd43c34f089d3a8ba6ad5919d532e0e5f1ebf08997ef13d8fc0feddc10c88b8e6f52b0bafb39cc14cd68629bba721adf01143ed955f5a95b3202231915e425ca8aebaf1eb9de3647fa95750711eefb2c9d9420dd0dfb01426a08fc88ab513967ec3ec5155a9b4e3c5c32f8b2e79954bb76d824f433dcd10b7c73f309b9f5392318a0f13bc064bdd84a29bc5971bf304d78fad7e1e3abcc7b3339e95bf1791e7b1a510a9cdebb30e2522e143c17f93670b7aa32988ae12e4662754d576dc35e11fa69da778a5ad86e52c20dd587b52f72fd21ef25fcbab44df60ca6b963f77b11f6386381fa2b1d286fbfd76bc556b3b05679df4c9fc71689c03a7349bb6aed88a22ca57e3add6a0422cd5787458a5fc90000f307b3c996d62a6461d9855858fe5da308ffa92370c7f32c33c29a771fde04dab7209c605e6fb0447efde7da74688999ff22e741821eb8d8ce5c55feb404d306e89085b4cbca2de4d5c17116c8c10d8b8e140a67622615c18ab56fb28f2c7367ae5f4b7ff5ed7db03fa6cafcc5d1c0609b86bb30e2516e9d562019a143a8f72aa6eceaa612b1edf0273a78132be9a61f096695c42eb1aafc826a19e2a4e29ef5e3b0006d71de82ef86af350352342857c3fe886a5dbdd085c7976ed2ff460736b3495c4f92a54a6bc1db241d663ac348a7784280478e2eb37d3b8f832def071e86c4d5ca8555a61fa9df3a107a7e7a2b1daddd8b84db1aadf3fd1033b40b56d0e0a8b2b177ffa2f603680564daed53666339aac675efbc57ce7134d4a63248a2cd3a4b542904f7506ae189c92e6ebe02f744b81cb5853414;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h395ea05334bee9f080016d90f233f06fcaaf55d05bd6f3a5e8a9aaf2fc931b929473255c80d94781311ecc624d57d4048966ee5c6b6cfb32bb2d499d8736c637a820c9826e393255d4d366a84cb5111030e79c2556cf9d27371f5e8a17d028b950ce89060829859e0dd457f78c326798f3fad26debec298a923b6e63a3579f8c9166106aa69b614597a507c7c365e6ac7a9108817c2bca3cf540e335bf0cffc96359204c14e230471e6eee283e5d056a6ab7d67d305a541cf63631277cd26562587d44dd432f637889a785663796445a0886d6d5e5fe2ea8b9f2be9990bf9ab6f244f65c45cb0f2dcbc7f1594d32ef18e2f6e650f29e066275dcd6f86fc426de83e3000440f41e9c3a5de873ec80b8f74f43bf2a7e6d4028e31e071340e669a3d3b2a22f347e84388366eb39aa3cef6b0ca2f556e0b1f7dd17408f01e5bce73b7fc2d8e7bfb6cff1bf7f6f93a8156ebfeb4d760cc4ba1c218f8541f7c810e0565e5904d6a99c0ec3393d5e8324b2fd162930bd12fdcef29b4ba8b30531682ab0f32aa7fc17d409d5fc8aa58d338a281bd7303ff95fc6ce47b894c03c90f6e499e90e5d805b9dd291a4a61290297474960c07032b1f45a499b145e8b8d90bf1d0d211be8e4de438ea92b191337cec3690f88138f82fa17e73e8b129a146a24cf369358431bbcc812910f79c6a5225b40f6ac7bb605727a829ef1e844b92f6f97a460e1ed343745e866f547d64e0ef31bf765876174bca8963f940ce83b24f2ceea51b66cf79ae613de8e9fc212bf5e5824c276cb3a17c34a6fec1004edfa95217ac5615ec33c1953fc82411c7c1339a6433af01a82e385faaf1a0dec2f4cb98a86c7c879c90285c017ade3e79ee9ff1a5f2b91e86a45b9806c7c447e800859ca0242598b7396102518c7074369cb4c0a31690c73e9770e1515611d6717794f40cf077c89192664b7c0fa85646481390b60e4b0761379ac39650ba1baf66f3ddeabff3cee51e0e2dd2315ad226ae0ab802173587872cabccb5e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h914a66389d018542927ece1e85d09b1dd3e4662e6ef1a71cc6e2f4203b911a374544d3e1c047708a9c1c9745f77deb6658997af94c68b7c36fd5e58ca0232342ac18c5f0eb4777d3e2100cc95794e4721172eb4516bf428aa26df8a4c47988619798bafdcfc57dccc83b41e3d4e09caf00045cea221d72966015d4b4c983176c85b3bef9cb5f0e453c6a9bdc9e90f07e6479e2a8a47a784990b2f1a444d8bebcaae33878eab232ef5e4377981ae9986ef9bc1d74e00aecabca930334844d07932096034b87f9753ab40b770a13600f8c30153923fc1e7b81ed6edc4710e81cad22982b7178318af95e40d69355fe50a2255210a637e1fc61d30d329d594bfc921979554e9a8f037a53621fc68c4671f711d0cb6e4a0fe0f249eb6a008792ac6fb969dd2fe4d05c0833ed31f6ab06e2e0f30e8477b50eba60ef6d19c91469e428f8129e4583ac7e333f3b34b9c7da2a2163acd9c56c5c78f62e527ddb0bb6892dc79385c6f6a4eec678e3f20065269b55f4f14c50a8ee15e3529610902ded0a4e9094fb71562bbc6da1e8d4391d73d1fc9af96f48633c11cc036147517840eec1046bd002f32ff385d19dd9241f93966eabe5570d2278f285bff09ef18f2f2048683e39264810d94c91d16274575c9699693095fc324825ce69a082b0db43ba04d09f2ea98142e6b75ad5bf748b70c82ffcb83a5ceff52594b4eca2f03b0f3ad66945646fcd364e920121281086f95ab9ba3c1a5c51160fceb81c6c3cb6cf5404b02defc906c25217272d43c26a0460887cdd6ca8c2177a295613c362473ed43a50fcb4e75d377929a85c2427ec49ba964407ec40ff04ce67d410b84b2a652b7cc2d88043072d73d5575f02939a397eb54a105013282a363c9c79b9c8b6f3cdf6758ee1deb548d90f67f8aa9066392f286f86b7a6dafa336b87e25f3bb5ffbb2bd9245de94ff31389911f8d7329d44de59599e84d7fda025167c650cb1f0bf03d0bf7c0f13cc864d1cafb0690189980ef28eecdfa52e53c6825;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hd643aaaec67ba3bbfa6e10ccb29f6acb0548cd3244ba6b9306fe12d219b6c2f3336d413c41711c4d0c33505a17d2db390e27296defe71e3e4dca3dc206b60b89f84753d16ab8afc0873ebf6aafeb63797de3b06f8b1658253ea37a74240ca132c7052e6a81859764fef5c5730aa27a86b750b3e2c63476dd46c1678d92467cd919b43a163ae36c0b6bcde910d38abba3fd7453e9099283995d2e6115cf5c34ae8df154e15e75175b3848e487098ce5e2650a706415497e011b5bb27894f5a8dba059ef0dec7d00da1199037df1a4a9c9b4e63059a52f1525d9e7537efe9a9b9b9f0334cfd854c93cd4545c640daae266ee2a129db10b8b6c86b9c1d32cf4d26008e63a5e47d5f67461c37dfd04e5ece6955ebbd24335365399f040224d7d821a386394594b9c08934b26557f1b325ab93e97e0ff6982bb6db62cb051e02a41b76ad7e99276fc95e3179d901fcba27a4fe0b360b5a09756378fef6390d0d7801f7c5025aa49808bf5b06c6f17f4f9ef48d9ff793a44e671bdbbea1acfb76f3e6a9de7514a0959e72905d9f774aee166f086927fa31650ee4598eddc4e007f578ea8b6bc766e57dcb2b83d36295c2498bd13d27a4aac740fb2c601bb1a35ae4fd80d0369dbed764162334d93c4190afa7db5218cbf3d5ac4c9a53e53330e5385e0ec16a9309ddd95f6c33d9b009fb4629ddf2c9e46a310bd7801adebb718d9fc594da789b44f57dd86a6677c526ebc6530fe6050d43664889dfbda828cd82698ec13ee8075a5ecea850163100a873586a1b73b45abc283fec164a702f3c66b53eeb6a1fa05d3c42bec3cb9914ad6346a91f28ef64b740e71926fc833a8d6c42aeb6f71c776c3f5a51fba96d17ffa63a490c868a12b67fa7479da585ed87726757e5c9e700f2cc40281a24fe48db76f8304e501268604fa032663d4c6f7dcdd8a7cd7616bfe61df50ef5487c7a65e2f5e592da2e3dce1742c5c3c679d474e3162f5dbddb51935e799ccf08ca1df09e248bf5651e5763a24d91d19;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h3dbfba1f58778a8d4316de0dc0787463ff53acbfc35a8728b9935c11907002e5c68518830d44119f6c921c2168d38d501067199bbe1abb6a47e52c0dad4152f5c36815f69942f54f7f9f69e1b5fcd3c401e7f8fb04a4c739b8912d16fef1df40ffb43f515c81c38788db1b8fad73e8da9f01eed5e199373d07b9b264705e7c1d6b55ae98b980bce08b874a6c78db13f24513fcffc580b56509fd58381d7650115cc9c7abcdf9383452a2efc27017eac4613e9eda4f1a6b72927308f5bcccc9d5bdeca7513a0c4cb41d32840ca71d37a6f65ab7fbc6772daa008779dad6ff605590db60a3c7255df9efef0cfc7a1fb914fbe1612168d128a7b05d40057318ecf7ed174ca57f7c2e4ecea07fd87e4bac2aab01f2a0ae4c40f158d1f85b3c033b83171fb03a1e4914cad98dc6a32ac057526ee569accb28850d17b45f765a55c6f84cb8e716e17053c95e486ce88cd920085c188f3432b22e6407942e3d23917581b7a8dcfbe680c89ae8020c9d18743e819d20ea5f47336c5b01ce88fe006b44c717249c1e9b64cb9ccd919c5648ce8e74adb49af81b4087804a0d0a529d9af184bc0bc3428ee0665d34d4e23e7602513b12b54469fd1f3b1f381eb29bfc598fdf3b2b52a16a9464ff23c1268e01e96967cc52acdcc47b1d0179524f3318b61f01c3e97b241ffb497ceefa83ad0fb75f186c7e3d01dc394def8074a82e64b5f176d2b92b0fa163bde11ea1224fbf52ca104cd3d6ec7f2cceb790f0fc3fb8479a68d2798c6294473860632b6109eae5b796e4dba7f08c7c554a45011d41bbf99170aedb852ae9e10a6562506950f789b1223885c1778c3603ed44da090866c1234097bee6c16df00a1f4fe800ba5658b99fcab97751385418e130491f2d53ea1644ddf139f3d50d8712f1c93832b69cec171ca397290a7d20b57de46226bd63ae6e26c831ebcaab1342f614f8f6b7c438452b4e89a4c0aaf38775cdf7a7fd5628096da8e815509a43794b89558703c7f1cc3119200bd32d233e04;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'he7e72ea6411f3294e74bf02ad13139a665a8097f3733335182ef4df4ab37a6f2076503cc22a0323c02c753652a0a7d17ec31f84b8b6c30bdab88a6002c1b89364a40733f7c137c3d0e9a3c53f75de1a6d734f7f33f9f1793f730a4bf1fef18f0692a075f095de085cb039232c29bd9106913845efcb5bf8d942bd5871fb06a74e661221eb96c92dd33219296bd6eac4c911f126580b9792a99781ecd0e252f55bed06b58c4566d6c7a68e404c70fcc85372f2b00f881bf3e0e214ddc6e5a831598405afaa978c34f540e2ab5cbac7cf54b602f13fb7f1021aa7f683a3c8ab2b4f0bfd6f2887df35de5d241e0ae5966c089c24df8337d2d36063c83fd3a722fa234e9cdcc0dfcb5d5bc9fb2e907d6c9259ea2bd72a953b6acfb2820d379ec4bb8825a21ad78549b61c67d014ec3ac7faaa55f672113536c2eb7d2212465bb11f104af52a24c5153d07d38a953640d642158175a5e57748ed5844c30f4e9494411067907170260ade7a5ff5b101da321c5a7be92bfd12e8c4fd70ebe2bde0ff76ba017841fbb44ba3bbdf23ecffdabedcc3d8d29179e9d71b62a4d6999ed43243665deed4901b6f834f285f577de0b1ca7e808bd6e759ffc7bdc748048ac38b3606a287b2f75c35a38d939a7f90691aad0eeebba593e515f6a88fe0cd5c2a2194e82a8ffb7c132941becd22fe1eeb04bab570c06a8a1fcaf5690753ecb5b0d2b809d19d164438f1b216b910da777d7810700d010abcb1766ee33147c8c2ab332a020c0407333c640ab94824133afe13bd821b7c045a8597bb12c6bc2b06cffb71ffada4afe202af58d567a548c7983659cadd186289793c090ea8d6f52ba3b6bd9c29173627f0ba0b877d6ead9fc3c851ae7d64834f06f9a1598451f973b854a3dea4ed08f9d74d492ceb6cc87ebbef8f416d83dfe8efedf2e48841c316e18925221edc0e84c21b31218fb3bfc4e48b03ebef71fe12a83b2ac5203e3381e6a3045c2d8d1b61d4cc3e75f0e61827a604ef95264227640bab95036;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'hc0126a736764d502831cb360bd659209403c14764b23ad9c9bc45c6a7947a31015d4dc7d7fd17f6a0d21017483e823369b50aeda3eb2d991c5a00b36921d9602b6ba8902bf6595ac95504b0d771de97289ba55c9c5c1f3c34f631182b2b3ccfccd3aa2ae4c9d0bcbc80cc152516f8457283a05d7259cafee65b43ea23b2d11d12a3a6ee1bf108d23aade28d2496d741881322117ef602d22c642c99523de7e6a00969a488a40ba4ba78f6d51615690252301a587c5be7dbc623b83efb01a71cee918f89b60d1e6fc719aa6098fd14c12acbeaeb17490aaa67ead4e5a6da88c171312dbfee966880a21c75f754b84359cf19d693e7a4511c90bd286219b3cf749bfc27e37e3e9f743b1b4d3906b3edca2c065c9638a171d928e9b551c7505339af5dee9d046aea448d465fa8e7283f0661a3af46cb1367e6561b5779b4831912330fdc44c02203e484f9b4283b98d380ed1ee719cc83e371d76e00a60b90631837a4ff686e9e02150277cadcedf84db9f2668f5b99a1d58240bba613a4e4e69777bf178b5fd0d6b3629990f9b7e2f1fa86165b1a32a75095565e99c3d9ad2f47a1415853f1da356a6023f0e2db6c46bf012a560268821a3acc8998286eb4f4df3d811a0fb6e827ee05b44c88d1d4ead8b05ce57be95180fa5d6a44342e13ed31db7929e9beb03b2e25e0f0f3cbe06dbf9f623d5c574e0421c7f0991443336c2043e4a54f333fd5132f91be0dfbdae8fec05d96a89bf020209d21d06f15503a3098e48867a3ff6aaea072a054e9013ff6e32c0ac4e3359f11c380ef9358ee5d1f75dde2a88c40fc5fd9400ed1447e4f79f3a29b7fd4e7eb83fc74871d2287355be85ec8e6cc0c3f6d54521b35789b11fff5190d63a2a76a1f919d93148ad6cf4e4bc6948327dae1d16c4a0ce68b98589c96ea24a9f059b5f3bbe9173c69f061e740662e981c22c63466a5f35af051fda20d6d7a1fe94262dee043d0221d888858015e63ae420be33986cbca0c7b05fc51c0e6a7cf6d2544a6995;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h6b0c2105ded53ea151944f1569f42426163fe3b114ffc47d0adb395770ee7da1c2a33e23cd4152f10cfd73dc3f34d481ef5edd8f59e30a749291395a984ad6ce6245ce6f59cf13fd089c20e39aa2604d9c3aa06b66074756c88ddd9734a75fc89960b903f07ac5af4a4905576521f8de2321c761d5fca1e0c36a4ca1f90b2357ece2b866b68de4878d872cc6da3695cbcab5cfbe41fc62cd4be8081136cec5411cc2d3b09859702da55a40858bf1dc09d69adf5fb4f83b6d2ab7a47fa51566fb747873bc3b65f43c8bc198b2a70a4c7bc6375fb995276567b4396b7295e319c4df90c6de742d9e7a1d86b3ac1efb26099eaae50b226d4aca0213d27a36b80f80e03f0c4727248ad95df15edb6e5de297735f3156f68dcdda7fecf4ac275792b23a54375c7f87c5c0626dc03712c00557b63e5d1c1ba2eaaa50c9c173dcbf1e0a29cd2ba4d6cf1d744b8bc74b9a08e388d3a7d366604a647211b5ffbec907fd6bbf4768af6cc28a57fec18a9dcaf749f5057fdde7f8310102d065243ea1a9aacc9266582a737d74e92d96d9cbe7338349cc2490c905d62b92dcfe3f7fcff7fadf82e19e500a65c9eb287dad656726e21f9885dfbc6a6abda709a66eb7f61db703996af86c83bca22e1390d3b34c3ae06b7376c78034e0571ee6c52ef614f6915c497d1ca0ee567e8c5957d5e40f26ed7cafbce211245cea26ac4b4f6d993bf7f726f37498eb11b1d2c7923d4ac62b89d8c713f253c3af1b7c5157e78dec536340362f0efadd2f01fb64dbe7b41afb1730921ac3cd26bc8018ea0d519f248bedbac74784089d8537e4d24d958b617229315e96aa0739cc2a3642026032299825fa24e795ee897c619ceb54efec7b68bf1e5b53c585d5ce2896327987d9009ad8247efdc67344891212c89093c45c2dcf6d982f91af5cf0bec81b3a8f026ce92df07105cecd069e5eaabece4d669566b0e91043da700a83400eed8d50e96f9073697bdf576f6cffa046536de02455134eaa2873ff03a8f5046f05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'ha3d036e18b3d144142573fdad07e8f9075b451fc6589fcdcca99db792635b795139f1e4a9bcfed77e31f7dd595006ef817f45db337cf0a7d7cd7270216ed08b1326a99789ac4007591aa23fa1b2f999d1fde72d41b6466b3394f4fe5a2c12e2d46c2d54a68167753ea7228116ae3418002ae4c41bc57de3a9c077dde946a3aed3de8c451d867e597d48cc0eb05147c335292b76110d4354a0a61a4ce7e7762eeffe7c461c8c2521e0c6d60d7063e0e54d6b6edeb639754e9fc9de9c0cbec3ba213c176b7ce41dea4d009b3687dd4c5670cdcce6166829a829e7969b048471dc002fc2b1eb3d11938e2164a8d65675c0079ff5fc8bfa8f0e09bbdb2aaa8debfe513143d3e0f169a0439614155f2b05787433100c93378a85eaf3a8b992f31ed3ec2e36e5349420caec8045e605e32777ae50ad073297f0ede4e4a85bd32b4a865f9ae6bb33638b21d68f6101011622f2c58c29776578f1e53c9899e9617c7b11e70e51903c718c92a5f59fe093959a45772d059a5c6b4b59ed572c52a6f3fa03e640fcd434e0d1c592336cfe1da1caf4f133b720d38a410a80651d093efefbacabc8faaa3adc1c594856959567efd4f48d1e4910bfcfe7e0f9b3e65c3cb4c5ae0ea258d995599e63baf617d090613ad721467ba8865e86e3eb3f6f2666d44aa0c29f6f1cec44c46a56fa80a51fdaa9e4bd574e987664f0d2da4b1040af6cb99e2e103cd537f43c14c2c474d4eb154035d95385be6798affe73f6da7f281392e7040b790d1de8c05f497029fb563e7c170c13e8131ed93de04286b4c6850aafc08680893c6801bf7d104e72573775f3408b2a9785e66aa783f1429c9576bb6c77d412ffe06db39f0efc4c02ff37cdc82a8afed4cc4533eafe4714d5aaac91aabe1184722f93fd5e3fd33078727444874b5dc3cc5a276a0d64c9c31b1803e25509889c0d571816f92507d9f81831ef99b88dc93e649d9efc5113c750fe041e21c8fd9693ca63436635ad62801aa72776097aa8839e8661c17abfe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5832'h69f3d28164bc2abc0c57cef3a02dcd137ffc9d2e29af60807d3eff51b4237283abfe1c4221ae0730550279f8cd48c4e5a1a7ab56283bb46d90537205dc151cec13b629892c6dcabb41d2f0e4b25c3e6f92c01a7be630b2df37f371fcef0c057742adfb4f9177ed2b1c9c4290208c5ed89091029162f0208b9b26c26c37cc20363a81d6500ce3e7f651c094b1c2bc1598307239768ec44ac158b04af52b574910785d054b47846fc55c1bdc9add472a0ef1b922feed8f5388299ab6dff65c973de70e1669067f871a1e30873a5cc58b21c8f19f66867e071826543068849e4e3bda438a9036d514824aa774adc3550f48561fc1ea800bf282ee5779181e9b87463376db2edd4f218ef440c88d09eef48c27dcc67621b155ddad2cfd8d79e2e620e29fd4f2a5e8edeb1260bc9cade17dc875f5f221a0a2c23b02bcc1db08fadacf2a0a8d7ae339a5bd3a97bbeeb0c8bcd8c8ec9030d760ccde158b5608e5bb4ec1e92578f354d7fde575a7f2f14ea74b7a5f0139ae9648666507613981216bb6fee089c95fb9086e917f0354bf560cb82942d756c54e7fab230d84f93f3ffaf9991061b8c884b866f69dc67c3ed4118cc3c37a22a63b5f42d9f1c6d87f3216c1c4a0e13f20cb016c88d16d8745d7edae8883cdae7e39efb45cb0a5c528e58625e536bca690e1cff307f438460833f4ec6216abaad72906d5362e29d017f007c68a4fd0dd164d9725739910e19f2156bb59516f3470971f32171fce7fecb0147e892a2b0c2230155f64429406d9002c9c5c86f359613536315797df7528e080492d40f301ca790222c1bc3e2143cbaab76fd1eed00a8f3fb966a75a3612398a59d65b828763708a40e3455dc85cda09985dd1cc9362806372a4c0d70759d91afec0719ed397fb6c6f73584ec4ee7d859809e2d627693ec65e34f429573975146ebb4066179a2f6d5fda14d1a08427310dac0e880ada6ad4f33b45a3e80ab4061d272468d7cb2be5bde7807a414fb58f00d0bbadb9853eedb79a08;
        #1
        $finish();
    end
endmodule
