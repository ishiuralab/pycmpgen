module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21);
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    compressor_CLA54_16 compressor_CLA54_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21));
    initial begin
        src0 <= 54'h0;
        src1 <= 54'h0;
        src2 <= 54'h0;
        src3 <= 54'h0;
        src4 <= 54'h0;
        src5 <= 54'h0;
        src6 <= 54'h0;
        src7 <= 54'h0;
        src8 <= 54'h0;
        src9 <= 54'h0;
        src10 <= 54'h0;
        src11 <= 54'h0;
        src12 <= 54'h0;
        src13 <= 54'h0;
        src14 <= 54'h0;
        src15 <= 54'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA54_16(
    input [53:0]src0,
    input [53:0]src1,
    input [53:0]src2,
    input [53:0]src3,
    input [53:0]src4,
    input [53:0]src5,
    input [53:0]src6,
    input [53:0]src7,
    input [53:0]src8,
    input [53:0]src9,
    input [53:0]src10,
    input [53:0]src11,
    input [53:0]src12,
    input [53:0]src13,
    input [53:0]src14,
    input [53:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [0:0] comp_out20;
    wire [1:0] comp_out21;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out21[1], 1'h0, comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      input wire [53:0] src12,
      input wire [53:0] src13,
      input wire [53:0] src14,
      input wire [53:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [0:0] dst20,
      output wire [1:0] dst21);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [53:0] stage0_12;
   wire [53:0] stage0_13;
   wire [53:0] stage0_14;
   wire [53:0] stage0_15;
   wire [13:0] stage1_0;
   wire [16:0] stage1_1;
   wire [22:0] stage1_2;
   wire [17:0] stage1_3;
   wire [34:0] stage1_4;
   wire [24:0] stage1_5;
   wire [18:0] stage1_6;
   wire [18:0] stage1_7;
   wire [25:0] stage1_8;
   wire [26:0] stage1_9;
   wire [18:0] stage1_10;
   wire [17:0] stage1_11;
   wire [25:0] stage1_12;
   wire [25:0] stage1_13;
   wire [17:0] stage1_14;
   wire [23:0] stage1_15;
   wire [16:0] stage1_16;
   wire [7:0] stage1_17;
   wire [7:0] stage2_0;
   wire [2:0] stage2_1;
   wire [7:0] stage2_2;
   wire [8:0] stage2_3;
   wire [11:0] stage2_4;
   wire [9:0] stage2_5;
   wire [11:0] stage2_6;
   wire [10:0] stage2_7;
   wire [7:0] stage2_8;
   wire [11:0] stage2_9;
   wire [12:0] stage2_10;
   wire [6:0] stage2_11;
   wire [8:0] stage2_12;
   wire [10:0] stage2_13;
   wire [8:0] stage2_14;
   wire [7:0] stage2_15;
   wire [9:0] stage2_16;
   wire [6:0] stage2_17;
   wire [2:0] stage2_18;
   wire [2:0] stage2_19;
   wire [0:0] stage2_20;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [1:0] stage3_2;
   wire [5:0] stage3_3;
   wire [3:0] stage3_4;
   wire [5:0] stage3_5;
   wire [2:0] stage3_6;
   wire [5:0] stage3_7;
   wire [4:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [2:0] stage3_14;
   wire [3:0] stage3_15;
   wire [5:0] stage3_16;
   wire [3:0] stage3_17;
   wire [3:0] stage3_18;
   wire [0:0] stage3_19;
   wire [0:0] stage3_20;
   wire [0:0] stage3_21;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [0:0] stage4_20;
   wire [1:0] stage4_21;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;
   assign dst21 = stage4_21;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1406_5 gpc8 (
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3]},
      {stage0_4[0]},
      {stage1_5[0],stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8]}
   );
   gpc1406_5 gpc9 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7]},
      {stage0_4[1]},
      {stage1_5[1],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[2],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[3],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[4],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[5],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[6],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[7],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[8],stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16]}
   );
   gpc615_5 gpc17 (
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], 1'b0},
      {stage0_4[2]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[0],stage1_5[9],stage1_4[17],stage1_3[17]}
   );
   gpc606_5 gpc18 (
      {stage0_4[3], stage0_4[4], stage0_4[5], stage0_4[6], stage0_4[7], stage0_4[8]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[1],stage1_5[10],stage1_4[18]}
   );
   gpc606_5 gpc19 (
      {stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[2],stage1_5[11],stage1_4[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19], stage0_4[20]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[3],stage1_5[12],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[4],stage1_5[13],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[5],stage1_5[14],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[6],stage1_5[15],stage1_4[23]}
   );
   gpc615_5 gpc24 (
      {stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43]},
      {stage0_5[6]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[7],stage1_5[16],stage1_4[24]}
   );
   gpc606_5 gpc25 (
      {stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[7],stage1_7[8],stage1_6[8],stage1_5[17]}
   );
   gpc606_5 gpc26 (
      {stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[8],stage1_7[9],stage1_6[9],stage1_5[18]}
   );
   gpc606_5 gpc27 (
      {stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[9],stage1_7[10],stage1_6[10],stage1_5[19]}
   );
   gpc606_5 gpc28 (
      {stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[10],stage1_7[11],stage1_6[11],stage1_5[20]}
   );
   gpc606_5 gpc29 (
      {stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[11],stage1_7[12],stage1_6[12],stage1_5[21]}
   );
   gpc606_5 gpc30 (
      {stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[12],stage1_7[13],stage1_6[13],stage1_5[22]}
   );
   gpc606_5 gpc31 (
      {stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[13],stage1_7[14],stage1_6[14],stage1_5[23]}
   );
   gpc615_5 gpc32 (
      {stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_6[42]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[14],stage1_7[15],stage1_6[15],stage1_5[24]}
   );
   gpc615_5 gpc33 (
      {stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage0_7[48]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[8],stage1_8[15],stage1_7[16],stage1_6[16]}
   );
   gpc615_5 gpc34 (
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52]},
      {stage0_7[49]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[9],stage1_8[16],stage1_7[17],stage1_6[17]}
   );
   gpc615_5 gpc35 (
      {stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53], 1'b0},
      {stage0_8[12]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[2],stage1_9[10],stage1_8[17],stage1_7[18]}
   );
   gpc606_5 gpc36 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[1],stage1_10[3],stage1_9[11],stage1_8[18]}
   );
   gpc615_5 gpc37 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_9[6]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[2],stage1_10[4],stage1_9[12],stage1_8[19]}
   );
   gpc615_5 gpc38 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28]},
      {stage0_9[7]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[3],stage1_10[5],stage1_9[13],stage1_8[20]}
   );
   gpc615_5 gpc39 (
      {stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_9[8]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[4],stage1_10[6],stage1_9[14],stage1_8[21]}
   );
   gpc615_5 gpc40 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38]},
      {stage0_9[9]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[5],stage1_10[7],stage1_9[15],stage1_8[22]}
   );
   gpc615_5 gpc41 (
      {stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_9[10]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[6],stage1_10[8],stage1_9[16],stage1_8[23]}
   );
   gpc615_5 gpc42 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_9[11]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[7],stage1_10[9],stage1_9[17],stage1_8[24]}
   );
   gpc615_5 gpc43 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_9[12]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[8],stage1_10[10],stage1_9[18],stage1_8[25]}
   );
   gpc606_5 gpc44 (
      {stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[8],stage1_11[9],stage1_10[11],stage1_9[19]}
   );
   gpc606_5 gpc45 (
      {stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[9],stage1_11[10],stage1_10[12],stage1_9[20]}
   );
   gpc615_5 gpc46 (
      {stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_10[48]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[10],stage1_11[11],stage1_10[13],stage1_9[21]}
   );
   gpc615_5 gpc47 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34]},
      {stage0_10[49]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[11],stage1_11[12],stage1_10[14],stage1_9[22]}
   );
   gpc615_5 gpc48 (
      {stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39]},
      {stage0_10[50]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[12],stage1_11[13],stage1_10[15],stage1_9[23]}
   );
   gpc615_5 gpc49 (
      {stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44]},
      {stage0_10[51]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[13],stage1_11[14],stage1_10[16],stage1_9[24]}
   );
   gpc615_5 gpc50 (
      {stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49]},
      {stage0_10[52]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[14],stage1_11[15],stage1_10[17],stage1_9[25]}
   );
   gpc615_5 gpc51 (
      {stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53], 1'b0},
      {stage0_10[53]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[15],stage1_11[16],stage1_10[18],stage1_9[26]}
   );
   gpc606_5 gpc52 (
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[0],stage1_13[8],stage1_12[16],stage1_11[17]}
   );
   gpc606_5 gpc53 (
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[1],stage1_13[9],stage1_12[17]}
   );
   gpc606_5 gpc54 (
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[2],stage1_13[10],stage1_12[18]}
   );
   gpc606_5 gpc55 (
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[3],stage1_13[11],stage1_12[19]}
   );
   gpc606_5 gpc56 (
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[4],stage1_13[12],stage1_12[20]}
   );
   gpc606_5 gpc57 (
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[5],stage1_14[5],stage1_13[13],stage1_12[21]}
   );
   gpc606_5 gpc58 (
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[6],stage1_14[6],stage1_13[14],stage1_12[22]}
   );
   gpc606_5 gpc59 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[7],stage1_14[7],stage1_13[15],stage1_12[23]}
   );
   gpc606_5 gpc60 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[8],stage1_14[8],stage1_13[16],stage1_12[24]}
   );
   gpc606_5 gpc61 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[9],stage1_14[9],stage1_13[17],stage1_12[25]}
   );
   gpc606_5 gpc62 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[9],stage1_15[10],stage1_14[10],stage1_13[18]}
   );
   gpc606_5 gpc63 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[10],stage1_15[11],stage1_14[11],stage1_13[19]}
   );
   gpc606_5 gpc64 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[11],stage1_15[12],stage1_14[12],stage1_13[20]}
   );
   gpc606_5 gpc65 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[12],stage1_15[13],stage1_14[13],stage1_13[21]}
   );
   gpc606_5 gpc66 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[13],stage1_15[14],stage1_14[14],stage1_13[22]}
   );
   gpc606_5 gpc67 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[14],stage1_15[15],stage1_14[15],stage1_13[23]}
   );
   gpc606_5 gpc68 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[15],stage1_15[16],stage1_14[16],stage1_13[24]}
   );
   gpc606_5 gpc69 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[16],stage1_15[17],stage1_14[17],stage1_13[25]}
   );
   gpc1_1 gpc70 (
      {stage0_0[48]},
      {stage1_0[8]}
   );
   gpc1_1 gpc71 (
      {stage0_0[49]},
      {stage1_0[9]}
   );
   gpc1_1 gpc72 (
      {stage0_0[50]},
      {stage1_0[10]}
   );
   gpc1_1 gpc73 (
      {stage0_0[51]},
      {stage1_0[11]}
   );
   gpc1_1 gpc74 (
      {stage0_0[52]},
      {stage1_0[12]}
   );
   gpc1_1 gpc75 (
      {stage0_0[53]},
      {stage1_0[13]}
   );
   gpc1_1 gpc76 (
      {stage0_2[48]},
      {stage1_2[17]}
   );
   gpc1_1 gpc77 (
      {stage0_2[49]},
      {stage1_2[18]}
   );
   gpc1_1 gpc78 (
      {stage0_2[50]},
      {stage1_2[19]}
   );
   gpc1_1 gpc79 (
      {stage0_2[51]},
      {stage1_2[20]}
   );
   gpc1_1 gpc80 (
      {stage0_2[52]},
      {stage1_2[21]}
   );
   gpc1_1 gpc81 (
      {stage0_2[53]},
      {stage1_2[22]}
   );
   gpc1_1 gpc82 (
      {stage0_4[44]},
      {stage1_4[25]}
   );
   gpc1_1 gpc83 (
      {stage0_4[45]},
      {stage1_4[26]}
   );
   gpc1_1 gpc84 (
      {stage0_4[46]},
      {stage1_4[27]}
   );
   gpc1_1 gpc85 (
      {stage0_4[47]},
      {stage1_4[28]}
   );
   gpc1_1 gpc86 (
      {stage0_4[48]},
      {stage1_4[29]}
   );
   gpc1_1 gpc87 (
      {stage0_4[49]},
      {stage1_4[30]}
   );
   gpc1_1 gpc88 (
      {stage0_4[50]},
      {stage1_4[31]}
   );
   gpc1_1 gpc89 (
      {stage0_4[51]},
      {stage1_4[32]}
   );
   gpc1_1 gpc90 (
      {stage0_4[52]},
      {stage1_4[33]}
   );
   gpc1_1 gpc91 (
      {stage0_4[53]},
      {stage1_4[34]}
   );
   gpc1_1 gpc92 (
      {stage0_6[53]},
      {stage1_6[18]}
   );
   gpc1_1 gpc93 (
      {stage0_15[48]},
      {stage1_15[18]}
   );
   gpc1_1 gpc94 (
      {stage0_15[49]},
      {stage1_15[19]}
   );
   gpc1_1 gpc95 (
      {stage0_15[50]},
      {stage1_15[20]}
   );
   gpc1_1 gpc96 (
      {stage0_15[51]},
      {stage1_15[21]}
   );
   gpc1_1 gpc97 (
      {stage0_15[52]},
      {stage1_15[22]}
   );
   gpc1_1 gpc98 (
      {stage0_15[53]},
      {stage1_15[23]}
   );
   gpc1163_5 gpc99 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc100 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc101 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], 1'b0},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc102 (
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[3],stage2_3[3],stage2_2[3]}
   );
   gpc606_5 gpc103 (
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc606_5 gpc104 (
      {stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc105 (
      {stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7]},
      {stage1_4[18]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[3],stage2_5[3],stage2_4[6],stage2_3[6]}
   );
   gpc615_5 gpc106 (
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage1_4[19]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[4],stage2_5[4],stage2_4[7],stage2_3[7]}
   );
   gpc615_5 gpc107 (
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage1_4[20]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[5],stage2_5[5],stage2_4[8],stage2_3[8]}
   );
   gpc207_4 gpc108 (
      {stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27]},
      {stage1_6[0], stage1_6[1]},
      {stage2_7[3],stage2_6[6],stage2_5[6],stage2_4[9]}
   );
   gpc606_5 gpc109 (
      {stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[0],stage2_7[4],stage2_6[7],stage2_5[7],stage2_4[10]}
   );
   gpc606_5 gpc110 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[5],stage2_6[8],stage2_5[8]}
   );
   gpc615_5 gpc111 (
      {stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage1_7[6]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[2],stage2_7[6],stage2_6[9]}
   );
   gpc615_5 gpc112 (
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage1_7[7]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[2],stage2_8[3],stage2_7[7],stage2_6[10]}
   );
   gpc615_5 gpc113 (
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_8[12]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[2],stage2_9[3],stage2_8[4],stage2_7[8]}
   );
   gpc615_5 gpc114 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage1_8[13]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[3],stage2_9[4],stage2_8[5],stage2_7[9]}
   );
   gpc606_5 gpc115 (
      {stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[2],stage2_10[4],stage2_9[5],stage2_8[6]}
   );
   gpc606_5 gpc116 (
      {stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[3],stage2_10[5],stage2_9[6],stage2_8[7]}
   );
   gpc606_5 gpc117 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[2],stage2_11[4],stage2_10[6],stage2_9[7]}
   );
   gpc606_5 gpc118 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[3],stage2_11[5],stage2_10[7],stage2_9[8]}
   );
   gpc1163_5 gpc119 (
      {stage1_10[12], stage1_10[13], stage1_10[14]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage1_12[0]},
      {stage1_13[0]},
      {stage2_14[0],stage2_13[2],stage2_12[4],stage2_11[6],stage2_10[8]}
   );
   gpc117_4 gpc120 (
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6], stage1_12[7]},
      {stage1_13[1]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[1],stage2_13[3],stage2_12[5]}
   );
   gpc606_5 gpc121 (
      {stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13]},
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage2_16[0],stage2_15[1],stage2_14[2],stage2_13[4],stage2_12[6]}
   );
   gpc606_5 gpc122 (
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19]},
      {stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12]},
      {stage2_16[1],stage2_15[2],stage2_14[3],stage2_13[5],stage2_12[7]}
   );
   gpc606_5 gpc123 (
      {stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25]},
      {stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], 1'b0},
      {stage2_16[2],stage2_15[3],stage2_14[4],stage2_13[6],stage2_12[8]}
   );
   gpc606_5 gpc124 (
      {stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[3],stage2_15[4],stage2_14[5],stage2_13[7]}
   );
   gpc606_5 gpc125 (
      {stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[4],stage2_15[5],stage2_14[6],stage2_13[8]}
   );
   gpc606_5 gpc126 (
      {stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17], stage1_13[18], stage1_13[19]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[5],stage2_15[6],stage2_14[7],stage2_13[9]}
   );
   gpc606_5 gpc127 (
      {stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[6],stage2_15[7],stage2_14[8],stage2_13[10]}
   );
   gpc117_4 gpc128 (
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage1_17[0]},
      {1'b0},
      {stage2_19[0],stage2_18[0],stage2_17[4],stage2_16[7]}
   );
   gpc117_4 gpc129 (
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12], stage1_16[13]},
      {stage1_17[1]},
      {1'b0},
      {stage2_19[1],stage2_18[1],stage2_17[5],stage2_16[8]}
   );
   gpc1163_5 gpc130 (
      {stage1_16[14], stage1_16[15], stage1_16[16]},
      {stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5], stage1_17[6], stage1_17[7]},
      {1'b0},
      {1'b0},
      {stage2_20[0],stage2_19[2],stage2_18[2],stage2_17[6],stage2_16[9]}
   );
   gpc1_1 gpc131 (
      {stage1_0[9]},
      {stage2_0[3]}
   );
   gpc1_1 gpc132 (
      {stage1_0[10]},
      {stage2_0[4]}
   );
   gpc1_1 gpc133 (
      {stage1_0[11]},
      {stage2_0[5]}
   );
   gpc1_1 gpc134 (
      {stage1_0[12]},
      {stage2_0[6]}
   );
   gpc1_1 gpc135 (
      {stage1_0[13]},
      {stage2_0[7]}
   );
   gpc1_1 gpc136 (
      {stage1_2[21]},
      {stage2_2[6]}
   );
   gpc1_1 gpc137 (
      {stage1_2[22]},
      {stage2_2[7]}
   );
   gpc1_1 gpc138 (
      {stage1_4[34]},
      {stage2_4[11]}
   );
   gpc1_1 gpc139 (
      {stage1_5[24]},
      {stage2_5[9]}
   );
   gpc1_1 gpc140 (
      {stage1_6[18]},
      {stage2_6[11]}
   );
   gpc1_1 gpc141 (
      {stage1_7[18]},
      {stage2_7[10]}
   );
   gpc1_1 gpc142 (
      {stage1_9[24]},
      {stage2_9[9]}
   );
   gpc1_1 gpc143 (
      {stage1_9[25]},
      {stage2_9[10]}
   );
   gpc1_1 gpc144 (
      {stage1_9[26]},
      {stage2_9[11]}
   );
   gpc1_1 gpc145 (
      {stage1_10[15]},
      {stage2_10[9]}
   );
   gpc1_1 gpc146 (
      {stage1_10[16]},
      {stage2_10[10]}
   );
   gpc1_1 gpc147 (
      {stage1_10[17]},
      {stage2_10[11]}
   );
   gpc1_1 gpc148 (
      {stage1_10[18]},
      {stage2_10[12]}
   );
   gpc207_4 gpc149 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6]},
      {stage2_2[0], stage2_2[1]},
      {stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc150 (
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7]},
      {stage2_3[0]},
      {stage2_4[0]},
      {stage3_5[0],stage3_4[0],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc615_5 gpc151 (
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage2_4[1]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[2]}
   );
   gpc615_5 gpc152 (
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage2_5[6]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[1],stage3_5[2],stage3_4[2]}
   );
   gpc615_5 gpc153 (
      {stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_5[7]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[2],stage3_6[2],stage3_5[3],stage3_4[3]}
   );
   gpc615_5 gpc154 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[3]}
   );
   gpc615_5 gpc155 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[4]}
   );
   gpc606_5 gpc156 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[2],stage3_9[2],stage3_8[4]}
   );
   gpc7_3 gpc157 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12]},
      {stage3_12[1],stage3_11[3],stage3_10[3]}
   );
   gpc606_5 gpc158 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[4]}
   );
   gpc1343_5 gpc159 (
      {stage2_12[0], stage2_12[1], stage2_12[2]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9]},
      {stage2_14[0], stage2_14[1], stage2_14[2]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[3]}
   );
   gpc615_5 gpc160 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7]},
      {stage2_13[10]},
      {stage2_14[3], stage2_14[4], stage2_14[5], stage2_14[6], stage2_14[7], stage2_14[8]},
      {stage3_16[1],stage3_15[2],stage3_14[2],stage3_13[2],stage3_12[4]}
   );
   gpc117_4 gpc161 (
      {stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6], stage2_15[7]},
      {stage2_16[0]},
      {stage2_17[0]},
      {stage3_18[0],stage3_17[0],stage3_16[2],stage3_15[3]}
   );
   gpc7_3 gpc162 (
      {stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6], stage2_16[7]},
      {stage3_18[1],stage3_17[1],stage3_16[3]}
   );
   gpc1325_5 gpc163 (
      {stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage2_18[0], stage2_18[1]},
      {stage2_19[0], stage2_19[1], stage2_19[2]},
      {stage2_20[0]},
      {stage3_21[0],stage3_20[0],stage3_19[0],stage3_18[2],stage3_17[2]}
   );
   gpc1_1 gpc164 (
      {stage2_0[7]},
      {stage3_0[1]}
   );
   gpc1_1 gpc165 (
      {stage2_3[6]},
      {stage3_3[3]}
   );
   gpc1_1 gpc166 (
      {stage2_3[7]},
      {stage3_3[4]}
   );
   gpc1_1 gpc167 (
      {stage2_3[8]},
      {stage3_3[5]}
   );
   gpc1_1 gpc168 (
      {stage2_5[8]},
      {stage3_5[4]}
   );
   gpc1_1 gpc169 (
      {stage2_5[9]},
      {stage3_5[5]}
   );
   gpc1_1 gpc170 (
      {stage2_7[10]},
      {stage3_7[5]}
   );
   gpc1_1 gpc171 (
      {stage2_11[6]},
      {stage3_11[5]}
   );
   gpc1_1 gpc172 (
      {stage2_12[8]},
      {stage3_12[5]}
   );
   gpc1_1 gpc173 (
      {stage2_16[8]},
      {stage3_16[4]}
   );
   gpc1_1 gpc174 (
      {stage2_16[9]},
      {stage3_16[5]}
   );
   gpc1_1 gpc175 (
      {stage2_17[6]},
      {stage3_17[3]}
   );
   gpc1_1 gpc176 (
      {stage2_18[2]},
      {stage3_18[3]}
   );
   gpc2135_5 gpc177 (
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4]},
      {stage3_4[0], stage3_4[1], stage3_4[2]},
      {stage3_5[0]},
      {stage3_6[0], stage3_6[1]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0]}
   );
   gpc615_5 gpc178 (
      {stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_6[2]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1]}
   );
   gpc135_4 gpc179 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1]}
   );
   gpc1163_5 gpc180 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc181 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], stage3_14[2]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc1163_5 gpc182 (
      {stage3_15[1], stage3_15[2], stage3_15[3]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage3_17[0]},
      {stage3_18[0]},
      {stage4_19[0],stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[1]}
   );
   gpc1163_5 gpc183 (
      {stage3_17[1], stage3_17[2], stage3_17[3]},
      {stage3_18[1], stage3_18[2], stage3_18[3], 1'b0, 1'b0, 1'b0},
      {stage3_19[0]},
      {stage3_20[0]},
      {stage4_21[0],stage4_20[0],stage4_19[1],stage4_18[1],stage4_17[1]}
   );
   gpc1_1 gpc184 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc185 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc186 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc187 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc188 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc189 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc190 (
      {stage3_3[5]},
      {stage4_3[1]}
   );
   gpc1_1 gpc191 (
      {stage3_4[3]},
      {stage4_4[1]}
   );
   gpc1_1 gpc192 (
      {stage3_21[0]},
      {stage4_21[1]}
   );
endmodule

module testbench();
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor_CLA54_16 compressor_CLA54_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hed2b37ad3e724c5ab9fb31a135c2ba3121ba5ce0fb53cf52f50eec4f6f80fc616e479c90bcd86c49949296f4ec6ef9183100069a916f981569e3e73b4860cdcfaaeb5d9f4998b18ad7f9b4a7bc8ff75ac0fd95ee10caa0f518d20c642553e012bb01a52b27db06ce0f7259ef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hcda0d53dfd686ef3da0a0d4e499f0a8d3ddd98c10a98ef963a7800a8a497b713d293765857d71f1593e7ea9673cd317147735fc757934f76c4fbd3712d1698a7a61e54bbf9528bebb58c0fedd33aaba65aa1d73502705909989bd911de41c27398212af2a8b5ab6f4a954d80;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h4c14d4df49ca24b387a0d0cc95091d4a09648ea08d7d6ab60d12af5443bd1b4086a4a14460ab3d0fb91574fef096f23e3cd1ece745e44fdd24ec68fb44760b4c59916c51efa386002cc7130ec717570c199ffca26664baa95b5cc014705853bb0d9150e35d765f7bed25d4c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'had087735dfc5bc4f2dca91cff6f037848b310e3630b253b3a2bbe329fd490df033585703a568cbce1de6440b1e1bda07e6c7b599fe78cebe0e6cf7409c841c97b7d6ebfb677e082c659f1bd228f98245932b98b8ee82615a2a7ed96b2c3de8a7c1bcfb666018536b2bcaa20f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hb11dd7e8e824ecb1366f591dd3bc2002871aa433fc0c9aef0dc73ff3d616859a75991127a39e994d48a430d534b30005b93eb255c3fe7bd730feb0d3a5a27a31410fe12a862748a96f1a3246c5258fec3fec5a707a15a24f18623d97fe97b513d5dc6997857a329b26cb6149;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h38d6f756e5bccb569f3ecf1c700c0b7c28566157db7e432ff39ce0ea31188eadc8ecc95a9dd4708d538e41a883dea5cfa6fcc49820e2f955080fcf58aad52507112e53699e12717516c385986a80b2e137854818d8504f141f9e9d97c050d39cc8eee1aec2efbe3fe2b300eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h2046313f9caa8b33556d4c9ae7d05fc56bd465218884bad92900d0d4641856dd6124c181c99d23ec6af37919ac0f55d1fadbc7d078141935788aae57a65fe621113a5f91a8527accd0b5e44c1b0208e331b966f693fee9a986469dba2ab2e4bbbac7d4ad68c6f416500ca0e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h4bc90ce54feccdc236355e4f5dec5aca1a434f578ac6b3e11fae43fdb05bc9b8fb335d616e44f283b120223f7db2450c7e16bd7a0d8c7af81550a337365c9fcddf6462876c70144c8eb4f99ec4b98729db68968297f882543ee8f8003eff94185f6f7a2200d26ad9dae61d4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hc77435fb05bd9cd59637f683a17b8f81a7e480b352b8d138de7d2af041742df136fddec190271d1287a52ff84940a1fc93909d1e4bdac9f9a34026fd84730a93dacc8198da78100c673ac87f546262308bd32d998bfce9a2abc339ec8e00aab711a60de8e27fe4e2a3ce6ba6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h11003fce4aea67787e4312f4f2039d44fc64299e6039509e05d29459c1d122ad1ca977c2f5e2412f9b94d09b6d7ad2212f3585cd2969629759a4632a1b444503bf6512d9dae2661a3a53be9ade7f7139ecd36635565d46d68d05194b45745437e9ccc470c7bac25c980baa05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h6ce9a8ff81b7a814fe35968da8e5fce1afcb8bd1e5159e691f8046cca129f1113709dc13216caf88832260869ef7f62bb25a31a3630bee0bc4fb572c9446b4ce6a2492f69dbb25f3688a6db4d24da599e0805d85e2f8deff480d4a294408921c760730716280b2cedabc79d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9aebd3124d743a40d768c191da233433b8158893b4a71343b86e5356f4119822c7f0ffa595e84e0c319e6ba5fa88e666ff127d74e23eb7e291a926a105268e9a473c065a912bd67749b3e1f80726b47b33f2c0e3df7980d8150bf10643b2c98c9b701a49bb7204ed62f0aa6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he23d52015736e14e80f3114292e1b93bcf183159531bc0bb0ed28c513edbee693b397e279b030f87864735daf281b5872e26e3fc99a8007727a716622a3c81dcb94643ae3a0752960a9249e4a490a302c34993fea20fc57b779093408a69ee83e3f16c37d6929b7f0384221d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf18c423d1a1d10c4309d4e175178ac4599ea11f5d2ef7aae2501c307e251cae58f3d7afcdae27e30e41de6178cc431e354488796fb3509feb3ebc0820e5028053dd976a7eed39d28327b6734499ee2f02be3cea577507b0cb2082920c2816054dac6f94b1065f25298cae8e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h24e74b6e7c8d8d2d8a7fef157725d30ca2c34f3b0f846ece2d93162fa1c8a129616d1081d5dc153896a49afa9af6fe5b279b70253581683730cf9c1952a67fac5422339cc4dc94cc36e64fa29b1f78ade1da968ac4fd63a8933eb079dcf983d08aeb967a51e1b80731377a8b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h87bd613dc30c55a183de569b270432443c59efd93e4d54b860bd70c40bb0c6d82872cedf6864964d52de1551554ee1b6dd14c2dab4c80b82ce55b8f8e6411d5b37c8a58726d0a1ba96f8aa0d2997d8f8043138e14baaa31b9fc961de56f1ad93af8474cdeddb14a376be5877;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h1a3e3aff12174ff49901a44f6e907198e599ad8f7f78aebe8e5270d09836c6c2c9b7e0ad18169ed21f75c9125345f19eb77256c8d25df313b48840660ef9d1208c85807fe655a73b4012b847f6a0ee52949156814023c9021de0265f04127a425796eb6e034d9a12f816a0c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h775bbf36f40ddb9f15291a24995f50494452e8182fcd8cabb7f6aacbf95621a10efde45266c17e58a6a4f05bc6bcf215912c4de5d5764ba24e1bd5ae69a82fc65fe251d8a67b0cf81e4a79a58e001cf0c5e6708037e2d66f958194b90af1cfcd471164d741c9b0e98c05fd0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hce7b57fa8b6cb2a66b71556be59944d4dfb9ab0898881d33d4ac20cb01675c72cb6743e1ceaa11c5300a562856b73d8c435cd6979f23e2520a71687e5582de839b674b23bfdb0311f4dfeee7061751f89df27cf85a47da10ac1bf7b2dc9bc3f5a9328f76dae9bda553a428b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h23833be80d382de5af742233e6be5d296544e2534bbc70a57a808be056b600c4f12e494b1484c8b0435e446e800baa42fa9663f02b6297f5ebfddf673c40719411231037849156f36451b49de2161f92cac06192e593f7567eeb4b0e6c85999568d0321ff49f400dc5375799;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd79d0adf33218d8bf98b1362b67537c5083a753326dfa0e77273d01006fa011fa4472347e9658b5b7ef3cb7de2ae313b67e61cf15a5f92c54ca2b79b66442b11b4eeccb7f0e7c6615122955af9a2839dd664b230e20f1d156e6c4bf42497e9555b6fd36d8f9b0cb97e451b14;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he513bf244a4ed4b0cebb733db7c4cc98d449cc0367877f028785a81926f9442e273bf53ee8322c141a5916f19acf72d5cb44915482879987a7eaa113eaf84c973fe24e8d2908620f89d8234b763402ee252ab2dfa5ddc17a6f7b05f977ed7a871b4043be8f299ba0b459bb76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha848e79a96b6f2d0d30af9c91316cbcbe92f68407a27edbec937e070101df01b1811acd68fd4fbe47070f92742a42d2a30088946b1456e7857f40d4105a63f3635f944a1be66508ce93a57c639bf82125769d18f64d00602708e4266c0736f07a3cb0d27ca282dcb391e638e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8df43d2c8e39362bc2462f8aaa252ab063cbc057933c5555fb32760b4167d55bf3253963b451c9c5d1b0d52a1f7b34bfb4bbce677edeb6140fbd78890155e27ee061fda4461d99d6268b335d59ad6a5bd9a77f910c94a274601b10dc9d3fc4dbc02104efd20bddcecdaf367;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h7c668ef6c13743bb4b88022579bd6644999acdefb7cef25a0bc256d9f24158f28f2cd844be22fbc8b95af834e21164ebc2a19f895e67ca4a357c4cd26eb76e78e1f279638ccdafcc0e653eb41d29fcbbff5d09fc652b9d8f7b92e50c7249a86738dde03942284fd4339cac22;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h51bab59092941ffeccf0807b4027fb8859a03ee85b1b0b84b8d5c1b4d81d88822805d1c9d34c812e17966e8630bde1ab175a06d94f77d0cce81d4abcf7b22f7d33e46bdda0fab5282fc90e2515ded66105821a7212a5b84554dc129c4c1465a7cc4b81ab7ce525cd3906a047;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h622196fb663747744d9a26af4713e14f2550f2bf25e4ca867c6a365abcd756ed1610060e7d0000f68d8ccfc2cfd8b006baaeb48c37465c5b7c5973e3b9b2500effa00015796c16113697270242178d07d2ff0cc806fed03a310e7caeb83beb6222f8d1bbc1932910cfa0edfc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h1ace88421e5e5933254e5e1dfd78a66941c131842e6d8aba1bb5e58b0e2bd0c6c928bd4cc0102972b2f82ef8118a818b5e44eacca9ff9caa27b6a8c490616ad200add8e03905875eb7c87511ea87e40488db3c4394cdd797ffa5f9500e705bdb0e4ac2075bcca03fe88ecdd4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h42db63d1c7ec725d54f1bd5e73cf5feb7452ca7702b86a0a568f6275404d5a2619c839086e1b672d1236c822c827f35a7927a51a6ce3183427ce668d0df54e66fbb00affe21304614dd5474a1c529dd3ec05ae31c337e6f371bc9dfc769ad689e143afcf00597e4c9a9ecd08;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hbfe26025b6cd003ad5a0de611262c5f68e9a77a9af3412ee0316e2f4024c7cc0dc083301d4c6367ea0858e63bd18dfdbc6d9841e5f8e62a39d75b8cc10f372c5f434bb780e23bbee2c81819bc443fbd45cab0c71a8880739e7e155215ed0e5f08dc0fa9dffd750cfc841fe46;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hae41d46fa72dbe7405b2eaef7b9e407f644d664fae93126af34ae628e72af9ac4ba2fef0da898c60c4777817419ab2814d9e4297681e3950c983613b92179a0bce25559b2dee74bea31ab4567ec518ad0b60e16ec994e5163fd3af4799e8e9281d531eb23b24b965c8e69805;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h4a93f6017155b1b6547b887b1d0383c3317546015c047391f18eb2575bcc4c9033bb06b640f4c9d84adeff90f9e4c783e9b4d474c01fb04c3bbb0cdb6605cae4059aa2b27ca863867c3dea6d6e1dc937930788fb811b942472b798afaa55440e7246d020005ac47705f5ce99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hceafe544188990559ea11187506b47d8be6d35322e34ca4583f163e9bbfad488c364d31071a5f43b9d0957646e8ce9ec03b3016423b943586d79a337b670d4bde73fc8fc44c5a414d7e1091fd9725cfccedca5443597d25df0a0363a2591c6fb28adec73ac3a610fa3b6c2e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h3dfa95c2c276255e4d6f6dd130a777ba51ee23143cd5a5038ab3864c2f1da31b3a5ed319856a1eb47d5b4ef5a1e42ffc3dd03d19e9f8b4bddd01bcc5122dd131fb4b0e9374b27d65e833796beb1f1601097a82b5260c96e5d30773539bec1e23b5505dec007f024306fe8787;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he4ad44a021ad8d4991379a6f4a3dcbec306d569fd55d05bbd76379252fb366d0f8ae67125cd7effa57e254b0d74f72e8432108dfc71e1f20bfa57681985466a2a4c109b1dca2769ef7c5e56f59b2c98b955c37b9da89ecabd17cac5759c2a659e60c0a52219620bb64f98bd5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h75c7b03ed8f42b9ad0de8880a04029975382126e4f9e5f2b86efaad102d0e628ce04767c7abbd334a05a4584c1dd717af993479cf83fd310ea41eee97e53652e2fa4fbefa94e97197381de32026cf85b8ce49abad76f77a47240d924f5be4c124444f7fdbbbcaf589c05cb9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h1394e29ba82800523cbab61b3b2c4a0360aca0c58c0912a58e6b62ef41ae61a991826f130d39a4b00455f02564ee42065a94e0ae408bc834cb45ac3cdd72ea47cd6ce2340145e7d8046fbdab8d09b6565eb135e3eaacb4cb73b3f8aefc99867a04761374aee8af9ff77d7bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd2822b9d2f311cc22e87f2242ca23b55ad7b8c49f64d4b13b92a19aa66b83b5a12e6beb055d5d18bdc8aa7868df038e2daba38c8a613f2fc379e53c98f716eaf5699493bcb18ccb022567287ba74aed1f375a628d3ea80e064d65ba5593d9f8072daabbac55d8cf08b97d2f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he8e375d3c7e948c769b127476af5dbd73decb9370649c2cc75d3888a39272517fc9f4d347722bad0f659c8c93963e0d45306be487fec2a4008e3ffb3ba770579e826e0b989c7e7da05c3de600a17f53a1b4f8e03932eb8b525046696f713b613111551036070886dc7a31c1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h16ba58a5cd924c31e39987f60c396d6635454618508dd9157ecc86a57e3dc3695736c6d9648aed3d11be98c52e0b911a96076a8933dcfd6fc9f20337dea20b8cab80e13b973d19116f046c4b1927f34c198678c8de01d0c3b219e64fb892b922f1ced0e9335cdc035e116d34;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h3d541dce60f76c59c15741b5d3f0ed4a40f647769173a011e0b4a98f310ab7713c345bf7d437d828619f79aece9ef10f3ee1b86635b90fc4688c82db4889ba11051369541f896de46398ff44176390de1d39381a403047c7001dbc6392b4de0fe18777da11956dc0e1f85df6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h3fc135d42347800689a986ac6e182582372377f1d79fb54b715936dc9f151e2de1e34d4be46f76bd54cb6179575eec97c0f72f6596aa5b4c3834b167b1c912a08d4b71b2c95d8f19fd4ced66ae98238c0a22b08750c9b4970b3d04ae1d7fb410a85cec8c7b824fa6f5b59e84;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h82d6d11f8c6471f915a7fdaeeaffebb4f3bd7ed194978c2b05e160a2370fd2a65b466e96a0e61796f097c8dde3509e59c33366563e690266b28739afce8f0ba4c7ba3f78ed777ce775365c2c15a6d6c565d5b9ae4eb869bde6810085c99c480cbfad2fd92abcbe8217fdfcaa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hcd86b492a212c3bbfad2f17736d50e40e5a000f420cec1f8654e0e11938144ece3d0f244fc604f18caf8b693edda2e8775eca055eefd59c458d8bce993d96442e82ffdb59d1353fcb806968a882e8ee5358bdbfa12659a80226c01540ab9154edbd00479132b3d41f7e4ea0d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h2525e2a74c0796cf671b326c771030f1d2e81beca3eb3ada44dd5de1a9263d6bf58a626494cabf5c121b771675b931d5cd91552c9bc36e2960922257cce97e0af78468289491d4648dfba4dc3467db59898055f2c9d4b2d4339a123a70d9b2a99c745e4c80444a62dcd7a592;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h7f2ee0173e640d7bed2f7fe2bd1feb70ba6c3ea37b81cf6c2915ee10e8c8ef3784987f7923e41b2ace42a67e26b50025b112f739076d3fba14198ff84caa1e4fa4ff8ac7a1f7c50e4984499d652a249388f4e21a5b50a3f15ef02cf9d23f875639ca5dcde5e7612aa142781c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'heb9ae4bf530df58191d3d0490f7ed1918cefc2ebf2dd7403bce75c535e92030eacfb294f6ce7d06d4cf9330d894ee9cbfdebdd32d272a46b3e850dccd93adb828c481234d76bf56460bbb64379f43bea718c731fbf4a7a9e43e1a286b5a4b45d950d4fbc2724315a98efa9da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h1d6f606d8a60b265929d95f7507843511612fa87dc398229f97117d9690919a29efda4860e8a508458b0c00a836a43a325c3008a3f92d24849f19a5e47903272c10b86e7ecf01b8a70d266e7399d566a478c30d7071c00f8b47b7f98d42579cf9edd94d76ee5bc19494dc74e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h76ca2bfe1bf134469b60393348c2dd7be416dc19c79576424b9566c6d8180fbc3b72e46e8e033e1512b05383a08dad87a3f643ca4a38d5dfe783aa53bdc254e6883f7d75f24872dfe3b481ac3c7aa22a2c55f7e5448a68c6513106e6fd69809ecd7d5d82cb901addad9b297b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hff006d94164c52a0923cb13eef61a510897cc0bff42f76ebbbc5a73221bd2c73c0d717b5dc28969104fde708bf57c4dce8bc91daea96280b4791e83de1f01d32dadc069ce1a3d862348dd9489cbbccaf9de5eae049320dca86856203cb1a3d463d43ecec6bc3fbabf04568db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h5e3f34d95e8daa2b0046516f5746c6073bcd1281137fb932e78b0aa7ed183aa51d9f50f52918736efc9ce2c9f32d626a2b9a4eeaa9cdd919b6611a9cec9ffd3a1673826461f4a45dd06759a030b255cf874b0eff7694b0b32b811726b47ff40ffc2908f1acf18f24f2b0cd48;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hbe0dcc94e2061ae56265cfff2e90986ac3cab84512d6a8abd9d481bd21a15827a2741bdcde63b091787aef23dd96fb105efda4395b443814580bad99d8098a14b8ec5e7d9a2e77a3a324555e8c3dc3b5aabd12e66e923f1eb46a5f633c9ace0682783692bb2bbe26337b5a35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd0a2c05f0245e152f115da3f0c8e097564d84492bac980d4a4d580f64069093a478d62d39535637a44f7a0ee8406ad7e276cd0b426ec1ab98f4f09854ce54898b8c0b3cf3285b3815dbcfbb1aca0968c6da08f20d815bc96617fec3cd6dfbdaaae3e1cdea529ac76c20522a5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h49810e4e2405a2bd0716540bc2cd66feaa8edd748afea952530f09a0411d518c5fb5a3f7af331890c29cc9ac761d425beeacf84a5d38aa55f1f9eaa3877cdf34eebda7d90331ec40f5b3e9c3bcf7cc702049d40e71886eb887ef14ef9d82fcf664e9c82e07df78b568397fb6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h5c136949fe6f46960922a8a6bfd0308138ceb4787ae7e31c7b398ea6be933824bb4c262d8bbb12cff58ab926dad52cca28061e602fe94e8510d3747cdde9db1cb981a5edb00b1dbdcf6a437291ce2023c52fa6e4f0de42bfd0820d695f0c2d346ccf957b76ecd6121757d566;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9a3afb57f8f56797a4a1367f22fb89fc3b98652e370789658b7f3368b36aeb147e351e1cf94eef02d6ee8fb565bc4be70ee4089e8cef99103cde726473fff2faac981228494e426bf7c1fec617b0539486cde0912644f514822dd98f34fe6ed48627c49ebc25608bf0443a8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hac6544d9a3cda6074ec0d212fab6d54928bccaaec5830074b9a6f079042c5d9b4705c92995e269dc020882ee5eb8cb240a7ea11b17c79632ed1e6d321f97ecb8bd1920a5b407807cb6ba96c6664b75887ef1fe7dbf6b5abe8cffa80c7191c28471c73df09ff7039db968729f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h37f0e90ae74c17b5e4f7b6d02b295ccbb39888070d7c2994ff7ed10118b2d8988b0179b6fd7fa36f7721298659120cc8e33d1414cc405434fb71db0c75c786f1d801c3362a0a96a33842e3306485e9b44cb8822f201ca9818b94c9863724d933cad05a0c21246f08bc1a69f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h1fe0bf3a659380b68c83778463372ed64edd1b63cc176e8a57648d689617b315919b63d0a8d7e5b164edad7467e0accfd2e3485afdc5a2f4a69cc4b898eb3e9662fe3f79a9ebe3c6e0f21aa4b8328b0e836ce79034df8991e2a6caf1217872f9d0f45b9242f90056a3b353ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9f77aac8d65a4765a94279b9be9ac4ab7b2e85e45ac7a71d18edd0477396ee450547814a9bb2fa46d7599b6d2b2a866afe2b077378a41b15002e29778023506828532600d371eeca3c9b796ae8496794332e5f4bb89a71e3c5f7b91e2fb7262cc39b5e882b4ce71fb2364507;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h7ad3a0a26b8b279f4fc64061e18bec829656fe0bb71f55aab5c74f93481221a5c8c144ada73ce67fc5f6d300cb0e35e6250016e1399be025462c2ab331b3a6393bf5e84bcfed520027ff6243432c094cbe6bb032d0af15b6e1e153b941b4ebeab3f782b934290d004e853e6c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h979c5e78e122b5e07b69c606a08d27619b3a3383b63bad70efc0100b7430f3233c3d73dba3ebd33dc1816f60d8f09ca0497a474b6ce92bfdb5c937c97501da5d5c0f5227e5c3c70c37e2f258df04b1276b02c0e490a4f840116460c186eb39231a11a13ffcb0286e6d39a111;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hdd0a4dfa0ad20b89b8e064e0c757bd987a838de8cb8144a2c23dab6940b3e8f3ba3895001d31f9857645476e16eec9c2bc0239c6d4ca9d9eb54e0964329e694446f476cb4e61d6603c7e15498d1747e80df16e1c008de0b97e62f85d25bb86df8cbcdf61ecd9e60d98d3efe3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h1735dc258c8129051988dc2bb1c1aba36100b2c3c17597c73c9ba14dbcf1aaa82029f7e5271b29f76423fda6703685ce9f405992c1421155794befbec6294740c619cc2299cbc924e55a9e2b333948e853cfad047f9c02f3e2c4bbda94c857105126fb213b2c9dc8f3443476;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8f948446d90cc48c84463379097dc1fd85f288a603603880763bc706bf05cd3eb6deafd59d93e377072b6462435c97e936e6744db81fae77c7530056e3224bf802b475bb1d848bae80015bfafd2dd1d4cd70d4732dcfba1048dff92b05b1bc054a1eabfaca12c3290f3e6021;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf6bd2ddf088c2c25125f2768ccef08b9c3ee78a54e8ba501ff956c1d129e6671994ec4e617270957b264800369bd62b85ef08a3bc6058d130f3676f654a0bc65036b2d5af0771914a51e874485e2caabe102aa152b0be584c6ab3992685950a1e76713e63955cadb80d60149;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h735cf64ac1a535b5a1fc72ac0f6cd84cc376db46bfb24f26428f18c3b67cc35606906a1df120f8727c517d67638ff20d831beb77d11a8d4541be9aae036154023ef602422b06cb5ee6f6ccabe5083085471bc67e52a8ba3a43c475144b265530d982feb9a1067df50dd6926b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd3b5a159ed3e5544527eafed8e07d16d709845bfef9f7d12440911afe615420bf9fda4b7dfd0c1f8dbeee6abdc41bfaed2e5754f9a90a65850f2846866e8d60c6329e09091aedf9ec1ecea2e221c582a11c47e52ada44a6713079f4de10e5c13a75980c592cbf405f4135fac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h894debb96b72677260a5fa6a7a1e9c39d413993e1c70b5bc472f99b012b6a236bb30291c2b9f796b03ab2b64003be1715cd1d68973431c2f9e379db9ca17356f48e72bd6e6a4db4f4f23fdd24950c66a4a93578648a6475a1678298dc614e43db0cd7b89b40d131eeec2cec8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h6ca1f7babb697d7553075476da306952369fbf9e8a892d33269c1b1dd7f5d3d5b3a8e741581dad8ab51c9386d5303a25dea32d0d0dbff025609a250b72c66d0a04e17951b866d21c0e9799a3cfb4212d758661043125819f66e63b873e7c62e7c6e5b801fb79649e495039f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hbccb556b0d296da5de49f2ab757d554769ded5776d2414cb2aee391d16e195342d763b7f2dccc146ccdad96b2b9281ccfd4aeaf31d25d372f7b2fcb2f79d375066d0e5dc3a0404c46cf583760f07c426a5a7fc7bbfceb42c257080b219c12abb75bd7b28ad14107778986f07;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd8edc51ffe90cba21b29e9c69d87087c09e0b349d8a18c1045b0d1272d6633c78e2c4c65313dbbb3931bff72f692f884048cd19c8703663725753a37bb8ddc70d493061da6c1d24c918a05bb20c3dc00bfe5931dc9af482c3577361b3c6b0f5eabc50452446ade356ffe6801;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h64e82cd4bd2e3bf55f9f32337025ec38eb919bcaeff57ddf0bb3b903eb522d73203aa7c269336c57b374b765f7b07e336befeb89998d161120b0100dd5202fc30a661ff4d502eb005e8af1d6bfa412b2a48504b2ad5b201bfe3d67d328df275b2898a6f86ac75e8bb0692316;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hdd55d3ec0deb71ad353c827385dc328d879684a2353ce2bb90eca6b8d5c0d069801a019c9347cbe4a5ac679ea14ff1fb9a843ec58b49a40554464bd58131ae48321891d93e2b380b93754b5f2f8d5175256e51a0664ec02a9ad1cfc34e6c30f9762fb3ca53d673b015255051;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd52e73dd1902686938ec454551baa1e60286f33ebdc33c3d0593d1bdc4dfc5b5abec5de6322b3a702a4050dc1bbb2eb5e3c6149ac5e9993071d3da43e77bff9f877426b21bd34f46581050c2db081515f3aaf6194d5da900853942337b18305c553c61786b96e07483c7f953;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h6bfa067017812836094757f35b19a2b48606ed70377936a1be908587fa255d70bcb5196ad7e0bb813493bfb806ded8eb58762b5047bf16d530157234135a522c59468dfe603d146221c332abe7d4fc97c94c28baf96dcda7c894828707e4a62d0d651351d0d2ffada5ebd6f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h48ac6e0fbc49d3744dec1393580aad659d849092036f8793ebee678171c36bf66f9080986d54edee6438af6f856f5785cfcbfd72425828de06124e5288cf44c20da95e0a39437a9cdfa256a777f8699ff68c42e4361175a2e8f0b65f056c02992050190c7a58de5c6c9007b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h31c0ed0fa1d459bc3bcabe3ead2039de971e72faa7662126db8fdca77a7ce0ec480622b3672d850b7d2f97eb49140be0f0d0bc1c0f93e043ae9a754e03a7cbf87fa2bdbda62ecf10f6af2eba27b80d9510fb10059ca5d6f078de7c378e0426e2d4fac1d1ec1beecae3ae4047;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8c86c0de1f3d699f74882bd205be5f0b774a261d995f68c7993be0c10fb8b42167baee8e59eeee01893bb8ce33ed540ece10d7a8ced7420b8135af10893eff145c4d01e42146d5e5a87463afa6de6ae015641cf63070e7b24c558a93330fe1e00ad9e4680645fa9cf62e0fef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h77a0af36f977c948f81e09016a751a06b07c63c535a60df61d2f6cfd5994f50ccdd448920b5941a5baa7e941e77dc6772c646daf8e1ec190d757ad9b05bf0df7ba07f27f655e94e6d437b373aed8147e750460d7e72361ec899560b1b73525f7714d4d55b38a3fb855a149ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hafae54c3763ea01da15e7c603af3a71b3d196ad7346621f666d83b1b3a44e71541488e7492db8af0fc9f5135ff27b84d12ebaec17d814092d8d2288a1df2edf106b6e6b37823a14586adc5f372a1b5b82d95b3f4e5617cde595bb6b1d999e1591391258f8d44159477e9618;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he6e1df845020f83e32c8cceace6d75c868920c650b31b250ca716253b83bb8f96761f08cc51b591c1f97fc4dd9f65b18d36b5f90c185bb42c98ed7d2298ba976dec2802420c2b7a71e397ea5bb41d9ec72e199a6fbba31060c17601281638468537a053e4eb002f8759306ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h95ccfdbc06c8bde634eae9c09464c47bd379415a57d182a25471c4202c8f4333e928106ccd601811698e27c59c4834b550883dd3da6b2edb21210774269042f8a5225b33724aaeaae82b11179143983b62ec1e9e05117cb1f30b4c3bd53eed4c3a8a6d5299bce586ef8a4ace;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h665cb63a6741122abbb409e379a939c5b6622f41b2351bc54dc357199d85c32811db606163148b39aec44f995d335ef14d69c436b2737c64864a83b7c609ce01808e932c7219d48eeaa785a2fbb5ea4f827b92e320afbfca39d07686dd9479432ada3356f2be7920d82b97cf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hebb92cb9f71ad318ae3d6483ff59bb134026a2fd760aa61e782f5e9ab4b021ef1851eaf7df1f6a1e6dab22fd58108c42501e9054714ef01023efa5d602a7dae58231833c88a1b8deef4121167313b09cd2d461f9afce79c8d51761b76f6448de3ccbd7b46b109df5eb74a149;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hc65512af8a6a74c1db300f5d74e2208f1d61b52d1daf0ecc285e6bed73e9175efc2304241166deece302b713ebe593198b6bf316bc33229eb1e9bbb5003face162a5987bee2796bb5918aa693d1bef4e3af647aadd182a05124b021cc45069042b140afbef0d7f37c1eecd94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h10d420406a2c0c901eaa779739f2aba318cbbd1141c04cc3f6072f5ff5a2b04f90287341150d539d83f5c26dc6eb1b27370e2c7802bc1ddff8d8654f11c920a35748a0bbe63f7f9baf803347b4f6d26f7e16c70d1e0862a2f656f83d99327f16461fe768191d35894a1f64f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h45b1f632d1ec94f0ab1e02dcf6c0efd3667d1195bf85d35e39fd6754325c9ca7a555281ee7e263495aa306894742f158e188f60e6c7e8baa0afc59476110fa6173e08c41e0bb91115ca0dbd559901884c613eb7b380bb2a00ff4a874f9bfca7d549d18c365c57d3a8112b53e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hb42fee90515d61394885b9d144aa70eccf27e24e1117c03ca0828926d75dfda45617cd0309d97172a05a2d09d8d084b304da8fbe1281e4e9e3e777fdc1e79888132f3c1d8048a2d082009848689d554bffc249c4d7a000ccdac65b4e0cdf163d204c057a6d5f71d3db0dc9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8d0a7a320cc7062bc7c17eff7e28d58df774ea4f3d2d42f07f865fa145c2a301ad73f2266280c5caca52da6557ca8de8271ab22af6a3c69e01728aa61d6a28d8fab876135b173aab83a497201d9b51e33924647eae00f03bebe198c4b2edb50a076f5551284ad5e44740eb69;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf5ebd5e6dd48a6652282172fd8fabc9d98e7f417510fed988691c0f4e2e203a1708dc63f0127aed1b689309332fbd6211bee08203f4b766c0dd4c17b089ccba5806c23c8a1a0d097821eef57d2959d5698ce2c415e811871185377e0f4baf835c82e1fb1c4bb9f47e49b899d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he317afb0b886a559177ffb2a73b32e4d9dd36c77fa8a784746b6755f09ebb0e45dd932510863c21836bb087de3af1b96821606d65e71545ceb55bb9feae2b9ac8ba0f81e3f6b4401d17f5843dfc712ac60b82d1b6e75f7a01429dc27d303f0e700090def1b2d66310aa8834;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hbc6a8fbd2d7be6e3ed67bbe50ef4f8344bc60505aa11f84759af5f0061cb3cad840e55738bcca598e936f30c960465597f1839e67f26322f9bbc4aa9eb5681d820b04aba650d02f2cfbbda05fb763e1eb7f5176cfb92c5748150ae77d26b2b82b60f146217fdad2e79739a60;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hcc340ceebdd1c1b45a018be1aa2e3a2bd582c3095c0896d74c35a824f486f6b30a155b46c80cdfbde6199f46be2768b396678fa8932821667f7830b37528ca20dd52b4d41e6bf2a4a30dec967208bf12ee926686787483068da5bdd8d600b26913f7944e735877d4e404451d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hfebf84176e44b95d0830e75a350a6492f74b10823a5b799b73a49763a52b67ca52c72def09a098bb7a0628016c701741707f2617ee60add9e5c2d6cbd20558b2347e0afb8b5096d5c71af59508b0ad6d0fa193faf7e2d335bf5d20ec4524fed4383eeebddff2541836c722c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h17490fd0612cf9a889a883a3d4e54300aaadb2e6ebb8784eba9e73bb1361f555439523ab123ee352614050d598732dcdd45b159c43eea5c2582ff90075076a0f3a29e8763bf5fa41b37991d31d0862143b790847d77dd8f3fd5c7e6b968e8519e10aff410dabbe6f783fabf3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hccfbd5b113c5525bf1f23bcc75d3c21cbdd7eb340d543d838833511bab01e35409a6d6dbf46bad443242393ccfbfaa780c3b4a0dc20dbea800c32c58eeb1f3f1e8e67cc6b8873c98d364d915bbdde7afa23cbb1879f044d1897cb19544ecbaaf6907c83bba4b4bc7d818e8b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8bee02253a4911b871b1b0467d49af38c56370bd225a07ae67fdf41d1d8d7d5907bf69c3d8da320fd0aa658e1a096351c5a99558ddad3d0bf1c2b557ff71abfa6465123df86ef2d8840649a565b6eba90033e93a5bb22710a3b74465a81508458a76baa8e5b360da7591581e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h76b5dc12330089c82ffe802b91e91fd01153dd5988ae04c096d3d7af1685c1c6c55465dfcbebc93976b440f3c4883fdc61c5175c4d0fd9520fad0a89d364da1b10417fd9160779587c94b35588b1831f6a094c4a62213de2b69f52927f6276bc7d9eeb8188256f35b18584f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9268417bd6c20a03f4350c758609edf8a65c775fafe0efca4634951a6c19a21169eff8a6edad41ee0d3e86b627fad65dd7e4d12f3d3da69d8143e39d9b3c46a6cc7ddc4e6fe4de6a5cb2b38341f1ff5b98854664473bc2a8acf5f0f26cfddc2ff026b33ef576de1c9e91f83f;
        #1
        $finish();
    end
endmodule
