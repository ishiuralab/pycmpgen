module testbench();
    reg [28:0] src0;
    reg [28:0] src1;
    reg [28:0] src2;
    reg [28:0] src3;
    reg [28:0] src4;
    reg [28:0] src5;
    reg [28:0] src6;
    reg [28:0] src7;
    reg [28:0] src8;
    reg [28:0] src9;
    reg [28:0] src10;
    reg [28:0] src11;
    reg [28:0] src12;
    reg [28:0] src13;
    reg [28:0] src14;
    reg [28:0] src15;
    reg [28:0] src16;
    reg [28:0] src17;
    reg [28:0] src18;
    reg [28:0] src19;
    reg [28:0] src20;
    reg [28:0] src21;
    reg [28:0] src22;
    reg [28:0] src23;
    reg [28:0] src24;
    reg [28:0] src25;
    reg [28:0] src26;
    reg [28:0] src27;
    reg [28:0] src28;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [33:0] srcsum;
    wire [33:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h156b83ed7b6823016782182fbefdd1f87df672b99123b86b8f22daa343a81b8aca71eb9ebd212ec429f1b198279dbeadeaa8333ad5d9273029938029435cc89b9017d66dac22465b856a2f7d462da616b859a570111a60e781b500f02d93fc34fb537ec978cb97edad3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15e2368048f5cf67269178c9f93c313001dd8b01979b4ae3743b2b89302b66669537bd690e4cae7e7bfc25e2c79299707cc938a651106873a1258828ffef9e1676eeac86f29bd529940ce79a410158025c96264399ac3b2b27b952016d2ab4c8165cb2010e837fc27ff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c6ef3a772da32202f627148234b458b4228ce9619f58f177c41a96561362d235ddd7950506c2e5bb8b9e55be86c665e752c2cda413d61c171877262443e3e22829989b5e22cc36467b9f256cd36012d152190a700a1f8ef1d603557ca261542b2fcaffadf48f07bd0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h131afe45832de4697884633c97c517439c9e109a2d27c24aceea1aa5d067709a8874a700e1e908bfe4fd93defa5bc218efcde040089801bf639e87e6ecaf6a21846c5c191e62e679e7454bcdba168a0f8997ee22aaae75519715a9da906a599d6fd81fdf74376e0b70b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4854d6dd29f2f5998fedd7dc04ca0bd2770367d793a4c3afb6f666118e27efd30dd3fcf9d38482e9e965033a124f1d975aad2ec8270cb8ef18ad0594b4297e89b8f5d5f60bba7f10d610f7e9b13461269a83a7381af856c8dbf2c427644bf4b7b5b4dc11b4635c6dd6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d6d06100f6f425316dd8b57b5d44ffc3aee5ffbd8d66b8b7e29983ed0f9965823d8d22f1ae9bb0308630d8f8d6d98ad6bf2a4717ef2f25f94c692c780c0f20a84fedf7c9ad04ce9697b2c398b08b39332e02a6e836ceef527627cb5d10dce258659cd2245f686628b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h606ef243618514b62aba5ccb51980162fb69481b0e7af75f0140546e3fd4d8892ea36b5e80e784d91360bd9fdae504716e59f4f75ca627ffe56985b730684380b809142519255ab0911ac1ac17391d562310f2f727000ec024899f1e681f89135573134be301af5999;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1805c84ebad2604b2b304d1e09e64c930f51f498f813256910df1254ee85cfe1eadd4f6d8d7f7ba259517caf6a15782280d510975534282bafcf1605335c4e079acd68f0cb57854adf3568db0c633ba5642a8d7f30cd0add8caecb229360b421d8a3de913657ac7f24c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h128700b211ce958c07548a86dbb48218f4d55c73854a7649933a1ae7f161799020a627d2595276cae31884096a7e6fde5a93e55e60e3661ceb8aadd542cac8927832a06b8ad73beac4a1dcd951deb75abbc35892e98fb4141356af1c076c6695ff2d086bc930b2b24cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc44b599bad97d1a05e9e202bc25831c7e5b006be568fab6b19d1f9895d2a126d20939edad1f16809cfb0c01676770a3194dcf699fc4f3731ec8d966015d16add6be577e82a3269798014bd3bdc7607575e08958b148f80e8375705f98fbb69c19fa91a2f65a613c7e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a7664c1678f630e93ffaee04e63d7dc7d34314d58227af61ed1a117c254a5b1aca47ada06c72f8e4336683105ed061c9b5832ded8872736c78bdbcf0ddd13c037335a4ca7800d244bbe4ba8b2e8e18ef453682e30bbdd44597f6b47fcd885e9e9436bf50e5fa23b578;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11bffaaf5f9cc23c1edc37e3468bbc1ca083e15ba1a353efeb358548e0af0a8c35cd831596086bcefc322962c3d577d4d06cbabd5d2ce15d811d8226067be2e5b1e00d41b7ed79e52b7fa5bf831295fd6088dbd82bec2883ef3e66a750a4cd4312de1fbef09fa570b9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac8955f929f049d259e72534b2a1e58303562645e1330eefa8d948587aefd7de79ee2180e5d360a7dc950632c542f9b1f3b4f699f9c3add165682fd7e3db3f97b1d61ae1d050e0aa61562d5147ad652bc1b86050c6b0ea28e4f1973efbb391ef5d3157cc2737d38a09;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc97945e323feb1810977d327874e1376d00c009507edc602998f34018a53d2c229b4b06b5448d71cebeb3292ff0a14e2c8372c5dc1f1ab0f0861b9e5b6e8bd49ec3cda437dd38c6d5f8b4b338bc2b58a2fc549f3321c7ab46bd52d0d387a5da497201cdd8e71d1ec8d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h151c8a6ce4267cf05c162cf87711b704b27e0ef3ec88c21a79a8d14a6545337d47ee485d7fc1db5134c7905c7e20829d838f856a53f7f1ded9eabce07205d1920ca7208d100bd515bac15139c6b0edac57a844f981c1decace884b54a6f4975b8681d2001d179618b8a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ce04aee554a4a7521ca8c463593aa8d0b8ad0a7ea4ee5a113711f9c030a556ebd057933bb7c2acf0c5fba30bce73a6531a62c23c48740578212eea90db9257d456f388984b75a8943efe7461ffac220366ff9785c7b9948488058011d2cebd12ad95e0e245d09ec71;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c755bbe3e5c7515d14a2d5e1df2babdc5599b680dc585287e253737f0a4af32b232636f7514c0334ab024432fab9e09f65660ff2686686c3e47a3028266d7336ff019fbec3097ca9318e758a095567331326c927062951c54b0905a8a82a0d79be1fcca0b1f72f5f7f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cfdc897f080b1816a3667eaf245d55c3eb6c716186ebed9f7ef12e650409899f11045b60b8756c942389101a91e15136c24fc3dc7899f084f33e2b039f49cab486b9c90929b846a64bc3ca9c88698e51b278c164a595f3964f5f4d5a17c788c6de40b513dd451062d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha50ff119279c5d451e9c1308d0121dd4a781fd98a1000bc1ad690970345738d6417828409073681f97fad61edbdc71899099a44e3125d93167d2bcef1376a376c95ad1d532108ac60b74e97645d92c1ab8dea74e9ed9cd2511d5eaa6e39874fa513ea6862933f200dd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he38d6132114a84adcc698aa13a4bd8c4cc811ad658ca9c8e314ce59038cc8cd5db078baea9511a63b5644b5d52aba87c721da9e1e344abda348485bb8b2127b3595cc541736c6e326559ed408322e92362cecdbc0c5e6da96eb4791f69dcd74d0da9492aacfea864cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcc6a30a9138667c05dda2d2eceea6b3a0e533d86e847de8d2c1063f0d359889cebac8cdf3318449187ce5a267e657c3d993db31ea3b4cfb558b937233c8986bccba72fdfc3894e9c4597ddeeebac4847d37bc0117e750dde14807157332daa93086016b05ea1ed3ed3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13c92c1fe675d56ede6c0f557277f08a8169f4ece33fbe22989f56febf09ca3f9664233e2186571d5581cdfbe634af724ffb953b0d6f14a833db2603c528126f18cb749e3d0a3e653e22aa276eac5d9d9004dee7d2f421412c291765977555b6d864fbec29a2a12086d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19bf34d9d0b910e3e03e13c88372575c421c38803b7d29237c0adc516e78e8023407574faa47bd2cac0406dd0d42dc8ab0b927bfdd7ddcd599e0a682b28a366694bdaac8d882a2a5e50c7d80836eb430469fe5813f7ca0135c6860edf8ba4b4c0a21ac05777e4b75808;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h193252562862aeb2f2d81c1653afebdd8b26eb98a8bf62b745ce9e0aae9ae8f2948240fcc4c9249b20af7304d4f44002b232142bcd34b668a913688c73a9955d3d07329f5572f9d62f2b956de6bbbf8b47792dc76e8881c50e8ad073d7ef7285fac8deecce1226e87a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7bc551474f7a2156029d6c3e2c6dba6b0647487c4cddce199e556f12c11371485164621dc3121a2ae2cb2985aa6b58d58b8860b4ebf4fd5f5b527b973b9c753c070ae8ddad5509a10586e81095f84f07aa4cfd530fad0ec63f7ca7204869ba758327c0913f26386fec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc4013e04a01b014eb1ba476cb6a200bce9586ad29e8500210c5e14d2644345a288fa635f49f5c93f4ea367646a99b2b94185c63091c4a6c4c09393d7d345e9e328a660c7359437200784af19e6d05d4eb3226e42b4d66a5a5e84dad5528863e03866575097bd15bf36;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h74e98465e9515a24f8597beb1753a7118f39d32018a151c0cdcec819d3fbfa15cbc427580639081aab9a682bcd6ab79d0fcfd1cb595693872ea1f1a6039c1d99d605c29cbee45eb58b5590df72ff2eb7f9d157bc215fb7bca86f62487b88ea26c3ac8f46b78ebc5beb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed02813e380a236d9b29d99fb3bd67a74f1a54c0ddfa1c7478cd5d598a4904883a48bf1d3045841f0b6f0f80de8bcaeb20eec2c3c6daf925e25aad2451eeda370a704157e1853201cb250731c05855ce2b70eeef506e5a16e396595b60d8399a23596ede0e5dc0b84a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb77a2ac873fc75aa40409e2feaaeb3585cfa9a08320ad5e78fabd64fbfb522495fd6304c6209eda0d9338dc4c86e3a269c1c6567057c05034345f157c7116f79a86316f77c97ae631acd02a1b40aca18c5cc720d6b634921cf9d1fc845eecf2510f45ed4e48952684;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5f1b27736d5d08ef6d54363f15a519ab1fe2578a561f53a44c3df23b1c09bb3388321779d6783a3ef3820b79f2766793a8cd56eb505b9947d2542e1202b046d021b236e333f6edf61a9b10a512530f3f561dcced2d328e9dc34dd1ea45018c7d67a4c31784f6ff503;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf84ef47af468612d9fcad3a7bc62510e35a2ac298b49bbebab139e83ca5eb42d16f014ca896c6cf1e40fd98474834b2928e86c9bdcb5012e1aa523d22ff905041e5179500f9dfdd286fbbe5e33d0576ddf0fade6b83163a7cd575bf2354154ef46476f856608d10485;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b1a38f2a6b81aad8a8c450a6b05b067d7e683085fb7008f05c177904e15e119badd2445c235f3eef056ba95f2220f7d01f6a120ca4b930d841ecaf1c02c37f8b6cfe75fbf062c8e4f4a4e3d4dd8e543e3994c08667ad255a2de22c3179290055bac0da9aa3bd92b58;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf09ad0b4bd56e3b8287c87b694449e5040724006a153ee5c07c11ceb30eb146a1e740d3b44fb68c370327324efc7b04f7e1c41d41e7697ffbe164e63081598e4565106b8187ba8944fd59507c207da1ab1b84f65bf63ac319ed1744ac98baec3b384b7fd080b3ea711;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h44a461f2a99cb86c606034ca4daba7d93f75eeb3c847af7b79c0cc2cf3f147875db98a48f9808b1dc586733d316c7617cc1b1b6962bfe347bfe22bc3d3e07d2eee642dd0ccad7f3af8addf0d715f25404acfdde0806a1362b9a463ced88872bbf3229a881815c4176a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18fded6f28c2d9c98767744753c5b6d6f4dab624f0e6bc064f93bfa0dae50ed64c9757bf7245ed0cfab2cbc7d1e1795b422e3c8c04c0857f42368e3b5264a8c872390fc7c2d3e976455fd9544e3e2badc7e949aac0e5f92edad6a1dcdd41af3501014dd6a329746fe65;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h162667fe2e224dd56b6f9e19f090588935480e98ffc6f439f96c6751da712e5e84fe0edaf4e64142f8a598726acb389bc00f5d5b6c693554e3e73cfee0cd2820b0b621d9df82993597417b055c71e179fc9b842f81fd9f12f469cdcda8352a523dae36a173d7c85cdc3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf489545cfd72fb33f6b027b9cc5f13dbe2e2342e2156aa0a5d2dd2dd29bf7a84cb0693a0e6cdc389fef1b8b466708b1fd2edbeb3b815be11d7b6207368d383a0223aa0cfe1857aca8806a2aab05bcab77425aad3296f680b2d72e3e8f432adcf0e3a802c651868a34;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h154713839711e5b0fabfcf5531058f080ab1d791e5729fb0bb4647846fc5239341d0926bf2c805b15a25c57cb76177a47c679b6d083e620fbcc1d9b4896c73ec2af6a964050b0fe4de8bebd7e971402f0aa9861b4c236de05a78f6e3b6f5fdc364ea1f9398f8a198056;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1397d1cc3091e18dccbfa4840839f9aa249cb0147262e9ca67c1f856a89467507df2150ee85b2f00a4b3496ffbbf4e89a64c3799786ae16e815ad0bf158627e21cfa866f159bdbe6360e2189046b2b3c378169c482473c9ab581f9358b0799a55a0674c898c2c88b94c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h110c2b78a1ad0cb43413d0baf263ef68239dc52f8fb3780f5d30181920500363f225ba7969b0896f6cd5a166a627a42c3492366985379c5e4d08f969a4950193517b48fde31bbf11c9bf93efc4acd273ecf50b0484392bb8f91bebe3007912a5ca81b9e2712fcd57208;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113d6182b153669ecb26c6f8be713c858666e3e74309fd8b9e52774a60e9cdd8ed900ec23bd6b91b133825f9a9566f5c1aab8bf4a133775028ca74ba72308ce3ff918c6a9efabb4d001e88cebc3d9820a1774f8eb7acb60dc7914da6379053f2ddc4270686882f9004b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1afe817f3506ee8a71fa526271f464aa9cd4b5c401fbab143fa814a5e44910f15fd9ec1e33d2f209d26f09a365c0f1dad9169cf4cbc42a1ca29c9748e4b3ee9de53d4110ebd54525ae2d17448dc11bbedb686b8962cdb76c95bc8a8094fbd147dc7acd32b8344abfc0e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h140e386e6872a57d0030c5028c9138ca051ef892fc42202889b5f55b6cb3950f8225a7c70c5ba8666fd9e29910cc9114200d435910f935a7ddbe276db3c53dd2cf7412d832182c4db6560890e0865f47509437ca759d3dc7810da315583e5de12ed6f880e0800a3c299;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf10a2b3e9bf1d01eb84d3a533c3a8e1444d3a59ee2a7247599bcbb2870e4d044e5467b3b41bc1b993a6f13d5d97f97dc75fa374535cee6f42dcacedea09cfcffa8bc6e9e4349663a6f4505f3bba913a763b43ad6674d503510a6ceb795631d538b1f5feecbcb48b34;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd95ef738a479b851d07ce4bf970a059c43320fde3162afe234ed39e21a6efe4f8e3d09314b7e60337a5c39d2aacfae5b65a39129573f05e2271daca50b9bc9c98ae733d27a24fec2d382e0d55b2d04a4f2fc04a292f5a7111602bf3a4427876b6531fc876ce7d0327e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c971b8a3f0b571d67ed71189cd2a0e7b2ec54a0dcd81dc03a7ad755dfed42739b2b058ba5cf2baddb9b29e938588ba0dc4cd84c358c238281d40afdd866304fdc0408a498b8f6f48bcc6f9fe7dc34bc5379e1d8dbd3fba51bbf58ca6a5b0d54a27a32443e29828ca69;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4318a920195cb90efbeec80aa30bdf9534087cebebe7adb1ddfd252700c70d4994f4b5dc246f6cb992d8f3b469e4adc327d5073484c841b812518bf43ddd43c18ba56b61aacc373e1d1db0ddd34d224261669b83d5186d94f6c21f4e9aceb1e9c22c0eb8b924de282f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf72fa377f0bd177f5defa20ed9922f7740aea5c9b496940c427cee1eb755b2252bcfc3e4f7c368de75fd610e32be430e1c0aa69a14aa5bae52111d656e901e0529039be09b10721875ab78cc6a6a7ca26eac23cbc7712bdae013be2d1134fdb32a91aa0df0f5af1f55;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f04ea659eddc91a4b5116435b65340030b8aeee7018dffb1ce7fc12fd4d8a7803e52c9cc5ee7eeea1e09d1786e5ac91d119f00e1ecb32ccf0f8d70c835ab4101d61d9083751cffe2169daccfc7bcd68ba80f16ec4fe5426a563c52f9c35679dad8f5258755b5b450f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5177ec800644c64ecc6190cad7d43f8d44e6bedf28ff43b141e327c55946fdb88e664c81061b3dac09e216b14f27502a7376b830cf57c59ff9e63257b70903394d186b6ac45c626e6baf0d9b957d3f9b72f73a354c9ab3afb5186b44e29a371857810025ecb6062526;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2f6772d6ac99bb6eae4eb577b6e606d38e6ffebed78410679ce7cd956f1f46a94f243ea9771f3bd51290750ee351780c05242215b7d115bde047f39d1f691a7691ce7a8a3f160976616f789184e88516fa6701f93a727272bbf46ee8a4ac7443298577ceb0c663dae5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcabac665bc7305717d06a161ff211252a940117b44b9d219978f0a340fe1e734b2950cae54f98778c90630800b2fe365a0a2450b0e40c9362ebb42c27177a266b9188a7432f437303fee1bfbd79148a91713e08251205b87d86ab93270291d6d28ae1b1060ced7fa84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc5f91acdaee5692fdec40e27f42103f7aa8c8a43859cd21b6f0265bb766967f750a09f9df62bfaad12eba1e596786b83851ca0755c4ba009f27cd24cded537c3d21d0b0d3222193d81352c07d6e6a9d1f659357d44282ee9e2573167a98357d7c025de18cfad322e10;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h56c5e581f92fd428273f5109015366dad3d4b0f7761f5d2de00be06fe6ae7b1d15a746a87ac0b8566350281aed5ceaca197b5429ef94108af4994fdedbc7221f57e4b5f0a2dc38001c1bc82f39fe8a30f5a7a77ada8ddbcb5408ea1e33ff7fe561af28283c6c2567d1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79f22abf5690b0584a55d1f721b2c5db559da3d0f7bbc2bb480633671b013e661915cf15cf4cf435c160dd36a45218040dcad1110a36aff5ddbc612b65521211e87f5c67867010223f744a75dde25cc8f2a963b313e9b11e340915f38cc638d1e167e3d145b28c58bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ddfa4f03559e7079eb36257d239033256a03e66dfae796c0fe2b5309575d147bf88f0fcfb49e6b795fddcfb5d2ab7941f5f2f839c3e96e1e947cd2cddc8a04271c8d6ccee5a8bee83381a9fa85db248fe3e99fea83c6e19069f4ed00af593b06a0741038408c95f11;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1263343dc2a4b0695eaa49e646ea29d11d1a6f1a6a90fda3b735fc5b0e1cb3d63f65100ab22d0d7bb13529d7dff693a25296f2ddd4dc31661801db093185699350e18c2021adcd0a58ca65152ab25e7541880171e94144640943ad7b8cf59c2c101849b591b14a203f8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c003aa791238de093473746dba69f064d89057094fbc86d00c0630d95bb4404a3d447b540e8d9254ea8582cc61f16c8f9144af4db91af8b10f3c1c3c8804537724fc8ec1fb8f388e377a8c851519555ef206e9a2476de04a23f54bfa2ee210e3e7f0c1fd37007659fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d985ea85d0ee67e858ff4298334648d936d0b525c3b3bd48d225036e65e50fa8251fdb16ca001b1f890c67a5014dfa8780cb857bf3aaac232d61899886f2802f3841d9f83bcdc428b5a01d92dc2050023b288749673ef3a41a1a310ff9493ca06a6cdf1c9c5edbd36c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hea005484e03482a4fac114c66ec18d244f8f6c62ec606d4bc8bde8117e46bb9c9aaae2635061654c037100520e89150627583d2edd4b080e7cc4eff6223377d5410638ec5805a5a0fcd11025d4fd814c20e4d3408c9f12bbd046ca71eb98864b603d32e11e1aee5974;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c348153214db2d459f9a440522abf87c82befc15cae8d76519874735cc8d18c4e721a6353329fee485d16890819f279f6f76ae41357c532ac252f2475b7b0f2860a0397220476149654027e253a2b22b0a1cea9f8c9c68886f6f6ec25aa342009ad1e51fc44da3d4ff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17fb3482d60a7736269f8c5b33fd7318f68db61f2a15620e1c7f6c8f0eb38e1f125a3a9287ebdf2dfefcfe4de1cb89b76f5ae2cbd5d59b11b61a0e1a87665fb8758196a34e808bec01c0d0750151013ed58b925304ce041580d909ee9c0a776357add8de2b3b0349e6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf07db734fa6ddbec41623b6e8147e2935055bfe1af5a686a3434931a59aefd05711a23e0571ae4ba9633c9091fec132db311b3f146dd2121570c356144144743702342136002e71ebcaf81431a3ad4d5384dffdb6712bdcd51c1df7a98e9af83ef1903212649b57c65;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b76e5edf7ee4733c46f3863a243a7f163003d5038426d49c55b8bf727440b83936e8f3eb2ce9c7dfe1781826d915dbbf04e2b1658bf2c182e08c14f40a4e18ed49c99a67152bdc460e8cd6ece2af8f852d28c49e095ff24e0eeed321db2342003c780d14b07b0825c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d76ac0630325cf626fb19a5dcfccd9c391f9fc9a90360cb5edd15066c8c8f12f8254f0d04e4ba792d5a8306b7ec21323d075fa411f4824b8a7c09a5945e086f0a027945907ec2c5b8ea5cb4481124a7a7af8436b37f42d30e0b452514497d6350ee48cf24e671adc13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10801202f2af59be22b59d9cf86fb782962d20abea3bf53ac9dbbcbc1d1bc190f2fbaf350e69d3f07af8d100c4d8750c47bd997c10ab6925a7cd8813470fe4308925d64364bcd797a7fbbb50096f7f7c2965a139cdd767d3a42b5650d595adfbf80757012a1d181e44f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11553f114f021f07a23d3951b69a81db7ea303ece59c0cc680e652c89e6dbed74f74fe4af02970566d68af0cf78badef81c6a26f278fb45e73876213ff11c0f4b9d866ef56e7a8f6171a95d729d67be8aff5a6787db3e26650c4093b9a1c1f598ce79b0ddf7ebb72609;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d90ef346ce2a71f24dc45db1d0595e5d2e9df1b7ff0dc99a0ba3fb5ad1dba48d745afdcdd1d0b452de11d053f63f3e749c97ee9a319a44a39c14a2943fb4ab67965e3bc267d8407f373be41fb9b07b4bb866afe1388a8fe743f8e536e24359bc4b1b435265a37e9ec6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15728375c79a3ef55697cf6413411b22203f2099f79c6ca62f6e039042979d9bc6072f22dc06dfcd4cd958ec35311960b54d9b547195792ac597073e9c20179a5405c2e695d1f9a3bf5982eb5350c467331d082bfa96a3b60c832ff7a563830edc830914257576e570;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ef178520f1a2b1429109dbde15d0d4ce1ae45be45070eec84b30732e723a94eef124bc5a63fc6b90f2ad02dfd0435ce320b7bc5326f47099956a7bbd1d34a7512b7dcad29b1a7be8dc6b0a4fccedb4c990eff7a605f9c3eda0866c2a40c5d5f8285abc1c0fbaf6f14;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc9dcc83a6c286002ab0f0c4da341e6082ac9feab8cce577ce313b290dc17eb9c52610a90c521701611a608c592ff268d61334aeb9dd49383daec37137c95c2fd53b46efaf74707f8d36fd3b51cc011a85c74a1f0d20f782e27968b663ad6c656a39f2a3add30e74fa2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1afb3b926a73d485a6860bb53152b9701da1a05f8e78a8bb74a3cbdb0fb6f21aec8930750d6c35777044d680b15b85c6a67f1d0808fba6cd86a7f7d6536b5b91d7c6d81bc27175c0a9ffeba84bfa759feaa71ab113b91ebaf6e509473f1663c790289f82f8634d20fc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heaa3113d391067032de4374ad5ffd821b4e2ba00d14a84234d41bd376deb3e7e3f19db6fbd1e8977f1843ed1ff2eaa6a8d68f954e79109f118c474bb557780a80ff6521c6c5c69b50febebf9e01afd9bdc5aa4eb1f07957c3c9fadd3a7e3f7468b0b97a42cd75e982d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a316e49e2c7579538d8cd2b725e47e220fe394f7a4eced7d7013b6cc832fdb687289c70ce7ba3a7caae8405ad0839e3d986eb684c0a1fb3edd51083a6bc53dc8f64b1b56fba09495227158f00f6deffeaec34d77949d767a1b30c40938a9eb114efa60158dcd12cdc0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2600649b32901e91bfa05ed94f981788a2f810ae1dd0201ee90ae71d3be0783025587ce516adfd6b81244c5319fb02744921053206d74d74364479aff82381d1c169f7d4ae35a9d44fdf07ed1386345578083a4df2f0c1bea90f5388bcbba1e1297cf3705c96964c9a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155c7ba8c52e81efd5a72e19b18d68f6605334084e298e7e9926427cf46a752cf777bab027b418e2f43a93bc2b9003df4d3cff98dc42cff141ecfe59b7b9128e87e088bd282b467bb40b79b1c997e28ab8b1672df39db9b159f7d8530efdbe09fee013a9427c11db48e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc7b0f962ccabac90f0036506bcbf746f6033b42cf27ad0a28099a807062811737819984ee8778a55efcc79eeb5f5713fb366d50cdeeb35912121c17450152fa0a0ee80ec3c8741ac04139be14b3459d30ade1eb4bbb2e2bf14d9cf9a704a6dd90e7a78cc91fa38d23;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c79170f721e51da8c1839814a2b45147ca21dc735d1f8c89af8a3e0d268a19d4cc57d580aec316ede7175ffd61f6fff2016607864a7b9481b0cb0b1b7d33f1e0e1110fa0cb1975288fd102bb4ab0aecf7c1be0c336cc11067cbcaa6e4db3bc585ccfdd8d6045ea865;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha82ce353f6b237d53ecd4c48a077118209cfad804ae69810867d3309e610e09558837db2ce85238851ffcb358a34b69281cba79cf585160418667b665a839035d5bf9d91e770e14930c388b2569a5c2b321f977ad32783541e532a6976ac007b6eeafc0b3de648e894;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3c419b126b5c4adfc659ddebdbac7a08b40b35d44c772ec855503e7ecc7c4ed66de92f29d2983038a56807a97d12a9b3ea3c5126976f5740c2b400760b1928569449bc70d2bd2ff9ca27a0197ec7dc6860723bc4b911bbaa56107a1fc9206c326ffb7bd226e377f081;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h176e0a2cb152f74df0728de6d33f43365a5bcdc2dc0f17d75685b2b20130fa5ffe9a350bd3762c473dc00ffd4a37eb8f3dd0759c57beb546a707e79939e22a7ec87bb641b36e93c0911da9c2ea2a32c8018092134385b120f2a5253d0a15cd079e0cdb339960b4cc347;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb457c5e5c7f2470e1e9ad8245f4ba0dfdf4f1c4f24a6c934d5f2621ef61abd186980a8df6a3f2b9c068f21fa9dc0963c6d4bdb43e259c00a470190361938401265180110c270c273db6348c44a8a4fc38dcb0c32773d8bf68daf6446086b7b6da970e9f20834ce47e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h180fa6c2c1914da956a6f806a2c43445871184a6acbc2e0bf6d2c46e536492ced945baf779f1c229f4912850d9188c9859269be415cb9615429e4e082bc72811105e56a4bf69887bcd87958ada3cace61026e2a85fbb8a410a0639fdd17c006f90ecd441926147db397;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c856850835f7980c4e171f471ad31776847cf30da5cdeef6bf928666244b58ac5822e50defe07eb1c925c508863dfd61eb0cb555807fb9d8f9714e5a3f204c4944905185efe786b56ffd9c8663e1ad653e9260b96128e19ce8e2c31c78482d0deca918440e2774a86;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h88c1d7a0e4bc47ad62011d68954bb3a47472bd7a48da9819ab084a87a4f0afd1fd78d257c160884ef878c587ccd8d5072c874b04c2a0e2a396fc00552097beae6f07d47b930161318bf740ba4aeeaab95cc5b94f32f051c17cdb464d5b7635dfd8c90ac551b836cff6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f7c83e3b914178f7731406a1ef6dbceb5c3b6f7602ffad418083475a2978a5922ac27f9c1a1df7a794f8852748c0bad8c2c5fa0db0b858b7fc06eb0ad50ddb3847d68c0063af256d65753bcb5d566c380be16ff37186a703608a92571253941c8b461e526f15100bf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h937df597d9144149ca93e1aa2e7142f00b07686a3634df5041839c3c7dd729d523b222b06cb801584cdbf62d188be0135fc8bb9da24bbad90d536f31d4694d726f878e8d79ddb289b10bdcc0848df3d788946681007830469e49ead881eb6e910814c66a051bab16f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb28710753f41b27be7a9cd2736f143e446e591ee7c822cef83d56cd7f0a00f45d93a868f5abd94cbeabe9f0c8c21be645b6ad4112c26d5ee921182971557f2fe868a21a09bf9ea71c04c51a6e9f4863e5a0d1f091a69efeec0048d080353039e5594c198528713ad84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hacd9cdc4621f8cba57e48de711fc3b5a4833709a77a9a803b329b40170c2e3e7deb756e591e4056824d88ba102270f88d56a6a32896acdd6999c480e2c052cf56db4b31c9bbd4c2c1b1c62af9c486c2d3f065a39a4fb8652201b92623f7ee3031b4f69442e59c0502e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hce2bbaff7eac949510cf03602fed8e021f0326e71711c794db57a3cdf3d5b20f5ce86271bac777f2851299049f72fdb2000ce790a88f3b8531c4b5ad6f7aede1c3cb95c56c2d747d4db70ce4a2c121f23a4ac320995704f7359d636dadfc26f377bbf1e7e08b7a3a00;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9cbe7d3676513a1e1ff556102dcf2af5eb3f52e0c8ac9c9a87926bd28526ca6627ba5eaaf0fb1f713cc6f837a7047ca6ff6a2e33cf5bbd5e4b41c9c7c9e0459d327b0224fe88c41d8d4680d6e63ce9e089a7b09b1edc4487f4339eb76feb7135ff9780e307dc5f8164;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf07275c9715d0abf3c492745385254d83c2f540d113d4b7a14bf4fdf92fde9b85aceb7050df50c63c607cdea190333e24135be626286ba6f54da19354bd60b60e90f924b1d9d29c22229266b2c8dd96cadfeb9bbd80d37e39049b26e8e9324ee1d34ddd8c5d88fec3a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1401d6f26b6e74532a491d76afc31d6a1538fa7b993e04d7683e099832302c6a23fbca05585bb464a1cee68d334bbc900da3b3518902337c8cefe13b9a6e76cc8754a01a5bb54ba90f61ada8cc0251469e7d9eb119f0191869384e3257d82ca938c7277f49a50e67f19;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h145af91cdda7d544aea86e02efbea30663955437d1582937c1b75e432e4aaf9423341798a326c61ad146420282358ed90b5032c0d9f1003c5487e8ded6d145f3a3a3c79cab97de43f6f762684e561edf32143f51ba915113f2262e0132ac025cb46d7a2662410bfc0b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd11509f275e1d22476a26729c8079457b8bbd4c56e0093bdbe2f6ab98c0a1f74b5f19b2bd6599b79425c82b1515d414a6fb97e109792623694ff6fc79e4c579f91f3d99a0ef387c30719a68c869035f4a521a01760052f694ebc79cc9d946dbaca85715beed0eb6712;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he412652079e11417913559b400670a0cf4d254a7bc5875aa1ca2c59ad84efb20061e908269c461ee50c33226856fa73efc58ed48589348a5ef56066a061531a3a6764d62cc50f48e7cb378b93650d66705588046484aea04007b0a5222a013d1636b1027f93312c801;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ad17c4ab23a0e356df94f8adf5a6ddfe8d779f45a4599a3af7c788acf07c8e41a68f0e8a02b7335799ccb45578301448180927fe27f02b4f9770aa79c1b8f1035cf435c9edc414d414a65a62406f53a398502fdfe6bc4dd16c75c3728a2edf0b985f4520a9ec14cf3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h168fffe1ba0bded6f5968c1c9020bdb1d0fae7a24a1bc0f5f08aa9ad4bf00fa354d26d1ba14a20ea6a98c394c69767edb99baad52f7353293cc0ed9547bd97ab4f1a5d79534a0bcf4e54bc395fa6152e4192f31604c069805196d84e1455fbdb0e04530588d643f9366;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdb77c5c95b5383d8744c6ee0affadc808eca6292e5e315cd5435d476cc6ed9d2ddf288f49354a921c710d1f4da69b8e14ce67acf8338d060713bebe6e46cfc7a7a3fa4368ce7e2dc5c9af93e3bc255e9f72b049c7eb8b961c34702a2f62ac99a774e875e5475ec973a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3317531147f39f8b23104155daa9076cccf3faf9032ace29c4b9e444d49648b31154f30018d42db12e3dc50f2a9fd00dc831eeab586bef5a300ba162e45fda4fdd2bcef588215c6b80e86ddf34fc71c0a25248b72a19eb740e5f8fcd594e74dd0ba214de1ccf85a3a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3760eb1982de6f832900374a56c9ecefeaeb0eb91c693350e96f8ba18eeaa81e35bd32daf1e7d9fa37718cdff01f2225d7f6cd9ec64a26ffd2cb766e7b5515626757a19dc6a9d3a0f88ee15ce84013754c98aea2917c1a5bdb28766542d440c402c18bf7cafa211c4a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13e5e0c749282c7394c0163f57e2f9995f441568bb75b2d4f11d883f6778a7ce4fc65687813643cdb6cf746745695da02ee6238bae5cbf2d0301256dc5bb4da1077ab4d1d6cd635a5d97efcf02e6b473baa038a7fe09bf0c8a8b80297af991b85b890e802951324915;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h359465dd6d1d1defc1104477820496c38fd0075b060cd6d41d0e11ecce5385cb2a3f119bfc33119dc0e2ef6c177b3f5bda34d59fe7c88c376c164e1e63720dd86d6e2ecf8dfe7e19701f853e04d46f1c798eb8f9ebfc5a233df9dfb7919601c616566c372dcbe19df8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1543fa381fdf33754e252e26adce1a8d51ce60bf25b9d9778027a2061b583c5c051933bebcd69a1794f7c1c58efe89686f71bc98973d6b2b64864f917b05aed53fdb06b940224f5d17f5efc43f179ba67c380ab5d91a32e63b9bdefe67bf5bbb6ef2358000d34a30655;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h153642d3ddf56d89ddb8f93549a26de76cef08447e5d7e898f2b1c2e8343407cad2ae6714db9288b188143684f46f01151f8623d025cc2807adc9f068cd018d9703efef63e9f3a3fa23d837a414a4ddf0c9186a37b1be35afa76934909c72b056ac986643be83fe764a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96dd637667dfecc8ed410aabac76e9b91295ea614f4850d79b241e3c4caffd1794ec58f9730b2fda12e61d69019cb7156bfa64254025a3c0a05240afee6d58c5c93d88180204cbcc84d54ecc0bbbef8d81cb7f8d3247e74847e3aad41f733ac74562ed0a68f53ce4d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he63a78149b90c430098f18c401bde15bd2f6d6df26b1c60d55b064c39eb1947bd9cf984fb22eb80379b887ee96c437701d50090cdef6992619623ff63199e203c68b7e8aa224b9ea9e7ea4c53b36d0a3ca1473ddf90a8aac31a8b5b3c1c70a1cd04799e41b4dcef563;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12eeb9f68b92d14ba9f1f84f693b4a8a5e5582e446a84583d4d55ed5555414efb68d840d4cb46a8ebcde54f2b273c06a32028f6db50d807e8f85906d3c9852b97275eccbc16ae336096e27f07df78c221e35a735a515b94871b84bee17779fb98a40f7b10e37f96b9dd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h92027d27fdf5bdf1f85f485718e780d87943e1c8fff9f86b074c72fa31488e8a90da50ac7bc4608835aad5c66227c6fd03a7a00f475a397a31af0bda7aae929d6ecc8dac0276a032c3566ad23ab14b794740f556458f9bc3029c1fbf93987863a5bad3199c58732efb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1134362b373288c3b72e8e1e7df9ffde5da66a9d64a91b12483b5cfd75be225a538a27daeecb1a472024fb4e6a9715ff2cff8fd372ef53fdc8d6210d9c3ba0c74a9064bceee07496b1b6b87d60bd56e7d0cf9e7d29b6b235e804a10885d67f8aa85bc0940cf88c1e3d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1612cf4cba1f9d3ce9b77a059632f499e94b498c38e73425ed5ae4db28548cabf173fd23dd800f154fc2ac157f29493688e8c6f447576fcadfb21c52e09fc7a79e6686d6d55bf6d32ba36c74de839ae51fb2e5016804880b8fa65c771230f9801196153c6b098e6123c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h433340f0faa5250ed8ff6c67c5f797e8a8103f65c4b64e778f04b4abbc39ffdff58dc22917638f59b72e3ef54ea33dfb087b1ac9bcc08d3334d06d13361a5e654f58a7688b1b082716699adf2775e0aa8613951ad04fa9942d628b8e8988a1938c8c424d713311e64b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11f6f652ebafcf2fe48ce37a74892b48878a9c4d2df68e99a28f6f466ba74e47d159b8bd61c3c1ed455ee475acb1a4a5f5534ba1bfbf6375558003b61a8a3d942f7759ef3071b06073933ddb25212469a3b6edc43603a0fc384afdb02db7c387e0ab8774ff5c19e5d53;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38c61c188125a7c349c72751890a811847653d0d55bef632d3a19d1136079648de14a32810a02992e794208b58269f8752141b63fecef73b22c17a94fc35b9b1c3d9fce63d1d6823a4c3cab3badc372e57da8aa20f714953d29cf0373801d46aa72a70f6ab7f37d015;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ad612daa579d7913b9b5824607f101d8b60e00ae22f081f29b546c2b663b1f69b274a5b395153865687965b884ec4d6013998f88d3cb548f009f77c3581ef20648a1fad148505b25c867c104768f24c6b7b1daf946093473340644e62d054caa9d5ab1137ee044164;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b36e16f47d66d27b6bde9dd152fd915b1c7de9b680763c6be8c20d0d2481acc9ddb742196aeac61da7cc731bb050b28e4ea21f526fc474eac267409a8c91b29062f63ed15e3bd8e556e51b3d3a65f73facba9c27562994117b20ff9e7565255f43d885a3b305787400;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bfb3ac0c0eb2b7df80d8170b64bcc7f41016de35c73609690edaf0d9307a17ab3fa5c6f9abd111854aa805b37f956e026204f2ac14d90efd85f25c37c3216c8b4e44347d7f4b9b0525700584895703ee31b69e82ec681cc0b302773e92dbbdab3f45cdbe02fa413206;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8ffc53f239368052e716b8f31b90eb59edf262a5a45489b179a6be4bd7d3cf4e0a3bb1acdae61c1763d761413b3c3abfbb0ec141562766109abbea9e46de413796c882079474c203a80f668ef6bce994cc40c0f7d9dfbceac70681f8ca4e1700303785a30d08e8b31;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5417abba1439ed9068fde6b887aaaa04c35086531d6f2ed89625d538709f0a0107e65ab20b23f61cf44afac73fc7358121238dc5ea2337d62ab098aa12db3e6b8dc7d4680519e3abc4100b8de46ca36181f6891ead37066f88227eec5d7f55ab9dca0d3e479b2f34be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d93050c9cbf74e13d4289230d0d55d50dc838346cf60f1b9c4ba83826463ffbd0137bff65e61bfb28609af2681ca3191752406673489438654d2ccca372a9c04bcb24264ebcce42163a4aa50d8c7a29f8d9b243bd8433c55913da31a414bffd81f4378fc18cbf86d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150ec04855adc9fcd21cd7c2cb941ad7c93c182f8b083e8003ffa3365c8d12474c6b04a4bb0ae2d5c2a114e0ebbbdfd9f4097b1b46be33e9a6206156849ddef684e17a725682050cc73eada8f269218c6fffa0b58741e29e48c076e0ae2d4de845cb6a07e3a3f27fa58;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a025a23eb4d826afad4102c30c63a4454193616f524a22eb2a6ef858ca54916d33943e3d5532b1e51ee4a5f90a1f8357391b2bda8f7fcb0e2f7a35b5cbf11af778aa10b1fccd1c568dc65d5b7dedda411e089c0ac77a74bcd28c1bb2f3a7d8c79fed5178a0f6281196;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b091635e38ae5500c0ed70c46b62f8b031eaea3340986532cdb5b212881f303b8ed1860d293c2b0505e1dd8dfa46a061533c7978a7069a642966f97734c4ef0b249662cbb7832a547eb05a4a082702f7a0ecc1842f121db0c3de34bf42bd19d5788db29b456a1eb527;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ddbf7eb14318138278a5a583983d5aeea4aa50dd82b66d3a9b4a18c0a5da46416f659c5799f87ca724677dcc60cae6173d0dfa62053d88d84a06e3644c7c7d8baf35b0f318d348ed4b55e659050ccaf0b338b055c4a7bd356f95e98ed32ec929e6cd79381540c8253f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1053f78eb899ea99591b56b6a5330c7ab90c8064ba468f213331e4c62874765eee985c0c41d886f9336c4c94113da8eee9c1d5c35534440547f401ac7195e18e251477d40e5a43a33766232d57365b9489f48eba5deea20ae127e3a9a16619567a585179d172e802a92;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha7983262d3ff52aaf955dfd07be0f1a980cd7783920a11870b8f431087c1c4c84a6adf9feab3db7698a1ddd4d50065027f305044c2f8a76dcb4704f75a10cb50cce4684bf3f8a574619199c92d770387336498e08bf7bc16367c54ecebbcc18263956574ff0f87c52a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c9522bed91a33483fdca824665b77abacfe9a5cf6f7be589f11b9506aaf3b5ca37bbcba1ae00d90e348c285be6776f0dbee3f638fa051f75cec2c1529f30301ccd70610a9416e13006cd15b552e77e5b1bfb09f18c11d797b6e06d75d8d696f89c697c7fb9cbf9b8bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38f7d253479613664daa4fed203fbcd36f0962a4b5d9292df50b7c5dae31c8020d9e30fa1827af14401e219acd5ed5d926f08b6fe6242ec5a07732c831fd35f5dd42d416e853b0c52bd42f8638673a2ab28bf5f5128d215178d9cf09754327d6e3566c1ca31ae58245;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2116dd25bc0f293011a35932e23be483409df8e5133657b28c25b4d8dac96a7988dfbac276624da4ec66b9b2bff4b41c546956c8452afa525cae8ca7fa0b38f866f4b465b86a0d2258dba2eee8156737dc877e2961b91bae774cc8fc624230070ecfd7567b6d78aaaf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112b153894ba556d106fb6ff40c0583290d5d7f9c4e269446fdd66b6cc27ead5a3eb223a872604bc8827c14be05ea5044086d2d5a89205fdf27ce2e7968ee441ee2d06646c1ee93cb2919188bd28d5382fc4a2f8e13a1a585812057a4879a8627dd2877f34f682db62d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10d5469d7c20c415297975a70b4dc031a8bbb566a0726d1dcfaf5cc823caccfa938d90121be539dbc91aaad70ffbfde3853da1fcc083743c6de1c3127c13e40dd8fbab0d73a16cbba91e55189e8bec47a2283cff4e5bd7b79e35eef6d8c9f456651e0f02d4e677be211;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcc6942da22d7f71f9fe94b556a0f8c024a03d734528291f6c7278a8d41854ebada3f57dcff77877070121863bd3eb292061b0adc0fa1ad6ef43d0a8e84d750329bc141f0842f94d41cba25ab232a622106b3896575a5fb5adb897f64117840e64e517184ec249c1b34;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5fedf9c32e9450d610b2664db0c426d31ccdeef08276fe3a08bbcbe80742bc17eb7beb2e49a3c8d507b6041de4e617419a848372f1aa4427e54141a20ac3542e53b24191e6dde7840bfd9da1f1d29765e1b2ed218c0792825a56dfc79e722c1368ed363b54d4db4370;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h182b5686b607dd518636312dff8c2fd6e0d09ba8eee2361e3cbd5d5081ce9062f8c52fea88f085222a0f5934fee4e88b7d779604e4edc9233202d9463b63623cf521a067e36bf5e3938bb25088d16a7e8f7a3787f099f0602e5eb31378184e6acac83be0d66c45a7d37;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b5e5a1921e9433a49cfaef1f88f6e1da80f3419ad2c5db67fc6b6dea8269d5fee1d9dc51157df5f7b362c955d6a0b015c44f9074771480d0ec64adbd9817c582e5097010dec1714c12fb9c8602420015dffa772b3fd7bb266061fbcbece637c5983a7c3c1c638ab5ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd3a985948740c011e42dddc7c7bd2ccb02cc4d0388e6dbee1036752b74273bc39bfd4731c4d4d9ac02b8bd2fd80853aec1db4b62e3b70c1f7dbeac9d2b48b200542d6591dfae10b26fc9351a586fac209bbad54710f3a54177e7066a4e037b698ad43641dfc50b753;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d4c89a4947cd6f3cee2541fcb9dc3f3d3a21c50449921ca52bfa221772b822f46bfb6b6b9e2fd931a74643ea90f7c2862b366e8a33087247d7f9342652ecbde176ca2ec9c7d395f24e99311c804868bdf32121a17b3f6788d9c1fb94f1983bc64133f88efbde7e232e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ab9ea071f526793accc8317e4aae3c6de480b680b46291660abb9d498ae42d138f195ba834b66b2906344ff8aeca50d53ac795e0532908d722c367a6d61923638fafccc9619961e9bf576a738981b4813ecc225bdd43d426107d38e1fd00bcae8227e3877ebc9a7c5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1878340361ae69971fd1f23690795e8df04a8c1c98a8e712bbaa433c7ec28b23548c23f30a61e51a34433993eab2fc46267881e46c57c4c35b01c83003e6766c36a834bd3708e5fae1d23cbc5041c323b6d32a69f27e374810c5b265ceba2e518c6a8dceedeec9e4832;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h124d8e956a70660fe9b02d750e1f986d41f27ac827dbefa89a010f63a69e239455362d944e38299b9b5e1496220d722f72cf0338527d1dfba72472fafe26ed28960dcddfc51462bd4a4f9db783bae6d79bb276d71da32b8b1b1f75d8512ecba20c48f0bd1c96a066a02;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2e09c5c4a0e823e2655606e0d6bafdf93a2439dffe60970d8627cc3ab917d753d8cb314c59bb5aff5c33547e93ccdfce0d4579074c60004691575e858c89c4ff7af50165eb245ebe7697c83a573fffab3ec1af1bd337d2d1e60ee7826a3ec8df0b07ab03d5beefa52f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3a35ff9f753ff023aa8ad14ecdbb342f6be063a83a206ef63d4f9bea304c21f93f94e5934c9d259292dcfd27814b85fe4c7c2ecb5e3a25b807163ba3f14dff76d61e46c34bd75c395f1b425e40a8239b79feba1731ee129b57651c24c5f7cd316ce984383775c68264;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbbddc3332b172f03c1eb8519f5e5f9b9acbac95bde8a559de3151d49aba73a080895b612f0b8e5823a01530b5ca61d881cedfca6a2b8a9cb98aa8b0497421b1368c760ae548568d47d3cf6f7c95e4f9f92c2d9556afe1c63eef4c1573deb7067f1e29eb891c9b0a06;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b942482d71456a027a9a92190030816f809a45ce28743ba10b0007108798f135dbfbf82190015a6138c967ec83f148e6c1210f6df3027784b3451520742eba7265b078a64890b2228d17696b9cf5052e290a63485a05192d201a6ec9cab61a2fb132150b5745f3a3b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1269b6affd55a77fe70e27f602b2dad9b6e548d697e7fc1b8e39e35c453a8de501d214a829d71bf40a6db5df29479697ca410f9ebc848407f639113351d72fc5c8a78f80848783e5b7429e37d5b3b49e24dbcdbc533074abd190a5ebced5f268a530d267c2b44b9cf1d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f03480555d87bb420136b4a290a6cccf8a06a4b272cd8e1e3084b0ece44756fc5a24f136d7ab8adf73dda581321257675fec57c977d6681e619b078cb9cf89c9a06d8b226e5499fd37a8168566de42227f39f7be5c71764ab42804cb2dfe1f3e15af5696949cdeb56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1809746b835a25f7910ee6e27dc49207c3439c6ca324d856f68a3e59940a9aa0dc4d977575d37029ab0544ed3016c1292c8237a10c3775928b976a0e967253a5d27ab5c14bbbbc60d13f73fe9efefb86c81f1c8aa9ec505dbc9405e8983182d3f6d7c286fe895971780;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfc59af5d5f9e0958b15e2d41622be916608ced7a3606cd6d87653b193296f95564101caeb07c2f5896464b29cee0b2eca3bc6f14f1c2e96afab429f20bfe3a3972d90b5ece55e769edbec5a46baddf64d6a067c99d70d4f77978bd4bfd681139d91123a1a3d6a3ec7d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14b0cd95987c5f901fecd919952a7ff51c089e55ee79c820811ba257e4852ba132120fc5635751c61612d3bd1465a5003f66f757735a81e20649812951012c24510ef9937d1d1c78de559e7374fbb7640f40906f96fb816c074b6e6eb8d75697e1f221e6ce56466bd0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12fa0385dc085150e6452af3963a36682bd4e65395bf0a788abcff63340bce9092c0f2894741f6647d0dac61ce50c4aecf7b72601c1da6dde74a645959741e4bddefb2881d006e982e7d38b1dfbf192efd839adef038f4f4f7a3c10fd3a9e0d17f90201ffb25e286dba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e69aadee35b6c4012c7d0d920093ec7df7da8a6d7a14210a12a1d0a06c7359269b07c4527fbf11b4be3dc23a66d65692b40d24eccb63ec32992bf1c4bd1c9a8115fd74482ff69a4134b79fbac9e84b8e0adc43d36371a33ca4a7162496f0b2780d1c65e7e8db1cd9d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h168b0148d9a19647a73a5e5953c51caf2945e66becf26cf0d3529f6fa2028b79151e59e57727a0de03320b5eb8343b506311c265db7bcd73c1d774131bb92fd0d0c341f59d3857d6ca875f51bcd0b470582b300479db0745c423fb9bf15a5893ff37992e4bc47fe34e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19ba53d5070749a724f1b5cbbdde9249d14189c576dc180aecddf11eeec9f2c6b08f7f9b342c68c7d941a85235d007773723c42b9580572cf902bdb1b75ccbff90cc647023b57bb0411f12a9c564bb620dcc30f2b46e95e3a9de7211ad97b473cc0881933a466b95922;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d931d3ae04bef4658477384d695ec048d0794299b5bfb27a0359eb3de17b250453bf737aa88a46888b748f2b2d8c1f89f3a19a3f8e8240cd6b29723f558e15ff244cc4f2e41629bd1a0d63fad411e7a56708689cd7e9ad23206e2716d4a6e5a2fe78ed78b4140ddacf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb4ad15ab18c2831653944388eed92ef2089a2d92622c9cab740b5c063d782e93f482c3cdad14f57286149261e8829cf5d4c1fbfb5dcf2eafb1bc40cc1378d594a60467e2cd044e184f8ca823fd2a0c2ebb58f67d4838402b8328b5289ef5dd7863b7cc1ae859ea1cd6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbb1d6c47056b8af27d97439aca90b28f61cf7caeab1f7749166995873cbc4ec127c4a322f642fabb95d410d048e2d2d69e1ae4e6598b67836b96a8fc50ccc3db2c6312e462941b1c3452236d6b87ecea589434f2d5de2ec3eaf1aba77f92e1aa55d04b7ebede25d0d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d313572f0a4aca8c71283cedff74def8cc3c96f6ba2e4f0383f84fe295fb6cba009308386627d9f3f7d2b83332cb5d4d42c85215e0018d4f57079c9b27f2b5ed2e4d9c87ed1f8f95750520dc587e0d881138bdbf5e0b19213d5c0d679c93823b2724f313aa0cf7386b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h64460f882828167e27e3d1df2a41c2f0cac29dd3b2c9560dbdda56627059488fe4f46078b978fc7928ac4f4d2e732338e1fe038b4c7f163e536c491c56e1b568abfdee7328ebed204d4af4e5456b0ef113dc884ef5e440b2c358d3691f34ca6fcca74d6686e2aa5572;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h858382dda00716928ba0470cc51c6ab9b108bd8f848b741d00671373554e3ad844c45333f7b2f3e95e02e1f40e12c691dfea472e107e6d662c4195dd3868bc9069f8af56c9e108c0f224156a25dfaf2377ef23e61607f1697246efff77387775ee6d2f7f474b030ea4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc04eecc61fea6c39fee78abf2530324544f569c7535193066ff5e7d00ef031c3874490b5ad2398132439b0074f6908e2af3fa6ffc2edc61802c01b02e1bfc08534ab1d33e647a68bf56c8848cb1a89981ebf679a4d1ba7b14206b5b3857cdfd1dae7e9a0a840e6086c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6959aaa9a8e2e88bb7a6a69587dfe8fe356a05f3d66769db81e313a1c1815259f49fc230b909b44ae835acffb2984074448f36f4b9a6934461abcd07207ce75ac32f37fd9e5db060c97540881b02b8984d1bb1030647a70a7dfdc151af41a6e73505895bd5e96fef74;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b5ba1df1ca0b7625f02661641115d88d3f07bad919eb4ca082a04d0504e518af066b6047da826a0a8a5c11dcabdb9524035c7109f96d585b36f8e92c52b668e22606e3c89f29cf9a995ddac542351cd4ba543b7970c62face57ead080d57311ca126bec15ae9aaafb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had4b60cb860a54c58ef6e82cb1334f1c8de1196cdd9c2063145cd20627281c9e8166bf29de5f6ca948296bbea2a69c8386961da82289bc98529f96fc32c6eeed9f837b170795af5a58a4c573265221f42d67e75436a05ae9ade0a96db51a4143028648e27b5624f201;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf03d4cb73445f7f7e57915dc5baf054feb365b894489a87cad368bcdf08bd26a14d0b0f0d1fc72b5f4c0020c57fe15f4819b0c808eec608ff4e30393ba5a7a73ce12e67f09d18abdad5f5993d44f14768e18910ab03e2c07a61b81762dc426fbe3b8be2833389172d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he4cb31b243e0dd7d307599a44beca6e33a0aabcb4b477a10df7cd61b4d6e88d1ad98601001823a3718a877cfd5b8e7a0aabfaeca8a02cc14c7223c1b19e43d4b45cc41ae3b66e55a9aafb5f30c2db6be40ade5229e800d53222d7f81e6973c44a206c59ccef4798407;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h782ab6d7a0bcaf2d2e2e4adfe9f999b2f51544fb8b1e82b8583b11778bf63e20013c436e2baecbfaedb1adb69cfa5a877feb58aff328f66a9a265ad6ce331e792d08896e218d2b49da7bdb0638d3c08dbbd01d9ed8ae1d7d431f300b5cb28c5a182f359e42d8a9ee1b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141e9d8396ef82fa44dcdcb5140c223080e26b0b7a21d29edae67c59a789f4c8ca4122e173b27fe540877eabc340704434fe33b0d196c473217df24327e23e5567cc79b9b8fbdea826b54cd34ae97336f4323337c02860dd11bc6a1d7e0138b845d3d6d47d37c47043d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c1e7b88211ad880212ca4051e5782424596447d67a5336a138a19eed6c268049e85a483e296618755610405179932242e02219669918466fc5b41449c82e287911c0fd5aa7f1708d30aaf21303dd656dfbcb81096612ad80f7577eecc2056b1b2551ba11ec9c580541;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b6f2a6cccd4a3e54488fe0aed1bb7927c370d68e3d32d9896d865c50adab072e2f30b1460458ffd23120b447e7b25cfb34f1b3128f148e503f8b061fa7c58dd27e8b1c4de30f9402b6e93bbe1b853db568640ab0578b1a5a8f0156c61dd442530f118c2658be46d8e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h164f7df5eaf1d74690ce1f5b49c61fb472e216d673b87e4ce1e539c59251f8a1725f53e37830b8452b42e89339c9776169e2950018fb13711c3d0a05395fd7a70b1d520fddb759a13e364f569ac8d46570ef504345301418cf5171a50dd5dcc91a770a6929c970a7f9f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf8c1a9f48b5e167e8fcab35a2964aaae20e9e08286f4f76346cb75201505f676ab0f99d7372fa5103a500adab5fc40795aa531ae187c491b30f4e1e1b4d134502c79c0c481adae28865de67f60a4f7b487eb70c61a530aa7c53a2f706723cd5791103d810040870151;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h455c5e88f48b6ab496317075ffb4d1f77fd4f04043f986c773352e6d037dc70d0522b10e68cb4b3bfb60a01ce173972b535eb7d60cd38ac6f3c14b526f6883e31abecce5f834dbc618b866f2a6893f8b0aab3534b2f4c276f36d044663a4fb85554f4f91182efc9c86;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a3127351e1e01c23c317ebd18d31d6e4fe57b75b32cc80dd9dbbe5544e934550cfd9ffcf745ea8579cb73c633cc93bc6eda5c28d46531be880c2aedd7be91b09daca781d65b3cd6c8c556a3da86711553d51567e5c88bfebb0baf2316b9afb9514ce82710b969c0ae8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h725af91a9199721f8c165c6457cb7ebfb99af1c532cb236fe9be775bf058f3fef454d2d7b66b1431894ccebda8fb8e6f3234775393534e1192aac94626a2a69b4a32ad85d7525c20165682462a7210c9bb4e486aee929d16b715b281d1ef60df910fcba28f05f0ea13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1162c9e27f979497481556c675741980834e65a016c5784dc02f5d4b150b5b159f866e7befa6b68e3bd790d6e457de9f93f0bc449ba1e27c547b62c7f48dbc2508be2c8d0bd6efb3d29a8f23e7ba6bd1b8aebc42c7bc6120e69b332677b48684c8d53091494f5bda79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e7de1357c72373c9aba2e8025f39e087d0730e408d6ecabfb4470686a42ec13059e2742c3de78f59af81e129fab949d7b07c8d8c75eac9be385c6f9654e20326ed005bc9d0804ef7764165ebbc5b825052a4993bf9eff5a562f139471d5cc2fcbc6669fdc60807b8fc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63d960e56113657fed007304e4327b85496f3a165d5e1814f4559ea177b65a59142ce989941a9b691285eadd961a2538dd4f03e3df38713f36e7b62a4555bb984e87eff7718bb38c4a08b293ee4a841194a671966064fb3b363bfcf565a9abffd36f9f4a540d53c783;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h180ef867dd6540179dec05b54273df14698f724e4eb5290dd48999aa983935ab2b485a63008aff5175fbab8bd05a158e5f43fd977730d6a1b7834dd2655816619d33901b0dacb9742368de987ea3140d28241c1ac133c8e6a8e37ac0b95c3524f25b2b2325ebd0196d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h32894802e2adb411ba4b0621350ca631d488fd89fe9ca46676353e0268e48f063bad6a54d591e594733c31e593d92d430a5d2815671cec7864ec1b74515e34c856a53bf1dd19156b3bcfeebf7173dec7934664e529284fcb14a3798ce617874710f0870ca7eaebb4a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15113faa6a0b2d79f4336606f7a3f79c1f2c6d8cf4dc49c719b40208c2aede28ee5591f5f4c0ef96d030f2ae9874fe7e0f4236080decb7ae7490992bbea5558c5c8b9cf69bbf42881f2f37af76b663aca00de82d61142fc4f08e1cd5bb7db0599b5f97c920d6940a77c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eba1ca9bfcb3c645581ceaf49a8d2b5b35b0e92804b64bb8c177fa2ef5619858a5f9f5de0c98adab637a36f556f613d843486c2dd5600b517a92b11a89ef8b4c206a7cd93c553dc23a3cf736f181bbea3e90165caae039cea7545466e6ea4ce292a10e926ee34d4ace;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h73c18f0fa69c97a1793c560fad9091909ed29dcc268d7618f92618b2d0b9957805b67acfed6dea51209b093fe7f52bb14cc18d88772b8c8fc6bce2b7e41560735926570778a2081bb6007643a0c109b0e459c8260753f26bed961803025aee36b5c2fe6d1a8ac8643a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b16788b42ce14052f0cb8e03c22a4049a4fd16d7b14d6b318edc02e539ff79db9ceeebfbad2853649bde3b4871babcd5c8c50f39fd0f3453de9e11fb1723a9507e9315e58ef79619a97e9602168f65fbd05a07e27f37ce3fc259f6e16d15a50c5cd1d966883cfa657;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he4b51700783c037cae3bde34d0f833a9b116f483426eeb45d1d10cbcdd112a07dcc3a6a7b1e6e1b168383a009442ad8c289e68f6707f3acdabbe1127681f76604e18914fd52bda3fcee95d9ce34f0dee2c8a2b124ffb5709e0277d99ab358d2a15f92465fd7d0fce7b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f6092f33be2e2abbddc0328bc5a9ad6ac45aa73f409db93cbfdc31a32eea2fbc32170e5b9f2c3840192a3dbf075c1563670e01a907ad07594a5ba628217a137dca0c18645d79edda996a0ce2cb40923302d86c4e96bf209845d4d8df1a662d78ae8f6b5dfaaf15759d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18551bc2a929dc2038a48a91bbfcd79b7c2922cda15cffe744e915c22a02608e2eae4517f78fbe2f8ae4b1af6339ba2dba7f7121db5c80498e6d4a4d63948c7f4787def31dddbc9e8c928989f31d783e9f59de20bbd9f64a96fc9720203bbce1b40aaaa4c96f7832e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc75cbb0b634969b6540e4815757d2995d435bf347dd6593b4490f33774eee853fa87818a906fe5962783e77508a37e75445083725b7cba9386809dedbe4b7fe8c19253e6e159b6ff4467e8d94f0b8ec21fe6039b2aabdba00746a983691588356541aa2772420214e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1befaabe2c98734ef140b0b40e06e02d5bc44c4f5d41af55e61d57b41a70743368b24aca74998506a79cc185fbdf142dec4475170a1d9b76ce8f5e9a0b5c8462564a4463bc1feeedb074f83914ca0e6b902d48504b0224efcda5990aeb985f342062d1ca889f439e818;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e70b918a5fff91cfa85eeb28ff99ead634b6ddde18f025a0b6f64dc94bf815254fd76a277c6f203f770b51a403fb2722bafb277a7a7a738f06d58ccf32cec6f4a9d3d1ca6b8ac4e60e63059b1b74e3a5b34e8919c079bd99f909322cd9865c8f16fc91e6d2a551db1a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee3c1caecb93e5c55cd9f4bacb8ea61a3db61b60b7e85b94f8a8c6a45bd45420487d3d6bb703234f9462926ebb424d00e6fb023375fc4dd8311c2efafe65c84579750a5d7c8da3d27b2aacb900561f34a4fc29bd896a6e824a3befb0674fea8a7ce90e03bec7d125d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142d17b30aac1f40dbe87e2926278d3d5c7da5d3870851ef08b298ebdaa69b9f9d1d95be002c4dfff86c21f787b6e7b631f89fe0a5044823570ba93bb14f6745923f18d4c2ebc4a226d09cfe6db5586c3e11058cbc0a96e8772c065d980ea4e25eef854065821f77217;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf52a2e5ee18b0caaae4b88fdf7da612316109a6de0b7b0255ec6fb1cd2baa35403dab8b2342f5131b8ab08e5b0eb5e52562f9206a4bc4b55c56445ce9ce82343f29b31d9b9419fe726a757add42dd6cd27aaed2db06fcdb47b45c5abb70aeb9b9a060d06c085261174;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8f29f4ae6e542f1d8d0b3c3714b256cfb48acda68762271641fdc4b5e1244be147fbe9e8d568c56eff04f8a117b54eeff1acfb3ac0e78b532af91df8451774574566ac8183d18101293b6d9201de29e40562a58daf9037d29b3183d078b57dcbae361e92424d6a0f62;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b04ee7ff2c45169e05492a6aa0ece8691234dbb91ebb3c6dda370fa607641ffd941fe95d82e41de299767971a4628d4e9b84add39c32b5f0f07e98e56c7a49e4cad4225ae7fcf6650e9730a58ddfefa2202447f419c9c913e360dccbf83f48a22ba59fa4585de11da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d9875561911c545087ba3a910b84ebc8aeea16ed11fbe2f2e4c0862667eaaa9a07c5652542862e1605e6dd4599e26ec2dc84d37e8045028f73badddfadcb60ee9a2a6922a51d2c9ad4c0053c176b5fc3e45ea69b0ded70f12dbe7f3c85d7c81991845154ae518a4cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h73023cbc48105c068f76a7bd4c12a59525a3df06d3a1c95ea9d0a10d10c4b938b0313805bb28c4ca8d730d537b6a5febe12f6dd4f11bab310d01f71102da831c61f6abaf9cbb633b47b138824463354feb1f7c591883f370d3a4adec97ffdff0402179679bde3d98e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h245119a16ca1723fb54fe2e57896764331fc84b1cda44652754e33b491a407743ea490ea69bfa252608ddbb1a7df0e335c41164a2efc5b60a371397c80be61047e235d30fc7eb2d044aa15137cdd6c24fd84b7de6f1345a6f0b0f33cd4a2d0173bb4fc3bf815d49300;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h99d2f5bda6e006b3df81ebd15b23659de855fa0d4b5dc65906c8e8dad7a1a689496535fcd2656e0598dbb189115e6628640bd026a20cdda6341ec71a7d8e6debe32aa8669715cd4d34eb4068fc21f428b09ec413f519031454ed4fac6df4b7392cbf7cd2c6476b9f98;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haedd422d1f7c5ca77e43e563cc7270d67ffd0caf4a853f767b3f06d5efd83eea9e0db8bf6cd9f701ca70ebeb66435f80430f1cca52bec6505300b58e31dce71c42348de0248184f01ffe85edb23af001b4b2c53961433014e50adc98cb4ea007663ca4d9ccdc4df6a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0dbab83403b9e6488c48c91cc446dd94046cc035a60927c435eaae3e0d51dfaf86d945e8d7f37d98d4009bd21db2609e7e286a53db0b3f8dc1cf3a3eee674a03cd0dc7488094f8c96e95931c78bfb59934bc3f96e14654f012a0f04635073b06ced45d72fd9146acf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h22a8dce952ebdd8053b2dd7e42e9fc3c11f7071aca933b38c522c39ba98c2f7cd499b4163a66fe8cf0d05fcc829e345931f917760f1abce8e7d4507f1b9291f52eaf5d5448f0d85428212c62d99f4997f2a1291709021e7760d6535d8b1c4d78b73174608137d0dfc8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha64b3b84a296f1bebdc3392bb6b40d7ce80ffbb8f39cdda467796ecce453f48cee3711c2ddfce85f345aaec9457db0f119a600b2a660c293d39cfc941568fb22085bd69ec007f5324958843c2903f12c34fadc2c3cfdf47c6d5473472fe866c82d52dec134196cc4b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h70e32693f6fc874a5a616e02e7957fbd95f1c5d966dd52d23f28c8fa9f5478d89203821c0a4180b749bb578465123932bf3648503407e425d929f231410ddf73cde3bcd1d010bd5374957a9c879079c22d345bd26010ea1d4d59e76fefcee0af76c38f3568c7d9fbc4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e5b1e9f2827442a0598cc7cc915edba9c9bb015321cdc030eee8116be0316e54d349067be7020374dd6ca6d5f07b68a686445dabba5863d6f1922feb4d1b0ad24657b1d75761c4ba003d49c9bab8112528d547618de09fb4cda0e9ae6ac72d52828f8688acf6ee17d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1979cdefbb811b6b407c8439e56ca3ca0dfa06ffb879337965e41d39004e1a5ba3260a97bdd394add32d429e8487f5c8bd0cb36ad58b75e48c040d2ee1db934d5c6ea6ced263ed4cd5052fbb2c67f15e42778a544368d810facb4dfb2f9aa31ffbdee04a7b20fcf5e0b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hacf566be805f3ab8ef0ba875216eaaa8b3f4212d2dc3012e5ce868ff34b7a367fc8d23ea0d34b879e585f70226c60a764949d577ceb4649ac4f2a35444caa8a29802217df1e1c6c4b13599d1e044d3567ac90e02253c6884d72453738843f85a91a60c03b99d375e77;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1890a42a2c8d083b6d60c1692b5345d0959ea98b691b6cbb1a4f968cf393e8fae4c1cb553b175bb4634c27486f22114df1207981053c940ea9f1787565239dea5c500abeceba5983bc524e6d0cf96bd284345ef0935e4061f7bfbd06606be1c7244b85c8605ad398cb4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h210bbac80720612af0eea0f8f435c513de8f1f96f1a504b07f8df202a48dc6cc256c6781547cd7473bd44ab28cc1a3fa0997481e1ad366f27607e8a3510c6527cf891eb9582889cb502de6c86976ff10e67d9a74a9feb5a0255cbe1aef92aec7621d7c5def16458d9c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h201e3311876a368cc0be5c0e0b7b625242e377371c803f6a1b17aa3b055e03f25b7880c4f51b02127ecd569d709d2b24f7d06879969aa8541487c3b29bcf60f45ac19297968cedd6111d93708be72e3ce11325a74b0aadc538441fcb8ccb7ababe1610a2c29e8a5f8e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19740f9a03b2b41caae22a5a1ccc09e6c3dfec1f08b39176a79778224af4c080a08ea17117619a66f0df14a72af89635efb20ad50462aeb14d697e7bfdb37494f75aa8d0ef9bcf4f5a1801932faa9bd8813d4fafbd61c68c24eb0c9aaa3559c3315bd6b1a34188d1155;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h102c1374438e8f13c86e4e36711116be192e6557acc7522255719e05a99120d8cc8f56d21942c3d886495d30866ac925d9428fbbbb1311bb282c050a2acbad70e3be9d5ac59d6fdfacdc1963dc6f830744561e8b82b38024e9b45e01bbca67415f3a7a4d3837fb72c89;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3435d45d11c06796aa667e412d95dcba03f18d1ea9fd999be4c3621ea177c86cdcf9af8afbdef3b3f37e7f4b5c27001b435881750a9be88dc514b86385f228b3f4a44a26c6369070a38114be72c8ef5ee51de0abcc16efec0584b2241af04a87e83eb0d48ea61a7532;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h572be30975a5fa457a0961679ae08d8d0a4d39092294bd76afd0b1ad471967dcfdb3e25af3a7d5dcf17900ccf9eecef17907fe4b7b9d66b37f891c12fe465de1cb126e706d1a2ce2020544549286e9bc719926684b02d7f158250ca0eb7fe57d04d7a4978faeaf55ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba85ac25cf02496cbb7d8dadaa4369f953fc1c8b21388e7ba5eacdbdd2db059ee642fa179e72e56338028d46b233bf17e0cb4ca92423aae9472cee98c89599d30769a62bc162b7f22b48c208bc12f98853774be1d9bde83f5bf9656cd5a54e324dc29693fbe68d62b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e25df305e43efb2c06e6efef98c42520f4e8ad7f1e86efc471455d0ab5c35e7f7895d3e4785dfc7a4cd9b00ba4e6d4e803c02254ce8c5651d93b3bee0ec26cf49c5e301ced79882d35cb11b49e38e9b19942a21aee27068b8efe2ff5ec6626f81845c1ec8355c4f303;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4c46e89bfc3b24bb9850365445538a83d87bfaa7acc0e3716259154cb7abda25edc2add8daa9c32ede1d412c5c0541a88bba8a3b91537b9338b4e513d326b3a57a6a261ef2219c419c09a7636088928f3e0f4cab44eb625b602d8fa7c14869462de897d8feccafc9d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h52165e1254badb50c718df9eff4d172f389a02abc2baa297e2a1e51fa9ca180442ce8880e1e5d58b7a67c43886e51381edf680d040f7339aaa976eecb0d5f92ab71c09a6ce0052c533976363dce26006b1a5b8a2d3b3854b46c688decaee4293cdeb18b9969288f66f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2140d137568ff8920da39f43e996d001160d5269da3519a805b36e8068ea659508a7b58377617fb4bda130e601b111ec37ac3611617024f79e5d9d9d1687579231ee0b38057a4607ee372ba39b212798d0ea0c528f433a4403fc8ac5b86f2f10008cb247bd572aec5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150fa7e2f817c0ba7f397616a1f9e08c45be4d5c66159f86d1bc5c5d7efa9d6e260e8dff557d1e6df12ef860a1eb3b6d71a9e3a1a44bb326e1a7e5fbfb3520129135dbe2356ee81e5af5c767dbd01363cfd3d557e54bb8f2a66044459aac9fb82f983bb0f1ae9512a52;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108e73b7072ac7efb4683a7207e14682c227f208fcedf62b14e23e6a98029c20469b387387e31670b5dc3fb3379b6107180dcfb2a7d8451e620426ac7c9768cb01387771d34b49c3d05839cfc8a607057bb0d49b1074cea9bdd8677240fdf04dd39057a663e534be61a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h405011fd92c43b0846a539082cad5b007a36a16ee7f1660156e74c164399e688f84751262addd03ad687d2fd228533ff42aecd1e164065da402c22a3f8141d089f8075f3ec48be93a827e30c977fd02c348213687633491ef0a1ad4f32d54f79a354a26913866d382f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9603e0793fcfd75a70caf16e2cb967510f42bd78fba3892406ab05f221635f6a3b3234e56d8b9d5d1095ededaab173591e27806a2989299b5cf66217309da696f69dc1aadc75773f457ae0d9b179bcadab4f29afb524fcca80d9e676c246fbc088b429966de0d4028;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa84a5af108bf2c8b2222b9ffcd448e075b1a8c2079163b64ce1494b3ef895a61343b987454465ac861b0790cbbaeab797f7ea3c08904308a503d3eac2dc2f56f36d4525caf629b1400b4d0bb81cb3ee5fce01f45c9588685e1bf702632f0115ea14cb1a390c325e05;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdb7a7c1086e7c6a6561d7f15873024e295a74eb253410bd84ec749be570765b188555f88f9ab3b5a8a8fc9e75b4b69f92af838b1aa94e0f39f8d17c6d2add0fe551ac426da2bcb92e7e8cba4a1cafecd00877c5dcb91f7d72f130c0f305ae96df79772efd1e7a12dff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a71eb00158e2471b112658fbfbdc39b09143fbce222daca5cda87ace321a763cd004c56cf5429dd545c82d409c468c099cded6b97cb2676959ab738e2c3dc534252293e1e252c7e65a4d9fe86bdf2b8c06c13641dd49933cf89f6418879bfa3e9f3d3232a598261b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5d90ce19a48e3601a63ccedd2c6a487838f36e30b87071ff72b48a38571e2b4fdbdb2e828cde308035028595bd225e5f1d9f92dbe17c6a26e2ad56b8af19b552c77c3b80aac3926ecd8b660f2b763e83c529d47a3e5ce5c2f1805e086607d8cb0d8cf116a2d31f2caa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6499f2ed0b67d003b03b964a6213f06fe2ad7eed1b097830916d10c1106f00564326c8cebbdb5ef87392e0b35edb54092ed1817f412d855b033f35861cbfe6e432bc73c98f7d8a8acc057f1f1a877a467b5ab8746d9f50d315ad1e6ae668b2d546f05d256a13e365a7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc1d733d774be67cac6706285d11e850736080fd6e075edfb0ee8e0ae36e2da2b635603ccfda0c499dfa656916e5a7c287ed4e40c7aab27c573f40fb8a70c497f75fc3de1e63e0d8ce7666784c8e8b1c533ec22a2f0cf29a9a294f44573f22941cdd5bf5ec4dca1512;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h72d8f747195bb4be9af5be3891530ab2804707bbe5c674f7b05d88abd5c8115c29f035e9b1a6c44489b37ceb1397426f43e94a56c0a3b15cd0a4e85769ab9c19438261ab2c5bc23bfa69cadc8f9c55aeaeffbd2f53f112298b17de9336a08384e642ab406e964e6516;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122c3eedbb10d185ec23085f32ffb8f805f6d4ffa21bb4d9fffcf60cd6bf8296cae2fdf8e3d36f4605071b707ec2f39dc82b422b49b124f63b962df3e9f058ef473fdb8c94f7d03ddee0b0bcfd9e0981f1af3d7c9295f7a82f94bc09cec9528b8999191dacf763c3f4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h178d9eff961ecaa34ee63dd6d53511e832fcfa6046895c2b9e817125f6c0528b23cf5c537a69814056e34c35cae55b9defcd450da848d27248a9b01ef842cf50786ddb464bf9e7e373afae534159df7c11b6c3622c02cee76bb4223399650654081c46856f31c71b8a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af417cdf47dd700352da480b2d8d843bf9cadb2dee3a81731152e4b63c7a67cfafa1deb486cd39d9b95c2229ef8f54cec72b52b97b47f37be01457c3a42e24d60587964cb84cad136db39ff1117e56162fc04f3314edd2ac6f32348334160075d9ed1a39dd2454921b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ecb02f494e056cfc5421a2c734afda579a115f71873ba2da8a3305ea9497bd1a267ab0367dc5c85de19727ae40453739890addd3122221d1ae72d28269be23bc131c233ea2c0f47507c27bbda879407673065b29fa9bf0b68d62f76e5d99ce74b4961f2692b34f6e64;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13a8f3e0d035956a2e585a4c99e9b0b77dd6e35697da12a09b193018a610accf1a3ada2b0fd4f3ffbe318b158ff06e1a2743d26203ea1b46c866387bfcc6486e1f3b1f00fb99734dbc2652f91d16deec9041444008a36776cc6e81fecfebefc658046b88cd95420f69d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67002a7870f415209a3ccf029882cf8a6da0cf5909a24958f25aaf0c8b3c34d01d9744cdfc7ca614ddc45ae189f2aeb573aebb8658bc5532c8b099359c9ff9bb5cb6afd5d3cef90597fe42e7a01a3d6e3a9602f559a1162900edcae1f25c2e86cea4066bb8639bdb7a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b9b7dc85a3cb8ac0114a976d2357aad4da95056ae4934e336f2b61a1d141411718d2f51724e9732c1a8eda61ca9af48d09fb68d708f8951f822c3c4c39c153f2b16cf9438850a3b984f904960c893fdccf180a6418eeb218d04c378e2d79ada0479aafba6368410498;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13c4b5f42a9384feff28a51b001dcfec1c1ea8b61ac551894733b4e7c8b369b79729235126aac6274aea4dd90fe92821cc3ff5ef8855fd217bfbf6e9c2066ed1d86ae4c2f00b00211dbaa7c64314286ffa9c2d98b47662a9cbd6697d2024c32daf8e2cefbf0d8b76c82;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eef6a876bb4b012300842e6fa64918bfe9d0c8d61881e2716f192d3481d46c746505a1bee0836d6cbd6756523b050987ce31d7f9499bf22c21cf592e0a4f8d83b5ae13c797661503d5e5b10e1d8674fd9df7f6e275c4f8efa78aa465f7e1d1ae192f47558d5f860b13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1083e6eab4c0788363ba52aa0937e7fd8b7631d83b46653fcecdaf76de9ce8f9a735a3ea231e6a8fc8e9cb2f76219f947b0db4edaf33253a6528364d224fc95a4d54993dac08f73e35b94511bd7b157d8df4ae767124e61be31f189c18571fc48ec263c00aacfadd9ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba2b34283107c9f0e21236ffe7e854ee8f5aab8add986c1170a3a3a08bea5b9a68e989a1e3be458751f11dd1c416b6708d9176d81eac63f4ece59ccf8b9449a2e43ae9d82818bd3735d883899d2c2b3ecfa9cc60272dee0bfd5fbf6f966d3e4198558ca7e748016d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4caf5d28e4329cef31fda43de9dfe7f375d79cbfa236d0e4dc58e133d695c2227bb8ebeff40b1ae4ab5c2db9f4969a8f3b9dee22b3f40940e047f4474bd2e42669f633f715f8693574f6d4b2581bfa5c3a72f3cb844047589be3c6ef0cb8c63f58b1f78df8681834d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf40fa960ae733a8c687aecc69dfd6bb301e6dc22d450eee3cb5c33d2b51b19d3c5ae1e52de6ef390ad99189340ba61a7ab0f1c8326e56897ad4e902ee3fba76e70e6c4c908f0ef0a620dc8e48fa263c7464b86a9c775cdfb326660fc74c71299f9896ea4e41afaae61;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h823624b0635bd6dfa7f567eb486af1866b891ec823af25a4e5c103475ae3ad2612cad927a3207cfa406a4f4632d7ef1bb1bf49b33d4f4ce7c21c600d593df367a1032e16cfa0e8b99d55be67e8eb5eed8e60a3ef513e9cd441b88743419192a62a6804789bfe8d67;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123ed9b0242e8388277e0774c977b24ab4da048fbcac1763605f59154a96edb7fc141c8da5f6fa0593eaa1037e1d7dc41cee1779afb7d2b0cd9cb9c6930f73da3382f9e53e81c96486ca629450005fd4ebf8e1f166b52393f01b16bb26e9c650aced20c8603a468ee6f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13536f97cd45e4325c5e6030f0ca08db595978120b19701f51aec78a6b20f71ea7a8b3f00f9cf5d84aac7e6f4bc4829be49c99fe337fb840e5a2f788eeda310aee14212f069d782611ac8000ded0d2974ddb3a07b9396cd458b73ba06b335599cbc6cbad30bf09a6fe3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d492ca128cbb1caa57d27f1b8e23eaed661be0f38866a52ebfc8f17f580bf124cd1af7d86c021c3cd14233009d56462758668e8c86dd63ce4f5c30844ba262a759a55b6dd96d67b37aa5ac8559cf2ccfd011f54d7524b24dfff881f817083172c25270c51421355e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d877a47fbfb7b0c91afda02e8742dbe0fc7652cbe852a90a866d9cc7828ae465aec64efec2b3614b4fb247e7d200bfc1dc1d6b76ed9a83dd1d00e46689ee40df0aa99a9b67bc906d0a3c196b7a2b5af9919be534eceda96c6a1eb836c2acb2e043fb486e8dfd27ac5c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e595b6f6a7e441e5d4420bd1fb6b6cdf45a53cab1b41bb3b52f5e44505591be49ba8204051f193a132972646493af18bbaf227b79dc61558de992d873db8bc554cb4026dc165ee88273da1ff73259dd9e2baf5c635e63c41d3cb56ce543fc83545f2e607ce5017bc9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc6ede55d878d2919952df0a68c3e5fd5e1b8afa7b392ac4214aa5ce98f51b4897ef965c800d8473003a87dc8cc9b122eab56ff623844c8b55aecebd1307b34695629fba76bdafdbdaec109cde186315b9b6c0436e5f5cc08f56639f3cf52e7f44c33568adef225193;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdb4254da7422b674b75e9fff399fd2677f72a6c5f0ce26bd0647c26302f3ca52c8e8dc101c271b21b3ef89b000fda1847229ed6723f59f0ac7354aa0b3e1a27cd95fd289cf1995f389aeb0795ccd4302dabf8c3831119b3fbcf73bdd2a43f7cd81f2e7a0df07acac6e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17e27a07ffeaf524ba52279613a8df22f96438d93b26ba325f3abfc0fd46a94a7761dec2de69e1b191286a85591e329018164faaeaf0a292702f84a9d72b0aff4e493009e749b419a9eced30e45bbbd83595aaaf19e69db9d84eff100d98929d3c3a2f4683effe3ef74;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hadf6bc48ba2dbbf7b2f7e73787b335bd954c3efaeae1e4c5a0dd268b141648d6c9388e0681e4192ac8c1dabf1e2790c9fb75353021fa5acafab8c3e53ee05397ba414eac95f118a681c276166b5e88ba08bc85b7785b8baa1bc22cd1a13945a2ec25fceecb29498601;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb904885e77baf8dd93f894c65b907b5a86c5bf9269670183ee7ed506d1e6e8d6d632fb696adc557a8afc65fdef8ebcad9fe7422a4e46607ed8199e3550926eea846e3f66174c5ead9f47cfb1121083c8c6dc912a90d98e2735309fc4fa7b64c35286b699934d3b8feb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28c9b2debd5fadcc23f6cbf683ec96f35e6641a882280101e8d88f7e923371b3b5b8d844f8884859ada09b59e0274f11cfd2aa4f04bb8b17e094f5926fc3e786404c1bbccb96a09322f7750540f0f6530f37427cdb877b4490ce965df0138dd18e44166edb12434d3f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15959b16d2d98285e2a103ea4128129cc1e5e1a0c1026e5b8f11b11f5554946e613111f170d69474dfdf5cf0beacf8a7a406dc5453f18bdc2da2652e2059ef30f827e7cde92f7cc49c000f9bd690fd7e62af49dceca57835d66bcf0ac05e485969f21580110b6b6f9d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d523bb0fd425ce14c72bbc8445dbfbd066de174ea1ee18f58a24ba9d9f0cda966525a38b57ee966b4e8399973d4c21aaecf3d2cfae59cdbcc79276f97c84f0548ebbb8525f2bbbbcb900204dfea8744dd8d589d01b122c620d05f5bb8342f076320146d2a85508dea3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13e155979d64c0c1dd9d15019342a963d16d60ba1f2c77324ec4043cffdfaab133bcea32442cd960ee86a4ccc7e45ea33ce962dc65fc7f9bcf99580499306e097b92d554acc35cc96f2b75764dbfa5bd57a08ddaf04c02f80e49d62c88a8835a62c7f1ce7c47ae25d9e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f38c6bf06e311b80a4f6aef9495d5157d66f2366c10af171b8784f7dbf6667767582f479193c84fd895676eb2dff16b29b86c0d485d08121648d69471e1751eee3fd443e715f058b8ceac40d800deb2d1220b232485bc8e20b19aa81a0b293430832f3c3aa833e68fc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h752ea928e12473555564091cf352019494f38c8b09a781bbf9956e0cb7e975a2929f01551a99bfbf9ca52dfe71d5b8cb33d60f305d4584c92d31c302b905191548667a90fbce2e5f7263ae6f507a24183808272084b02448cf1c0695e92811ffab54a8e3c8c0ccfd0e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8bbb7e2c9bf411c7dc5478b0b52450ccfc3cecb173ab14cfca21dae118a0b6ee8781745d556c784c9134d5f9f427e85f8d2cec9a8502a3b4451f057904a7adbf994dc5463c7650de8397f447ebd44ca7816c4d4202fdb200e4e19cc814d24884982a8010e36aad81fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd4f7b02f99c6c815150a97b58796b95d1943a38294c1e3616d568349266ddf5533c33ecfd6f374256dab9e270cd910aee5ea17dbf74881b067e73e25917f706c96b01faab6863366aa9f86f630d64f737d9bbf4b28568693cf85006fdcbaf758af8b228cbfb0f33c0a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he527634d59e3c212549ccf40a977997c66df0054e7b0bf2fe67598dfca293d38c24b827a4c068e72033eee28faed1f4780d87e4aa367c143d3cd6eb8ba1fc876141947ef22a27d5273a47064bdb8f550ce504b96c8ca49a4abf448667532f49e6876efde47c7a3015c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf067e28de9040e283c44489e2818601537d4c31074c7cf6ec9641cb33c87809f5d52c29a23877f4290ae1be2f1896bc60bd0534a2189a5daa3237b2ff05d51239283c527f4b24c4261731e5cafba6993120c3c69dfb2b5a738b1dfaa0522625c34fb12eac3441faaea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5a22493c9d2f178780ee857fcf4ab8b5b93bcbba4a578297e6a6cc68cdf76099b89ee231ed892fc4adfba9cdf4fea9e0d7c687eaaf8e3bc05ee7b529f2c89841a32d0215b993e962aa20df0799167a3ed0379bdb9b656251b3fb00e5a0b9e298fe492647143e622b61;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h105299e8fa2305c129ee2ec4d5e50668b103ef79edf42dfcef798dcaa74fe76b2e6ad64c6a5f574eb5cf9a60051d9119603c08183759de0c08095a11d01d44da66bd1968a5deb858f60c6b0225634a785e3227fbd74eaff970b7ede359212d3e06324b205db7acaa61a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c577847b0323b9919cb9970ed2b02f086eee3d44ef863ab5864293508c56444f04666b009fb2159e8e53226af1980502961483548834cd90cf9a2f511c23b9092da8add7a42205ba36e5d205fa1a8d5154b24d698f1b5caecd51b4691b55225d04874c8246f709f1e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c690db6ffbafba261ef0802893b32e62abe4637c2f4e6f846ac70227ff596ca244777a29f84580adfcb7ca65c1476e9e6fb2b3d45d9fd15fd86c8151533e1ef9b72f5476499a0eed0403a51fcd35e862bd5054ce631cdd6890752cbae038295c7ef4da2dbe77b2aae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h361a77dcc4eb94260373eedd7e360c14341440f83bcb851b7f34999cbc7a8e79049e56de5811672c8d49aeaefc2986027d4d03c0bfcadffa3852fd1a7d98df0cc97c51dea7b1673cf7fba3d78a83c317576c0c354eb29b51202751d3384aefa86c49d79b7e9f5ee316;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d86a0e42ff5b2967c6625dc189b14fdc0e3b4368a933178d1860d9311fd1c2cbf5c8964e7bfd695e3ed955dad9f7aac091771e052e66fb3557340aedf6d6aeb3d9e6176b0ff3f3d0bc941b51ccb521088519d9851355976c7441b2d3e4d5d0cfd0cdd05658fe8b190;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h48009c7f5d2db3e60152c19f2bb87863ec2904c44cf4ce9c2237ae929ea0dde54fd8a6472231b4964118d3f078b84b0a489155a35bde98fb6427752ce2f90de8c3190f3c2c81838f8da6a3d4ac843490bc9d51c7297885dc0cd2ad5abf45165cf092c51ae34b189581;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19d959ce42587a5a41f46d77884c5baff5c698481c085bfaed55337b33b81022f0f203a437a05b73d6994aef99a7b320f44214cf81d76f1e5953baa363bf6c3bb7f9b30a994a60185129400de5bbd2d424501ff50227b693028888896cdc3df24937dad4e31476508c5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da3afc3eec03905bc5e98631b4b9dcb81ddb19bd750a653e7bf95456f02b5d5c9875245c7a1bf15247c1728d593d8881f07402f5dfe3ba3bbf90f7dc02493138186b99a71d4e8e284231fffbc1109d5b2769cd581ec9f874b5e8a30b2251c8b9fb835c76b68fa14fe7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15b00d8c551f9de8ce005c65d8758eab7e4f5d07ba5a0057ee8db09123aaab6272e9ef2a29f7dd5af19a1d502476a0354b2787cfe4519956b7715e1a6d77376ef45a00f175d9ca562707361b24d40d2c834d7a81ee1b2303a0bd37df9845fb9cd133936d21cc13a4a8c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h166f04b97f0ab952d2a538306e6b28b2456b9832036a30009100e453ce74e766a84cf16046577aa3bf191c0f18794e4908fff2c04150a9571e5f8252497abf45e3a8cde9168e3c51cd5cd6027b21d7b6f2e6a26f2c2e0dbbafdb88b3ebbaa4531b08a26bfaad6cfc4ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h173fc228fe948da4df8d36e8770758b91b2e3459e00ec2a97513b0595557ace1829c50848aa8401ffe00e236ed62642a3cf90272c80db00d61f7589ea7752a2a1b5f3cbc118b063331997647e82e410ad81692383a7eb87df9b5751d8d9752142d5fb2706163d1ef628;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h188dcd359e51341185d3cacc9d218dc139cfd6d6b86168892e1e08926c2a3c104cc71bf428a9af48d6dd4ada0080764d3f5b644400c557a43b235a21d288768a8b71fe30f9fcc2103a4ebbe3052681ed9ae668d98e00ef53c0928abfc05c44636a196db352b66673a6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h33ec3c38421a3ac7ddd291029c51f8f1c0c777e6b2b48c70487eefe52870f24396d0b19a097840c2f19a39dde643770fb8a48f967626bbd4784b3565871c2fc8ae62637dcb3a5f48e50ca608a3b995e128e8b395e6012e6440ee28d18027dea569a242e3bcb5a826c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h103c02ce4f43933abca7dff1196645990af7ed75a93a2aa08c77dbcc591639e2ff6a88ba2261667f822d8e131a3acc3444a7fe1f21ca1c7b0462639981f13c3d8d6f2c67ddd0ba6f31d142725c8224350e91d99bf426b9ddb589e71d9292498beee7a3be04a98e41380;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3325102b39fe2f848bcc83e9cae5c56eeeccc2774b515f45522dc07c3b790d5953934c384f7ea20a9001111bf70fcd0e462151db7d601427376f428061c62e0b4aa745bd34f2038a9b108757fb3f5ed40d2b94ae88c933d5b0e42b930993e8c7d3ded7c902b1df918f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2e1dd0c2de2752a7a73776c41da816f214f6369218e2e2260b1d5135c584023fc86141e069a46a1011d30969dc2da0dc5b0c5a9864aa002444d8c2384f3a3cdc241f2d6c10104568f3e32393a1bead95671bc1e65c9ac7faca7e96134d410de3f483e96f85058ffc68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf433952a0263bae1210da796992f17eaca50e7e4504f5d61a37499002c1b2d78556891574fcf5e66d343a99b61de17242d1dd5626d63dc75dc928c7e01ddfdc2b6ffbf1f48c8eed83739f9a65346a6e771bd5f99234096fd738a6275238d27f707257fb4e46cd97353;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2263d7863300c49a4eaa83855c7ca553eb5626e74c9f56dd1656b6b84ca2181379aab42b84ed78b344b136909d8425283fc5f1601f5127b8b49e5513f13c9da8273fc526cf1bf2cb16ec92e30f7d46f372297119d42dcbae2d853c7d4f85c289b0d35bc47660febfca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e1c5552da28b640f92f4eadfafb059a469611ca4bf5ceb69d81431cce430562787885fdc8ca907980335e1f01c5ee91c05a8519bf8fa5011d85f41a44df017c4d382f6f0a5190f106b22fc9276d40fe11a52b2180407904215e90ab752d2e0a29ae5099a9104e8eccb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2d1ce0930c7c77f91216c9ead46a914ccf3fc7a39fc1a8601766ad85ea60003fc64087018439a6efb8b87e1ae7e79cd73a9ea4adc252db64c41e37b3d5d8571f12cf0f9d6bb548ce4dc06eff1bb78416ed798855c9460213abf7d4d8cd79957b49b9a1a7cd1f5c0856;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c44885c11c86e9b40123261b037e417033fe09eccfb564b90562d6e22efff1b46c679dd395c122e5c608d81e71d044ad15526e7f856db797ce9319d52b1e6da42057ba785442fc3c3ae1dc884b485a82dc4ca244b404bf7bb537f1759bd4003f57bbedc8f827d9c46c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe57e78a454f5bf296409a5e4f9336cdaf22cc7bb98e7c51497e1586bd29d19fec8b7498abe43bcf0d8bb1f47a6c982e0e933601a1b77e616915fd20379240b54193adc47b84c81c7d0640d4efb63f1f08059e5a38a6fcd91be9fed27301e99eabc0a2d21af08005f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae36b56b31c8450ca0edaf232fcc56998311cd134fedaff5e651b27e50abd3db3b48eef191c22215945869d9086cd8433aaf30093066b88a609aedde260f77d23bb739ffd8054cf7ad9c06fca067c78d3df3f619357e5903ecaf3ebb9b25415d0b333518fdfc1ccdf3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he2e2bef72b8c5157184f6c5d47026787c9bcbaf31b64eba34ce673de27fccef36775ea68c033396196ef1e2f7c8d3f580fdae4d327926cc9f769a9a2f937d5ac808522d5a58061b5d7cc29d3bfe46ed297eaa08de5d201638370a45b4bba5a5de909fe81e5b4ab82c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83cb952ef1d4e3f1ad2cdfc4cd390fa2fb4bec9fb03bc385cd470e2455db461128c9ad9c9dfe05dcd17113ebb88ce8dc0ac065ace23dcf69867b5caca55111ed4820cfdc4af31fdd6935e303bc935b242a143eb9186f8bb537d4d75d569ccf71c7cf2d1107ce67f9e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bb6da446313535943be18ea6a1a5f2ba7c73f8178fea2970fd025a68e76ede7cfb8303866c73ebfec0639933311d241a816a7e5b4b45961de116619b3e09cd555345daffb994543d23ad5d23c79607b170c006c59afaac36678c5823f70f8c6c1e1a68b61ccfd7397f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf8d27420c7af83db69623c89885ee977793e38ee1a4a7d1c883b7c3a57b33432c18675fef882d02006e182925ce2ed42d5b0b39d05ba0be39a3d77e4b46d1767e7d96cf78dd75f3466e01ff28347ef4b119404283d3d6e95751d6a0ba253e5e38ccdbdedd3efdf39;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2710ae634c542a9d4b48717e4ea0c73c3867a4bc8c929c34548891242c87c740fe754cc43299d4f60ce4b6569ab256781702c3f51d70a2d833fa8f66e1c20e6192b1b1d39fa057de17bcdaae21827d82d52569e549b0191c5bbf0fac1d0b91201e8933f832c13209b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1afbbbd4eebd44f2174dbe26e5751075a0ca288815140036ef85a6ee77e85069d98a6d03b0c22895f8819e7f2172c5457e479dfc40bc737f492e7025f45c08bcfd26a5a198a8b9b6f45acb143d911f1ab5fd555fda22f17a8f5013d7e9c32abf732401157d655058b1d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha5df3aae05c445f3eee961f0a14211309c94fc040f6528d68443d5b2c1da418e11aa4eb545b4b819fe63545aca9326d899697fd2f9ecbcda1c35d17f25ea79bea95c32971d6c52e3ca8383332223df5ba7badc1fca454b620c92015d91998145a4110a235238dc78bf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heb1b03c064f8f62b0874fe6806390f21ad5a4dbebf6d8c7d132b6c69cd647777a1b4377c0cea04b0dcee6be4efe3d408bd93277eff65f3ac16bb41a2e44d9e81cb5a79185f4d792af61ae2c9ad6f4677de512dc9a363aed24cbb16a0a13adef49a3287f91f72297839;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbb2a21ff497a0fc7989532832b3d87059ba21ce562fdf3648fbbae23642bb1425abdb62a952c7a2f12012891e13624c8f1b3ab47d7f1f72fe83e6a8f23a8c51e262ef63dc72a8e9659a29bf8092fe9ed878c7c2a2478eb2270978cf1d5df41c87992bc170a3dfe8cba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6169f35b7a227cfe851513d6913a8fc62af8194e355dd7d4e527342eb3ec829941698eaae1f789e2c17e1b81a25fde88784aeb90c552059e876da688256f82e590608a6ba55f166f3993ea95d8db4e2830860dccd9e4061075b40f7c4e68931590d0b9b36fd8b2f90d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1de27af017e41e00830d7cd58d76b3779e35783772a93856f591b32da44f50c62a128b0ab53d10777868c98e1b9022f28108ae38f52f267b179137dca6d8091a6d0a9e9ca2939b262eee281fb88d8b6e1ad42ace9e2e55c77440cf02118183bedd3309ae00a6f21e557;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h943464b7d048c7a8109cfd98f9cbefecc2c9b84b2397f3ac78d6c3157aca9ed69c1e84bba556c75c5970dd63dfa01a5cd002b25793150153adf082b9bbd91ea37dd0be389bea483b3d1ca0d6aa3d492cd9f0e1f44c6d1585cad02080993b4c814b867f37edbdcb0f22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h77ebd2ddbbd7272d1eea01ccb0dcdb7bb939e4f681e8a147c34a607d6dc9ffca8f8c2d49995db7f26cf491e0cc171ba414efdbcc1b58584e52b1292bcffc960a0f333b681f77661ea9c19f0531a7c617e117f65ffc99c0adc1a7feae868a08c1fca7ce2479db584101;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11851f1e095e449596a0ada0e827178c8471cc02d2325b3d37ea8fdc14a226e793d5f1aace461a765417f3b2616ae100e24b816987aaf3b47bfedd2aeca451881c347f48717b81f4a6251dac9dae55a24cff02aa8576e31d605349e7587057cb0543cdeb8e77f386215;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a283b61baff07ec95dec8c93d2ffd98fd6906b4227959f132d2b6b1b3885fca4859bf4c056fa61317f16eb10cb2166662cfb8e53f5bfb54d95fcc67d0dbd84e24a0c35415403dfc2ae2b163454b8addff832fb32015aac2dc216d07372f34bfdeb9e9936fbb1132ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc3ba71d91eef7ae8ff3a413e471a4a381143b1b7cd9edd11ce3fe9b409b7944b40feaca835acb74ced4f75b0f645bd56b72a3f0d3a4e9b1d78d1388c947c17856e4e24ec594bdcf15c9099b39d8a71492f5dc6e1e3d825df0f280c4114edb730244355d72b35bb4af5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h54b07d2f64a92077e1762cbb7465030a7c79dea85998119392997de496c35151fec7f5a0bfd935668d5baffb8532dc184a15028fd64bda86fdda4937352814f5ca79758f2d92d55d7d0f8df6871f8c3eda396d061d6ab69e66141cc17adf39127c0500ca587da6b674;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1454423ba4fd63706e64c586de61f4ef74dbcbf42ae69ca02d94a25c0f438a63d022c5032381e4b31688dec7f6ef7dde049791fa2a04c3767de468e6a4abc78c9b56ced0d2e7bab03b5f1b6b1ae32fdbc99d90af6f8896fa3b60d96e8043875ad53ea1d7c9459206e93;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8f31e990516ec079d95454ecb42bc0f064d932cf72cce529575ddb2adb56acffde9c4deacd2c3d58f0d53b874eeb14609a5874ffd5a36f8db177f0153fdbf6aa17d56a9cf9fc52c18463d2a511c702f18203cfa9d63c7373745622feee729e0dd8d2e8650ad289a68d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfe0bbd0acf909d7ae7af4437be35f87a8d79424f83c9b881e337b4308b6bafe6b97eb332fe377f5480485c5155fb0b1741133ab60eee46277d6f0b889f49911fa25eebd1898e1f18ccb24711cd89cd0414e6e0d4e94f494be07ae2b24e7a4bbe2010745e37b7926926;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd22d6c353ffe91b46dc81c77d5f537b1e97a627e1ad6a4ae08502742b001cfeb519be6c93cce9153c8e1439163573d92cc3f6bf745a6818fcc42235cab3510610a73af084c4ab0709cb67d3467df003a774b7ae3cba6b21f9a0b804c1f60b99d8e26955ce54b33cb4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h418c6c812dd90e462ba37c8d22fa8a41efa36d4aaf0391bc18e904f70dd5dce153fa80a289dbf3b8901cd7d30a520ff30e75c8b3c2c2e6c821056f27d93d3d4a24741c0513d673bc3ae31ee178ea1409ddb09adcb86e4d76f69cfbdad55ea8bde9bb524b2ee3365b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb741af6f8e2f01f59af91a765490a8916335574b107ea20a71f4075f8a8599d65784b8fecd4c2c726fe604b5a19441d0da02c2c21270e33e08b2e8b27239ad24df0146d8c46ac84d819f6a8a92effe598ade2cc6148b12fb6cca1970bdf293dfb5ed3eeb7e8aa1c66;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba08577cab37441e79e68fbe172b1252edcef2937609f1e15a54c0d262f6ede7bf8809335c45473cdd3bb3d705465759abfa77989470bd37bbe5d2d1a3eaa9f1fa6f169664f312769c2e27b96109d03d3305b2be1e656b49c921b98a736cb4d13b44765aa716a19837;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha23e7bd030b0dcd58b558388123747c14395f2d2b8f69b5762e39b783b645e72fb30005c4831851c3afc1a3e2ce3585757bc7c85171f99a22f116ae51028e3326831fd61dcd196224edc3911e42d6b181ccc1289f6e9ab520ca0164cf5a5ed83b7d7251567f51f8f2e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd905b5f7de879dbd44bf23509d9ac4bcf93adea3288a0964a3c9863b874198c6523ba53c84fcb12130f223b038d2d8781107a7d4640158990785f63f7d9ca662f2f5fc85223e4f9aa28cbed9ce98a5a1be6b7325284cebffd3ff37176854ccc4fb4d9dba693444a5e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19824666186b15d898d845fe120094b866d11e4696486f3690559140e6b7b272556e6e833cd6a393e9cfbe893c312469adad49924fd894b3d9a84b5b32f4a085df07e53f968fe0a48713bcf4e7b1a4b029366220ac302439a01822ee82046c20429455342a27b3a6564;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7226ed57d0c4fc06768deaca5d8cb43bc122631be2aaa7303d3e4c656fd8fcbc7c9e8d62ed17b516ce9f71f0f00453ac8eb90a11a982405ddfcf5cdc4159d92d132662adb357e8b4eaf6489992908b91ff38266fdb419433c85e4cef09c16a5ef58b256d3a9cf50f54;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd24b192b9bfff001571da861e0d89a98ba249a224295ae0c2ced3e37d759c4c0ef7ed7c589b2a156c53c3b9e2e9a4214833408ef71c5e106bbd59425cf420d18c14a0ef10814ae8d52f89c6a9fef88ab842a0b4e1b9de6d8928e377b13a12ebd8ab96c2b8eccb2855c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c9a2b686b457b072117b9a2ed71823008e99a8f1cbe84abdaf1c4f8542c659c7516d4438ae97831b5ceb796a1e7b30d456366bb5f550264a64d9dd515c857e1a7334716b79999b3da31fa99a2e3adc02dddcc1da1ed4b2b45dbe5fba4edf0e68b9865f45b05c2ac203;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f7200cfd929b9fdf431b00bbb82aae401508a900cd3d1107103b9f687dc7f2ae630a484a7b7e1b89dff100b015b6e16ef814aea688788eb649c9fa85e082f47588879c7cfdc50b56192edd15918b0942f34b089f0aebb3bb214aac4604d25a34829f3a8ce90c2631c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3db4e8471a49c7023e71b0f69d7fb2eac0cb0f39ff741e38758494bc898ec086764de8aa99b7272981ff81dd6ad95713a00db53901a184be1ee6a98c660368684d77ad3bf6922dcbdd7c876dbf3f7d6c5236445b76e6c39abe696a6fa34da45bcd0af4531362dda613;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12e52342ef8041ee7ea1298229cc81d10372a4bb9ab734241e3719529ce36aefb7d76cc625d64418d20f30e094d0c305b0281bdbac1f0ec190ef5ca72217242c1d36cbe44b9d6b9f0cc8a13ffa86cc77121519a29469c6c56de939afc9f887da57c3682b4a13d23bcb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e7fbb8dccfd36c8897b4be5cd6d009fc26f5d6f7d9b2afac240820a71edad0845dde2c4555118932d68fcd74b5bf476bf36b3200e885f659d882dae249d666502566bde7d261f75974a18c56f837dd5cb79787eb7bd334a2ecf816265bbaf2873c8e7152ca204e5f45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175ec09165161c5426f3433b8f84e12bd6287066d20fe8720578aee5604d8285c45da37e4e3c4dbd3168f863e75ea951f7f0a73d803f65cf4ff057f7800a933a2dd9578ac71460dba85129a2fe56945ea70b2010ef19259ad166dd9ab389ae5d2c0e826f6a48ba48360;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a50711d580f7dca1e7a0c6f50b561be97fce36f53c9f17fc732751203062ad4533e7bfbe5e798301646a2e075b0019c006e9f17785cfb69476dc7db94b77c672991bc95034534e8cce6fa6da95dd4f1538ed191a5f886ad152390ad9760182bdd224af8926855538a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h169995acf9db6e549c7b8bdae387aa5af32fc896e6a2afe821128fb672cfa7a17c2433f6199e8fb6104d5fe818d2544c81fbe20f5d4cbc2be09f41291d5e6b7eecccf85cf569cf283f0e811df33a73b00c9b461e10b8cd1945e520a65eb5564eb57164b224c8005cbcb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b02cc34ef74c265790bdf265fda19588e2ed15044ac9af963acef9fbf2abc06470f357e47677ae853ff534fbc8bbe869ae2570e2a8acd842bed2351734d2e62c63d999bdff6837e92b6f32f54d6bf18ef0985d69df25b091b07f3fe1935927f3b8f7c6ec5de0093fcb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2649ce2bcba93010c7beb5ab08587ac5d156de7967e43084f3747c7499ecbd4469eaf06e064ef06a3e9ffb009ccfc947c9c576eb9ac44aefb1b9e24569849aa6f58444b4690845e66735c03b32b84e4644d2e84a417896923e3a4f1cdd089b8ad7736b868f3f49c75b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1066657b91e27e8bc951875c416b33980370aec4a23bfcea28d2862bd619a28706ae30295d18c1efa7fa95a5e0e07e931a235c30dbb0d3ac5844d7f5b40b54c99bbde773c9110ac5d2263d4667cb9c7cd1b93e34f4100b1c38f71f2dccecb454e32faa87dcb54df4d14;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17300a4c593b7a8b939f0784a0775c76bb2f64b03fd782a1c0f94c44ea77473c97e2ce2accc12b1a090f4cc1051a1e15cba316d664fd14298903771389862e3d5eb8360b0fca5b8153cb4b0894a750b1cc308ca19a8b524b0812bfff3c29cc99c3bde3dd3b65c8f0770;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h81f10e628a89e2c47e9fbfd99853356edb597d5af1f101c1cb73add9ac686308caae8c2b4268713eb6cb8320e706c4dbf72da9f1b1c95e03acde7e6e36194334579f452251fb2df67d081594a9d9ae95c12c6a6ed26c353b920c9dd835c565c477b3e32e019d34fb6a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e7074648ea5188b16644030a2167d5dd0571bad629a24ba835438ac25426c032c72ac9e682f9ad5cf50c9c0a116833d41605a92bffb739340a48cf671c597502864f0eb9fc893d395c78efeb70d0f981be35f9635cc2e72e60a914cbb7514fe6a37b959a0a60c0bdf4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha2e2fa9ec4f60867c00883526c567202340bafdd945ad0d389b8c1cafb4464bd9e6d6e2ec44b93840079077e190748db74740af947a28f91365422dedd9092e278d9f507b7c7e70f5cd7c6f52c0524f3c6fb2a5eb73598fa2b60492d3929a598444cf85143b3bd1b91;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfd0c612427713653df725437bedf8060a6e639fc41f07a5bd753647aac3c3e786e22103efa95c9ebc09a7613ffe4f252e6ef9fca8f87b43dd678a9d768d51369c9df87652768f0e950e47fb7b6903d45b3f4beb1535722abe5d9eac0cc83815a3618435353aa1c901;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h344daa3ab127eab825d8ce157ee59bb90ad2edd1c8ab01b2ee0d7acff079efb59be9ccc6ec5c0d3498debeafd6cd682faf61983bba794cc3523cabbdab0744438e1ba01d25cd6ce25716225abfb2eaed23c6539352641089219b47483911c8f6b512038d9c89d07be0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he048503152ffe8249bcf5f1fe8acb8d6e3042ed3e9d2e41af1ebbc504722416beef395c64cf4a0c211a34b677a619a5cc79647f530f5cf753887597da33b146b79682987f39b66fad68d821bdb69077abb94327b5de9e2f92ba4592d900f4e224da9e5e06229cb7554;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3dc2b623ccb2f19d37fc4b3eb0be7adea481010297a2a6731f5f5eed2bedc6eaa37c09e8b60fd6790dd7f6c1b07383f622c5204d007f42ddcd2c57c984f7e0eb846deaba61556023ce4c35cd46e7b51622fcd4795ee187acd278e9cf974bf67684e72bade435ad0898;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1341702b9b8804db56cf71e74442b873dc56ad3753ff7d169cf3a3bd989106334cb904f6b14376f03082589be6e82e83d09b611c6940e6ba2450c22ab68b021da1665b5112d20b7d965e1671c857a4fe26a87894a54b5bc123aac0eccc4267ec624dca90d3bac477b1d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf03f0f1031de1381ec6d5517457879afd261b727c1a10c06c84d6de00d7acf20291c61c2f900446526ccbc06ff858c8987b4a47e6fb1c51d969f08d4470739c82080d5e8394254ae3e170e318c6b692b88d72eeab5842d18633d0a121c6173f2c627d2b3ab879cd455;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fa0ff6d9034f91ad5bbf94d693e5f0a64f588839899e0778f1163c2a9cf5d9883855fc53cc8b77cbb9f46b09ff1433eac6786cd6f45a1f903295eb2deff19cb1770d8d878f545c14187e27af30fa0f62c39bcaffe8e926708c095458881e35a2caafe86d36203f65;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he53a41ac02f573f9d8628aa8080fff6814c63b6ae174206d31d05455b76bb950bafe4cddf421c7d5934acbda1b0f4542f008b4d15dfad7580e1a306bd78c2802ca0508a614c01f042cddfeef932ae31bae7018079708da7c6f890ab2952cf79fba6c2d74dc7ff676a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d4173e83fd8ff03572d55fe692751bd6eebb65d61fb1583b73aed25ebab4b4f8864d1799f1bf95b8c90d05e228aa9388fe8d826dac6e0404d043f29dc699fc1c39e29be8e369d06ec2fe5b5ca56af7fbd4e50e8731b85982ffcd51e7ef9b7cc5d77cf583faca5c503;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8478a0fb349674b7476961a6c7870c5d7de0e85cba2cbd1f06d58c7a1a983ae56dac0b3135be0be75ff9aac977e0d2bb239124df0176c808c769fff099020069c59f319e11ff7d340897b0d63d715779fbc5d38352cd15f1e3865200148ea4a4c5c22bcb47ef9da820;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf9cee0ac4e858b3f9026592977fdb314da270e4f74c68ec295db1fad753007ba4d07f4e68a791b6441897f5d5781ceb90815d9a0d0673739ef65529f6677044e19341298b809a198fd27fb732f4b4bfcf23f91983efcbab5657badac75458e0539c2f66798393d4847;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a5b79c410a89eb0500380deccea5157a561b79a9a92a898c27b2538227db5893eaea7f933adac1128f1ef2746ee7d4cbf79aa62dd9e388e0f4a3e631fefa24b4e85815a855d97b843dc1f91f580bbdb92a72b7fb956fbd928c30694ab9bfff8fcee956bb37527b50e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1508c9db8e68260ce20ffcbeea6b98d8911ae71c96b9e4961baa23803796080872799c79e6f0cf2aaabc062c2d55f76b74e4d1ceb636abd3c79bfce936911e43e80db986c8238955868b9bfe6c82fe62ca50ed3d1791d3a2b64a6d455845557097b52c67ea8297da833;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h107bcea9c7294716f7b0818a95acdbacd7c48375e79fcb95de43d3186bc1d6b73bcd46aad342120796dc671aa77ac59b762b2e6b91973d74fff47a0479e5d2e63e40d9f0c28505b6bd5db571aa49351cd63386a4c357ba5612d06014e4bc6ff2266ecc1fc93a159dcbe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2883c2746e41c83c94d120c6caac82d1b5a2bc8f33df2fdf1cce5c15d39984fae36951de1fb28a2054ba3c8797672a4535b09c6b32d6d755381c107d8a0ec14a4889c31accb7cc863125b30f7c2e89535064413811fa85dfefdc9e64a70069137ed0d44ecf46c35ecd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed694978a74fcf31d59bb421b961968ca1ade5dbfd412fb53fb3f362806f7d01e87da6d237dad74b40cb5ef8d96b0821d72c6e096b8a76479942ae2d159cc2402d66d0ea8fa72638328411823a7454eb391b6467b3194557684d156a990e02facb6a94f4375131ac27;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c49434b0bb81d0190ad8668544596d381e7ac4970cdccf799db976b5293ce03accbf54d6185b4b137aae6dce212d90b32b375977d314d25e687ebb53f96f6ba131a120bb9ab8d5d53c7e2d5a7ea838aa58e8c3eedbc8cdabb4132b346760eaa5ec245811030c49dbac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'habbbda0c6dd43164cee7dde9f7cebd4df96eb05837939610057622243cd4d0a2c804139df9d80e89bcb8317a05a5c8413936c2291c7d19e828a8246d63cae9fcf7edbdbac634de4a8f68915ea05e8e5c8741646ffd18a86991d194b4c46e6350a43572fc8e32d0aa0b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59485c123d3345649078ab0541b7ab2906dec7f904ada91e93b49b388c6484b1b9f883cd133c77ad37ee6c0a511f0bf7e033e31110587c6698cce6756e56f67fbc5d78046e542a96dea93278acfb090df652c1a7a2b3b6e5811e8c973e78ea69e0f85ada58b01f7ea6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8a2df72f189258fc06b2a2d6f6b75ea0c1e8111a79ff3b21e2950c59bb3ad333f1d1100609024ab749f86790d27456759d1286db4dcd8f00272365ee05bac658c69550bb410f109d19c371fee545cf25f1f24f200e08ee4d9de1b28097391b54b14812c16d3f423365;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4bd0c5f0ea25a0ae2dbc9d6ac892e5aa814bc54453d3e465ae8369230e7b8dc2edd712281782cd65703608a8ecf2cda0d6e2ff559047478f10524f534d2ee3bb11334512b2868a45900f8660e8cb488fd1e283bce4df8ea70144f562d2de8612491c0b10ccffa61fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd99379589f82b09799745c0ffc6fd01c81f29927be3d775646304ffa2059c61842369887907f05a139d97b03316e5f2e2b0c07eb60171b46cf7d8c7aeda6f776e3c1d9db57a6a9cdbae5fc4ed06f52a7a09c83583fa8a0037351a00cacadf2f925c98bb47c0d740df;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h44de72702f005c30d2388434e43bf3b690d1b80a08d488a280adef0ad5771805d4e6244bca3fc78bc5afe31937eef3774d2fdcfc68d443636c53d3bdcb81d577011f9f4f7079b3affff9a6f35831e6bf46f347aaaac256fe17344c612bd9b8ced13423a039e4c67a67;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h172234b4873752f627d1144c50808a876ac9748bdf7cf521c5d4ebe1f794c9042631e060191f8ee718b1df3d50d23d1c680400caa7f2d388e732fa2e7ce3c74d6d18d6217946209bf089d7d32b1cbc6a3a12e5102ace77d71b5a2971b72b4ed426f2a62589752b293ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb40a2999a29e4567ba1fabd502d098af67e2227cb28f2e69d868e4754ed31bbec5290db07985cfabeef61f1f3a0dcc1cb7b56f020fd0449255f6e97fdbeb200092849e53459db9b4ce08414f7070241275d8923cd1204560e8a6c24fd70349193e78f582b78e2c7812;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38261136822c9a9108ac3741da072b18c438ddce17f842513cbff9c773cd3582ea42780c4c4f08ce497ef2799a8485f1f7e5b7987e453d59a04c3b0835b79a4ee7d175eae67b88e08f31ddd43591ab94401485bfe87f8b9ef3e6eb5e10ffac8e6ccd6eb61ae2e707a7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e2630f74d8e44cb90b82f91ef40a103b2275439d83c6798ae5fa00e0026a642fe3742ea8a9efb79b1435c21272f7e203cb60b336929e668574e8e88e3020b0e73d8ca03afe86abb8f13a3f41ca344b7a704dba455d695b1b5a814ec95d94a92b79b6fad4ff9c06e90;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h154e6b248146042906d006f336a353f5349417336f25ae268d15fa2a00c96f92fd90069ec281d7e4088d68ec0777db9d16173fa9f7461ebb664a210e34681517eb2a039babafe4b04febf7988814f65c4e6d1758c04280efa6d455eecbd4f8a9661216805f5c6ead013;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15fc462911f7b0f34f102c8a6ec31ec1dcfcc3ada7a6b431605e43ee469eb3908677529d07d74712cb152f819fe302e2e252f5aa0ac6b40bac70e63b2d5b08bfb1b27436851f33f1ae2c8317c8743966e89a259bce78520b492c36988288c3aafeb6a7e7929d55171a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11a136e43f0747781f62ddd3d32c60c0b1be403740ac086062b716e9f62949b1c771ba1dd255d905f21ef835d44aa7e3bb60264827418ffaf0100b92db690c490056ab5212ecb6441d8abb476b4a100b2766f4dbd4b7c6d667b7aee18cc60ac1965e68992851365419c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h77160220231d44c87d7ec9bd47efc3e67720b85c33f82990fd03babe934f99c77846e5c9f605f84b26345fafbba933a12c521ab3ea1008414a42c0bf7fc5040633288f5532cbc4a640303096a4cc6f40a5fb6937eec4bf34512dafd2f20ca4283a2f8c83a82106d679;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8f58478014d94b2bb2226c1282c907fa5ec9ab3ee74ca71c1fbd6c53e14fdd39679ab57e7e19cd621df65daf71ef5a35e41af5643681c1ad1f58c0f9d36b07bacef9101f57438d300c92bfc5760928805e205d5dc353a71e379ccf0b039d3b85f3ce48222c81f1202b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17462155fe1d731776264ecbb065adaec71cab72f73685041d6d5ddacc6a8c1d62f7f85369f1e8a6b9097fec3baa662d928294c0067278cde4d695c421298ab98763ed6c85eddb3d7e02696826d41b276e755b93c1e657883aa9c60c8ca62f3d90cd15c0ca0c888131f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c322fda8ee01d126051a7b2e18614d31193d248f97a38792e4912002fc84faf256a84b6306fe6308aca607d12c2155f6eef250d03b0d7d26037327cdf0e49cfc80a2619f1028aef27866f8f136e99b26998dc51b30b2a36e8bde10b8ee593bbce0dbf99dd813cee481;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2084897e02059de74d8ca0d33b568666eb549db1498a3cd9c22e1d9cdd1978777e3d7aa37e8afdf89aa0b2e98c2dcb42261187e4ff6ed50e24aab7dbb050c2bd472f0c6225840f1dd4e5965a7ec15f6761df4f68a0ac825f9dd35bb23f126d33ed27eedd729ceb1d46;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1897e04a52c6fc52d66221906c21ea0cee09ee55f4d6b0190f397a2ecd218a672bb42208ceef80249711b9358b4fdc9dc6bf066b9825559126375fd83e6f514aad4e64a83d4c13519f7de909f40a140166138ac1f10f7efcb17f90340a3be510563f7db291a4012cbc0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a1e6aac812264287716ea6191d39cc5a51bcab0f4ebe68b7b402141f8944587d36357931928a48be38906e2470b6f166d1e571e2047dd25feda825681edc7a20da1cfbd0142220c9208bc9754300c81a17835de072f77f581cc062242c257204f42ac13a0a2210595b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b101d2713038831e3b6d1d9849e062d5a8ada82940a3e68c06c21fa0eb8c43ceebff2e3465948d55a74ec1ad554379ebd77b783e0d98661eaf180f3f992546129869c2c7feec4ee488e537d9b861442e2e81cc003e268e2860f49dea51f81d9380ae8a50989e170846;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e7f19d4a74f161efc405316c9f1b132f1dd41c33828b7778e57cbf048568d2c550ed2b4d9ee8b5bfc5ff66d8fcd4235d5056c0a85160ec7d948d37341274815ef42e709848185de91e97016ae96821bad627502564e20af4dd6d0fc019d6638339877a00cf3bd0d896;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c1a37af36e1a7fac15f927050e8f115a5238e1e38e75c0a02a2dcfc78b096328e3f65c745bb164068828cd9fc0ceadf42a13b99ce0a513632d282b0521ca54ccf36bb3bb7cce1f1ada07d13c941792de92053dafd25b3ccd3d2baaa63c43cfdd1682580f27717fbb23;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h80b281ae9df85fcbe43a943cf299d5605728958755ad15f2e69f69bcccba9a211328916c3331c1e4959816615d6f3f577214e3c6f3a3663e5ddbb4778687bc9623d27ced1e83902d38d3d90b2379dafb6215a08834687f78b64a5328e8413b2226dd6a5cf224dd2ff4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9cd462fdeb0591de103c715ebf8a9b79373657992009c14e217a9b0c3c51f90e816e06cb58157a75b9e18b8c2333a674854c4531a01b5481349d514f2a97d9208f8f3687ca31b65c5203012a67fa07f201b1f1adaad3083ec244db6665afb4afc859f366793ce810a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cababdd511af0bf3f98bd1bba8b739a9bb02f2a11280cc22f351a6703bbe8764573e57f9eb738e28c4c741f4b206daaf2726e316ff50046785aa56d93e23ff5dcec869690d2ad936cbbb94dcc94e8c56daf8d84c8d598a863249ac721424cb06d1cb439acf1d141598;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c895a4fb5ef899aa059576f7042a004060457d2af866868e2574b5560b01a0404906db0762692c7edee906d29183a33c7bfa510c06b80b70204d0ae0052dfab85439157308e559853b7677f1f3d984d4f49c0b617d785810a56b79221f16312300f72649da7f7f244;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd6186803f5a76c2d55461c3d03274ccd99b513bb285a80d83fbfb366a0e6ace36002b1ff1f5717f4a9162f750f4019c681e35c73041fdba5e3129dd99c800566387a712ccb2916d39ad99bd3e0556345b8e412c18b6c89ec6953b1b7a9bd7cc91c1ec42c1dfcdd7cbf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dfdbe532cbf4fb732c03f07c722c8ceb759931a3ad6daeb1ead5ac79222d0dce34f659b374f844eb9f11a906700bc3a2bda986666f6d96740727ccf811bdfdacfcdc5080cdd576f32bcdd91cd0dce1d4296b7c418face07e4337a097458b5c85f5e3399ec881a1f49f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167e2791f8f3f7879bc7a2ba6b99a6bd9d71a9dccbb1052fada29ce681e065ee2a006c2995087aaa2fba11bb890e57d42e137aa4a8e284a5e3f2ef95410ce2ab0ed4070f9450644e4afd282934333bfbc33ccf1475011687d7d94c473f52cfdd33dcc8eb4a89cdb2726;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76b1c72783782dcd0f3d9937135b273ed3847246b7a7c68f59cee507c7e8907e732919c2fb33ddd37cd748e9f4f3b84d8caf7bbb7ae25c34c340c399df9f40347a8cb0f5c13d30c91e53aa918bda4b6d0bd195d07796702f2afd95c4783d2b7771dd0ccccb384f08ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd494f673bd547c915d0847a991f93479802ba39de7488e8a49e3728d54a4638095f708ab10931394c66fce3d58abe26d2f0e8d1dade7c54ff9c468a89cb837bc7a5881f4741a5f44c103306bc84a9d752d3abe9c1b141881316e40e32fdbb5fb27c88e5ede77912acc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1acadf0b67dc19c798839fc4c398a4da1512cbe17b044ef5e4b87a26715093686049dfe3f96d5d372e661580a2e719e7a0e0dec94153c5d922c8d95441a9f67f8c0949bc48775d18e64df2d88bf5fbbf9da1a9faf504d26523543c4290476dba576f9b069756fb58f69;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ccdd68b5cf3d1085738ef0730bee25848dd667e5fb823ed1647d7420ecf57af0768bf3fda12432362da4c9299ce0cf10ca47138ad99ac7089e26134fc87d4d04df39ce1d22200dd21070bf7952ea5d4bc9909a5920965ce9a39d54b11c5cfb1c8050acb2cad792044;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfc2cf6ab4ac5b685e361a7a02e8a0e86bb647fef2255a5b4cd36fb77c99e60412c023d085f174655044047255dbb57751fa676d53caeaa4766eeab513a2f26f899e74ee56233bd858ba1ebb991a37b7417b4f4680ed76eb37e806e5eaa6d4f1cb0ef4611dee8155c13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc2a55b902fde9a95bc31baaed7af1aac19117989a551cb07ef4a605fda2b787fdbb629f14b2034b280a6bdae5dd33181c65566928a69da46dbe51764add62fb3eefc7bf86f8490d1b86d9482df7f3617d2eec5779670af2d87e73e3fcde0fac75b1c921feeacba2bcb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbc2e3174b26a8c5007db0bf3a75ba144f28504e64cf5acb246591279a2eae6efb9c90632806e46b921bd11f676ca864903996922a05b196393a5459170f1c4bfb8b427dc2659dd848cf1045fb7b85a3a54f02b0c92ca475f5f6eff3ad5d105b483cb355a07a4840082;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16e18b9e27d0d287ffac6a4343debf3131cbac8a8531444ac0366c269bcde1429e11017fe01a50b91d4290d18b0ba7d2034cbb2b489bb20cc635dfa43b88625131cf68478226ff422b30d13bcd1215f0d6a15754870e84a94f2aba213ad67d3ec62739062be8884fc8a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h168c5fc7161955ce347407203826dc760353470c2eea7f67c95211460fff489288ea0bd3a26ff5a86d61d75d3e23b8498538259366c2f363ed8404243e0c57bcf77bc62ba773ffcfae17a9e5ef6f11382e771a897494ea5a0761530d61b8646501cd16edb2231454709;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h107e7d27c27866ffde78b344b27856ae71c8249ae8110b9df0470fc4d9af46a54218bf90243db8b7fd357eb5ee430920970fb7ad2a569e1ef881433d04c8d30844ddec2ee879512fe1f8a6390b582ff2c0f81076610f49d9abb2711c7fb406074a66624e1fceab1f4c9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f0ed03179936be2176c0b44a9123b50c473bbba6e5c6b592558ddf32c10ee28f31bc68852c8cd6cfb6862b72fd5ded0aad7c558005b0f8bbb86313f2c3a7b950b1cce0aecc8e5b97365af2dc65feb1e1d0fafe17ca64dd72994cfa046c154f472346729c5e7faba1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h81a2dd65ca880e90fae8193906a8f7ef668571c9217e113e4bc948fa871f650c805c99a132e5f22c016e671ca866825aac5122be2fe6bd5f812d4b14a13cc4010426d44531bd1f2ed47e3b8a15494fb8eb0064902e197de5e03c15aa326700469214d1be618b00070b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h550118ea3401c4f7694d601c4cd0427f117ec0e05e8bf749589e8f29d0fdcb463682c1c7b0bf8bb02d1d67dc685a7c82b6fae19ba44ccb17484aa9da0c5149ebaeec2de5fe9f356b65ed564f23e94fd2dbec7b8d8cf1342505447d808efc26399dcdf9daba40c8dee2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed6cc9bdfe6d3f8a6ee6cd17e7515ee0e01bb14887032814c0d5094bf82b44c56828a5137a9cf0f42cfe2854526c9a3898726cce3f2581902fb453fc204c14bb4cf8d4e747c813b2593fe75874a48c91520366285c753db242b74fef1afc4fda01df1ad3992cfc6f18;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h22190a0ec9ec1fa99b1490dbffdfdcf6ef8a5e13a295b08d00a593846203f2d64957f914c6a6f029f5a1a0ba7157ebd0d133bcb068a66f39362f16067b438801d50bd61badc1fc36baad828d7ce59d204f258f8fd86b063faea0f7b0fd01188d1fa83301e55d785964;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b35999af27b751e56f993efcff800a512896a29c25a87a9fc7c8c1a79372fb91bafb2f1ba7bc8c6150d654f66313376f2077b83cd8cd65b241326e6af3a40e67e75683bd70aef52d73c63a409b200b7234aaea69eefae8f77c182933c224fab03106860ac46f6872be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h774a82bc03614da1e74eb46c16fc030d7dbe0610fd681debea045c5eb5de09a4fb88f59805044cca1b5590515a1c2b209871b2cca04cbf13d0cbc9c727b59504ae92fc369f489ae109ce2306109b649d218584eec8d0d1d63743b7dbcdea3e6dbf2dea854da4f0d830;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he6a867c94800a9390d4fd88f22d38fad06602fb1c6e42eda764f7cb4d19b8736d2ec27145bf1a596c704e7ff03a46d33f4862eeafbdaa8583bd79e8a03a4e84457340ea41bf234fca3bd399e732a09de6fc946132b30f29d3d888c7358651fbd4031f550f4a1fdce3e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha314aaabc5da89c2d95c27a779021f73ef58e94dbdf5c96fac2437b8f652ba69562572bd0b9cb2bf37d2d4a11a2de3a9295df3d96672fe8a426c315cdf8e3456f5f14f46031431234489fec5dc01820e7f5fba8e9e041e839c016a2b85ea515ed31e31f389294a76a3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ce79627bf96f001d77207ed0cf0828f6494f6687e4c393456243e140c4044a04e8e977042964f7934b6dff9937c475f2a8f7e1a59bc02eb0676a334ef8423abcd28bc965fad0b6273fade00513ab60932cbbd225a0f71d5442920e70cc9f3ee08564b874f2121478;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1413c20da1fec79076f717a5281f71c2c3d3ebe58b27c328141f0af92a5b902da88f825e401200663b4b58cfbcc427c6779f0a90af783bcdfd9e2a9832ea8a9aac4a18ba03e126f874d4f1484af0cbbcb3772c4752ba75eb8a7e01b0cc80d560cdc88049d4cd3056209;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h92ab26cda1859cfbc3ac97a77346b84c0f9d34f27c522576a16718513953c9f14a2e07c32d049ea44c907f83b181930944f4a0c84bafd87f5e3268111a557e404610333d28062681e8d9adecd59a1eac14ae1f803f24e965c32532c4991ee63833f2ecdcca7308e3fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c64bde46a37ea27955169cbcb9c87ba32c2f8a28fc185250c54b1fc2c9c38efc86fd609ee580ef5410b3320330e99a71be9510a05adb88ae867d98bd3987e264a429fa3defdf3f41935782035e565c35c4472e33cba758fd93a0acf36c08be180e8abfe5fbbb27bf71;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9760809cebc8f08198229e6fa669694cca5a635182169c3021409f19c79aaed04b1db7ad99cb24cb7acafa9bf860b95d516125dbb57e48ec955da0efd975dc402db86f61c62e17e93ac1c121207bf3a654170d368853748a5107797939923986ac5b387a755f31139;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb02e217c6e2dd45ad0b3a4e63e5d76e2a138d14b5b276f37927f1baf1a50cd03f9c632d4bdd98ec643b516a672b2f6c451b4989a415128b3af239f333246e6166680a09e076a01690710593c151b290313f87950cb04745afa40b25b7490815c9105a0df3c54fdaae1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bfa432fd1892984867727050494e4950a3679e9d9686a295a3240756dca0e8e5725ab98b945e9c607121284e1c3c2a3ebd9cb22b9a1c26baad32f980a8f13e40bd7ca55a06ffe0ad5d54ace0334c6a991e7c3789a4ae324a83e20047f8946a9b5efe42b1676870003c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18eff96b5bdef872892e388bcb177f17e847a512ae263c90bc6bf5687839ee646f9d4fbfab5c1f672fb88329aba4fab723a73fdd5e73a5536d2c2f1730fcbf2fe3367ff709ad43ac3bf3fd8e67b4acc264410d4bb16e26cf4d366d02ce86721be55044697bc43e36305;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15bbaf7a5d4fb73b38f3d8a15161cb59f9ffb5384fcaf84ff74383b9cb0b631dff24a28c544f70c64baca90ef43e067e9ecb399ab3e4cb93807dcb9c0de885d0ebc1f0e1f78fc61f3eb2062cedf8cbd7c991025346154ceb822489ceccb3a9d3ca42b72bf375819bf72;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ae21c9d6f446a39b6a752fd902778d6826b2d5239aa0c011a52768dc7b177ad1d3970ecf5d4996f6dca6b1d5fa9b59c46ff456f657540ed41bdd2f5a1a4c08dc5638222ac108e4a2d8e9caa83dc82319c03ccc4ad77cb2a1a0fa1523ea1f3c70ccba2badea903d87e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h135a3ec688e660334fdf9a80c8b898c56f275137e6c109364c518c1411f6261d9b4bb6af7315bef9c9c7d614e639fad3fdc5d65090b9cf58317c000e1f9833d2cc5dd7b11e3a105b8665eee2ce60e2caab3abd18185f2368e21e15c2c1d4920bb82a845fc85a5f7f005;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b60ebbc434f8d01e8ffbb9bad41f8dabd726d6d91c70775b8ee421c7c7d0502aa8f79da497b12e7244da4eafddc7eddd33a08d98294eabb87aa18f998601f9f8fdee8b95c0304d704e2a9ec889abe46a09ecd74cb58fa1b0543748b0b0c4f3f888a672612575d9adb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h351e3bd78b071eb04cd3b628448716f356fc3902d79283625aa851efb01da030db4db6d965c762a826b71d96e25a6c53e43677e6cdbb36fa9e8fd1958f166f183ae2c67d910d928b9ac2ea38517d4254419f249d30b06024d77263d836abcfdb210bf8362ce689a81a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4fe2436defa770e03accaa736dcb4c0757f63927ba5a7b5e9d9ee34dfc93e3e58e9e919066222f9d3c49630d9428a3948b823d4583288a87201d54f76caa3a6b04c6e68c97c9e1d0c1ff2c1ed96e0dda82e000b1a43ac2f57a09b7165ca0d54427a983b5c5932c43aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc835a7a3f988454011316838b3eea98902b07ca2ba4be1b4853265cc3f8ba9a433f86f3377680a57fe38369d418d3890d475e4b830c5ec31a3d2d7545bffec85224b4caec5dc5b8f526a0db9fc88195ed0657913e3523a44cc72567beff4e0013ac9015144876e7246;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4c35e2523e6f1d048c8af9eeed6925716dfc1bafed5c49ba07687bdbaf8994e4027e358f421a261b2c5343da99aa8bce48248510c0e4377f8f60bcfb0337aa64a1ffd3e40582ec63387baeadc6cbda34a5bf1dd93ef7f59e66dd897fcd401474e2b290f399788d3f5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc51473523f62056d5c97265f5a6cde91406d6428f6885e114f5f1c69a40f74444daf68cd475edd1ac3bc78312f1a6e6bdd13b72bb0e4ba63f7686e1d9247beb6d45697e75546ac7a107caf3d2b162eebd82cc51489460f3687f1a99ab7464c5838691a7be2c854cff4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15daee3de466d555f07499cebbc4c8c3e3d7dee11749f4425cbd80dc4c86810c633743e579202159a2591b9d97839825ffb0ebff0bf3af0e647e5bc7d4c99eee87b0b069b05aaa9d962f764ac22bba18ab62a6a1c88f8dd7a4d1430e1049943260dd3663391c73ccaa4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hffc6b494ff7571b5df9da4114f9ef278c57442797188075a4be37f027f456aedc718b61d8f9d4d1972fc628e5c0ebc34627dc3bae33813acb500d9ba53563f75bbe1b2db058f96d6a11211a12f49ea5a7029bd8b68eb36fae6e0a169669fd56d925ae64fddc50b580;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h324e57fd06de85eeae4efecf740081fe648b3996307295963ae995cccec8dc8a0fe95a109d4485f5ccc7501fa7c1885a8c42f5fb80045fd8063989eaf5f248e896a676504520aef73be8acf5be5056fa73913ebd38c17673c608f0599c2a78ebc80b1c2b253688408;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7997a2fdf56885f9e3a1290d57c00aa363f8f168ecac33b3bf6a3312fdb0e9716429cf8a24dcb2dbccdaed3f5588d26608a090e347234cb614d17b421d521528a1d360328bf321324d7ad92ac27bc5a7bac90102f956a457acc96231afee64bd0fcd7c975f8b63082c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14b3edfc2a51d0581a065af6ab3de71b872559fdba377cf4b34a2230aaa9b47d1492c63e1eb7c337bade7753d47975ebf0ab1a98d7daca5ad36c6f62f45dee308c92877edf0b7e455cbe317f6cc11849d588deb8ec99206febc8b4e4176e8060ec172d10665e9247d4b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc85fded50732c5625d6f596b2de870c1033b2af2656048b878a0bde70beb3f599bbf844df4a2f6a91f32995988e2e83609320572ef0a17c01f0c1b2c9d62f7a33f2191a6eab234f1128edefe3361bae26d86661bfd69cfc24fe0967b5dfb22599e03b610dc34fb1d5f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hffcb3dd12181d3ad83571e12a9de2f585cd7f6c6db18094c403bc6ea8d304e180815d552c5129da313c52156c06cb3091e70d871b2d02c5565b35a765384872a47cdfbb3daf0e9ac162339ab8ffd377bb8350fc28e06582d349061afee737b8db36278e80ca26f4f23;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fa136baa884c1ca2eaa7e96c469ae5d9ead089bf58797f041e892f96a11a44c4fbbac0d9b9737754235fb89d3d709e72cf5b24024f1b57e488f8bac0ecbe6bdd0453fb191802161883b65cfa5ae50eb0f73c7d402593bb3f5581dfeaf96b6b3fc010afd5858e62245b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1225ad0c52e4d5a128025ca51e708b8f383b28de21e7239355a7e2d5326180c2e2e4e23dcd12ea2795a3c9de927ab2ec5fac4fdb8287ecbdef13116dfe7d5bb1705ec0da21823bcdb87e2bc66a54b454513ec4f86c6adfbcf30f9fe4f86194e6f72ca0cf53d59106eee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hda4db8d62126034019c8191d7a4397a41ecaf4f008912b73c2315d43cdfd93c7db8b8d7eb0b6580a5f889a2c60baa39132c8f12aa6da888f1c1da63b5a099d7c1cb232974a71aef96cdfcacf17ddb5f4d31c4241cb81729eb73c2430afe4aae3b98a8af8423795ddbc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67e636744279e444f3e7322ad8e33c408ffbee5a31483324e75c7c8faee8258652787ca75fa53188e855ca645a79fe5c8bf24786efce574e3d41203f6b8352fce901811fde71b674e8ae1a65d6e71ccb4c99d766dfe150dab150362e481b7899477a37e21a16d8514a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h55fd70bbc137dcc6bbd5c93c25163ff09395fdf207d72ddbf643f4681aa245e28cb049b215c049f3b3919e18982f05319e5f223c0784cc53feb919763ba3ea76965840f64d108a2da4a52adc49fb7406a5cca4b88d074a6945945213e13d58fef50fe3dfd0f62a3ec8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ea50967f96985ab9c4fd53fd5e173d550f352c2cb9f43278183868e5973b1ef24dede925f0a4a3f90a4559fbb7c3b33b1c0350073544045f02cf215bc80c8a68cf1e2adf11ce1c565f07d65da6c72195f74b6832bcdbba68b6b4040c0e3bfb74ff1c3857dd83471aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63c999a1eaaeb2b96c0cec12e8dbcb18f492353fb630944218c321dd8963442a4c683afdf8c5401267eb509ce708f9a00d3262f61a5ae2a0167172267d8c236548274cab2319efdd56a40355997396dc2352621fd35be828ab9a52a42704ae456e31b1cf9830875bae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h172aa91a590a88228265d3016e79db6523dbe9acca2d0013c455f1eb2d9b315479502a007ad2d5ee7a74bea2b4c83b460e9947ba7863780b3da82af2744f1f617122922eafee6c1e41d4f8d6b1eb6f1a1277c94029ca77569067317fb64f6799bbe69b838c113cbcb73;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2970553869d5c6531996222851629f55c92989972ce924388edfff34ae73bdc0adc071a658b41d0f0b5704c5fac010b52a64c9658cf5a52e607b19341104725496a6486a3bc521a9ef6c7fb2771171bd83d5a66d1c2bae43958351564fce8be38f166b11082effb2ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd78f5a8bdd7c13aa1bb4e1074a299ec62ee3cf11e609c97b1479364f9dbcb762d9001784aa32ed8a16d4b0eb953d4f46a7a6cc5143f83f873fb2a809840882ed1d976268ddbf8190f1975d3dcef06bdd862c12d1ce46512cac0adbdca672a986f5f3d4d6d9ca8d6317;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd35c415bc33cb5d4578cb8f85d3f7a3a6b6aff8c9a1a1231c492a34e74af802a3533efa9ecd3b57bbb6aa2a9c57edd35faa1bb061362039598b97656133266f89c9049ef04afcfca29ca95dd8ed004ee3c92e8416d0752629acabfa59f3bcffc7a1f832b00f6e61b4f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fbf2d21f3f017e8c2f01cf38f17b20ebcbc4f11d587c94b5451f323ca9da630dc92e00ec50fd567a4a699a132baad3a188fc227b1ae5dd0c1abd05aba075bdbfcea86ec4f43dba296aa6db7d096f305ab233e56c56742912600f5ff939cdc9019bfdb3a8cff5cb2c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfb2615b313499683d9faae5e67e9fb6fb597f2fa2d926319a4de08051690aae2a34258769dd64266f555d64b2674eaac0f52fcb6cf17c9f0b72cb2235cc631341a052088b7427981bf26eebf823bdfa3a5b1d37fb0466feee337c03a60f27bac57c814a5f3913c5003;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d10a73930f4d4b64dfcaa73043400e578900a5cbe3425527a4a530ad973c2260777c2c513c9ce628514b84ea3037d0487f442cce79687c883f9d6874c15ea5e6986d1192d30ebb0bdcbeef06fd5268849646a428eec4d834279da38487771a4041551dfa2e7ed19e8a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h147142d61d7df0c18638545ce1e48bbd3e62bd4a1625eb22bd6b854c59d342e868d2ccc08a7af422ee7111d78759ad8220ad08d30433e9fd6e3152e9b5c1cab091bb3073e5bd9dc476736f9627afeed32b504d14945abe7aea11f567318ff01a21fb26b8c43e7e5dbf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c99d7de75556d871241a1c273af34f263cc62fb6f54bb518a14def306c0d85a4b97c5b2fb8e20686615b2d4d685e66c625f6d82421e42b56cd74c936bc4314abc8a4650d2eb7e09007db81fa581bb55084e95c39eda870333dd22b2a35b4676cf1209337997f53d43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e4c99ec333739d857711e016375426dcfc33ce13e789816e2296673de3ccfa2ece8b095531e8289df36cbb3d61f96aa7963d7dfb9fb96679875fe858e900ea97ced12ef1bce3d9715e869b556576c04dc948d2d57ad6e0ffdf194d7574e1d015cdb1a6a3e5abcf6e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc18253edb50f5f61fabefa3a88f6fcb8e74ccb25d1a46f5bdc286eec06ab73ba184a5478f14f619bf2744c41ba6383d3a6e14ffd279b0b0f5529a31e5b0cde312c4978b2eca881bfca16bc2a8d74866b48a42cd4f3a4938fdbf244d872ecdfa892e449c50122d70e1c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hca1a74ddf05c494d7312e0b39ab16a343def8bd674934b5ec07593b4c0b0a6fdd4defe93481edb56c8633e6eb38ff3183ce14bc09d7f2bd67f45c5b6540d85f26605e1a24438a5fc8931d83c18b8de0fd6834ca77868fc2e3b42a22e6abec6a80c7ebcae8ea01d62da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1776827121eb61d43c48babf59d54b87231e1f8ce9ac0c9fc2d704ae5f51c5ed87971e46cba99508faec4e4a008c2e108574c694ae408783f42ba1239b913468fabc866f7b135c4e0a6a0ef1e5826843bfe52e576f88d19691e3dcd175f048ee4e263db142ddbc20ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb40fcdd8cdce08986694d055ac9bac6d5908a2ea716c5f7c8398d69324fee33ff9d2825bf1addb799fa39e3d87ee56113ec772ee4c8a0cfcbc70c37e496192c31fd57f551def7cb29039c7e0a5ea1532bd9021d28831e3d5f1d60d80deaa96442778b1fa2a40ca1217;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h876ba9410167d7d5da7c31278854f63fca58f81af4180d1383df5906d46c2e22534dbcac7c250900f888b97ea99543008ca9eb102847c4bd1f1b9994620a7b11149352545bbd1bc8191e0dab13166e47cfa79259acad8934a979d35c2d5050e1dda73adda6e57f215;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4b0bc6d70739fe2f05a89665bb394f60b3c403527b6d45744efb12d2bad0a7f16a79ecca44201a8ab3972354e507783a2546bdb795fe7d9bc6407ef4cf2478c2228850759e22f72a76e48c58c1cb33d508aee1a925622c6b00151f1e9f53338d07f42c7cd4de5c8b76;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h74b60a224d9fe96ed19c7fa27042fd0f6de0486319f7baca3854e479d1c5b7f413aa7ca5ad96aa57c27786e89b8af81f15f51ead96ca448dd64d7b7ba8ccc776ff8316d67c5bb7bdd865d20c56fbd61705104e79fc029a81b694cc28dd0f000f42b5a2c6dc2772e861;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ce6663ebd031101b2e6b2b1301a30e804ab59138060d87a949fd302cafcfae6951f191a5c6c93710f1c9a0ca4baad694bca652462c8e9f23e8704684aa39ea5bc08d29cf0ff5b1378b6c32fcbfe52aff72ef2b78c80ca94d13b199fc9152847e1ca8450258a074f4c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f1676b81e052e05c7092521d3d4319e4fd6e0bebfb2dbeca0f6ba6efab9226c161aa3b9f57fd79a4b7c3eb1c6789e906363889a9907aaa68c2254433d9618f61a495a807609044d4ca76926357be172c62a35f1e58a71dd8b5c2b66c81f6dc67b27758c9ab5c4efa68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e3546918770fa5b7021db6d68d4aea8a837e31d7189b7f07ff08e80f274ac3f4e8cdccba069f4a52f90dbba06c2d0e60535ca4d69c7ba4f0db41c8fb7113ae01edc14f82738fc73bd3adea3c731f5f7753f5c5dd1750d90bcbc27d8dd56c16ea05c7a92a9ae4181d87;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12caa6385e82cdd732002c68b4eaa047715a28f106e3cbe7ab90b9083ae626c7746f310d306641a5727a15fcea8168059b0fd7163e6165ad55d768976b9931ee8ff45d15224671151fd9648267fe6096cb13a2881a1d427c7bb1a39f88cea889e420e020d42a2435625;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c8820d2e92779f36a635f1ec74c9c700e27cb9a0c495f806cfa4f9abbb1ec9d6b6071b963ce0566acb3fb4ded3d2800e6caf39d7d46b4031321286b2b52cc87707580077403fdd1fed82c9f240f1e7ce195f3026bd6430710bd724d8e48bd9858c42965456f583b62d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17e7e4a68ceb714a529e953940a8e4a1e5b62712352e6ae3beb55084e88da2045fce1101a70c90ccfb07879df62121cfb12d1fb48024d8e196eb7e07c9156df8650ae7b96baa7e7b798649ba1abc11844700f9d0159b56ddfff490773f524165e14825f1b61e5f33b7f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h680432f70cb7ced09af429b35ae0849cdcc91994b45a6d3223d88a2a25668d08431cd606d45905691b90393a3815150472c0b52616b0b840dd64f95812c0b66208f0abbfec369f535993428c28f1d1735041e206d7e61b954a4a96b8ff3d21b11f71198140b9d3fb40;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h74ff31bc26715ddc4f702479da71f1ccab7195075ba8faf34b02c930865af25d0c916f8980898710abec8f436d9302a5fc650ff1b8a9c042c034fe313b397e3a98952d2622555b16d3994e8903d56411bfb40a97e921dc819cc7864b8f1727bb054e841ed604eb2e98;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7724c8519cd61a664e443157e4be115a9c3e9405f74c545b1a6c1436a51336335fd8f60e65d7802a32db5e8ca5cbba3805aa270f6fa9a1b7a2d8c27aad117005b2da9c0d5bae23a5a46517cb1b3c4aeaf9545c013c86cf81cc701dea0a9457709b9e41145a320dff0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb4d4357bef3a6e67ab698b985e40d5acd52ec37dd59a1e4ec9e111f97fcb884b5eafdbd9825f12f1027477c8b32fe2df1724a6c4797c0607eed16c1b2894cab8d3b9841076168cb54afcfb08f5cdc3745ff7f75acde316c825d43dc030c0dd4968398984ec12feb51b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1897938fe74d8d553ff66a42d4086e335c1573c0bf038ad1a29587b8c5052e7ec28de9626f53c2fbc26d4e3952f6dccd7274e4aa6c753471387e2bcde126e6cf996011114b11f785f72a060edfcef69553888a0326fd79eb92a081725b224eb14c3c34ed4af5c89547a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1435e07e593011f20d1e63f15ef850d532ac35f7437de355f6562fbb09f53d52e4bf79e2599f1f1343001af1a656c237d322a51044ed58ca7b8a5d82515e2d4acf396180b403147b07492d2833274528b546f34f492085d3d2fdeec7bf9ef3b81abbf7627dc3e23dae8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha149f098693c3f098bd483ffb6f0dc900159cc5cd00cf94d8fe74856f0aa6cdf39b74e882299623c4dd0a131d8d6a1c153ff81fa32ee257becf5a3dbbdcaa60d57dc55383c54bb5458443093cc0224bd7c9afebe356b12f2cbff2400fc2729f7e465b6c1912dc2588f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18c3bf79b378d49c38101f7b79e0d5d00715da6f3f61faf36054c60b67ea4278dd527701dfe5072006d987b9bb90580930fd0ff9bfb0d99b4616cf3e7dd6488104ef962f94eb57ad1eb08ae7d354d5183de0bc69fc847046667acda39cf9b37e25ec2867f84c2dea4b4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4137b3e7205f9a33ea35296849fc0e2f2251d85ad8d892cf02eaf80545b34e0d6ae59559c194691d4a171293f71120d54cfbe9cdf86eb9977c275c3a246d4bf3ceb074f99fe07d84c71d0056aeb73e30d5548b0ad4ce30e1ed6e76b7bbd2a46c05618703b6108031f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163a57c2aa83dc1496a598223ce7b979a57cc3eb20207da53fb3189d273ba1c95ee19f5b522144fc62abf203f34f6a9c9d0afd5cf9a5e82d9b2223bbd4e15457e1fe4180cc59b09777151b791356db01ad6c78d300af0b2725af0cc98c4449d5d50e49ebe1723fdfd97;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h193c97b13d58794b07b338b9604bd8052fe7f4349935e108e82a50f50f39cb8d8a9bd5df2d08b02905be3aa77fef55cc942a56f9a0f1dda0e5c3d9c6c83ad6b867fa5809b667ccf1e58f043e89914a6f0281fefe38171ea19d00303564aaafaddae082a6293b4daf21;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79dae6c2ffcacdb595688bb873afb613bfc77678e21f2a5c4d980b589a240a0ab0d45add72e3eaa85d48c258625b83c9085dcbcce3a54fb89c1ec7bf0f61e8085b6c8dbbf8fe2ddcf116ba22ee422df53e593f85d63e527833d1a7192e77ce28351583cbf1c3259f0f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123f893de54d34563571616f58672c74079f7331e848e78a14367bcc38b84cae06b59604615e2b888a096dd23006e13a18e263e1387fd8689e635f5b3f3749ae57ce9d9519c7a177fe7f34d1d67194bb854a3c20fdef8bc450d04543304deb9b72bdb19e841c5a1edc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h145859ae51feaecf251876afad033fc383b12ba1d1dd4c463394c7f02c150cc857e484a44e48cbc6c101d1801f11db5d374c179a057ecae1e40cc034d02319e71aab1b201e941c9a98c0fe6f7182a8d36468b9ddedfe6bd768202259d13a6ee9fd995816f318ed02250;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he11bff71236fefc0e251b3ee518295f94b81efeaf308a2d9017a85e9db22a13457bb98b1ba0213cefe99ae4b6a0dfad3277f7cd31f016451fd7ab05c2a8338ec187be4f4d34fe55e88007b889e2522a4232f9200cd26944e04569c8ff8c6e403d95d5d9b1a3cc1673b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14744780d7f0743d60797cc65699040437711d25d8cdae46abe81066ea8eccb89c1e3b9be7ed132b7bab079c909cbab11ddbec1266a7884b86deecfad26a0a89029532b850f8b255e7b7078ca24ca40ac5de71e4e88a93df70d60202a913a431b66d1dc25d9510f6636;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b2bf63336d753a20f36b00bc47c78af3e3198912956c5fcb15b1479e3fe8d738e7aa3a3bef6fb6aa91fc630abe83d2a71a28c9ce565126c8d54cbbddc9e38cfc8711b82d9bd17d2b9f01f79fd7a9f7c5de6695d18a3634471ceff6402cab145f7c589aa1d1f5159bb6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8703b08dce778f24cd43a3df45941c34a6f601904dbcc0927437572d2e85f33f5007e174ba39932630dae0f6690a9f58b5ea247e0c32518e7e97f0126be3aabd49f71cbc374cd99821e786a6c1b27b64cef03601e0cb8dcd48eebb10621fc00cd70b4f2de5f8e3f56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h26bece424a48a537277b55245fd0dbd66e3489702b7d49a7ab1ce36f13fce1f03fd2d9eda58fc1d42b375ec4e8d8b8e35f9ccdf9b2bb2e537426adecf489ceb243fbe27e1ae7c6ee8cba0cc23cea19aa2d0f94a3cef7fb575310925a49dc00b4feb4bccf84eedba146;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16d6a25becba9c54168920e20b0851fabb17830681af9a0eb31f56cdab0168a96c906da2c6ed537ea80fef6f89bd010a3f0dd2342f65e8855ae07157d0b4dca3912940954bf38cf6948720c9496c853b6a6ce689c569aa966bd75dbeaf1956babc6f798de92c83e8049;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19b1774d7524491d968c7e71d9a371e95647a5de52ef271b59f6cc92f28c22edb810b0b87787b1d09192af1f99ab780f04c651b7bdd3e34b9ed9f9b03a1ce7c5310e69005457040d38779632d3a92a00ea5cd2baa8ddc8b27afd15f899f3117910dc0a06d834a605508;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db526fdec8cb566c734eb940a8e7c6723a31f21e5083b062a7a86abd99f480fea36b0a6705846abb5102d65d126bb9857d3511661c1a5704dc3c5f73f251b0145ba22cb7b40243baaaa6b9aafed222a73fca7072f49bb07389758e102812a5a132a30d2254d0f875d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf9c0793f55837b1840d196f5af62bb703237ddfed1ed14c0dc167bea0257c3c0562d8db07b10d3f8fad63d403b12abd6e8ee18ce5310ad1243eb61e434eae9aacb46121329b47da3556845f45328514ab6d2255245e6949f1effab063a54acabc39784d89570a7e8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h128b156ba99ffdd87761f5de49c7bc12662336724a397869adf08c5b150c6ab9f9efbda4bebab01278a6ed6d8410bef0438f5e1ea0647740af165345b060dd284556f8966d4bfd4bd2a01050142a5ddf8b0587faf1390a2cba67c95632e440e6f8ed2da937e6b69ed27;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h917827a5344d9e213fbd2b3e15c8427ec1a63e8abc191a12b1b010cbb44624c355828574e69abda9fa248518af93b86594d864617178a2b8978bb2bb3cfc273b4092320ab87de8c4cd9b0719f24ad063b5b1a382b1c91e4ebac9b42ffba0a14e03810b42bec74767d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h114d4cf4a69e1d22d87556f23f0694c490644fc3598c1a37c22c5b370cff0757da896ce003855bde09c5d90036c4dd137887dd40bd2e32e9a0bbe039cb92b74fe14ca1ae20f5de0c75bca3c6b7118cd70bb69d1667ebb3956a1b1d996cce9b251d0513cb62952a869fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b544ff8cc847a147c9920cbf3ecf9caa7c9841dbc6d4ba8ad30c19e62c1f7041180720374bc54ba1521daabcb4cbc11e5e2ca27550d98258a5ff3981458c1ecaa7b887b143d63956f65881254b54b7b274a1943728c713ce73d0faa31eb77a8256fd0dabef4350348;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h166f8570422958141c335151fc72ebd3be4753a77131dc24bbe384e1fc79bf0748134077c326055e971bcb808f1e949d7fed0c9927ff929a9ad8b7d1a1c42e49426120ae4e837c8c103ce01dd44835660fdc61cf17e69bcabb5c720ce9bff8ab204383eb4c33728c5f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd8b7c5593bc301d0859986f4c1f3e23b3b7ee7368d2d27b05559599977c3b3df26afb7492057d85b61834169b4bc7e5fe54c24f4e19435749bb058245df72bba0d190e2587fb69e6d939268aa26b59a72e0e30a420e78a1c748f0903e78e00fd2841dc449222f53f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134aaff3f66414392d6269cf2cce51daba5b27a3a1c83f22f6dc8b8f7e7bf7f38d5664d526c47f658b3521faac89951e3bf721f529a519a97a98fccb46f711ec1118d45b5266b1df6ace2ea489f93d264dd67de95ae99a9db841827bf17039acb6105b51186e15c1f96;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ad41905159d2c34aaf5c7b80dc0418c6e12f773a9ca99badfc9552a1bd0eab3a01e8e22125075c73ae6719907c59d83f3c8eff621dfa66abace824170d711b1b5aae8646cf65a9108e99fc4de2aa697450573ca271d6dde0e47f8f6557d87478231553dbc829e3cdd8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1727a6d7a8ba89ce01b069c0c52736f28bbbc9105aa8ebc0007a15122e603a83d1055f821304b0c110521a86152f56f8792ac87cdc7aa83de813691a0878e9046e62c462435e7c85f423a6c893fcd77bf7f38dae51fdf690d92d881421c35f84cb955623efb76ebb73f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e990983daafcdf7851ceae93157acb174bcbdc89470c062eca88865f2b6aaf0adac3f7065c1c5522b055b446ff8f7d8417aeda883811f05ceba9b27b6aea7ebc311439474aed10652a0804e6adfbac0cd012eec4edc7f99500db6899cc060d5088755b451a10dcd2b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae09e5ec7559c2a71533a2aea8d4b6b3da9ece6c7436c29340f33c764aa19f362e3fecdf4d2af7703e084328612cd043f35d1daa880b7b009f8a11b2223178fdee6ef91527c3168a2e176d22f7fcb509c7e52e0710735f76c3d951302d68190c3a506853aa0f373b3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5a86ace7d85c216550502c2d9c765ed202e38bb7809446b4dec5695041e39cad74838d25699f61c9a96ae86584092fee7aceada66ac1578239304f4d163b9ef47a2866c07950d3c81d82e73e5aeca3ca75c572503db8461ae254f84299ba38f01b67871f3eac6218c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5405667ba8f3c3ae9aa96f2dcff242e164b57e950589e7cf16381544bf70a833fdeb9ce8e6f11686a86c66b46ac3803435bb6f1bfb23d18831493924d7b3f9045629e9a487cd073556068d300887c8eb689f4d98c9bbdff803c008d98a2554a8af2fb9899bb8b9054;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f99ca0ed30cc53a3dcd014acd53790b9027baf2f90c768b9a5fe3a96ea752bd356ad807381fd5c60e4895eb2ea509bbca874df910855ecb0cfc8661b7d0b0d6d667c52feb809c2dc8f75bb3c893353762cc9b9538cdd74f5ee496a0acc01c622040a38280ab524817b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27833f1ecc1993764ef4a6dabd6c13be71f7f74b431508ac5434fc53aa2c03e153bbae9192d164683a022c7b8cc00536b0e0e1ea7bc0357c3209ca7453bac163acae99030237ed1fecd351eb7dd2cea06094f8d98770958771dc01c62e0f13205f1c7d232b504338a3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e44fedf229bb484b1df48c72c967675ff7b7110a70918350797941a60d8798f40a85659afbbe0ee40f0ea86c95d357d52d9dd22a5f35f4f4c372c7e3c34d507c799edd75f350dcbaf5951cb1d2c619087cb584bb3ce5d39102ee72b58080d772bd0cda2b19bd1d665;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h236188e161ca116babf1f0ee0a6448862e6a751d5cf46991c627161b0180ae50a188e3e896c68f2df207913f934dab92681dbbd2032b18fbad4bfc5c2a3db521c30a69209f3c6ec563e81885a37f703a0138ceb5ac4f5a45b9a1d2ea03d3cbb17605c591addf449daa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ee10277bdbbc601fed1d5ba682a04b8d7346c48caa22e524e6cde175d218dc4db7082e15a1e176d0d7b3c3235c9c169b8cc51223bfb7f98e69900e368faa553dad9ba808a9073fb6c89b152d0f0c8d75cb577abcdc9a037c0a71b25a9b5face7aaff44a7e4dee25fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14b0039891f56acfdc77f3400488c44dfe08da3571bf5a9c6b20536d33a1449c175ab847eca86fe4009ff0bd612d52d7b1f67cc8caec1e5cf608476f9b55a22029d78eaa9a5f188333bf66c25ac119d7db50ae2ce3625c3d3fcf0bf133080823f5c965c034441410c31;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9faef6aadd26e3580057662b82c1fa18abb95fe541c172c8ecdab85cf4ecd2463abc108922be77bae333d95f193b943d973cce9a09378b21209f0e407c9786977f273e12aeabea92313cf117a38f51c6305f531d37be01be47198357e10a4cd2c46290b6207029d04b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc92b09fe0d93718871ed3a96852e49ab2da1a682e0235003ff72002a5a7f9ee15b7020af59bf443e3dcfe86f99c90d7bad3f082915222ffb3585b2b465aa48a8a635cc39dc632a91084da1ec3190735d0e4cc440e9be15fcde48800f31c325ff9872745b9e85d36c0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5feda0da71460c811e788c23a702334e126c509866206732eac083691b262ac1c5856927faf4699c3e29d67506df96b0aaec4b770afa957a6b8fc7a32caa777ed04873ae257e48cd4da94e1ba84d5a9fa35a681d2f5fda39b28efbf150d758c0c20a19e7b1abccc862;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf1fd0d68ab3880203d77caea4eca23adbcb63b7571ec5f7c9cf7c48b4def3ef89adb318ae95fe183ffcc2fde620690f21ae8bdc4149c5427d05de4b98c2035ad872f65230ea52001299fa22fc68112118449ff7c37c659c90144d44810a7a631df19c3dcbd103d392;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he94e551c64091b8052ed2b7ee60e0de1cbd2f466833bcb4e8abd443bc748780891ef2db3c383f35647204741c4d6acf0c5e7f9022b72d5ee4837ecf9123e768322fcd9dbf9ebed563691181c252dc0d6360c24ba6c130a97e916c767252887677d85814e8094b27d03;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b68e7b2f797a19fbb3c7dbf181e7274d162e65d0ee41297e4b0513ab230d976bdebaf2d1fce7f4b7b329492e5a6a40d7402704197a2c73e4c68b25530ff5e198d52b1504b0bc70914b1cfa821dab74c840fdb01f2680dc48ec16f2a51745767ccb34426a5f0c327c1c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b788185c42b05474700ecc8685278e04d56880c70e5624308bd26d1dba3653e9d7a78637a3af5a7ba02b5a12d800c58092c44b2451776c18ea42c5568c29381afb4a52a271db90f960121bf2f68e509375d707124fc70d9c8770872930c668db93380777a7a175e00;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c2a08ed19cdb46637f03216fe30e66a572c6f1ac67d704bb223bbc9efe268d1116e0f6c66d13a85e655c9847aa293d17304e97fb9a83a6b3e36139e876250342ee8323024d06be28774a16f0224e8d8a57a73f836ab641885b2ee0d166faa58950c238a6324b5e3fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c0c0da1d77b45242d60ffaadee315bf45f21824c1f2d077e413222a442021f0ef8fb58df2bf5fe7d9736c866b34c3e3f60b8fe0f2345b067af10306151f86532f12b0faa9dd403cf53501b311d4066d1e5a14e3390eafd3561ddbcb2d4af82b6e24b4799efc5b1187c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee13291df59ea2288aab840a8a9e13719facee7210e144d9e3f87f2015a734cdd7d5ef03f4ffb630542d28957b1464f7394f4cf192ffda3abd580e890df7ab231fe97c49dde4a3b18efcf8bf95e6f3b4abdf5a5218113a6fc6f65c35e97862f0005f3976c19c0c3a41;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ea89628702ea7ca74ebf5476b6a7888d14fdc4aeda12f1203c4ec0109978ee1ca4775a79ba4e4838e0874cc2ae9ddf36d66b44cf098a35de7f90457102277414cf1b52def6e5117a30ebe0490816e1a16479b7a93035811a8d9f78faa11da1bb87dbb00998230852;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h580cccd1f899ac065d7de0c9b05598f52afff8c7f2f7bde2b6c06a90dacf5254b9d86cd2995fc0490a7ee9c3305583363acef8d0a366ce3b0bb8bc72cfe33cc038faba2a8d9152e2329700eb2986ccc9bd96bd135ef4cbf9db7edab67a5fb241b178a1a57d0c95a6c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b5062b10b8aa6d0c084b665a047d5773430bdf3faa88435fbbdef6fbfdae56db51f160bff926692041ea6c85fdae16b52872c6d204a3389c6d8c7fd9a6425802008953c269fe05ab02cd403df9fef523735246b7e84091bb49d3eb44fa4c57953ee907f26923b285fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h151e30dfdc4c9db62bb1475070276fffb216820620b3d4f12ad6d28387fe5c81b9fed5d9f23a6c8c4faadfb2280e3a329cb27c12d4076191a5840d83051188a368813da462eec65e97f111477b5ff18eb801d47f3405b21c2f22ed34c0df7b0723948e296c99296ab93;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1f3a3a188dd383f90b855b085ce37f31770172334122a9e678cbdb3be7c983f24badb7404560fc4a1527b6d13fde4cde5f7aa3ae385cc7fabc656e89de57b49611df58f36338058f8a1974094e67d69a6345284c89a4a2de3b9817a789559610d318f624e6a52ccc2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f521e7886995e46524c03d5b175375288f28db38f98bbc6394c75db706e77ff393869a6401a9f2368f6030c4437af5aa06af75956ac65750619b269d07e8ce37a88558201208e5345e4043fa5b6f89b4169a8674b85086e01d3825a93cba693bf776931595f4eac86;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16874e5d0b558df36553e6dbe6aa9ad9eba258863f41b64de1ae37844a497feb1ffde0c72cb1f24b5c3a972430326d92fcfa697b4bf1c48e906215a65c51354671560a35c4145c15341681adab82eda93ec1e5d45c2c58a487e9bcb34ba4e773e0c3dacaf34245ab7f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3c236412518413eb7a4e656c2a63bcd6345a59732cb0e8e6596cd9a2ff8371ac3689bba9d7c40aa9d9b283005326e2b15031d330e4ba30097dabf63d902a9d81071bd78eb898db355100691bade6756de6ee2cb3764cce1f864be9455e83e5cebf622048b8d068ddf4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18de9fc3e3c04674bff9ff6b35434a99816734f84ef82853a4a94a886bb025b1e46fc0909748e64714f5b65d95d372a48180a2c317a7afe59018a245c73068473a846f2955499b05bb77af095bc9c90fbb6d972882f2474180d3b24d01bf0cda2efd74365c7a4c1e76d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1302019f4506cd0e3fb9a70b83ddb05ac0fac9350555ca7e283e29479144e17eb9caa1a3e0664f3feb33264b3cfbad6b14ddafa769aa15deb1f7a15938479212702888b9437da7172f4ddf75b3037966c5d9ee4031acf3750316c5927eba93780ce295ef862b3f7ba9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fc0b59baebbb049120ead7d912bf088bef4c41a54f02eab0c89b8a75b82856653af9481e8279711ed3e1238eb52fb7f12e532ff8b4f2c6a44ad74d869aae8addb862a7238fb51603baaeb0321aadac0b6795009fc1fc1917420b985235504d3198b9bcf61a2332cf40;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e1c0952933a8e1c20536881cd6b262ce53d2626fe15b948a0ba012453f8cc4bd2933da8119f836937fa8e65f73398452667b87640c7b6c8e960ab6c8f5de68b50cb6255a63fc418f94f0fd35d794645466cbc4318e58363f3c6c3d63fff73c48b25f2aa19870df4857;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c1d7812eebda4570971bfa7df66d1fb50f29a3ec52cc64c53030b6b07c3a4d0062492766aac2c14d91a9faa95d76c3a4ddc48fe02a9d02e96b856ef5ccddac0e1bcef366026cb8285696a2a5c328cda3571614c5c68d6a502b803843cbf7bcc1bf4b911ba8462091d1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c0ea28699724b723cd886db22edd57f357ba3b35ebe46a939a7a975ce58a3c1c8b4bdc0ed4ae4c710d126baf8a6884a5204990348f43c54ee92072843f9d936c3272de3366782c2e38e24ff554f412644d2c6add71c40797e9e13b34d3902fe88b1a12da2a1fe152cb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8bf3d062f8309d3697dd9cb35d9e82b2dfcc9c6cae2bfdeca66e0a2f0edfee08e92f3907f43e96803ce7cdafef77766e28a4782566949618cc3773df3c49d351f3b52041af8b2da1a7d97776b4e5e94529b4d16c9076d74ffc30fec6ffd92411028cfd78f5472a325c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1785b2f74cda0cf435a6df978eb67bf52c88b326c52822147e34a5df683e80293f941ea9c836d3b447f7aec81070f62b50db3ad751224522a999dc852be73e540a621bbcd224c3e28b260f61f3d332c0457c1952836810206df1ec6cabdef15ff08ccc02f43010956c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e3450f9d2fa69b7c9753c1b01ed46ac51d0b8b71ecb18230e42eedec764188aea7ced5d8584b1ae986bc8abaafa70bb6d683e79e759f3ea8ea97f7ccc7901ebee67ff000f2d378eddd83c1c55203a9ad2c6c5b39de0859c0256c013d27c2a42edcc52d9916a84b791;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62a7b7f34b7a4789904153bde76191894c6204fe2756733f9161d6f5c655943a7985cc03fdda553552a77d29cd35ca1674900ebd63b561e7dfc40f46213b01a85d7fd86764f99db942284aa15e995b48772bcddcb58f66bb95efb3f7bafe1c7e8b0d75631fa663c28c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96576d4afb75b38b49c2e8f7f582cfd329e85ffb5951875f2bad3007be69b7b2075f162d6b33a3e6f59af62b680c28c7628a96a3eff1dd674e1d3ca102b381d1a8265ae6533a8d89626bec158534e5b301caf93d4b749a03461ee31719cc139c8a9941646df2b04ad7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha3beddfbb7efe496398258ccaf3a97249708ebd529433796743c29f83e5dc664aee8db3cccc6bd1cffe8b7c14a51db601e55793ab074d0b651bfcacdff91a312ace96486ab8bbfe2a666c5ad0cb81c9a330774eff701a0f74c3338c45fb193d6c91805b933814128af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d63e4fb3ca0dc8d5a226822d74f73ea6d37114f26093c8e6ea62db464abacfc99f3492b5dc9a876bc547ac483541b4543d34a02bd4527c7e16d3cd748253bd374d50b019f87173e6ba3baa2d74d868f7b4765503b0e99f4cde5ead31e06f04a6e0b6cddb03157d16e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb358f4ca2ce80aa5d5046199da6326b1039657b5484188d2453a50313959eccc7543bfd0070fda904a926ece8805db9be8ebcffaa94fb1b37bf2f9e3eba3c7f09e2a3ba616711e60bfab13569264857defbc59d0c6dbc11ec811cedb5457be7e43b4412a9102030e90;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d79f84268e2d75d3254a61e563c0b3f3cab77e0d8017da08182b758811d7dcb5d740e790927a7391adc1553122fb2a357a72cce07e93043629204e4961c60ec3f99db7b0e61cd5dc0c731f73315efd707aa11b84cbb53a22af582af185d36945e1166c3c2ecf3e32a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1250b32958e17cad6cfee66dc8a0a1013f1f8d13a4c27204d54a9901d1f4f581a4b450f8ce5afa96cb8959c575eeffccb9ca313ecd982bd10d1cc31f3bc6d71a503c3908b19a698afa1ee4e1e692201c9c3adbcf1602aaa27ebe52785809b1bde5589d55bcc23b935cb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2e407b4a84b33f843536d7981c79bfa23a92cded065c210a5b26089f92cd48dac9a8b27ae208b0685f083442d6c521f251e9a96827b75d155844f5fe2832e8dadbad5bd9ca95fe3ee8ae15696264feaf5d4e72b270c2f8c4951a642a847b0c178c6764c3824d39e511;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he0cf970c887ae305117c18704b901e2dd5ccfbb1a62e1bfea7449aa757496a0ecbab297f98df9b383ad9e08a3b39f22126f2949b532c6eccf2a98f168a69aff293e109671a38ebf6a64d46ffffba57fa26646bf8fe47bac6d0ed9abfbc29c78a555e4a957e69ac1b54;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b184d0b00680bd3809c65e6e00b8f26c38b578aabadae6410006943274dc135e3f8887079d9d04f6abf608c11313cc676e4cc75204938cbeb318804d7777e60d676e368791902585cfb79ec893940ea0251bf068c15158fc8e09315200b3f18829e2ae525c7a76c6b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f74f6dfb6c380ce3b0bb9e8131840dd8bc44314490b36020acaa1f80c649f2b3ef83c9e72dfbc36bbc36dc0933b4edd22317790ea16b174c43dc51189d65eb22140625d2a7ebb44f4e27f1d621441a9a4e0362ed2e19c42443a7e2a1d0fce5c51c6017f0617e3bab59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13d7b75351fdd4315488c26e7a3f76f80010d6a88389b7f94d404f7dbcae0f7ac4475715bb465eb76ed9c8ae24c1cd1332166fcbfb1240698a056ad0bc8ba4f8c483aaac4a32476b523a65ef9597be736ea7081ebdae4d5ad3511b63994e903d32b875f71cc47ef0697;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9603275a0c08d89d708e1a259d817f623367cdb2cc1038420ffec35c4fb3d54cf435eef73df453d4a3d97007e49f42675740d57aba45eb1b176a0467b5462e7a46f0649cab4b06343adb85fc9048675b85cb43de6b4e0f1ee14ba9d9cf01f029ef6d21976fb9df4a59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f44f3a5bcaef7dfc67b15e086ebf9a519d2807c860b2fa93a46f7bb9f4ba6b8654537d724fd909636a4bf39a1dcb7478e888a855f6e04fc31a1c50d219a86087faf45e3c9c5b63e4abc6fa6e44957422a7d601167e9cb39096ea39ea454be5b1663da20e4e14526c40;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc6e20087369a3d89c1ef48a98e649f8182521cef25c95eb7f7bbf2f2d68ce33ec9c39e7ffe2868910aa533f3e268ebeef3077e5411ba7c3fa48ed049ed1c3fe3df5a212204008b113ec93085c242813071a9e81f0dbb17993e8148b731831a18752e6beff7236ac38;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he641f17a5b293a543cb3e99dbf8fd55ba47f89ca434973b8c577395bcbc62a5ff940becde5a306aedbd902ca55ab1d04836e0ce7923eee93efd3ccaf1936894f0a949f8748488b453d42b5889cf7584e4a9158a1391433d621f6316a418025c28ca578d968d3f270c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4855bebb6333142a5f64da070d5b98698af272a45ec1f07db2ace9a7c3588ac386438269335ba7ad10f8ef6bc2de5deeedb4dc374d05da87635dfacd929aa297f929e3e66983b48747999ea65b5c15b39cd28047debe7f426d5762ca71f17c2d4645d1d54f978e02c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h193f3b58f9ea51ab7afbd682eee71b9e30285cceb1e1724781aef7c0a63ce2720ef8fdbf34517e9c5043ea574da1d8b35b922fa602ff1d52cf1c6a5078ff92705b861b469c6e8e4d1eda3d73f021a594366a49347a9de94ba5b911050c3653b400bd0840a5df6fb96fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc67d7f7782fe0f22bfbbee4760f64172ee9536ac2460a65b8d2d6e4177b84feefa6f3b11c8cc656c0a02592715a5bfe477e112bdb49bf17e7c22177608066a4215a6988accc03396df00cdf9fb3827017e5ffcb000ad497c6b2242b2cc0664783d280f20a9681a9cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19907b4b8e8378cddf2284f4fbdb2a65c0948c5c238a0ad972533b6b97deb3e006dc231163d5d887c2024a92d2791e911837feb8944fad7cf6a0cc39ddab04ddcb7b20068bcbcd323097dc9e8594a406d4b5f2d1c77184a35b4515e1e62b62ff82a229b1b797a6dd0f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2b99d98773e31cb7226a5d8d8999111947b8f5ff33a12722d9e36badf59da123edd3cdd2e82700f76ab57f9702253e76b8158c84f81a1d0ba6f7f5e866d1273147a2a9445e04511e39d3ffee66c98e2d8e34b608eebf8cd6f955f609256386c60cbe4cb9cf07add2f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba2bad35f140bb9b15d66687ff1237e75adfc701aadfa05e95f17270e56aa31edb62c99fa1bb4ab59790b0095f22941cb63db93c38c413b22a0b1932ef218ae6a56452da6c21b9ea8d95df7326e1cb01dde0acbc7233d8e3b8889055c6ddcd1f804f7caf7fbc98f4f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e59dee5464cf12d5131d3e13dc1bf1df8f682b589fd11b7a72d71bc7d22ab30f694f55d7a6311a44d76ec2d324856ec5934fdd952bd5caeed10a60e21fcf45514360287c195b88dce1b90a7d295d4425b93cd5fc07bfd74794746ab5ce17905dfc8a626e0784820855;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a03a56352b11eed57202ed66eae6dfbb086f0fbe82ee49e589694a038162339679d48c368c16975225b7e052e8c46cae47dd1d990f3d37e8c5c6aa251d847fc2a7240ba410d3975971d6c92d2925407d7f353a6a57ffb29fde196be3e691c4afbcb442ba44203b1e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183d2828ae22982bc4565787228c8d678da5802fa47d1f7d6c4441682ad6b56073acd8fe819796fa7aa988757a090257455df3eb80cbaa28558568523143489895ed943b0dceb9913ef740a9fda0cbde9dca5a9be491e565e362bbace72777a40b2cedf3a4020a238f7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b5c9628af95af8a0042672e127c86d549b410f714efa913fc3b87ea1af8fd2b9f6e39992dd06d358817a54e7e33966488526e548a9658281680ae2f2bfbd53bd7d4fa88fb0b786a229ce5bddd7246ad4a96077f1133a6fa7c2aec3317f01cbe656d198787d16bf926e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1933fe5eee6a7da7b51f07f168143356e036b7d87e9b15bb83d5fff0188448ec26c5b58fa2be5e15d3a8e7dd1c3b511d9c95126fc58b72388eeff98bf4146dff847e8a8ce58b9b98ff2ceb24de9adeaa5bb80296335c18a930b3457e1742871abbe2a968a8ba3870e8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b03f3bf537a323405325c2e192916ff03b1e041045e0df361ac4543e38ec6613df3b68aa9f3be30508a62e26025590ee747962a5e9b0c07dc364e0c3aaccd1138a5c96f189e4fee1c17ada87d432336f08cb3916a420867ebe58da126d8bd78905858e50f9d54bdf3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1970c01a5c8be7613a132d60eedb48199bbecfb657ead107b531531912594c8f31fb6e1e4be67f13ee2197e4e41b9e28caeb993f23759ade63dc16a0784e39dc8714dc73dd40518165a7e33a5d6f92bf1511ddbfab6244ef03e35104604caa2a15db30d171fd9230ad5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb17cd71dae730f378318c70d445964f7d54d24ba18ee00366b4696df158747539c73ca57ea747c9652abd1c77a3aee7f226c91f139e57afe95741b6373cb737146ee4a50f1ff04e3260c3650c0ea6585e1040902ea72fa61590fe0d520a24aad72fdf0540f31488d6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1322b5c89fd828cc16422c5c2e26011600ac713cb4181ebf25bfdcab934c584e057ce3ea1cf30d39d7cd7d53e30e850080d514e9b9a59d2113412b95fff45eedc68a3f651dbb2597cde5060385cb67b7d67af3c0050e64667bb2ce11a14b02ebc76b7f4cb3cdb34d0d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8fbbaf34e8c75baad1eddbadc5f8bf6bfdc6f94e3a9505ea36ef880387af42cafc247256bb1fef276e10d018933bcb7e8e38117dd1481a425f79ce5a63e563e5e0b1239552e3e4637fad8e4caa8a5679e231ef1373f9ac6f2dfb8397643b0745b5a3842a3d51febb33;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2f1414f5023b2f515ab170b7a93253439d38223cf2ff854af2ca483799b6cc81a300c55e37fef6d239774c8cae0eef5cefb36651d809358e137592cc64db2e67bbb2ce4406a48c792d79e12db8969b687201368cb393281b0a97c8f9d813712d14f295f6dfa23971;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bf525d2f3ff8df44c6cdb3719b8625e223faea54e0cbe364b584bfc02831668b8a776b5545fc25e8207907b8a141ccd79cbb19f16ca3b4e88a3ee18e3c6b1add87894cabf9385aa7139b66dfedfbc272b25d5e0eab755145c2a7b7f400e4d244f1f8d8e681c86a9f2b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb98436d89d1a49258019318a54434f8645a1d17bb51336a96a6492d9f561f9f5f14ebce19311244efb5eccea931c0ca2933f9be7573b5ff60c4f58a431d249ca18399a58c55fc1be8615ef75d4733904cc829d57f7d8c271ad97d1c6617b2cf1cb24889551fd088cae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a57aa3facbc25f7ea15a457eb72fc43c7ae374515be9583a85fa1c452916b7bfcb436bc5dbea80c2c8ca6383544e004d4f9649c56f9079fc87144a6cdea4890f7328e58decf872e0cab3d8215f5827208f3172647a1525299c081e365bdb457e7575388a5ecead085e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha90bd962661d7f1616b1cb02aa5802b68cbc2091ba82dc15e3e9f94a9b9356656c1d94fbfbee22d5868b9f95c8e25317d56da22b84e5d3978aa328a166b25f77d4ac4d04b45cd26a0e31ad13e9a0c91b46e67691af507f395f4d8d53762f0256bcd5bff0fcb473a815;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc626b0775924183fe33cbafb7d78432553505b34a4d8d35c8c892aa735ca22a000942fea7f25d8541a1657a2bd22bc843adcf1d8825f4a80c707316d00f23e258e768e1ab5a816eab6ad448152c7e710ce46265f2fa4a2064caa0c8f4aa25a905a54aa7a218c74f99a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h174110999afc8f918cec541a469cffdcdfd10675a533b3168297b4325156ef0e1fdea09f4ae25d66eb7e6f9ee8ee7a779ec09edb3786a39147561f88c8aa2962d45d21111e758b35e775a503c4b174033098783062c101f260f99241afd92a29f519c8b8107bd5622f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ae66e892b65989082cfa43c4225add787100c7f1c93b5b3dd1005a8b00558cdfac938c8e8508f67042582213aa6631cf7ffc267caa5aaa5c0b8393e37d8250f5b17b3dde3200c6bb86c63173a64e17d14b5990b1b2f8cb57d013e0d4cede1f55dbb750bb6cf9564060;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16fd0279bdd8081c33d5a5691113019a5d7471e221bd104eadc5dfcda0e035f795b5c39a3cc895186865a938c5acf78c7cb14b5eef2adb92ce76152572330017cac3f09b8905d797772ff99e6476fec85c29a570b2c1c889f136b4d1dd52e4d9c7af80b1146334d485c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7094356d22042e6dd65988279bc018fafa4f41a31d93105bf3ee47c6ff008fcbb62f1bafe1f370f3803d1537611189ed6b603ac359f8e2b63a460908ba8c3d970eda2edd327daa1e6144f928219559c6653c53c07225f58b819810e418972e53e4c57259967871bb9e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed09d7bb5325447fde783d7b139a265c826eff630299008a97ab4ec5f95b54e43ac0603d8a1f64c70809a050ee7fad380c85b7d65f270df25b289b0eb57882a144ce88fb2a19bd3c8d181d2f91dc86619653cb7df909dd0719e76d377902894ec3522b991cb90c72cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h152bf60e2ed1de06d387629d72f95818cf8c605e3b9d006a56ab27e857c6a2a35038e2a253dcf32b5d8fbf571b6f13d2116724af7df79d09a2a06a6b0dcd2641a8f5f32f06f12dd7f7098fadbfacef4e07e8761a2b9f8bfe59d5f94deae16576e0f5e5b7a7f930176d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc02d61b44c59b1f8c3742c13cd0b69d5ff693fc9623c3a22c2fe850ccabe093d0d08aebf94844f3b82b4ad1f42a1e54e1b8929303988a164c552f6854d7af79dfd6fe15eb6de7bab44af45af5be1bf84fe5298acf740c92e4e2c2626f7b2f25dce7df4996594bc1fd2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h178320038f0d7b900bc965e9d3e1d0090b54d3644dc724ce9972372cdf38db3f98b2284b7178073694e1daf45b3d4e6df94a90dd3c5381729c39b05fc5c0a3800d4a788be0a55fa887d7fbbbef599c68828ddca6663e4871e9c2ae369405b2d9243c646cd7461ccfc1b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h185b31319f32893f63647c5e1e21e7e99774c558903cc0f1754ba7f726e64d870e3d5856445312c1537b5e8c4bea27bef19c16d8d7bc88ba8a1b7e43c3213d43ca6801bbf264067fc0deecc79630f064a0c07be6069ca5586d8a79b2118d20e96e002e60a6b3f31ddc1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d279be41b25c18a10cd908ec259f5e17184d2fd3161462aecdad1a43ced23908d5b3649f7bd8b3c2e2534ef9b63a3ef24b0ed987645eaa95ab7bcfc1fc46050c21e6929c3225218168b7a109bbda02d3344e944e7f7816ac4f2eef9c745cbc3385b35e662a46697c8a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1817b2db67c209e3a09acb25f9e006d72a1522580de47768830d0c728eb777df4558afa6a484bc5999f3774d82cfaa7a35293916cc95549f5f1bd1f790664d30cc216c9749a2e98a42492bb92a96cf1fc05a724d07bac8baa63b48b829b3a8da09ff94ff0e9002910cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59a0c7d5d9cf772490e850313b12c21477f2e54acbe9271aa66e99f2bb734fb411989abeefd04f86830a43087c24928271645f4ae509bff4063bf1c905dd817bb49bf7a4175915270d501fdab036096264b5e1c42e51cc3601a18eab0f61947126676c60d82b0c9759;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd3b64fb1d800caab7da8e15487c7269276ca1bd224042ffca4a03ff528f50090c3a3a48664ec07dee2e1e334c4eee38f2d64f3c7c511572a7bc531c221092ad07a3980141383a8c77f2a1f92376eddd1f09d060cbb0d934763fb501ad063a36928e6244bc42ae65b23;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h393b40967d08bbd645e317367f544a8be3057daf6891c9b07f9923c2994b98848b9ac17f7dbe3354561a785015bc7f79675e408c5d04822f3b22bcf314fe98546122756ef5bdad68c6ac63187c68ce6dcbe8f91a44aee298b921f1133cb2c31ac1aec793da5bdcf8f8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4a529897993ff9777b9a95f9092e75dcf4246d6cdef422a30d97a6498bb9aa7f78d767bcb7ec135e6db1a25e5993527b965443e9ed35c29c56116f3904f0c661e9f8e25690560f4901ddd91bf7d06ec63f1925b82e8b9039cae8131dcb2b74427d599a4dab12b81cea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb43e1310eb256b9c93ae5da8995bdf67cd7e6f0e1f701d1c3b3a41feb3a315432431e75758072e8e588bd308c6330acb482e2caad57989c7f502c9b946beac1ce40717e6ce0c532cf919326df24f3c4a2ef8554ecaa0d4dae9642aa1d981479aa98ce66eea508b178a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1794f8cb14c6a448238681bc32d4d9ac7492a777f219f26a2ff95cef50e1836900bc4a256cde5777dca927a41acbf60d216020fb6a69463a5f9fe9cb745d8f4849f85ab6476eb1d780b43a234d8f7f3a898bbba4ca852758d46e6af5869601eeaf06e199078d1acd53b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1215a4e4e3af2d0508e8541a1c07a6dea85ef9d783e215febaa776a744443e3f4a8a91abe62897f4c80b91f1255a9c4dcd6e9431cd3e4765866f05212e674f28933a5aa5b952f3dd6f509d2e6bc23c1d30fa72c188f8377cea64fa798629da173f3a3b0f29f73d1ed17;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha79dc9dfc6e71455cc787684c4c2a5cf7714ff3b37fb916ec89dc9f67d2d79cc3c706134ec45ef83a510499ffe30307c72079cdd23ab1a8c1cf88797f1ebc0cd32463de0147f391b595e9cc0ff9ebd7d402a860b0b2095746827b309420c248d8fee3b3f66c524ff3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha280edb3425ffd6a4fbd24f6f96b77a38326832eab285d47f1bcb131904c3d661fb8afad71a1c917cfebe43eccf350300e63d4f9039bd68df6a380c94afdbbe2c6b583ddffc4ea832c94b9a0ef9096bae9a54c03f8fc9b4ebf51be4033f7889e78b57385bd61d85f0d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c8ba50c8a876bd490e73d5bcf5d2e0a335b3a69a39ccf19d00ca46c9dea9e5af53ee28ea99cdd81d96f43ab6947a19640a4dacaba502fc84669b152d4101f97a852811affe3f359a578986b55db503fea03b775f1ce30853abbfc4583f28fd099ba4789e2ad92ac2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c92def2f5b0d983cd9f9d6cb4d43f5cd708a620dc21233eebef67dcee9ce3d6f43414a51eae31ef662a2d3ee7e46ab6dfcc961cc6fb11978ccb5ae00838c1cbab3d7586be5b195683888f75cee32c496847f18e3606728135b6c1c5aafe9a04923ad962d41c8a5572;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1849e57a690c9205ca17ceca3fafaabde48079ff53e0f8bca25599132abc874e7c2e78820410832eae74319227406fa46c9043f667f8232d0f0f4d6619810fde5c21bcb9b8f902372d291945c65c8af3ef45611788edfa6f6beb0a5755c3aeeb2f01b9d66c54af6e5e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdbf78d909edb84b492709c43e54264353cdbb226d522958d109efdfcc42db3261df62aaf54e9d08738cbf6683cb3b60ad7ec6be4a95495f4f7bcfe618181514933656ecad3f2ac78d827b8b2ce012e270358c078f0417c513b0a5b33f55055ab6d779871a917ac3111;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2b1325a3ce4477a3d339808af1fa553479f7be066fa1e97fdab7b1625caf46677d76457d9109704a82f9b853511d2960dbf51f7a8953db0d7d8c651a1f3865b97ee1fbae0e6eba02921e2807d321e37e451ebd35eff44c936975d291d8cac51949f334437074a4869e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d213a125700860de8ce7ac198d9c9596bb302053c057ebcb1c64cb6592ca266361f10ec32d1aea59836a8a7f5425235a3538b34edd32490cb89f4f40b4cb2f1f30dfd95ece4896e1c94d6461b79503531fa1553d326e66af9cdfc3f9c54572fcadaabca9384fcb8ca0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h104d935758027512ebe5f1ae236963ef313fbfb181a3a16aa053aafe9904f6959e251bba78ba31f867fe78b3e19a3cd7f4d0758e930ccc101a16f6e5ab3993d4c9016433eed029d278f3875b72cd97082a75e52c58a5b924a48201c7a93d773d0c6e1d61e59ea7f8fe2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c08c55667370396e915ec7000fa7faf9dc542a54b5401a918efd565cc109616d00f974ad6b383a32f391c9c57dfe3701f219cfe5f7864c6460b2a9fef8ff6655bfa708783bdb8db5bf68499937a298c4b199628cdd43b0615fae2c977b6ac45af29ebf4d98e815ff3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b3af43163111b8d9ea239e1ce8aa749cd097ab9dcf7e98f48370d93c51fd8ea5d895994a9deda9a1c271e994abb58fef21486fc73c78be53ef40bb2ee1ca46a7094ff5a68e06a09a450f08f4fd79116e000899601aea86cf8ecd69432633d2af1e205799f3065d82f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dca080b5cc3a72690da168fe4deb9890531ce1c054d3a240f0aa63a3921baf73571cf6aa5864b90143d6f04c361d7ec4eb64ac27a818be23e15d9b0e314737827cb54f15d855e281659954dd5b8e102e836f67ec0b98a3c7f924c5ab0ca10970b351c22a8734b23dec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc4db2a51ab75655a487e7b77b64d67437927fd79a8afcfd935f9f709d2c56650f7c4a5ae8d04082d5f74a7d26300e24d930e1713d87b10b51fd9ea0ccbd56ca62dfd8edbdcfe8e996adc5802b22747e07a0bc7e48f3daeb3a46a19595a1ab4a37a1311a3545a5ce97d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fc412c8e4fd38cd00902d03a44a282c726650df7bd760788b0de5397726ca439a694f666a96d31d3149b2b8e203a72c4a5c8ed2713e2f10155bfa09d69a46c9451e482843f702cc1c4bc21793fd4d6641563175d2422130f303f43e978d10929dab91ca84e8d8b0245;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ed4ac8c9172ccf5d95366029e5f89e5e1d1516f587e6d12127ad48da3e650795a18c8d67bfedf2af4c185899897c3afdcf54128042c924f8f0f16b8d0a42cf1e1e50d7689f28f22de19a580efce1a12757782374c3491f37a0a99a2ec0ef5c084d85104b86448157a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8082b2840dc3ac8b004e05e04401b74078f9c94db193f62f8ff824024c249625e6415c6118eb11d48628e04992ee93dcaa28b0c26a2c98bd41d5e04dfd5c43ce15e7b5bfa9ae11facbb02dcd03a42732942510c30c950ceb3091c5b409b7e49905de6c366b5be49495;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h160a6918e6e3caf166db56a0f3398233508e97fe5ee22f863435279810432dc816884a61e14c01dfa4aff111d541c2154dd320a36163becbfdbaa7a5d1ea161badc245c98db5f5ed089fd4b0eb4737629742565fb7bf000e1bfe2a0300eed45376163b1c46e8c5b3a99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2da827dd77c7b2544b694abf05db89193c3a9cf6b48e58391c74bed0fadeebb504c4ba1a06acc3c647035e8ec98246d9eb94b089db164e82c9bbe92086f478cb93f52189f0027b6d073db608c571302bc6bd0e7fb397ec757829d05d66583ecce885741c3070d0913f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9565945ed89bc5d5609b3a283f37f6a762428ae0da6cc8daee127d74ce5670d9d2fc57614eadda254ccb84e35ec9e7a3b2d9f20150140a27b30bc1d0647c01b079adadf429f1594f5cd49632f3893856fe8bf77663b8f16907ba837d00c3976cf6ba7e79e2d58d0c61;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c2339491dece2881f09ea8e963caf247c5aff43cdacbda0692e09253e7c63fd5ecc04ad1750d361676ba58a50e13f8268236a552f80ff5e857c4e94902e630a0e38e6665e45104f606064c7c1e6f58238ccbcb9ea42e0ea2f58e22e6de15cff69b7379913b476ec14b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be8b23993f0ee07d6517e84cda5ab110dab4779ee8f2f33c91864661aa5e6798f7e45eb927edc7c3b2ad7ae546779ffd4ce6302074b41382b46e18b3723ba5d9e650707b599edbd31917e05cca803f59dae208b5d4f825df615845818779d79cb1f4db44778f41501e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2d4fbb155e164c18abd159ad94302534e9c79a67262d09ac5e7535a1ecaba95a537461f5485c147332a56a95f8d1bb4a7d6af330ec8283736a11b1a659b56cfea6b74764df43665452525b9d5774dcdb1d6785fd30970d5569c8746cd69ef3d4fc720258c939dd107;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd5716e10bd5290a5a82cca34031e55ab5443745cd13c9093f45c01d8d6b0d1119aa6628f5446a32e893bb8ef586d898e65af7c53e28ce695dce0a2d30091201b43bbebbc7be7479cb1c73a4c964f7a9dc92e4f43246758c9893abf7f8bafe9256ecbf1bece4b57dc70;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9fb42c68a92d500d2a2777629dc48880b5a1082a0d9d9475438b4d993c0c54734ab5c9d5bff07213ed38db701006baaa2a47d1e6feb0470c7efa4ed2484552098c4e401fd1906445d8ba9e42c0e425d5b039df1ef08d5c5b7c7acd7cfece9fd6417dc3a1e9bb62e55b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6bf74862b0860a99790e0df3905b31d873593ff466233fc39078152229388d19e09d1260b2be748ec73f52ccea8a5e5ac479ef9cbd92d2412a22b3c9d59872a2febf631c3c9d1f3de97f19947071c2a2540929b937dfccafee865c77c0b6fa3418e963aa6361eaf54;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haee3b9a5c83c2f9135a1a08d7ef53d75fa3a158a098491ca1f0281f4039ba25cb90a5f50ad9943f0bdbbe1086d46a632ce205006666b1d79330924108549970c2c036ac11860f26e429038bcfc9854ad3524b949bd1fe002c1ba7e58c569505819e3487fed20d31353;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h462325922defe1ff0dec8b9f68e27f65304e657eb175a16024f7aad07c056f2de9c91717c902662e4b8f3f4d22a6e71a3b3c2370bcd3311a2cf4d931da534253331a91df4fd4838a778fc1eaa24b7bc249623448d6ea512bba7f5ce6e6ab7be2842c4b0cc2fec0ae4d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16431028c22c5602864239e164b5eee6ea2d3ada307b6f35fb94e54e0ba49c7f795b6c432a0f68484063a27b7280166e3c9ff5520e251d136340f6031daaa952071508505d37543b068a69b2fd04287580809f278b8a2729b20ddeb98ac7d6987848978abcaf6e2241c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7c2e2bc579e6232fd3767757f838734b66d05e57ae6e0d926e42cd017b7871fb4f46d932d1f02377a6cdcfdee7391bccd4d6c6c83e07129caa471c18a88ccff41a39a9a9d6bef05fb4576ef5d7a444f984d57e519a0cb1518913f5926c65cff358b3df468d24ba0c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f51c7222ea08c54163ddb91e88a52287accc0dbb8b2efa2290333240b08973f6886c040b25f3153b7fb79ba0b4e580d25862cc85cabc825f8e23f97c1588b2d4badb05d0411f7fc2b03269e81539bc70a5267e1f496c99c3c9feffd2aef04f45047de0b51c16948c6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10da4b2b548b09b9654e7c41c11baea4a72967a708617946f0f57757d984af3cddb0b68f17f6966b546989ab965a9ca6e070414cb5a1b60a49f964ecd6c875cde73867e9fc5483973888a5667e9dfa696c12d7859215a8b5b6eaa9473eb9ebf2b94071a0e1c9d2598a9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b556bfe6fcb0309972ef918613f1e51a289473f45e54df35b12507077bd5105721207313ab7bbd795f7a59175c31530364ad85bffef2680dd5f0a8979dc6caea87a4807e1df86595871ac7702c3ff213a42ee68bb28bdc0434b16a77934a9e0c082e350f20b1514989;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1930b668571c3d133363bab2fb7cd11eef98f55d99e8bd55a4244634d26d6503dba6bbf07291169ea19e5bf917cdd606191d45425786cc4ee5be13022299bd8051d6a4cf665025529135193aaa08da59f8a6072486cd39a241a815cd0e2c746cbe31eed2dafd2382a4a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f0a03781ace6ad6b1452c102f933fedd20c38d79bd2a0c7fa0aec5e249d004b54cb6fcf9f5c6c4cfb06bf2f828880feeb17ae2e8caccff48d716bb7c3a3ddee109cf2e104a3c4e02e3221c84fcc62b08ad34bca9a57fc0021967ebbb2679cb2f074b6af9171ae35352;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d1ace529538b0a170bf351659966cf3efad550f6bf8d261ed44cc1a3eb2afd6d60c3ed0a5c29233fbf4d87fcdb44e6ec8ba91797ae4dddda3edfdb4bf2eaff901c5b33ea6cb1abb6414c08f23f429ef76aef146ae1e8ce448f5368c1ecbd7b683a61b83cef716e9151;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a9554ff9d05b2208f629192026bdde662585312190c848442013d20ad40b7db75809e25af239a5b4614b7ab8efcc26c2c6ac351d30c8e34097f649dc254847db61c8aab97a1b267c16f9c1ee886982fa1f671550694daa0c30423858a5a04492f2301bbc8eec7d07b4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8dbef88979fd79e3e9d3597517e9452d6a5dc24782fe4266294ed61b480d9f51a90928dcf3f1313ebe3c7066ee44ba9c256951328fccdbe922d1797f4273de57c572589df1d22092c2c44e73d92ccf753ea6be59426d855fb29766eafcc8910ef1a0d43f05573e999;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h616e376a7ff2b74cda7cf61f9de2ec867107fce4b56a0effbe2824a94c98da0ad78cfd1ca050b91c487106e5b400ab8df1e7811fe413ec77fc3fe0152f777432f44ad84783302d62b890b2d823fc681d6e61dbb086e2b6f45761fa2801989b6ba1740496f59da5cd6e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19b90c889b58a7ba74e2ade087d99a4d731fec184c764fc24ae19aa1110d6a7b1131c53858186fe0a3dd32fb741d602bdf0d1fdf265706ed9635a5b25ceeaad71f6beb843588fef92156468a27735d66ff7cd8f3343ae143471ecc9ae5fef8f047005dd12594ffea6ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc22d0e613f59c0687cf0ef8a67f236093e65c6e1ec7ce46e74edd7f996a1c7a16bd7421edec6b6dbada258b6b62f85f719b09a9e016ccacbf9039405f36148bcf13da02ddf4072531353fde666c712a307391993ee2437f106117f057d2512690716d03bbebc70b33b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e83921b3605f96c0aca039329af7e614329f4169b47ffa9a7dd5f275cce6ea39131e735234e77345e5c7c9d1ebcb251a94ca9b7140cda025d09bc81b4cfd4de09f8c3ef5ae3d87151a08442b375959119cbc98a08ca7ffc6446802316b195b8df9c277723414ada39b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb9a8008cb5576c722eb5f4168112079aff3841d6f89363da0ea9445e7a309358158c032c7b698ce43ef3d59539f626a34a1c10e840ed867f35702dc34cb6c347635d8b23a06afb733d17865537c18a97c411e286415778666f08220f141c8b33b16b5f5c08ac3397ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d6cc5e538a625327143a425906024cb8a3fb3338cce68e25c2f1cdec911025d680e4bcc95d3588587909bea6dd9f9b4384477dd768a23e79ae0aa880e31e1bf5d4f5176ce5a0675881ea504c884fe11ff1250fa07ceaebb7031d435a6c189cf699c7b03d8358f637ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12b62d6279e454534607a1616490a97b1d3e63d39cfeeceab3580874b2b805865404d803c780d55781db92d0f93100eb308d03c596e089c970439e0d4e5194dc113864720aa9ab7428db76cfb420e2fe0d081c9a54bb4d78fa62cec42ce70cda7cee0b9df6aa3d3408f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb5edb3dfa3df249fbfe358efa5e98d71f51c790d866b4ee60f5b84509395a5d1fd32e0f9f12f45bea82e28400c993ea56f5860ee777ee5a2c350a9d5241fb5070b058b3cb45c559e31fc59c484b6d33d40b2cda4661211b56bd0a0b95bc3cc4dafdabdb55f5a655a65;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcba9d09666a65f925f784f3db569fd9146f7eca6b1ad74026e5b92d3abded242ba9a66d1e7b70147c7d36a3433c99739f0e56f5f915d9a5e671f67f32ba9e1963a827373d63399c857e40bc2e7f901f7bcf86dd02c16aff1b1c28be01816c53b7a382f1ead8890738c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14e9b6252be24cad1503da212bf7caf67f6caa3bf7e10b7a1baed0f0d4e1304f16812cf20c39f4cda8e58113f3059552ada73cbf06ad877eb38375dec6c12652415170690a1a7f1e5904b7770a0316970afa3d3d5c59d89a9d2afb29c95e96ec9d39fea5b12345f83ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h168437336c55ecf6f7e7d7b8bea66e9134ef9131e51eceaef62fcd64a4a1bc098653af24f1614ba408261fac7346150d94c22a929a168adcefbbdbc041b4e7d1c66f286e22e898c9abb965390c588547eb68e9de5f2bf49c27bd23bdb38bc7dc758e5dcec1ab596d0d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h41bcf07c255986f4ee60dc5653c5b3a027cd9ce04b6dc017d31ea509205d1360e6368d53e5312f1182a21630580d155b18fef534c3a96199523f5d0439d4c055d54568e6e6069306337c85767f5dc86313956bd748a67d96e22e7b7294cf057092b8991818195b34c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h30e4962dfaf978686a036e2a92c2601bb459d9c3511ec19ce0cae024db14f72fbad5eabd7c61dfa22226401522cf0ddcf9fbf1d5df21d5de00b13ee5385e0a70dc7b62fd0db0f14e8775a303ff9168f59ed6c48b04bc5d346e998fdbd60c63a2d5f1296aa3cd5d9f66;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h103565012e200d5f43c7df6bf3e67a0beb9a743f9d7c825c7ec3bf2a976781ba91a5e8b01783825081087df12b7e80905156d40a2df8c26418769e441398947f2353652cbcc873d046dbc95cdf9df82ccf8561829e848b08e1c32586a6458c67b4a1ec05e7dd67789a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f3d32a5dcdac09a57d956da86032b44ca736cc6e34056374a96dc2d9d675f787f8d6474a676cad3121b4978d4154db255af2f7bb4ae14b57c96b2c51b5dae99fa66cd28b870cb75a41576e87e8c5cd9530f17fff2bcf12fe96581fa6f5ee4871c0a1df23edacc779e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1018c5f799a078aed379b68f19217d7d320c6e04433cb38820a9e2ebe4d564241697306bdaa8d8a173f7df9f7ec70d1d6ab481e2da9fdbec82f49ffc1e6b5c455bc339112dd80e0f3915bfd80ac0aec0495177059970f10b8d8a040563bf09a96c52c84882124299fd0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1107cc0835600a02526b53e24dbc06bffbc6b8511e26157432a70056087211230a83167ae82365ae386c641c8adb62e1827d443e2963236936a781ba3b657623d5b605bb6b5d287668768a491ac27660ca5653176e51d9d8e6c15ada9350fce0967105002bc4b05454a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14cab25d388fa7b1e8cdc7a9a33a6f5eccce49ea4e3e568cb17c3823a4b16f085ae7e6b4bea8bef576953c59eebe59c3199c9a9f358ff3da445ef7449a5d6320de4253788a1746bcbbfe1143aef8d5c017cf08b410b812a850e097bb387a4d292e256d7f1d300eeb0e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be71246017f8e6f12235dcada3fd2f20dd7c7340d8b1a5e548daea1e92fa22d44f578a6eb7232bf950eb9c8e465ca0bdd86d8f1791bd0806c0edd72b69601aa82f5a2574a6cb5fa7fa14c60babcc4c76cbd32481e25661662ac8587c136e539d513c8db781db9264b1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11bfccbccb4491aab28a2c1d0c3a6383dd8b1d7f41e9bde3a9b85eddef17aec6d75133c3ed1fe44f3fde2d8da3fc36b3a099100082d125663500c93e66242835a3ab388d342b378f4db206de0cf94861cbae10658b8f21807296bca2b95dc2b415456fc90496df7ebd5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a6f01a66db32b45cc9f38d96321b918f50593a959618b5f081b641fd3e8c0910bb268dbbeb754bc62d7a6425339797bd9a0c239cb6265dd71aee21983ea89eced8fe8499220ace3b433917f1727b5aff12ba51d583784fb8b1702ea59450f7bb3ed1c2422fc9232857;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h99835028e630037eeed196a4f2dd9ad9767d20ddb854b3ecbc527e2ae965f5ac64cceee6d7993ced2466b2088d7e99908c57702dbbf0217f32f2cee62ac93c78d72b8438d5f1f4dfb588ad95ef277f432b92a34b4c663398042f1dddd1b3978954b8ed082d8d8dcd56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h33bd1e473d460d9feeeade3c6ede65b4b09caf6124f887195575286639701d6eca50799306285625a6c3d54becd95981441baf0d2ed63a2639e6c9315f029f8466eaeaf70dad5d6d8e69da473839114778fc8f88c5562636fe9e0c6a2b553a05233b2531fafb092941;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c80fdcc876cf908abcadfc81ed1ab03a7f2e8c1cff8698a11432260162314a82262c10afbe9880cc0aad15cafb19b6ac5d3b7800fdfa61971df3013f1997d2394e52121b292369ae49092a5392851aad51c7c3201fdd13a04634fa00696b3193f24e52637f4ba2f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h71d9e9468c8d20bfd2d8f9a0e8d175d86dce7067320d1f93ad7890b10ed40052a87d36be10ce4961573feb5eaea0a4eb9f6fd0827a283c6e387e537e872d94248de39769875d2ea44bf20fb35e6abee5e4e7ca1fb9d0fc179e667d1a8ac87606058e18640023826685;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h159ee6357ca8313a1843a54ddc04f92d3f79b02da5144c2d225ccc7526ee8939f831b0f5b8dc30439fd3d0e30d909c2ba73f6f199a216b7a0b2eef829913d56bb6e18eb7f0117ee391836d4fa675a6247345e9b7b840989dbbdeeb553dbdb23ec2b4a8500eef3c5b86f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c923572879a82a365e5fb7ca6291b8a894c166973a18d1c0da2f7b2be3720fbb2d432b569ab498c76f128a6c558105a3ce506c55ec68c2196a18591ef78f654368efb861f04d8aada1c537e4970850231342a1f16ee91ffc65d6eb6f697db992c38d77cc2d513168e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16fc84f05d4a2f886ab717ab74090612c15164fd487698e49e868c04ab135f6f69600f85f5b1e9f8bb40ae251c9dfd036dc4efb4fa4d67880b7b4388b5efc1cd0baf6c102b0e76e3e159a90dfd3c4ae1e12ce08b6b3c24962d1db2a3e9365c3a07bfee2476e8ea9a1c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc8ca1af2af0925848603b39c55db48432f82e5e3c8c37bd5ee6b519ce0884a52d58280c7cc174a3f5612a1e2d835e11cb49d349fa2e871b43976d521a0195158637dd14572cba0cc005687149d4060581c694706e574d438b3c2b48611303be7e88712593d7bf7127;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197dc143f533b0525bf60394ff9c0cdfe2c45058f8715c3569e804c2341cb5106286efe82cad3f442a77ce62ae7beb99a536a01dd19c35010e30bf38f587bc3bbd56ad9a1c4deaa313e68300cdbb839fcaa5d672c2b6a0ab828fd3ce1d16852e34f59c0f17ec588a8ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14cdef26ceedcd763b6385aad0ca24e49c266d1b573fa6ff2f2d8a7d2eece61eeb6d61efe090eb361b1aaf88708d20c8792ad686306c7e01efe0a99e166d4fedd455de1b5ba491e112103406096381ee575c85274b0bef179f534083ac9aefb4f32d402bc8cadf0c341;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h637322ed6459c70e3ff1059042bf5836680d1592de59562dcc6e9cb94e11126d29200a2d9511255e92184fc07c0a2fbdf36ff7a3d61c4530d97557679ea0589fc109e0c4b8cccf5b1d5795152056507b041d38e90abdefa6abefeff953a10c092ab4b245661a52ba5a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1741804c3db6ea072f477c6d0151084618c6890364a8e0df5419dd9aeedf02bbdd2bc4ec8c175508422053f692795c062073b03130209591821779a9cedba3bfafaa28fabc868023fba2833401f0db0fc5525bc15aa52e3aa1373395103f3337c0fc5ca44a739ed1828;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd6b6ff25ab16a8ddf4e0edc48b46ce1625b9440d5b852609fa72bf2c50792eb419417d37c137b6d2402455e49509bf0d0d6dc59b027fc71b502d37e60479c78ba6389bf9e93c1729025e63452d22897a04a512c0a5034ea82377b9ca331d5c27e4a575f0673379a257;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2aa1e5bf6426350730351f48307b385453aa42706a096f42d1370b70d2f47916507d5b9687d2d44754eb2196f7bf2b70f525ff79025a06e932edfa6d3a6d1d35e22230d5fc73e1ad968900716a03413b6beb72f3ee12c5c5778c6b2c18bef52fc93fe8d7e6c5856b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19cc85c755fe3928116338301a77cc9147ab4d05f7720dba3d36c95f48aa5d9e87a29522e3e1cf8f3faf46aace9a82d25f4a453ac4afcef37f2e9b073ad87aed802633c7bc202870ed2d1a933097470b3e5bb9108df29985166eec462008cffb9a819f1cb84e0bd0ef2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hede1accd38ec01e94465ac478a227d21fe8a8e049ae019b924e5c4e57fd498d7c6ce4d2ebedb1624215ddde6c12ccb9a1b2c4e236298425ec2b23dd3a10db934af73dc2e5a64d2bc47dea386c7562f5ad36c440b84ba1e5d4e01ac6edcce88cd07c12078f613b5db8f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2e81730970bdf57c5f5abf235e53be2078c95b3a15e3464c19c746e71324d7e122bc5fdf6366573a117180a838cb50cd15991d6b31f651fbd9c1182eddf706f9806139dc3046dcb76923d9e9724e4accf0832f22a349c5001b9ebfa991e8ccb4863b03f85d44621e9a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd53c3c9f9a3d9a088cb1631cf098779b6e2473ade830423413d7dcc39794303de7c4ebdfb59a16349489b4ba360ebc7dc851fe1cf3ebee58d0f7eb4403e0fa64ae87a5eb50f52095027ab971023894884f1181d31010030b7b8dc8ee209124fed1651781d3b55a044d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4cb60a57bda7e09bc31e2b1e8f241228392f4c2871033a7cce0313b7213764fb1e5853683715932a96b1d80c0731f5791c1abaa468256cae1028a39fadfd5d500a9d03da06f06ab420afa59ddf1836bb5a92352f8a7efa951f8f2880bc569ef56af2529e785b83eb25;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h893e10c528617abdf997213204593756b9c9e6eeea76bc74f37f99d35e560c32f33c5031821acf35430ee57e24c440077786aad24c668ede4cb307964f5a794933e9de89b0f289bbde048f0037ab16fc6fe1ba33bb2702ecfb42d8309698b95a0a19ce481507dfdc22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h57ab6f1e047a0c380f4638043959efdaaf1ee446814ed7e6109c0286d15e9121aefb3f085d28d6f6409f55c0e111265c56d353402cc34deb61005ae522fa103deacdd1d88cc88bf57dbdd1b0acf437b8f0f35f5021ca496e941ac23df0c04ef627412710093f78a677;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8bdf6a6ea039d4d4c43fffbc6500b4f9cde762968ed5ac8c47ebcb4a38c88854721f1314a7d164f122349fe0965731238bd7713bb47e90348530eb7235217fecbf167dddb946f7732f9672a4c9a52dad4a1a3362a7e69c74e65acf91c9fa940740df98b70f491ebaa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a2acab18db46369e276b929e8075a30f3aef9523486a171be058b5eed49446d39eed02178f2fb674a3af711ac4e72b68f04455348e82d35b7794e1df88764ec2d57d7b2d4ea1faad97d035ec8024b995449bac56f6c0d6a130cd4b8c9ce0121c8630a2b2e9437be879;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a85d9db98ca1eb901d329fc7c05c94db0d05eefb15a2aae9d741a6fb1a1087602938c835e3cee5933e2eeebcdb9a6b97165afbf327efa02ab078f8c9be4482279c10188820b0be15ed6e3039aeb7360094854857e8579e014d70d16bd55e2facfeedce61d8941c3b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc73bda47a1469edde7a101aec0d38bc2c96c67a7749ba817a465324a695576cc012f1fe02507c37b9a7ea0411fdca640cdab09624e6663f48fb4f705db2109b72e191e1a8f135ffb29d609a6b2c7d4739497299591da07c3e44c4807eee7d8a6e400fc0de1f938b0c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d347c14efe91c136c3593049b220b020c857a293398b375dd58048110239066246e488ff5665d57ffbe5d7998a5c16731ca377680d6a965087c2ec3335cd5a5acde9244ea29ebb35558e3aecb90ffa632ccbfc8c4105fecc4d0a012186d6cf8881ca3c48ce6db9bd0e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h81daecba8a251ba3599f21a03a283c112a1b348fbe3d640c951c6d8ed67968a5ff1c60aa8ca29f58b8dbb0df46a5ba738b488ae83c683e63d73c015d2ea4fb17ce4fa1acee42af62e83547098be8a003eb6b76d60f8ba40a1baf74a7ed31a3edc1a48057bdfcc3fd75;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde4f7f960b862e45bf36fab8d6bfdf0a01d7627d7bdad41d3d4eac60f0cb91be86effa7a45ac4a0ea228b808e6b01a17dc992cdbb2353e332ab59b37a260b17816499248c2be1ac8d0558e53ba0dcd1932d53fac3391abf9ba665acd59a2a13d3e9582929b1b17df66;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0b1aebe0eda58cf324f333173786a98fcadba2be89dc97c06991b43abaa04d0df462cd9f344f5964cc1f1b5f952bf310635eb3ede8cda2669b5f2e635181b58d9f5eeb3aba60884e1dab9265b787e3b7960602c6c4ce2087490ed5f536a3726b57b1c1597da960332;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h172699659215b2921c1ed34e162546603ed75638a699d863c590af50c02d7bcdcc608fad7e9db81a0e0102ad20160fb1d5724105131740bca2c87a547ca32b4bc254277aacb5779d8cd4832154c38f97d9fcd00b2d115a329a9795b8963283efe117ad671b1bc23b13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183c0ed929a954d7a082f76205765ef109131313e364b3f62a63bbe2c6710a03bddf616137bd946a74f89b0c12cbc00de60dab2555ad688c8ca06585849d6fbdd115437cd988a41d9e1ac1634b115beb7b89a488529e9c941263526a062ec2a505e81d1b617941f28bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14aaf9d1ca7102b78b1e421c84c576d6388ee23a5663ca23c222fc2efaf71d0b0cfb0e0d761744e707f6eeb2790462c60c3d979df4c3a2aa9cc9f7566f7f48ce71dd6b6b47543eb59fcefc4d3b7406fc382bc389bf686ab17fea61cf15c61ead179d9d1406d1fefbce3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13415495beb23f38fea7247ed922d22ee6eb3e77b5233a659de5a8fa0b5a12152bca00c0c713efea5a1ee04bc54799e9539fbf4b817bf894f9e5658175e38f2a72bd1271744ae91853faf658b3ebb8e92396cc347e43436cbf9a809c3b4869955ef4213dbf872378f54;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ff2b27a516dc8481c7601b42623f8fb34e19834d717ad3ebb2acdc3463ec3057c164299743d16d7d507ce7961d60c261cce9e48c16bbe6ae787cfbb66f8374af2fabcf311d60ca7d4d016a9df3fa8b49197d00ad0e97fc9a1703526ab4588817cbe9482c3ff9c03ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf35e0acd85369b0833264888c5cac09641b789d6701c05314a7dab68af788fb83d9886c29d26f850757dcdaa5423ef15652648492b08788f7e66391cac6165a085da446eb6d3219c731dd18454b567ed44ced5b2f4c79fa4af354d0f176a9a0029c1d032ba4a834c99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h72857ed21278a6018906b9010968171abc1fa66049742fe92ba98bf033fcd8bd719f8feb0ae18c05b5ef5f8b67bce2e65b268c003101ec3abcf3bb5db80b07c844b9c7d2b158ce70299ee45bb498150f60935169f280c4c0163008f9cf1dbae1a470bd771f19c9ba96;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f18954f8c75793d18c72520d4995c40375a5d129e3f5483867cb7950d63b926720eaddb2d444249b2ab498cdac0ecd0792e5f9f180b58a2554b0df1fe10c28b5fc76658dbc422fff82f596c6eda5706c05edce8657825e75e20540702d96ef3e586f5234e295793f8b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d0c958f59db11662e09e1555c3da39290f96184d5e6dcd874501267fc936bc65ea47e197c661f9981850e1a0760f894f8d601990f64474eb8fb34c2f4bda368e3b46b389a6dab0243745adaac7cdc94902f1073a1d648c292fff551e0df64e8ea6ed0c6aad93a8f11c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1118b8acfd745e691bee7f9f1aa77772e49ca0fc7f91d6e2ab57531abd2aafe39819e5d6f695c44b3dd1082b5cb6234a21ac2a7ed26a3089388a98ac7b4ced8bb2040d776c3415a94bcdb0b0fc63af0c2588b0e0e46e5c08bcfafc3078f1b4f89b4740e99e102c2aba5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1672a9225091387e2d1fcb17b88b7c7700c6acd02474f0d0a681dd9cb9526cd4e86df348d1b14973d4a96de983f0514a6db7a42849a234e6852ec8ba9d14850efd08ff593f211c9914d3eb4fc995e2ba053c85e37abd6de4f53869a47a559cacb7c2c775363132ecde5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfa59e03def6ef25d995567aa064eac5faedde21a3fdd4056d9a0640dd35aea302ff3d70b3abbb83814d4302502970c6185c88d501649e8434b1bb666b0587e6839dc5684732d6c5828b2c71a6379b801f33510a8cf6452914ff6905a3c2057ea58008830062c209499;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6dfe1da49be1ef1c9bf0b951c1b12963d98fb860aa7d8ff46070b7040db06fc2d150a425ba5d499971cadb46f9a90e27565ebd9122eae62184a923b4196e5f0d166ef0cbe0218a091e707e3adeaac1a4589ac00d21cf8497b38cb759888e734eb25d4ca4cf2c45d6f8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1417df6fe14f5ce44fa7c8d10e602101f7219fe5f5911fc4de36aaa54b8461acbea77b893447c4510ddae8044ef4ee1a2b89475a2b8ace42be82f97a8989928514991f2d1ecc115033f28e7fa91e6a07643500f17e4cdcdaa04e6643b62d884f719220ac04b203fdbde;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h138abfea18ec9c49658027cfb24810413a419e6654d47ebbdc575ba54af63da3c9306c5a57aa0d9306f9a0c247696fd5122d9e9136e888d83d9c3034a3b15ac5ca36c469a80b569fc3370c45296092463d4c0b2201bb53d2ea68986a7cc696229400ddc61479f7f0f38;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3a82da06e9961cc9a5a598eb8d01c7730f7b0b33d2950ca9db0500f55870b8ef040a5364b152fef398e4a1a4e228e4630d39171de7445836c9e58ca7dfb26036d799034a3faa36778d23b89e9304680fe7e245721e4201ad216f9196ab495aabf0f4a2c31abb206fbe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he4d40266d86b642a4930362dc6f2894c87c449cf41729724cfc1bb833db8d070c8aa7f4d177e014e7ec39a0db689d04adb16c4240ad927afdf9ad409ff2f9eff51e9f9e067a585c18f5a5e9a341424ac755a6c4d0f06d416590c34b2ae7d307d2a337234d2ac7bbdf7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf9bf6014d9ceaed3529dfdb3744f787197e1642e2b711711ac537e2c95e1fa74b2e045d90359a1c940e292b2923d2a1e26150618e2141a329e9bd049fbe66c4b3bcdae7c15dae6900d136f77ba39dfb18fe5a39cb88db743ef4ed01b9c20c834ae80a89dbaa185bf23;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h143cec82b10bc8f276fc32ec6edde06cdf9cd2403a5215ca75a07dcee28b75bb2c80f1fdab987094a81c80f1b7d999826be8ff9df9a77a460f6cf6701ad9d6a22398984dcde8ddb7f53c52eef91b0f1ed85ed7fd5ff100f3e089553a238c436464b5c8fb06acaa8b0d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he803eccd331811267db19a160178aed0b370e8a80fbf93f156223c758b65433bd812b577d6f05ce90829f58bb855709c6cd763121d4cdb30165ea1412e7d1c7db9792d8773bd71d912ddc4a912b199e03e6bdf9d2bd2f39fa0d8b208747855621ad8e41b80a83c6cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e18b3fd9e2e5c7b015626ba5f26a5f1039562a6e0cc754926ca73da691b023ab86f5b6552d1923be6d9fe6a9f73e2171c68110d3fa32cf7343a3f3aa7d477d83e930738f32db6c632117b982705bdf66e9b62bf1b34adcc3c42b63ecf0a64dfd7564e9c4e776490db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde5e50f049d5ce2c92e82277a40e4becb8e3471471c7fb5d69450bacebc9ecbb4484e7e5c9107406b4d7c00d39b7e0bc9e5205cb9b9baff80b058c6013aa0d974a8bdec45f9e21752daca36e7af4c76babf28ee3fe3388acdf18b9c3296bfcce693d069fa316537a5a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he1f783b5df6285238e1db62ab0c7de6c59c951537a31eeb726de58420ba14e9b581f6243edbb016a300223363532ce570dbbacb5c6b05138efe0a35b004f11fe6bb8999efb8693d8f93976874f4c018f96360abaf0ca8da03d411061dc573c7362758907a482f69f1e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11e710ed33e325920321c69bdc92bff7ad33dbb4c167bb5369fe5ec0335e73bd96becad863c30c6306a1c4beaaaec311b42c5753072d0ba7e670fd885ff623012677cdcd01fb2c5d38bd0b4f42521fe21eeb27069ac00635524d39f6dad5df9d358d47ba4fbc54ec2f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1384d99b16900b3d24344b7334a8dbd3053e604f70f34ecee9975814c62724f5d13e0df884a686144067fca46b197da84fa09b587f23c1c698b279d326bf2322c8ed773c7b26f18b72942deefee8db374668c77da4450e672df640c096e1351bd246fd68df9aeabe077;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hefd6f4e36d66be0ad534d611f44a37ad61377476c71029996bd0dd071175be6734a843770ba8df87adf42292c7dc7acf998b8c1d912a31d5a6f1344071256861d991f50f756e963ab439ef87212543172756eac3f3840f7a444560c2158483ef1014da36996edfb3f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h715335a8a7611dc146bb3cb749624c6c6dff695bec8c8ce9da622be613b0331573bd1d17d7a017a3535de005a71e7304bd1de858fe411dab8bd2ee032825172acee282e6914f073944a954ae1e7e815f0e836f9588150cf7ffc5978820295720ddb337bf3d2b67a9da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e636b7c72625c90939c1dbb8cfb26ea16f5a4510df2815070253048abbf2c98e672fcfbfb0876c355dc095f6411cb9f4e106cd469b3c6d8faea6d17562dc2cb85619cc8d272d1ccee66f9bdbc33c2cb8801874310eaa9279d3e920409b5f257d8cbba957af57496fe6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h181bed1e1f8bbc0c29001d16bf7d16865c19f6762da086cdbbfdabdc8add52b728a2ff14f0fa27ec16af1f9a5912920c8a9d7be944ab23c863c87916a9647d473fef102dbf2be30d09d78aee0bffdb5fa847810c8a98cce2c5d0c0b051e2fdb4c7d8be02fa581ea0687;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fda8d755833b14a5e1189da62dc7cd52ed110fa1c90869576d9160e6101d7d6476c482f13a720d502313a3dafa331e2a56648f8054bbceeabe6c31ac93c6f44817f4373217020ea857c08f661067b3ea583e7ec08da8c74bff046cf3e78633877e9723fd8a5e6fb1b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf026f98fccb7a1f704c4bc2c60d35ccc6bab5d91d6b32fc12e5e9296e4219c5b31e3189309ccb747710e0f623a26cac25f773fb161665151d0b3a2e2a05c871e8c8733bb600606c5aa983f3922aa3860386143919ac2e709386db92f5d99aabfabe184a31984eb848;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19792790ef29dacb13317e4895544df7d957900c70a615513963f03f8e2e91bc40741a115e25e5d8b7bac8ab08390e80f2472dc03e9b15701b83b9bcf17efa37e754206da1109a9e47f297df079babef129165b3a61988cb7f62c9b4bf2841e435daa57a7f328fbf15b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3bd6281899b285320e8d1fb1e24a2827e027e69b82496290c86c4db89f530c4ac3b07d184f0962bb28d027039a70b75d1410016ec3b8af0ebd446f8dc2f7701115dc3f3b0f890fd03825c6dd88a2f9bfc1d3b9e41960ae2d00d7bd8053c6d7264227702cec7baf1e53;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h832e0eaadfbae6a86ddd7104518a732c3691aa22789562daba8ca4fff16f2ab46a15f651b9ff1b3e2436fcc830a6f6bf00d6ad7fffad77cdae976560d10ca355242101a6f8752415bd953b16bffcd2875492e243b965f7e78b436f3165a06c7a7df69ebb744ab2ee13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ef0df7cba68074ea981cd9ee24cae67cbb20142acf5efc50114d5ac4a43c248675d2cd163c6d4631c9fa74dfc74319521bc4b9ba8c00a7614a23c47dad18d4791207b666d078e434c77c127f3dbeca828d3566a30a4007c4349441dd97e528a1f19ec913311c8a2f92;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hddd29040bbf8978d0e96e8c5aeaafd689f3e508e2f85949cc785352681633e75ad33e30a1b340a5488da8c07763540d5fbe20a895bf23c8b682b9001f491dd6aa0214ef95f69e5492efa142da4eaae8fc93ad041ae07be82dab7a6974cddeb71d3b4eb255062acafe7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h86887fe05da34e7a8e02c5e049b43267e7872fe18ff0f5c97adf620e95254a7d08637b5b498bd784f4a5972a5dff53a96d6089ac06ad48039e9b93caf2e08436e588ab0404f2a8e330ec823c6a49797713309f8cb9a189f8fb23747b283aefdf6ae0f5ef4a81719a76;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be4cc0a1083be5b57f03f3e6e4ec960dc90c2738d95e62fe329e045321058ddc0ecefabb5e3c1080e9e4030786d6290d87ce2ae9de8e2d830bdd33152c7523656163280d9bca036b7c13817fd774380866d2c825209953e4f70431deff7898725fe41fb466069a53d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18617cd0b1de58dc8530ebeb4fdf8c7cb42c8862ef627893b1ec11697f5c30a615f22ea007f860aeefbaf3ddb78baf3de1639d4fd67817081c65eded780c14dfc46c1aff274a4343e833be3334b7ff4e48cacdadbfd2d76bfe775df3fa67fc66126bd3dd446d19f45a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h169473673792610f3c54a594c1d7750c3e536acf06d40612e7446d275efa0b61933f5fe58c48ee33cadc19fe97d08a6773aeeb2c1bde487d6c54129e64e05526cd412bc7ac5cf271677adadc1bd0704831dce0c119f8b27911b3f6bb72726471e9ab0b4124e60007d88;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a5817b1b660d56b99d106fabe9e0522046dae7fdf9d6a945a9dadfd42c286d151edf828116ad9498c40c2fa3d6bbaf370e5ff8afd1d1c57479314c88d23d2d02b83e24e3ac37d47f32c16799b83d0ff8dce618b13176584531ce917eab6ed3bf267adffee2d35def1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15128d8b9823ef8b44c718a494815430fc671ebe00a65e99fcdd26b98e46a386dae94bc3267eeae6ab3d061034b57498288726a6794d75b22037ddf128738dc393f3a7e818f38d022753e26bc4845ad7af6bf3605b95dd014f2d14ef8a7da827ef5b10400192e6762db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfad6ba429ba9d10ee5c98bf31cab377d55ec8edb54e60bbcbe75aba99b9ee1f062398ee48f9aaa8edc5d622e578ded2fef1fb92590157799ee84c8f546f51d067d8547da7c5eb8af71756e1f9f849fb76e5e57c363a0211b1c60f167fae790ee3d1b55812947cb6b65;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed06e98410936019615340158f1f46ff2ee701156e8e1cf068e551a00dd6fe8282879342532f2d087da821a8cd94a64108dbc32f4cb47b6e9252a606c426d86cb77f3b404a105820fc263dd83d8ad39af52fd41d7f923db5d19c5320808fb8b9f258f4ba8b38cb0569;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f1c229d06ec7dfd2a4b78699fe91da3f952d81e365f1b672b2e90aae5e4e7b70a1d6c130260e9ddc39693da93c1f200031141da9947c543fe960b505282ab009aa6928bb66360b2346ef77430a37f7edd9f9f6199aa771d723e15fe37dcb96ef9aa5bb58150cb4ceff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h129d3ecd576ee39d0f12416ef3361ca34553fc8f90e4a2c36a4a8b80f451c6c23915948cdf90858e3aa80085c4019bf6d0750a7dfdff942ded1ebc2c755853207903860bcd9b7aea0fd92ef459d653f18e3009eca8f14c59a2e1deb85b3c771b740e87a19151cdc5d79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e0b3b4f8c53e6231a54e96a4858db17b567cb16d5436919ed7c9c8535625b73cdaef0a72e70365a27dc13b0c41955f3ffbc0d010cf86420e3cf90abe8e3d0e1656cba88cca36dcc7307f51680ae2067d0a39fd138b3e4e1f7b8838d9374f1afc44e7f5d4dd2c8b8f5c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a56e4ae823b8433c4a885e7c7a196a7c81dfe765ce4b6659a73383054abcf6888ddf8bf98c58206694a8737ff7c298264e208bb0fce442d47a50ff19644529a3b1a9b31567f7778ea30e4ba31dd11b204677349595d8a5f64e85ed292e460d913b67e77e3bdf428cd0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8b6fcbd80a92144309dd34e9f1262a1e3496dad5bd5e2e7e27453fa9b8fb6a9ea3d364668a5bb25ab8856f92d1d119a116be6eff83761f6175a9b1f6db22c61ebf73eb5fd4c07d8b78e230574ed11b0f1eec31bc7a2775d20738699c2a0203261dd03f72910203b4a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6b0469eaf4cb78f033630c725f7094a0206899b6f56e7bd5f7e684ed8fb560e4f347dbfbc01673c210f31d9bf052ef407e0b129b165830e3dcc476d9c59175bed813aca25e151712f7477036afb8caf055f9bdc1d6bac44c4a470eb15a37727c10026bb1b493c0e4e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1b7c6949ca69a07691f5fe5de64c4925ca58c9d75d125564d4de30b528232bf80b8bd476bf43c3e57b652b4bb552d93ec3ea07512e67bddd57fd156082a65d9dec76553cdee2ac70d244ffe6a2125d6c00294091a5401af699a47cc1e94accec206960faa77ff2996;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1006d23317d5c503f274842cfd1211c186ebd8b2c20d6652dac5aa8aabe4842f897b4c146933d13dcc3950c2a86810b727020fa9875035adcb3aa4e343184e18d4ce3b09b96d12cfab65249ba1b680f73edba7d8b60c08f31861e316d936f6f89a670efc914c89aaad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba1f2d840ba6cca244f521d2fe1ef8db7863c33b15e356cf92bcdf42b8b58c11b4fcc5c24d81debe2e92b55b231bb55d45ae785e5b5af8204c4f55dae809d87fa99a67bf06d8577daab8509a8c98f3e30445d22047672cda3b114834b8bc57413329188067b47cbec3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd1e1e4ff4ab1921debeb6a042dcefe628774e9643f30649c7bc152a08405a929315793cb6e7cd840b6735cb5dec053b9153b1b983a971951a9cab7ab448fdf0300a8f8e742a52ccbf7e842daaa055b054f9c1f5a73764147e124c632e745e894ccb8fa9f25f9fea85;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c6e690e7911f115cdcce948ccca2e59df9b5c11d7f904eda086c5569443a80290d91e090504a49abbc6d1b058ec92b971e0265eeeb0fee0ce8d3c42b85a5ce53f0450860f12cc2717dee70de651a10ab71a8a03d913f6f65cf2ff970ddd082b04c60ad903ca9c7e23c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a600b5a7f014e90619166641fd7b499179bbca28a19cecff5374b3ad880fbf459d7e8749f4158b27fc91e9c5e9685a3d47605129d52689f548970882aff10a53e46c31ad6969f00c03ffcb9c0e8bdc64d57b43039f279a81a47adcd0bf97ef9b484f7040a4308dcf6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb2a26f063887bd52791e9145b175c479c1b555e0027b4fa1f4bb5b24dafaa68bbe19a1e0e4cc97247b92b67c8697b713466e1663600e0092d1d3259cd625cc1c4b3853f942f91268a0433fbadc8ab936130f4770b767d8f61cbd039f50c2ba76634e802ce31ebbb0a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd85b926cbe108c477dfde5b73731716c9af6e7a1242c3f6d8e4070aa5c12d38ec1dfdadd1ad1b9aa560dfefeddffc142064bf03ca5217b1d4d534955420efb6d2548a05e4c84730853ada73c5e123519a76d90cb5cb0943b954651c072e2e86eed9be941f9745d1b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e15102878fbeefc59a2eb887a735752c00895ef990f683f7035380103f9212f1045345fbdbce3c78bea95d326be7dc8afb64d56ed517b959bf0134571d87b0818511c540c46ad8dda7a8b00fc5fb27397f00d5aec1317cb7cfd39586da7f6f50c688961ac9e85b1715;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c92da1aa742f0ae87a633bfad61444779a21dd2cd167c15366cbdb071e9c6e6a91e7eadf9c75468939d482eefa8f585edad52942f7bcf009ad83d30fc71d971c66c295eb9ec5388fa2988303a92021983d9118bab1d64471728ed2312f24f4e7783591e98dc21e2959;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18923f376f7401857f36398e1de8b7391dc03665dea8ec19da274acfe1585a50ebccb94514cfe13ccae37f88c224cead1ce382cadc2e43c5139bb384fc55f129b26e1297e2eec24a214c21fcb171000571b61539c76d3284b75bff0e7670eb0c29e0ceb9957a0bd440d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha8cdec9a54e108d86d7b30a0965637be268b1ae37ad1853fa981db1be257f50a2fc430c5f3a9e678aa7cb860deb627a87f2413d38aa7a0f27e3ce96438b953bbfd3c08b9870166cfe67eec62d8c337feca75287a351cd24e63f66a68fa8c1d2425bed53b636c8472f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11a8126849ba178f96920ec246d00b49f27ad38df0992a2c7dcf95d14c6e57aaadfc2faba2d81681dc50cc45b9c8da463cb3856fd39329564d7f4562edc6ef3aac2bbcea472d263476c8369ead3786e8e451928a3e4e27fc662b1bb2eba2c2673c47f6728d8959b433d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12f1671260d25860011ea8485a08888a151f04a14a549c6134527cee80096ad4a0bfe0c7667ee60a5274efdc56c1e9b7473d3d3026e7e5b3b35c85d738caa7dd84dfb67100a8c1ff965b5820f6c7c0551de5bea23c14456e220c3432d83fa928302b675fe24fc6fc776;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155baafd5ede5c4dde5b6cc3509f027814a4b93d82cbe1cd1d0e9abec2edf22b36792e2c7d85b46da0c3711e7ee68f0e5f99415a594bb4fe80245223f166b8f18edd6e08eacf5e2ec61ce7e8a8b06ed199ff99b1071d69db1e555d118298392f37a184999d8b0c57c31;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1707116ee071cf7cb379b1ef87b54333a241eb0f299d74254e690fe1b993d53989c9be9197145effaf91b1ca19d22394e329a2c1604ead8a24f177f4e5f75e9ee591dec5603fd958640f6a6f1a45df2e3b342b4523b0f99ce9fada9e80c90cc1d4c9a5e3b8033a90322;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10d19c9e56bffd21b096960109dcf769e24da519970908b5b4257433e455a50a57ea6eabf35fcb43cf4c0e0b792a1b5af7ca4a368bf39f4bd67408bf1382a6455a01e9caee50378b4c907eb9595ca6a47f4d5525d770b6b1bb9ac1773a0f336a7377ffd95e3ac646c4c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c7251b8dc42da89670cedc57230edcff87209a3b0315a5524d19e1e61befd9ce2555ff64565c097edc0e5d9034c4bf0e8f9f90e08dab170504939a82647165d6199aaf6073216a5c83c50f21ef78d07db67a9a6c22de52249f9015bb088546bad9de32b6ca43b83a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5296f5f04e9b12b590d8da9c446fadde0f8198ed73bc9bf5fce7b747e602f55c01ecf261a56747d44d5d553e3e96d614adaffa1cc7a588e390bb3dd106c4c11dc544da1b2b2f1e5a561b84f2ea2dfbaf0293fe3f77262225ec8b59ee698278bd9efcb505e77b51cc3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3f0b4ab8bc8d62472cf007777ae964f90f07d6d81bef8e40b845598b1edbb905be8fb48f90e62fa6c7ecc1d5c69466c9177d73b462ae2a5fe17ea669aef7de81dd4778fffae40be7b04d3af1dd1ab67dbaac95e5da3472d5cc2de91f79dfc1f890328fed33129f8b19;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144115ca73e1fa27baef73232254d798357b5cae24ed386727a726fdc2ab457500d2b13cbe53a44107d258fc5beff7f106bc88f8e506e0d78655b24a333c275d13db5264fc7621764152a1a0de48b5b38c3c63d9bca0d30d1024ffae485edb1d41baa4e6650e6bb60fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1c2b6078e409e3a9539cd7ea4df580d65224893ff42f5e80ce6fe5e8825bb2e9616ae83d8de32c4a1ca69fbf270bbe27ff8b26cf57739ee8375a0a387734505feb94dddbfde26f2f0818fa2f94fd2bc3fa755446e9f6924f1348b383a0a42540331350771604bb91c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79f6473a079c8a2293b51fabfd74d6d2d01b49a8cc017d374ad142a07d5fca48871ad356f65101f0fcd07ae9f54c9754ec8d64b3cc5b9e3eb16945eb4aae8087cce8a99f4b0bf7de691268d9a5ff1cd4b0e4d6da64955d963a2556d609356335398714dd6d9aeddac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3067fdbc9c97f746be7e160efb2dc9d454f4412046525cf9c259bf0396f56ccb670c1a2de82cab4ab34b82fd8678a9656b71a119f5e95c5ff7db3e2cb941fe8a5d096e2002efee2ccafbee3801e2a056a831f8b41f904752aa60e92bed2cdb46578f77ee5b909bcdd9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a364e883b7b2007e0891e50a0bef7fcf06531e25193455f731b09544f10f2217a2cb09469b513a667494f03715a04c7964d94fc2991dd1b6b855ff33665c25593b37628108ea454e4a8beefd66537f00ea3706eec1ed9bf0ab3aa865f44d6750abcc184284cb6ef5a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd6a1026ccc049a67c2d3192727e61f35cedf4b3e21d2ba313ec9bc13adcf752df51c8fe52627989f6beaee1453821459d5cad8dd926f37a0b75dc7d9049839998ac3761d8a7ca6af5a9a9382fdb3edae3b93ccc24e7eb439e00bd901ca419ec73e2f720c76aea691de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc995b45b9b704759797cf3bb9ae6606f471e266407a982a3adba6ad8bbfc7c4a74930694bce4ff00577237269e96db248c269e058a5f82d96c0bcf5f32b56f46bff669924df3f84dc6345c95081b16de43eae60a4242a1e244f0497c89b491b72ddd2de519ea224754;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10030a135378ba52da9a2b68f9ea2d59a9119ed3f437c5786a88a70eaa8dd4471a38b4a4bff1d5ee421c1305f70dd8b5489ef59663e9beb7a2d48e65a333f101de605d6c8e744d77c42e03899079870f62daee3e63f473d9a57c2082dd14f4627607062948baa75c9d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a87f8772934ce5f6a15b93d6259887daad183769034f0e1fe190850b9c9eedd64e34cda4a69eb5b3910e10c0c2d1d8ff0edc2f545fe7d9a8c9fd15545af30a56ef7ce476430e7be7688a11c56e6f87ce00ff317e493218c7df9a448e4b72155e05017a92fa61fd671d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3a531ecc8003c6edbe1b35087f4bce065fcbe9843a7db17d13311d16019477f6edc2a6f79d292e4d3704ff6bccca0ba5a52e9c5e2439288a8d40ad13e5c909518922b1d8d86492464dca0fbdb64d003487e58f54dcea8821b970e5aeb274c98f05b1df852928b61148;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf38aa6a1bdc53497bc23ff1d454a86993bd7fd007a373ce073612660dcc0f5d9c44f07cf72811b5befcfad0cb9d29ce0ab13dd744d623ec8fa1663e8a3aeb9bf7259792b26f5bdf58b87f7767c780376dc7e183847f0d9f3162a394f75db843847f63c076877b16033;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9ea627c09fdcdd829b23b17ea5e3d15773eb2c11b836633e86dd6107b68ebe6199bdb7d93b457cf34b678470802ef00bd5ae17ec00ea582ad54290366446acce5d2a17ab296dee82e96fee663784a9f192f0deea085e5622f21c0a6592b8037a4de6a51f214c02e522;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1239b33896ece798772a4a2fa359e1bd21f9b06e0e2345f1cc050f3f8c7e403f227e9c629cc35ac5259aaff28dc4d4fb73d644792150597b0c2953ec4af5a49a16d973bebcf94e9f0c0b12d6df13297ea91512fa19cf1b144f17e5bd492ee2295f31bd5f50a9220ec3c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf24cb743f1abc08acfbd9b8ad481e7f298c178ace44e8a0aa5f1ebcbdea77ff89bc1d71c4dbd902b6631e60ef5f3f60aca60d199e27660c522b259afe312d7deb8ce87a9fd163eee05cc2549e84fd066046181fba8631add95ddd0ea0feef5fee2e5ff8c8395f13d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hedae44c7ddb38394db6137f8500a0919cd801a57782c9d85a8a3f725930aa71581566bb4d667a743bc9b4a7b3d2798887174cc10bcb8d96d29cc3b4fae209d2c41924dfea00e3b47424addcfa9a205b029235a3a72929fdd1c692041f35b1a340b632b1deff70b93d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c509c1e8b57f492505a7152994b173e1bc2dc52d978f523f609d896f8a2db24031611dbf249aafcf00f1fa2cb72d2e1a42ffd892de044884fb1dcf4f85390487745452854b788396d0efaff544471fc0f8f8eff93c042318e434c57642b6edfb81acbf08a3ee45b301;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b17662c9e82c0f24818b97fe2ae3e54397b6261c2e10cf5069db5b1be7d6c1d14077b04ef40542af4d2f5f2185f8647d3778f882eaebb2dc404b2295fc7ae4ca0372052fb54aa03c9aa34c8ca8050f78da8b77db61e81e05b6d9b139d558c559c88b1b69009dba99c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a1a18fdd58769fd3a835d1a29eba36f7a0c8e8fc9857d3edb7c6aab63339a948930196d9ca68525c834bd8788daaf8d959a5dba275ab8643bc0e98e3b030fb803a3e80458fc06dc0af8608559c0c935771955c991d26cfdb35ef0c97b16fd7a5bcabb82345e6de1e8b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5a4aec2de0011272883a1ce9e50106ed2df0ebbd120693b157414d02f0232c18fe360b01a20e0b4e9009219f5a4081b6049346ecd5417d8209146fd19dc77b3347d4d72f42dd4eb96e3323c936cb9d4c231ce341b1f3f5710bb49316e3edf0906db5dab7a8874132be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c46c96005b304fe08b38e4cb291e98302ef6f106a12b9ae6eb85afb5087aa3bead9749ed665801278c91d2f566bb1e408dedfc535c22d29f8a82fec2412c37e272e9bde4a2ff045acd41c7ce035abce54ec22d030e2f3dface7d59b104803bd60396dd81d1b2c2b90;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h170b9f16d253f44b16df01de88b08741eb64742a3586f9b9fbae45459ede5134b2d04f8cd151c258d07a692231bec7b270895d71aae7f075f745a2f0ba8ea83425e8ffa7f6573f58fa7d9581aa3e3a2cee529e71c63b70e9abae80425bf9793432cef24650a122d61ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cce92df36ed2e194707edd7beefd65622ecd7e1f8815ffd1e1cf68155b77559270cc618731ee5e7a3a0cfebef8b8be1d91462ab6a1d06c619227cf360af00d7ef4473a85f6f731f625676ad9124c5e67798c5ca3ae106aed71a9db41678081a3f46769e10655aa2944;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12e56bfb8652d4876523c460f3512f3edecdb321b3fae0a4d364b430ccf931cf19a8d533bf1593c9271105574110270940fa438616e60a103f8f7d3765742ebcc988aa16c7795c81be5371d97d7f9172658ce18c2206dd001014aae5997a830bd6da2048c66e7bc9378;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h88344cc59146f34efcb072f0c440c1d1f24092974f939c02dbbc5a8ae51a12b06e0004ec0fdabbc690dfa948f3382220dd200f93bc99ba481ba1aa2e4004b3361927619bf425811697d25950ef7f2edf51281e23ddcbfab3aa53dab8c1a094fe54118eb7ee3b212c1d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf750916fa46b392b981d68a5e99a9967b225b7df27b16581cc46f373fcbb4001ee5e7fc98028aa96e5676b9150eb2e92f756b206978ae024d92b978432a1f90d783265caa972a8a4a5bee6e3e01a34e571365d96dbf0ae7082ac56d8b32e67f8f9da2d0f83e858bb3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17be89be696370d89089ce31b3a095f5ec91800f34374662b0313c94df752982009373d13065b06953e548e1a0139158b9a037270ccaa088bd591e999d60bcdab91888de0fd97470ddafc6ca0f44043bc18eb694ae33df87578e919e4a3801d3944deb9391d7007a02f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116077f5e7ac2d61cdd32af8133c2527f1ef2d0b1f4354ebdd3b74e21d7b3f6d2985ced99e8836d4127e1ad2d54db6548d5707f530e79bba4a25ff8b80164fba27ff751ebf411b283981d270908acf9666399903f95448226b43a73f832df8de74dc6ff14445c1de9fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bc259d70863ca34fe8867965493f4879bd3ad1eb44fb7ce068ed218429fae2340aa145af0d99166fd8e0c83387360b7e9271361624d7e4775ae89a75b510a229572b5a6471a2728836611dfdd813b4c46c36335fb26d37da87853db677a4b5e42eb02518292755b736;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2f5b8e6c399e45042cecf5d1b30f60e9641f5e97503b62f2f0b20ea899963f3f0c32a5860635a37dbaaa67309eae01f7687e4e476d1af4faec572eb1e680074a10a0ed6b68a8a7a11abbb919a560a352f9ceb840eaa8f9850675ce6760c88ae8526bd932264ca28430;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b11b14e23b9ade1d1efb9335402b6841654d23265ee0dbaa06fc26693a2276fe2e0b816385a3f9e54a3e3e6b1db8aa3f322e8a5e53660c3eea43dbd137ce3ee13af99a0e002b46d9d21e402ff8e3037d27e4e8586e9a8352ad5216372ec01737f7f878d22d1c486734;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f8625ec87b85a89b30b365d66035b99de42e40e3b270daf2284865b8bbfc4d0f229a5637cb7508b8b8e8ebf3c7b3b228b759394a19c91185fea097c80307b35669de1fbbd833a746b07332196de3be64bbb21eccfc94b924cd12626c9fca3c5fcef00e096a87cc10a7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1655e7d4fbe7899eeb0e0ae2755f917b56f8dfb5ad9c14eaee78262db6b6959c8894cdd8cf65c529f38e4279dc1c479afc43f4309106cab7f4fed7ee00e0635a3abc9b427fe6733bbc697f1de29bd506eec25e59d53861f758619e3a7da3788f6f9cd9cdc1e11d1269c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15182fbf52886c38cf5d90f6c2d6b8e68bb3cf5d1b6c66c595cca8fefb4d03b7f34e6d7557c7906e316689a6f12d90db99a181e4637df53ce5b4c80b1273e499a5197fd7c41183e8bff64995905e12032af0a5c4a2424894dc02799015962a4d55d520e78a75a1ead1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1397c7696295baf5860886fd1d4e09dfde8c0530fc285eb6397604bab69ca876a7113ef84cc6d51a0594f791cb1f60c9a1fdbd9584ec60ab6c1a5f4ed5b293111c75bdb90f48e3daa2a842a5e513070f183a235c3d13ef0bbfad291303c0f1b28dfe7c748170657a4ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h190aa21d602938af6699b147ca1d784e26348b6b9d058c66734a687c03935b8b8a1fab96b1c3c35ba62d050805a8e96e02ec7dac0f3a731749733b38eaac2347f188a0b564b835d6bb19f8a87dc0656778f2f1f299e02f0d31b85883e6fabb50fa0c1ccd18bdd838c6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha37e590e69636b8e7b9d85ad386abddfe0c0434946ebfa99d184d521f16751179eac82b15450c457785940170786b98a76229df829dfcffb19a9d71dc25e39c304f760b7945903cd03d3eb74c3aeab5d1e7aa70cf61548ee7fba7341b00ed97a1f8917c37398af6cc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167081e7a6659fef37db4d6385643f701f13ac5d4b6afc1ffd2a277abbb019f8d83062cb62844b9496dffbc9cb10a7250edefd23154341ed3a4e4f0c874ad70ca06a3315dcfec8f416aa18c618ee858e5d94e5a40658d7f1cb91ea036da757f09094d76cd55eea9220e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd7a10b06d2f29e74e98a5e7c522cbd94cf4086cdcfea3233461cd703d4daeacc72a11d9ff9e5e82df5f84f8954585d8ad504598864cb740efd43d4d5810b0dd9e655d1b5dfcd5931db5cfc609cd7de7d30036dad2af0fa234f9474d36df7d2aae452cbc323bd3008ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc0300617bfa1ba86c7908732d46bc3cc789e07481c10e4a3a3adfe00e6be90f655acc12a179a4fa9914ff8d8ddeacaa65af48589ac468327b2c6d65a27f402d02caeb10474c6d836868f4689aeff7dfb7b4f232c97b8f9e71dbcee92994d5e448ff997523d2b93665a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1885fdc44084afa950940ef525275fb9a223493aaf342533d5f1c096495c5262104d527930c155880d1d128cf1aa96b8409a8ce907ad3f37bbc9393e829d861c429b84201c3261bfb46cac0d04bc0ef6ee8cefd8669a8962d7b8e90564160a419ef105aa880357fedff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8cc1698d5a883eda07c650d852c6db2cc23ecb03d9392a03f43db9df05b94c053a6d73377ac9162c5abbc37aa5a38c055fe396fb61fd30b9bcf1268bf36bb9dd7fd53c411a02861e90d828938aeba865e92d26885b48a1ec3aafb2275a797d7f61f998d9696e984a08;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d53b2fee4eca49ef1f2cae192eb752d871eb73de97084b6820d8169fed323e977c600f700ab96b94f326898f7267facd815c57293cb9949ed16bbf8da3f8e613794285001270e045838e206601c3bdc9529c96a21f8e870c8b592a54b4a506fc2c13f1b8b386189dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h73488304411b1a9bbef64360adffa73f0f591955a21cd1344bc8337767a5a601192786352da113377c24fec56ff61b1b3fcb1620a8d4ca3423be5cbeb51993968b7224a1d1051bda0f3139902a9bbb588dc7eb5cbe16d63e8a48ec1efead519bb78f5967df2c885774;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h74eb1c30c8035c5a0c33b2f723d650467e28e707f71f3547415262d6b22c76c6983b1469660fa0d244cbe4eb6f02ecf73c0fe6e85bf0f932060ac5edd4077ba32de4b10d481b0d568fbf15ce6d400dc6282e8008456687b15cdd2d6d716b03c563c250d4e771e9c20e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b5f4fddadf1ed981e628cc04b05672d65f5ee2d0ef08b0675c0f314325e1cb6f0b1d77578c9f8197f1f5641d4eeefc64e5efec8a0659f801b032a9e86df56885aac83fbee6d491d113b178ad3c171cbb62d2dd0ea8b60ce958f2e3e0e344d82ccecde5c1977425e46d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d053408d433a9efe2c96d2224ca74f92e8693d2020c5f6b8f30b801e42dbe84332818439fa821941a8d34470a23c3150bade0647d348aff2dbb5c71ca3e577dccd0ca8388ab5aae42f8307609572d202a969be91118dd5abf40766cff66ec5d2b8066f676a6ed3b34;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he98d796762a3d0811e20d2aec85559b1e0434beecabfbd51c380a13ea3bc1651639de5620c0a5a43c037a45ad99e4c75d1db689b2ffc85a326bcdc02d74ace55c04141f0cffd5e2d9b6fd482160d65eb771c1c65aa327e378e6f5bc741797f88733c5fc55cc38a2767;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f4d361a4e4267feeef24f2494d587b1ccb147c0691184fdd06e22b3c458736840212d563fd1ad8a4b4f4326821129d8db7abe5864e67d6074654a28306886016ccc441c3d915d8e83d06389212f1d9f49c4d935030375c82d631908013ec89bf8057ea9bdb53ff2cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf8813638ef0533f947e802eccbe83c6dfd0b99f4e03ee7c784ee91e3055744086dd8f34f44eac17d6399f7e0227b796165add0e4b7ad6190fa985d602aca7abacac165b60aa23b31467cab8d43ce4889e71b45f589a6639d806b1465f469ca4b001adeedd326e78958;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h33c9471f7a86098cb0b86e205fdfaee4f4e92ddfe1706b2f01a8cfdd15ce6e2e1808afb8a1d960193f78c022f254a17babaf07ebd442be1325e56acf366a3faabae8560855abe64f31993336724865a32071c952d6b36f6431f9990460a6b512704e0e8c9d42fe4f4c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10499673de83e9005c52e003682d49182364d5322286e4051547e4aebb1ce867d4c9c93846dae46f0bffa3ea742c98d7ededf83eaa2a37fceb276caa71848d3849a90526ab94f38160e77eb4ce848aa066d34efc9eaa4d2503f705d0f48c502f3de2b0ee14b0f39ac51;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be83d04c94332416cc71059731b13775c8b19a246cc22948382f1a7a1ce2d67f9880bb626346f758b84b3cb1e756ebdf3d0b377e124ffa5d671cb51d74b4635ece026cf61148955725e5c90a18eb8946969df1f7e18d0315bcb9e2a753fc5b4d218ede631f8ee30ec6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd8e57cd125b813d6707165cddf587181a5e703a04ded63e3a8e27bd255a6ce1f5a0fd5c214a00cb9ad21c8c7ee23785e21985f66f8426126d395a28beb958a425be5bac0e40d6761e163945476d2d0c91ac9792f5ea7be082f11636db6a138cdf7190d9ddb0361f2c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10be46bf9df30427830586bd2f402b59798acbde0959819b7e2351892796e3734f59181da0c9c11e2738d795958aa553d6592a441f793d9b9a8237bc059f7a3454a030454416e582d5d6789d6dba324528f089293e1ad54752d6c3ae3ccd94d902d9e1d4b6c8e82f9a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec9a1ad289d81c8960c7822f223bef8ac751a03b9cf0769a4ac64eed166217ccc216580a7860f917e6b931feecec29fc23f4c477f38fdcf7c7942943b6bb4499502d1d56378808329660a86d7788d01b4cff965448cf45ad00554c36123673486d94f6e8f6eb96c7e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5fca599c710537cec7bc685d6fccd48d42e19520c0ab9cec71fe78069399452e970ae48b4a8beea2fd566efd487a8578e69a9010a8157512dca005cc2cf29d7cde1dcf2d5c29fd2d409110909dc17cadaaf0be5b358170d4815f5355560d491a81e203d4f746c930a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h52b1d2f064118a140735c84e50a580d746512d68a12aa6215208ed685d2d512eebf548330e3d5840d7de86e462671bf425ae8a8ccddfd6a6ea6848e889ff276dae704f05d9a487a4b12e6ed13bdeb225a823062e9f82377fb17ae668de390aae4d64fcc4f721b2730f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf8fce9e4fd20f8f67424995d1863ec7f430354dd558608e77c10ee9c330e14cd139303fdae17a3be6b5ebb7f2d3d139ebcf5c3d35a8099421662322e4263334589b4d85a5f36d5343e6a39ad560186b83af9e75901fabb51b8b461f77cddd84c4cc91e0b32ff1c3757;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bb8111581d8c1c13ac790d111f1c275ed63503a3f88e72442db51fdb204bc06590fff6e88a17ef4272c037cf912ccff89e904d7e786ed91576547d9226c248c2944f6bd732a1d4fe9781d724e226793daca357d877e43966b9f15587cd7b6861c588ed861f292b4ed6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1493c27af6d218643d7df7d253138a84de6e25ea9cb3bed3f5c3ea32cfbc45a64c74a439713a88d71d1056528230902d3315e9f518979c5bb23b99155b54b7e32b7270dbb1cdd92b20bf9f19d4d21fbd3180e6bb19b5e30ccba74bd9a132cf81d30f0a92af081287ca3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5bd9376e81511406b2dae87132a8567766d9d3ee4d03555e7a98b88d77d72ae768215d311227099281119d3aaebd6f467701ca1756a6391833d9a00302df6d6070fca326d103ad5c7c503e772f1a30927683b80ebe509e2db94b402fe82d531e2c1398202a70013ade;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h182bd262ee2c0871c8371a0de422fa73fd6ab3c61c02c70f7802f48926406f9b7669d08ada5741c7c83000950d0f7b53d9a9f77bd6c905a02ca52e78c0919bfa19577a813511b9c68831631a9345d21f064f47aa29a4fe52758e1fd7c39edcc391ff0028c6c8d2ed78;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12492fc372b9bb7ec15f1c65aa3c96cce7ff6b8b169c78446976e83da59ea50f2ea29300375031d425ff2023d6199cd8e0d1d3a148dbd91bf38e18f7e04db4e85e9f7b563b57efe5529b7c922d79d26094d0c4c97595ee2cca1ee917cead795884a7f0acc9fc3caafa0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17be331a54c9a20586d195572cb55ebfe728188992e74efe53238d9ce76c096839fa84de8e1f6cd6b31a0cb8de2c7fe95cf2fbca48dda75ec2cd85631397280943c466e0ea3e588a853c0347144097b113c2f20c2ef314115ee5931eb351e4bf2ea3edd79e369a69006;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf3c6d8c2749a11e9d93f82ccc06d98784a981e38dc17b07fe7965a05729d1e32c55c5ef3740a383ce8dc11c7b94edbb924fbd2c5c879dd53fe6e948e96f2540716d0561491501e7026448610f9064971228738364af59a3335835d80a27fd5c0ba277ebefc6082acaa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf9b7484234583a5df2d0e2ccaf4ae025d8e22f89f6c70fab8248717bc453b62483a3dd339c76ecfade7869a5f872525b81617ab76f3335d502dcddcf8a3a573ff164f9db5523725a97b007c256c7f2b7a7c06d89c21a4f73cdef19a6bae68c004982749ce3141c020b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1547c58bdf8d0e55ad7c5fc5bf54c9a56ff6404cec3c0b745064aebdf89564f72fd1a6dc13c39e14028e9bf54663bd4a851117b031cc11ccf7de16162a14162380679fc20f202d239000941bd39178469ba31d5a2f1756e4753a01cd9e6d8e237fbad9e8b3c3e5d93a7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c4d061af1f727f84b406b7b77e318aee5bc2d504510e6036ed843e280de961188e3d5a99bc56f8001a3af3daabd7015c7df82c606b0b734b15a8a05744d0ec3fddf939e7d7e818e931fa8bf48471f9ee23281611e9bb8d6bef02d0b94f98655b6f75b2c026bc25f8e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17007dd199fde903b1c3589512642748bc5f2ad1884c73424a3c72bb2d529a22ca14de8393903e8b2a5fd6ad9da8227f0bfcbac6f5722183b6802eca3f8c634f6c34409605322746c38a6f6688b2f9edbc364cc5cdda5816b216b9712057b89a4cc5617da9d6d9ed52a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb53e97f1401795cc779c051cd007fd26cd2a0e405740386d73a780a7e3ade3cfdbae5486a62982b4cfe86e45fbd7f45850996ceb425ebb11be853ddb73ad3341a5bb3c0c495dd2b774d9a43077f982779916120270a7b05e767cd30133e5ab3fbe130dd90af92176e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ee4029caf9b17ed3340b38ac7a7baa93833f8f4035849c4e9be54acae947a19242633e00357c77b74fa2e1d36f73ab86d53df207181d171b10f6ce92b0c5472b637a4657ee8dd11f0c4e2f293f010c1c26fe22f605d562811ac7f36f9f2255d9f27fde26918f4abe7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17a764090d08ee259529baa2016dc93dc8ccad78917e451a5ccef11c8544b5c820f184e972aceb0cf3623f7bb1bdebfdd8b28e0066263b4a8b3494049623eb8c58fc2cfaff92453a25ba2c84ab3c108ac2e8c5204d9e6372fd1a4cb0de4ccd5a7b2854d36952967cc65;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h135a32b01d4cdec789a3133a1383c8a4e1616b11eeecc7971aecbff0454f76cd0db18eb64c8e645c078068091020df4ff03b7c2d3a80269d31ad1f20d03653e2666925a456e7643b29ccfc4b9d415cce764a9035cf3548603bae7414ce0fc486a7d063d0cf2e0f1933d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101102b1f49be96192b60e7d1111dc5df0a13c43b01c9d7dd597cb981816ceda5d6e46de2428237596a4d154d93fc34f01caf6d1c2ca0a1193701c1d3fc9bc21c29ef3fd55ce48bc4c6ea4de855c678e92d05be00542e59f88265292ee41a293d0508d52830cf85d36;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1211b0415fa18e01b0cd3d7bade41f3121c90ca5f553184b3de8e88f5a072bda9053f54b1a74601e7fc224965b83e5b6636e534487d6d0a0037a1d7ab2ee0089a8b3e7041728911a8d7b85c484e60bca30201e703d4756f4a7cae20c65f237b5f821a92e13ed4710195;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b415b9dfe3a76adfe8f0ad5520637ed513ba3d42f9b61b3fd9fa061f8f517886d144df837e8e7400906a1d484fa6a9702ca569239b67871adb623fa314e7ca2435276dbc9c9d9e5fb3c55e2910851f1ae1dce01868a94bb4221b371a410308dd9a30070c962bfe97d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1158bf563afafadb4019ce26ee6692bcd0cd063b0c8133d207a6e7d7c83193536b75623dae6dfba4aabb917f5d96be73c740775fc2f745827047eb468d41718d3666dcff08675e1217436032858a9ef5129778540544c4d35d65daa627edf63985ef691d90f7561edd0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h89044bb135073517f963aa7fb74585b0b336d172208d3303077ac58d421299b0464a89ceb10f101cbcff0b721f2c57db9339172eb27bddd6688d67974e2fef6544cb8a55085bd4a51326f85ccade1359cc96b980c6912f2e961f902c0c90163bd9ae76801a2a9c09b1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h646ba1113f3c2fe2be0ecf28cc4af538068a1ff30995b42ea405398f74e9d05d34fce6b3c7828ffc6630aea0d855172888c67afcd02c307b510a0a471d2659bef1496227a2fa08fcf385058ca6f668956f54d273835251806fbd821fb51c73e45267fd2abe7ad20c5c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5011f0fa7850d9588013a7ba7680b082bdb10067fe461db0b093f860251d352a7229fd3398331fad3b4d14ad97585d9747153dc8adbe0f92d08cd0c2ef0e762d21d7210bc1259427117366b7609dea585a04afa92ff02330bdef636a8c86e6f34eb7d346b06df9ced0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a2e9998ee677e1f02dc9606670e84b916e68fe897b7a4bc4c9162c65e318d7488ceeba397dbe40215a964a80e78b8fd770b0ee6daec0c3dcf6d66db5d07e83bb2ee83a7f2b59123b83cab90a50933d4dd5549c30db0cf7a4e60fd67f59b36b6ff55f3824e47127b06;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113b70e28a7064a8e0b56e2b93cf76d75836e6193e70b23efe93f9f844868f99f8769666f5f3d80a0f4837afa68842cdd71b5c8154cf918ede4ff371e4792d9102ae36cdf5fdcd360bb80c35c45d13ffbeb6727ff6b8344f8b4ffe55d4a4807ded8eff92f735ed7ba35;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14b1c038175ab1c03902ed49591c7126efaba42a12b4b58780d607c2390d2d456411884d2f86958e8fde60b619ec46b7fdcab74d040a02f9806e0180b30438ab8e77bf9776ed3d34deb0ab343f616c902897c9dea2ea27eaffc76344284404ca66978aefacdb6b10ab1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h20a83a875a1c45267df284a750f0885dfe1a7c5e759a4bd4019561b5e48b561e916f3f325f8932b302b09517c596ee6504d81fdbd19628187ede6e2a32406bd3fd46c7c8255dc785b8f71be718f40a911357fcecc14bf6e8583b08b85d27ac0c3ea8465ddc23fddd8b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14f5bfcc95c3dedaf03e48a8c19bcc843b11ffe6f9f82a52820fb059d4cb55e225af46df7a3052acaf16b7c7d461e57df01225f6e56aede372753788d8c5a820920e0ef8af7ffa4869750ba88c8345a28202d3cf91084d1798aad385e8a1e050048d315a8ca7bbd5624;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eda744d18bcc62efe13eb29f6a060a18c90e1e9866b59c121d33adcb416fe6e4afb1e67a370707ceada71c4464021329071509e3df3e6cf336e70485d157784c86abf29222ee87b179b257d31ea557ed738f48e3dbd87e5f2fc69b8db9b3eb7b152ec998b3db39883b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha8616be9efc1838ad1bc905b0cfd9ae81838985dae3ff112a56b5b056409e237f06a84dc7e58ee35fc3e93e04cee31fcf34c0078c181f3b01a9fe403b1c123aff88b0b6ff028ce98c3b7a21260306a4fcc360fa37940541e342dfa40873fd8897dcd4d4ae3293ce912;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf26efb45e13ab3a1ffaf8b6a91a4a95f367d46999b12acee7be1f5929c990e1bb4ec8d767bd621d68dfcfc23636770707808e72e3ef3e614a43ac81a234262530ab1f14d3f3e7079e64ef34162bb9f04a430c48c62318d746e5f8fefab14d44fa74546d95f3792e737;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1590dffb0b760e97726f75dd8965d967c52b77f80c6f7cbdd3783b9a09545b9ae0127f829e0619dd1907336e4254137271b64b967f23f17785b5040422fdd3cf109dcc5a001561bfa530c23fcc45a0785a6a9d9ed81dda68a5a42f0247f02f0e1f8bbe9c93571d2e88;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdcbdc4f51eeb1f62db8ec8d586d12ffe611451352a4e890d0810d0568e457add28cba7259d72f09f705cd4a174f10829f13fd920978b48ade0452901545002e6dfb1dfdbf6a85f26ed49181d6f704de0d2a5ee73f4fc763c211af07d2ac5d424ca0b27f89d3a5ba38f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0336718542872493bbd36f34e9a4a58ac540618460545351fc25ab339bbf355f5fa0341f2b238e275b183f601216fa57d5a442eee0be115cebcec24616a24f5e179027d67a6bfe78b95f70846af0239e45259184fadaf7c191c0c67304ed9fa9a489ee4c7efb60ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfeeb3db768bb04a496ff7a959252287b35a87cfb9837efff08e13b865b263329ce028b04bf3ac88a623802d3ed9c066513b8e670544f703eeb0a8cb773317915c64ad7422a5ff1a4cdcb68f67bbf8dade50a6a0edc8b1bbb8e421104853f372d68b73efb7403e65ef9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde9c3db1d7f340e211fef921d88a36ab3335a6c66f381cf2cff8e7c0b83519125e5a4914638f93c608fe418b0a5f51ae827bc7ba702f93458ce78c62f9f6dfe73170ec0bc3aed8d87fd91c6e6c4250220c5e3a868ef842f4ee78dd10d78d0ef68d941baafd5fb8e543;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1932122fae07420ce61f5bd68cf59a7841b950f57b16576ea9aa2525e57c210e326ad2192eb49d398e80fb6206ecf47e595e19efc7857c13da142a3cc2bd5cf0e86851bf7efaa9eee2e5b6abd5992ad95aca944842177dc699521ef26dece8dd0cc607df3c34eced67f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h275b4712d1132fedf0f29f1a8dbf5ebbaaec247e9672984043dba7fbf41e0b67ffe480c76109234da487bec0a9a0201006e3764e631948a5ab7dab44eb39517afb7dbb9a0b7abfc5c0c3223e85056ba5c88d583c462e81d210bb2c244bd165046ee23106231d25d814;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28ef496dda6316208fcac0c78948acd32647f3d711715e9767a4f0c6e48e8ed88b4b562b9c98721792c01ac43a53879b966bdca9344661319955d73d94d6ef27ab876e3dbaaa8d77fc09a117a3e44dcf415fd9ca9e92d0e595eaa6cc64810d670102071a9dc0be0320;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h25bcf04d0dfa9acb5770c0616b1870d35a9144dabb6965ee158c73e7ca4334ada1449d9bad39c6bc5b48952f6e70c9ad704a69b4136706eb1312e70ab814c9a3cbded114d5fe8c006b96d3c841dd3ff7a5f425fee4ecb43f239db21067f18b253be1a940e41f9ac109;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h180c59f979a5cad1697e177928d0b50cad2181e24d8ed18480cd0abaa140c88dd2956d0a4ce023a7288c688d28a6f21f9b2ea9a7c10c8f82a5ab596eb3151ee5620ee4fc9c13503202a71cbea772e4435803e6b202d7aeb1c234b97c10d32fa79a8cc77ddbedea4d526;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f6b2c328bf3a29832ba523cde529354839fce4626f0a22e42e770a0674e657f6c72ba722ff3b4eb95dc21935be7b6f698d128dc8745e101010a8e0e1f63075e022707078c23b236e5f69c65f898d0059e9ed7ce0a1ac05803cda6c25a92b757cbc6cc6aae7f419f365;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he96fed8be7af433f5e8e0555f3603fb081ecadfb5747559e024c0ca8327d62cb5d195c52b111b6850dcd710ea79cbada962d89c5c48734b85a8ab3fcf5f1dbba3b531b313b34f72f535d3988c523e9e9356a1a307201d4f4a121fd3cd9a690cc2f45f193ba9a6d7171;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h91fe1e56d1d01a2aedc623e2e5aabdd04085c2224d2f0f0deae61158445f188b26cb1c8f16f02458fad23ba3c35515c362312cc1a67c173cab26b89cff98ddc60f11d3265a1d10aa4b3550bd9a414e66483a4fb1a9258c5d0d91e03bde37ef43db4da6a7d5196206d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heac411b743669d146a30125fe0d8875fa8a01ff727c191ba779b4a5c68a40f7943c134dd31e9d56f86b4e78e92be5d2d7d60da843555da4a23f80ecd6d1a065c109c16c64d4724800e0446fa2ccf2fdd57fb903851855fed0d86a1472e14ecf0d798302925414be412;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h40450703504d938d314cf4a13927d9a0224bc5b1d57793453eb4dac444c2b2edbf6465b2933ccd8ac738d53082ef7007ce505a80c08875363cc07a98382d2c356d4c346519aa3904db132bd0f63607918838c57e74f77ab16216151310003066c32c6dba7642e5cbc8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5212304277842d306c52352e0709965a5a80c33cdbcecae988749c7eaf6bbc08e49e2fb9eb1121f0d0cce540f9df777706ff6ac8f0be9aa8571083d33ce9aa0e1329928f7971fb64fa4e892ee8e21e67f134f95350aee5f95077a2f37e248ccec0f01b0ad17b2bb58f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c110b670529d2439c4e1b18023dfee995fc95540ad36b0600ab4a7f2c36320005b9674965b7aad33ac0361a8f611a65d5857b019d8a06ddf8615fc017cf0d183753662b4b5b0e3ee93fc176096a0c4b52551a5d87f45e405437d2fd47dff578079d2fa7f9ce9ee89d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5c3b6abd53fa66e1579591681d599a149b3d7e34f12ae5f31ffc86115fc04b0992e807d570e867577bb9a7ab40b0650b3c668ed47316d483419e4a053acd9b2efea802a4aca4069b526732c6f36446bdb0780b54d57070f87d9f9dfb1d35691034f807b3d1616e57e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2d201db17fca022622115e21be682cd7b967a2d87c4cbfa73adc15b45cd0ea197c302577087a8a5bc0f7d28851e2e9c931e31859154351d2fd1d38c5778a5c8e8befe564a958f2312b8d038a530c710b87f5ab822b78b582033e0ef2cabe059320f0a48ef53617a4bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h110953b7349d78a16477c65b7979a82f824f343de0cebf05f3cdd55f67c29494e5f1fae2f8375c5f96480dc2eb6cc8a6df4ccc578e23277620b58995e5a01c299c4833591e39288f9bb5655cbfcbcf7b7d0e4f02a57aad8e2af537b238675ff7145034727e8b4f02cb9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16743abf25d1da5c9c0a979479bed4bdd7d13f1f8e32940e73d6e1ad669015dfd72ed1c84f3e7892c4b20fd7331bb0a46d1fc8b02d1ead8a07113e63633a33e5acd39abfc9a69645cd89f92ea6d998900979829dab82739f439a013b21d55e7a1e425054481a9b72c86;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hce686c4a5ec0c52b08184f4264e42d00af079bf7874b0f76fd17e3148cecb2b8521e0a29f8646edfa19124e8a3d11fa03b11f80f380839ea25f676b9d495cccf6fa1479154dc7190f57ac9cf2dbbb098434b493d401e5c9f0f97a38f8715317842ee19bd11a5decaff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc2fd1787d52a8ee7271c2bf9fac0af5dea016b364899d9110883b7bb54e4498ee6704d813239cc944adc6e2993c5b875bad78d2ea8699dac33344cfef5a7cf7cc450a735530882e76ea9a725452632a938f50805a2a38f1e16809237576475e44cc3fbefd494e7f66e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9be1e59e7b043c8412802247ed1b6827910e77f7f45736a89cff79745a6f41350a3a0bec2f38cd418bcd3336476027dd7c200f9d90ce81405ffcaac44da3d40cd467d261f405f4faca62f64e7b3333401cad20a94a700c83a4d265acd78f70d0c5016e2390e12bfbf5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18923bf38f2e4d2f811ca690ba9ced6133051cdf36eb0aac286fcf6c904debd08b239fa0eae6e81935ef558c361b9d5233f5e4c611b2dc533943c7c457c6ab9e532e9e719f459d06c77a537ccdfd212cd7f293e741cbb403daeeedcce1da30ca92cd680eb92be014228;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf110edbc5098a5894cc320d9b33a38a14c7ae5c18276c2886763cffbf07ca26ad492259d116a82c26f56a94aca9ab58178aa5718c04be094273c1bb3d9b45dc96cd66f62ebaf16fd628d5324d6210f7454857037936aaf4183247cdda85396a079ce10904f9571a9e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c73f719769ba1b38a40628a368745f5c6651886f22e6279e82e98ff41910114510c644213bf9bc52a48e6faeb767b4f58d80fa852ca01df73451a92bc1c6d7dccbfcd5998988f2d5566eb4080b18e1f0cf9cb5172a747912b00ab3464bd14599d6e5bbfb73b81e7495;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1244b13c5726d2471ffe216a17eabd2208d6baa3a80dae73cbd5d75e6a6f3d6375656e693df0a1d8606248908b42cab80faa59991dd82fb1440789b1dd8a2eb117efdb0d86bb3d3eafd81e992849ed9c7e11c258fcf8de30cf68e06b7e469e102957aec90c2c497063d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12829c6db236035b3819b8302deded28b95df6ef5f82e44694fdb8d2266ab69072b57ddd050f994d56d6dee383892c63da741da9c028dd0d295c4ca6eaeb00bfd5566dfa057bc8e718f6e7f864a0fb1b6f7a3493cae56a2ec6fb00f31f7b913c2549719e65c59890258;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h682cad236ed74b284fa609c1f398dc45077cbca93b30ed4a8701ecf7ff91bc1bb313fed388fe9459579f1b976ba2ab6864780d60ea40eb14c4ae7a1a87c7a9e8ddbfe31e6c0d2d16b386c6b3df9946a5202af578354f7aa1225742446e1ca28a9767cc8b3baa607172;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he6474f6dc38829f7e42bdfcf4056e5a2b98db50ca13b71779623082caef11103f66670d70615ffe9465195042f26494f4f807100b4bf5160dedf94716fa314e5c359585f76d2e5b8b72e9a5391097633436dad282c04e8980788e7a7f8c8774ad7f77b2a184b10f330;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19ee4564a8e48df42f78befebf12af38a88cd34dec0e7698359ffae16754a474eeadb399ecc389fe91e87c67a7c56cd8d8172cec350226aba896c91293daa40f8db403749fceaa9b65bfdcdb6dbe044d39e46be8e06bcaaeea9ec042dea52ca18d8b6efde37e7cce82a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1870da8fe9c978faa38a89085a7925c491a0e9cbc96a0a7d9d3222b93ea4b63e77155601b5b42dd3a2a0dcd899d957123c30e8cd1b1f343b660659731acaa0b6592b1f966e5a26429f74f67c2751087730bd06413973f3527496261cac2a422afef19ae1b20048b748b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161a635196689fc2822d8ef23e67a13543ca62c5fa17f203ffa1755683779b2f3b6b6c89b78bd1e4b423556b69ddc0e737fe85d3c864f15429a67df23f7ffb700232401c38d112607d6b63d2dc1deb00db74f6473ca42c72dce5c82a4b088ff93a56a45a1dabd24dbc3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc07a787e77133d0fba5aaef86a6fb25aa658a9bf6e22476953c33c4eb41bf8e7e7c23c25b0850fb28c4e8489c52a1b5e3c36838899e9b3603762682214e69c81874637232b45749ea8b4f184cc2c06bb6b4eed7808de796cee592c75a382f4b37e99bd3be6a4e5db3d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h139018ed5bf45fc4328cf516fd02344daa0a213080c7c91d069ad4931e7a00baeaf37ab7c66fab6d53b1f111636dadf447c654e09dacf82fdf8fdd49252f3b9f0be732ca6be65a9bbf6dd2d68118609675bcf752d59ff7489aadd198f48c9b28b1f85db0795942996e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c5fc091d5d042da76dfb8c9dad591255726e1d719d31c9eccab260f36aa5706c24d013a49b48da3d06f7fbc52a6e996ea594c3d4aa329bb385651d0f0e0d2fb7ba6e1e19f2829572c9e4fa2fff386e1b38cc8f1429fb51b28374dbf6cd866d26a498730c5ea991e78;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h44766b5f1dfd59846cc46af1c354bbe9bd49f2578cb29ad2951fa7d17a071ef305055768a320155f2be5857886d9391058a97c23b881508c45969262afae28bff41b0ac19c62b1f84512a4e7c5cc1b95078b06fbc9461c40a0b4878c8311cbe58a32fed5d8afd81ba3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19fe36e71679c1728dc79f794a64fe72fd082658c9d521fd8c538984a65ef2664823b034ee636c4dafb81730bb1e0c6fbfd8189c56ec8d23be23f0e2151c71217a089cef994833c4b35019228acd4f3b65eda6836249ed44f0df0dfe35781ec2b2ac9e5b56ad7479c55;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he933c5679fee163579b828187ecc802d089695b8fcec16eef49388269664d1f6e51e113640c548aef10c4e66f60b763da475ff75a37e8b0c72d4f60e9158a0b0d186c0bcc3be9654d8f131c913c16f5e11e2ee4c0d5a4d482d893c3f63f3002cb5df56f0021e31718f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d58e97750809c92a9519a1679fbcf97f2a46dd58599b8e54e2b76482b97b8012be963123f86b5096a5a6a34c01a5291c09791cd617a54546d26b99c230193925e8509b988adcfcfbe6b30017f42a0aca53aad5d38e70b345c3ad994aeaf5d66513ad68e8ad6998445f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dcbf05c851621c910b1bf3e88e9c5a5f18e8d783ee50bcb79bb505cf6d9291ea887240f02ca56ce3febe16a4fc4dfe515ccfbc29ab2f015c0a47e391c22b2c81b070d03ebf3da81ceaaec49ae20edbea7e059bd5f48eab3fc2aceaf10f6c9830e19f88607a1ecd1d2d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b36689fd297bf7d3c2e9c719165b37b5a991ec6c1badbabf0f46b22b30b4d1aed487d9d547205f88022642864de8c5ccfa03214931ff3076dfed729cd11b4579943cd6bf1985cffd24bfa63104756feb92b7004d671e658ca7010f3f930da763f49337838b3054b52;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h138434fd5883b7397f2fe8548b6542a69ee6d238e2592b6b6eaafe612b6fd4ef78d7f3a091cec01e96ee51bf8b6111216f144d291e128cb787a75187663eab50c42d6a6275a63672222d262d0317005222878ff90d319b1cd28747e87ad13b402d91ca9ca676c713eb7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h104a2c1493bdd9582a656b526a9490318a192e36c745dda6e19826092b87463aafd40f007fddbe207cc3a7b186cd540d28b5bbff1e6411b94559b89703e98007144b7ba9c86f6068c4c6580d78aff3dc872747fbdd37ed0a16670ce47630b6de8f61680bbb061a0d21d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf895f4aa4679249490acaaad14e2f9dcfaaf2e022f221e63a763f467e71ded25112b9b6456a2fe8dd86c4c2d48eae2b340b3a61ad4932de7629a14b6dad37f233b97e074202595f7beac11f2bb125e137ed53864a2e47ae76814c30efb0c03d901da89ebc2b57749e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ace7384e15f7951867974726f7f569e52c7880022f8230f9f44b196fe59b03d7a7a1b98a3a32a7ab4f320dd184eefab2a066bfe8b4f936187ca34a893209c9ad88831dcedea72d2c46fcb7f58c38d573d55db39db1f8380e5ceabd4522100ca8116e3dacce3e829cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h129975041a4539c6eccad14c84bca3307e8ae44caa5d6acdd31c492e530696e738cc6d54c477ae4d36028cc0910235630236274626312570c6c40d0633156334c6e92269a7d33b04aa70fa9151cb0ca110999b6797b74e74dcf76a65904ba68c8adaa6466ecfd0498d5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1afb7da3ac8979dffda4ac78c85085b2a02d85228430da520aeba9e9c003c4dc36baca93d76344d1830deefa5b465c820f786d6a323d2d9dafffeae06113ce95155a3ba26c71a09f7f3059fa49f06a34621d5b69bb8c8a5c9dd2e60b483404eb08aa16d2c25de9cd8fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ab47677cfed12415d8d87cea31188804d4c1003c1ef16a2a64e57eedab6b792ef774b836c4fa5a776ffb9f03cb972623d4271197e4deb540ff5ebda7c396ef04fd669eccba5a493beec030a1e9a42f9ad93224b7b2ab1ca1d48d15bf3db62a4168ca4dfdbada790f6e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f4de7a4d8a960045376b1301c4deac52288f63432ef410c8ff248b5555adbdf701ce5501140ec4f970569a37c58c74b8c2eee45caeda8d37d3c4f3cb2bdb101fc428598de0b76aa3d556604e35b8097ef4c17565a3d0e33216b8c25b4cbe96c154d4df824718c0144d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f64c4dfd007b790119313d97a76fffadce1d8a0d0eb601ef33ead313f3b135b06b2b0d9869f28843acbf15084a83953626610c0cbff6facdf97e9dd945d994bb95729989be03e2ef1ecc9243b079c492693a0f5dc8d9b308e6315870dc84821ee114a9c2dd3e9f802;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5de57f464b974488d8f3fd455700d396b2e0f191c109f326a6898bcdc3a528f75ceeffc437211d62e7445ca35568879a0fdb091992040e0c011d8fef6b940f4855708173fac3064718e7233b234d41cead14a192c58a0c4e8d2ae55344c6e156f91d819c6d3b0bb1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5808a1f6fd56a32d2a3c1ed9bfd4aca6e0717771835959f94c3f16559d623e1c0820a389ba358f6502e7b76c09d36112d3bb158a3ec54e4ab17f8fef426783f3604e6ccb2c68c16064912aced3cb707b83d9235d47ef2457acbce34460cf8ad4f5e08db705026f412f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h171ef0681cc079f81ff50d318f930a663814ada2fd138ba611dd0952fb954752802887a303b9a3e7daaffa2dc6f25dd8ea00b0eb0ff3baff63c54fb5ae9525e1d8039880602d84bd52099131b1f96c3123e17eeded47b6875f54328c029645d8885fb7bcd2472431129;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108c5f5d5325483a084357f2863ff6f656bb1cea789401b28be45790bdc7bbb05ea3ac17697de760cbbd416412a9624e67f319c3c4577c6d142fe53cede545bf6eeceb73909100698fe3a3863da518f14a3c62cb6d75520f1409b2f60f7f9de4c6a13a857f67fb49fc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he4d665d618cc82561ed831b42e58d167a2b247db2686e335f4bfcd347a2b1e08b91195cf17f89cd1d4d9dd41da2f41764a33460df7adc2b8089d161eac963234b1dff4836c6de7871fa91d65d7fbedf03644c2e77b4da0ff0ba27ad009c4a34c49bf947538c38f5c4f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1abb0b55ea48b31c5090497ffab02d16e82bc047027329e25bba3d3c841a6ca7052c1072b03577d0bdb356daf3c940ca07b5069cbb376ecb8c8b74e681671cac2404ff61d7da26b524178a855c29982c134ffabeec7d625192bec003ea84998c0a1d787006d2681645c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfa06d96922b2cfbe2366620f88ac8d735b3b2f9f46ee4dbfd8f6aadca6f5acfc816b027c727a5b982c02f58fcf5165d695346242a9a6835474f4b32074fa716ebb98188f74156845c294a42de522094f56ec2f70581764f7f2be8a683c120a8a27ec9c1d4f6ffbd85b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f0ecf5cba8d50d3a5d56ddb789dfa75fd4b7e24737a4958e814192f624ae5df96915d955e82b4554798a91c16da0d72e7ee21722b03a8db922ef87dc5affbcd5b35366359030d44f36835dd8c99759371195fba7b73d99b2633aa9d14552396ea7ea85b2a6709c8a52;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1567e1d017615a0599cf2e4035edac1b55e550e616694d9da8b44fa78626a0ecbf27c5d4b4122795832ffd0611f0378c0beab10fa731b09c182870b11be784e448e5c8681cde67467b33f287add8c3b1ccc9d777e87abcd2ebb5c73293061128561925a239f3b2b90c2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7dfa570ea57b3c080c0a91efbd9ead298f4a14e35a2fc196caec488cc2155737a9ee638d56d33350f5fa4b50b6be4b6d61a41e63777971387f81260d1cc4ff44b1ee10db0786e6d585d74ef842d212b7ebfe1e463ad36593dc852e401423f2bc7fb7de9c3beb5250d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9ad5d69a927d484dc5bd3df1abc505103c4b22cd5f7077d1ebc14d4e8e4d23db0668278a38bbded7f4f7bd935f8ba91ce968f32a058cabc217173e68d9b281d70a6791ac94d5046871d87131b9b07bbbc43c2b3ef4330a7383ba28067ee4aed64cf791593716a173c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1100b971724ee1b76ee7cad6934feb5ee271767c0663373fbc10f3b82552c986908a21ab607b71732fd8c5c59ad5968c6426cc8b607dc28f0490dc07ce0ec8a09b09c5543c44bb8fc33f632a602d8c321c1e98442c97cf582045dfb3d91b0805af39b621a956a463802;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h205ce381a30ed608119046da4293f9504a55a3b05799e4efabfd5e4f1b76db8e4550d5ec174e1a313de20eecff59eeeac2c026a4ead4829afad7d11f2efb6caaa81081446bdd8df688b2f3878fab334cf11d07e6598576517d9f93dafd4a2dfc1bf709c52553cc8e6d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d482d3deb5537cc55d28d9469f61b4654a93329dc436c54dfc39286da723de33e7e357211cd65349f532321ae73bc250a3a3a49ae0567ec4a9da1b15e2a1a923a8ecf310098aff06a5e6445981ec6d27b05401d1bfe252acddb885c82ef9ab6b0f7b9b7174652acf5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c2b2f2ada25526f12d0896fc0fc0555375bd0e24fcd9be0eacace8fad7ad8ecf6e35638dd48ac7e67409351554fde53266a6dd660eceb0456d5ebaf44912bdb06c5f4c0cb20dd357e4edd43a2babe572497926aea4fc674dfb1883f920c63cb6ee4c6b0b9358e6dfab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b7d4e03be7e0ff2f910ce67720079ffab0db612c190a0de7eb7b66f86c0d8f16ef5304ebc349ae747fa2d3121951f110ea2a09dabae67166483790dd7ed1585c772d6ac96a1f1789179b037740b1499e9581dc5711495a35628082b608dab70ffb07266409e033ccff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90c9d850fb253e734d24c431244c9ef6358ba1e188142cec5e5dbd541243bcf663b15f1bfecac245f5721433fc69f2d803af530d690661c3779faed16918fad7b89f443d575689cf191c5c76b471c136772d0c9bd5a575f60235dcb07d4bce9099ea3cac128c9e4e9f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8b23b11b263567a1bdd63abc52bdf09802e90c28ef2eaadcf8051050b55a1488f8a352b4aa85536d69299e543ad724b7c0bbbbf21b0250aa2a2b05e61ba347dbd616c4dc287bf4519828ad3d4a41b48df479b6557f6711e3bfc27f6fa9dd00f92a8d493d4ac1fed3f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19b3e1d98bc27463891047419976333cc998a6ffd68c4bb8625ea8bbb8a8af964fd43e91744518969cfbd05b0cf73c34e609cf45797ed16d2f46e3584134bc6d3ec20beedbc5ddb55ac7b4dc836cfb997485d4f18ce2aefd5ac6254a9c2094e26d24d933a48acc25934;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6db20877fc9ae823f2b772529a523f6e0835ea95475c3a0d713f230dee9a97801aedf8df762d38113d51894a5a131db13f8d154b47fc6f457787946d730f2911dabdf1c7e33c83b1cb23dfae2d31025ca3575d4a51c38df8497977d75594ef2cd8fd3470bdbf093945;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed6612517d7210cb32e52db6a938accce0b375582524982cb1280607815684b5676019ced70e91d24c13b6ba58e0e26fdbf10a73d1670b985cb6f7ba956863762843509aa460c3a338d912a10c1a16c2b80abd7be46b8d4f335c5703efdc7b489ed48ad5195e495477;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc79e93e027e308f42d70a93b20e761bab52dc4fc0c9f4e18e4f5da89993d4c1aef5526b458e5626fc512685bc35f0e426e8ff6b6656be0915514f4672cf7f776182736f544b507acad7556c0d696dd42aa5a270a914ccfd8fc0de4d4079c434ba09543bc2d0a76cf2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he3a1c25c68be3f0fd1da3bade41184f9dcf9711e98ef8824a2fce58404182773ef76a7c33d306b45c11117dbb3ca56964cc9a0f50b67573a212687ca6d5d210597b68a0ae7f7b87e8ef9b2c60fcc3a077354ba54a8d8b57f043827798aeee035610cabe92cb56534e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h928d99dd18ae981ea839960e5fb780ffb87d78894372ecccb3029b2404254db95c90ddb040c64ad75130492a2b13940bc591bea30dab128db4d88053c6a274ca152194de429d2148522d3ee0678dd3bc61afb860812cd9fa4c2966eb2cf77dca233d2003ace70c5d83;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5d0beaed15eebff220ef8c2d7ce0d9d32678bf94a212645a49103461d1734d53006b8aef50ea2ff51ad36b2ef3dcf822983c80da4f7ae8922bc555a6345dcb0be828183d6868635447034dcb192783963ec28d32523122c57ff9630c840eb11895abc8cf4a9353e407;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8e56b5b15ede1bd827bb9aff1aecf4ad0424f2a3ce8c7d690f0fe54f992d9419d574e12ddfbdfd74786081fc28a9d715d90c69d2a55109421e25d2ba204e1043d1c51a7c24c2c8678f3696d5591be00929e6ad2ef0e0338cabc320fdb74714f5714e679a12dc3570c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14de22cce9c18f0c9e10a5ec40a8cab63fb3de184972bf580d6503899a944c4a5343012e78b55dbf498db78e950f26c88ac9fde8e4e5bbfef8bb0320beab9c51bf7be3542d5e530c9fbc265042a5cdd6fcc1447e52adb0c06b1409f7139cec8af44d868faae9ab518b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ebed448158628c44260c5e8dd151d1f5a49929f54a468455e3351b01909da127a56fdfca5cd9e9442049c8fc42f7af35dae2a8faf2927c31b96c01144ffe44a54e70d8c22ae9a3519ff9c7acebe5cc6b2036693d1a22e1307f18cc451cd8cb82acd522f1c551b528a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc882b17e55c0a445bdf33b8774a1883f41432493e660568e3517b2e57261cda9cd9eba344ffc251127a8bc8013f868886c4834ea5a8ea57a9639141d1c3b738ec6cf51e54089221bbbf4ca215d529393a9aa55d09e8f63cbc782e75769ed85eb70e2b9b4154873c72d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc065252bc97e1f50a7e060aca8fc84b6de24cd39f40529a4be165b3c00ad5f8f1ad91d00f4c78e597188a4bc59b30cfb16497a6fcaee629f461897e0e40a0f960add1a91fef134eaa9f2aa03ce3ff0d746e3b8d719ebb39ad1a26c2bfaa3433eaae6b3ffa0bb7e0039;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc78224af7f8a9adb74dbda43b0abc0df7ba750c1bde40a2720fc61df3b07d6cd83bf99de91cbfb19f8bff867c67e9790da99a306e7ea07409b31114db1863f48195115413144211b97e7a4a80ce859968edf197048a7c2174c23ee845e050a6b838fe231d92b28a79a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8a310efa464b52733cacfe41cb268e7f699c70e061e49e470a830708668bae72a34e3fe45ddc958fb8d8df77c47af9d6b6f086832421095b61409663dcd7c92cf4748c800743bb8db01cde9d3a082d1476ce2a46beee68bda06f9b645be3fab0d63a604f1f36808031;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dd4500e74a917e3adf362cf5d6dd4daee340a1f5a5dc34f7a3f2f6cf045001f842b0d73943b76d44b5ab440cf650f98f14e8d0af8a154c1547cb3050561dec6dc139964b9b609e441626ede7da78aa88069ce22100916f1177cb22e3e27e68b8f0a5f7a558a2c7aa37;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hda6f0bc08a8b8e225bc7e3fb685f464c5d6d25e05857c54a8ee42f1814b9c8a7fef8c859d432e77997ce8c88af1349080b57fd9dbf2b899daa444aa86e7c64d2a5d30b82e6c96d384c9cacc0e66c0f7d54323a825babed3a251611da68415383ca799d58001fc7c29a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h92fb867f6b06b6804bcbcdb7c9486c4814e1cd1c9e8800edd650c05221b7bb92bfbcfb48a7508bf992ad66dac99bf0cd443b5e698026d838537b2e858c76e16b1b9a13cd8380639657f38b6737d9bc2e8daf1e2a7a076207d9ffb75997999f764d9bf44b779b1f8643;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h99e922eda391f190cdef1bb4e15b151b74c6ac53adf7776b6c1bb1d3d293f7fd96cbe87aa844528a44b533af57b6104052aafa5f9073ce697760612a01964b05e0ead76d319cbe70405f9716846affc159a91a24f502bdd157196d91339365e14cb55ae3a51d01cea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he22214528791bb3845eb134d76578a1a93d65307f08a06ea674ef58f7f1b2b716028c89e4707eae119b275ae2cdb515572554080cd60a1688680e8e0a897be63c8aa98af9c57826742b9b03ecea1d5395d1a3f41415764276a02171f3706e89338dc2d0abe3419c900;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c28e3d0d6e34777a81aa19e62ab1481112f454f48637cc966d3fd9f09872bd30c410aeddca17d06c0417acee0492dfad15555c9f6b03a16ba4e668598e4a38bd12fb9a678cd34b97527ce4f5163520e3fbb7e2381880fc356bae366f96199cedbefa4fbc0ee5ba0cab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d1470425777607fa11843c4f2605f62493902c700cb89d6469ce4d0ccf1d556f6c81c6b6bfa3d9fe4cd473a73064cb576f7fa59b9d34b8b7a5edc3e035e6ddfb2c29ac5cfc375610c7ed4cc9ec7daef7735dcd7fa68c925f2ebc4816620f53c2e69c5c3a23582c1c0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b37dd7483b872b5bda583a2582927f2b1af0c0c692d42eacfa59f9eb63a408b3cc10bf5a78608b659bfc99beaedc1162acc8a0f7b42ad0dc60248916e9a6b755d736c4f7025ed4cab65f49d42fe7f56ae8968ce2c6fb332bcb6a67e91fedfbfb2b288b1d46deb2e4e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h368b551bf58c0a67f94e974f2173793565ab5bb970865993a6c1258b1d644ef36c17cc57598b6683d1c609b213694f7464fec8785137f005007f7b090e78366ff0182fcc6d6491d5c4261af1c6aa7c8acec47deb94ffd14fe92f306681069b5381931cddc19b88f6a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb95ede526ba70a7ece2a99cdfe0f414dac05358f66a5ce884b4aa2530ddb628ee552e430dbe5524bb255c973f289e72859647cd892704e2270a777fce2fab2c44b85d02682239c035f3f6a59a88583fa0d214d093bcbd4696d1a43dbeabf57c270c223c59c49cb890;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2d02f524a743b3597f1c9041cb9398ea4e2db6f7d3cf3de9f6b52a93cb6722fcf24a9a6e7c123b8c96c92bc2d9b9405ae081815be50abd6fb863a00c3f11a2b16aa3a32cab55ca8a6c2e4f4abbe0eb14fe6ccb5b5f6f722c3d1c347c09dd7648d425fb09b52758c05e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h184b10939a90b0f577295118d047bcc95cae38246fc49661f3ccf5afd918627564c83d0f46fc5b2cf12b3ceb9b05e23ee77cb83422c6c0dbc6a97731bc6c6932cc8bc5114815bd5dc4d35d98b894fcd83c8a3cb8686abf1c0bbaead3801efc9a925a94fe37c2f69b85d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h642a0cca87009c0a30b04a42767a841c2cc1568b11efd9a3e688b771f4a99dc04113391508791e1eae727c491663b075d14ac226f5b2e2135ca1ce6996a693c352a1c2301fe81a7b031c77f2509d6f2dab970266c94c5b1d917ee048a96e3c1e505d72afaeac885d42;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d6fd54de980ff966788e0802d1b1404210c1d4c4df012582847a0164e431c60c4d57babf4b91d0c1346eb351878dee49b471507c92ec08e6187230e2bc2347ef5232b7bab7716134af52993b54fb95e2cfdc7199ad7949f3957b61c9232d879268aed0eeafbf92827;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h294736c1a23de06f5b8397249ba34e5f7f5fa3e6b34b5bde77549ad06e39c34c94e89fdfa47a3985d4def3b08e8a57270004232da5815f448a54e703a5afda8116efd70bcc78fc39517878de88888d71af4ef286801620d2c79386e96c9bdadb1d0dc935bc2ef72757;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd4d6c69e9521487656633a711c1b710cdb81c2201e0bf124c2e60b4595e44330eeaf13f5b85dd1d32498fa11d960268c9fbc52ce2acabcbe1b6b4aa0741551b34b2b4c9808541af8ab861e7eb3506064e9b0da83b5b3c0b208ae48834426d6649e00d5c5881f349bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1e3a1be9837ff967b46a343aa6b640f1789a22cf505853ad26ae3b7ab650f426a2c6c21ea8eb56d761143b115391a5f260a593c9fc89ec98e3fb7a5b17cc93c0d51036fe55f86431c1df4bd7613da2ba21e4ce3ae4915e05b15d9b1371020332ffb4b8f3d1029842b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h558b241460262537e524718e7c555dd64b7b0ca5988055b57543873ba03588162cdfd75eb070e1cb541270a6c521f12a392a7778097044e7f092e13643c3dc03b342b6f9e6bb761f8b8807d4dbc2046a39e5df57178bdd460184c5f6ea09a8eee621c5624338cedcec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h280f582121a0e298038ed234c4885af139f8b6d0dbf4d8c06e780b770527362983658474defdeb249152d9ecbf315483017cd66c476f6e298ddfda6ce16a05a92755a7e3206245506836cf35bf9590ff94ebc4c0c134eba280a701500caa5014b68877a6d1b5469e57;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2107eb7532bc0e0d86dd3f34921da2c9204d8cac872d7b61560520c172ecbd8f43c0c4cdbfe44a994df7892699a22e5540dd86cf89bb61126708d3fe394d1b12171cc1fea3f8b8d304bc98f77bf572dbb58d8cfae56f2a7f28bfc867bc89c6a0e364def35635e9b6a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdec0763a26f0a97034fe6c8fb84ec747e647ca079bfdb4172d25f522405779424809a350b41d434a6015b8beb7ef1cdd56ce1fa053671c2afc7237aa4cb73f13e96616352c61f7a1242255fe30401c49c644e875c4b27d66f811a05412b5e1fa1b343ae5494e82de73;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17ddece271bd1e04699adbb53089143c81624055470f37a6cfc00b030c366240d293d454bcd875c7f1386b92ee72e8563485be70a43a895ba5645c08ecb52ccabee78d7aef331ab11a0ea122d0458880d6c5564cceb730da270b82f6732ab87e1f1686e66431efcbf60;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbc028c102bf04e138c50b68189abf8c869fafccb5732b335bb68d35fd9840380db3aa01c3a6d8b55c84b5d81c21bf6ed54ca18542c6a5da8774f63dbdc246150281208dfe46a854c8c58a704d8392652b95f194ee3460a8d5c856f46bb6719dec7ec692e036e676eb9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15e13136866edc93f0f2ca8d8d22c645dafdfc2b50b78630d29529b4248b62942211565d9d1fad5934573dd243ad76903295eb90eb1d583ddfe86e642ef0849af87a46600185370403a8c90fe6e625eda12a707f32b37eef941f3d00deda65c4493a5e1a4853f423111;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec7a1df751cfebcd3787c6c000c2ba2b9ec30501477dcef11c4071a73fca3fbe01043edcf1f76b0fc01ac3e11ec02580d6227421e2901de4f917660695c9506d35bae22561016bb04b7a9f9941fc59acc20b6668b063ca5a7bcaae5edf50f5a0b15e2e167b87724539;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3a6e7f59b711d319b942bc7508c950fe0014793b2e93053a733a9d51b2ee144f90c33ec7ddfd0416d4a1a3debbb02dab3605fad3186d50f21295ca71897a00b70e35d9b552ad8a1b2928b82d166db40ba4fed188a56dacec53644b7d8394970c9ce43c4107ada9a473;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17dc5e649736ab572754b7bd32d857b05f10d184b33a8768a7222874cec6746a364fc5298fd67e66371bf70472cbfe83b539ad70b450f9913f02bfb305a7df0d154b8d4241912622a5b22cb32263d736230fa55a11978647048746fe16f782e1636e7f5aaf05477848f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13d6edeffd104324b66c72317edb8c84a6dabb2a9bcc645ad40ab36d7aa36de1d4d087991614aca8fb45311c08823e26c6c8d34fd16cecc07c512467f884513ae80d976b61ee8e577676bf99dd8e68114b518974a091dfbb9005a5f55eb88a6f7b07358191e0fb8bcd2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1628288a604f4af607b3e5c2f89774641c9077c66cf8709c8851235598f02b35cc277b8a7a877e2025c1a827a6e78f457cd91227ea95fe90c895470e620c463e0d86332c6d7e97ddbe2ed20b3b640d5069943def9906aa320e40e0593952b87b5a3a3151e83c139c257;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc633574979739ee7c3746e30d1728b9668d3a3003bc54fab416d53ce3e7ecdba2717b76a8865d916996fe5dfa391c444d09dce41f2c2d496d90432ff3657cedfafc164294a7664ca0c561812a3d096b6ef8dd8fcb86a22a8c6269f89f24d275f8fdbf39fc29de286ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed47a94fb85002c6147cdeffdfc2ed30ebd127f238a1764d6f1c60dada28217e2a2f3cd3e1be30592f06bdd624c4818869c4c5e872298c45e449508c40ee89592c679734f17fe52a6b7375caf10a12d16f07615cd50ace37c740bf7b8d883837a0f9ff567c2b51a925;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h172835269028d425c3e96e3e2293a73344deee44bc49efa752850ef07f44dd5fa87b3e84ccd32974f5c2e52ed98890eab26234b75d0dd5dad6c37e96e09c2c99bd8440c7db9d837ea10f388078367ac81bd5dad0963398c314cc6eaf7ab1bb47342ba13f0296edba719;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb36ca791aaf6595b52b13aee8ef66551fa266e13a493ce2b2fd9e68520e3d1cb35e1dce6984c7e0c5a35f1fb53ae5ab8cb3e0883e6e73bd844b0554356e5529b8c4a8e1be25a3e03428e9e2220f51f2f1e4bcc60c7e7cd304a87311ba1ef985f34601c8f408062dba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ec774200387f56113e627f14208940e1391bb96b8763b46da33b6aae6f34b83569099d0961322d222a6c5f3c779e7460b6857108847d545fc1d1dbd2dbc0ab44970855157cdb4c321eded32e3bcd33f3e8809843c21d2d8e931c0be43edb9a8388043fe3ad2fa16b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffa3a0e1193b58ee65e8b263ba9694875f79957fbcd6e1f5badbe49591d6ed4c51e1568a72c9bb0654a086bfd1459bf26b05d40bea33398f54a2f8915b436e4ce84bb8d4d33347a3e76a8d378205369d8e3b60496fab23b630e0f99ab47854458db2689e7bfb038d68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14f6c2e3969877f1f1b9411b5050f9f1138514d9a294383f99fbc8e8a712d3686f5b54085964089db68ce74a587ba8006fb77f4c66035aece58dc1d9d9c430fc8395056a86786e871d2d8cc03f0f223fb616f1ad1614abe6f5ef70824a81e84fb8709c94151a4c706d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10ce44d1248cb9a598bddb910fe78847d0f9292854112087b802d768d12509ea50d9454cf755f26314410d253bfd846eb2211dc912ced93acf7d6273f738a0b0edc12871d0a5747440b4fb5cc4eefcd831458e63ca036b4d40eb85dd1e481da93039281ad810df7bed4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h663a982cc83b35ebfc5a5e0a4744f112f1008dc223158634e7b9505d060ca000ff43339a6033352f28ad5174bc74e6c2936cbec533e66394a04126a288a084baa4b9d0183bbbbe75fb17bc0f70e93fc11a8ec20e898962427a2f2feb84f13a7ee9514330df7bed5ec2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4987fac0d2230eb385f195164353081350796cf7e162162aaf6336fdbc695a443c285f01b88cdb2984d5132dbea18a4467c23e769fff057ceaf1981ddbbbaae75e311f81b850a28bdbd1dd9fbac38203a0acf0f6c0e0bf00d872172843d6439ac64411b19c6451e85e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h124be4ee48c52f8aaa1423a87e218086d31be52ca37d59fefa3eb0690ce2f42dc0979182be087f1cae7983faa7fb729fb91b32b4ca87244f471405acb0fbbeaceed081d45f8813b3bed261370313e2b0968b5a21e1fd14ce9124d285fff4ba159d327a4e62300e39a4e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h162841bb9b2d262140993e0d23029fa357779d5be7693980b6e0d9c6ac10d38b94db379333376c2363f1e6e377f19fd907cd223460918f240f6778d7425d34e3ebd647b4ac86799f3bc297bedc8dce07c4fb58f993824e9bb3223ee6cd661eebb7d42fb91012d3be040;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h159aa33b1569287d87fee6f6c5c694b6538a7f7b417dd8b5cd01ae0f33d9a397a15618b7e0f98b69b423948454a97372e13cce1a241a52a67548c59b27a3c42fd0a0625984ca286bb8099c8cc9d090da1c6d175c6e6a4b5b8cdc76a11f21b4acd7f05ca4d4ca6b1d640;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a176a988ed5331c0f62633942e11dfa5dd85e6c60fdec79c8ba93dcb4b5cd5fb078cc330d2189c805ac42ba181307f40a6b05dd568103bc8a1aa2491e353930269f5ded40ef4a6dbf0a26d0714da8c417d4da936dc59c2baf9b762ba055de023528c46dab552fb7d03;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c379ca08c34215a3cd71c9d81dcbe89251e85984a51eb7f05ec077dce2243ffb30d305f56e2fe287475158366ee68ef41a225525e804589abd6856f45fab857ee7e9b510d48b4f5a28cfa5ee30b1917bf354bebfff7a331fdca7b878e2d306df105b9554599336e21;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d14c5fc4d29da1b50fa17b1cc7f765cbc8740e8321d906db52dd66fae352ac97f38b63ca4d23c4564a2bf15afe7b68ac30932acf0246b9aeeb8387dccac88bd081a43e8c76b763ed4699d7016a3ad9702d9436a9f5a87d56aee6ffbdcd732e84ec5851f9fd33e4ab3e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h94a18d41b6dc2597e5b9c46b7379939b22b549f1517daf07ecc8b5d0ff96a7272430f650db4f2c66b6089dd1175021159f693cb5ea49479dd4c8517a7d895f18070e0cebc071a866931bbb38d5f7d8e5b217eb15e1b93c3c69b758527bb69674d7f154fda9123b2ac8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d7626cbb5b613a1bec271d84e6aeef0b1c87df5b54b4a5d64c98ff9901963961a696421ed0c2bc49bd913fb4f6fb24052a527daf720211487f0a0c2b2f66cd2aa7b78237e86985ac46c6d79f53dbdeecee7d2b43f42c854a5d30c31b27d67f2622a153f10f105a5a4e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b7426032274f2d46bf08997ddcf5eec456811ea755651705ce60d35a288a48feee14e3828d07cc9ab4ec62d1cb9b06b6d935df4b8b102936c888ac7e8c2b7d18d736f52e0e88449fe45c129263d9cb73713542df444e7966b6a45cdaab4d4894c9ee6ff43bd5056a1e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14608befd51c9799334a9f6007073b64fcf54689f0fc2b434119e44a3ec633256572d73e7059191fd5b8fa52ca1bfeb31e4d06850fa7036fa4bda90e8623f13080b424bd521ba4d57e4fa4651cf916141b9df2d474f8c413d69c533a3a5cdb6f7b8dff168da7e8b79cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h449477056693ae559cedd08d53b244491be2e3a464a0a5abe10f777a356575a1daeec5134ee1c698d3ceb0a18492bad14741e559f743abec73ecb13b18808d2f0aa508cb02aa97e50eae1ac1800c864d77369ae65d01b77155ddbd1d406401ab9d79f11ebced88588d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h69e3230a4fb75f74d2d4094a3313810fd0f4c3322abc6424cc1fa179eed4effc12e94c16a1edeef5dda0a397d78f1ea4c84ececca3bbd956429a4598f6ec9e6a643008ae92608b9f4225167a466d451e5ba1efeacb2efba15648b1b8aa8957c3d4d17844c10fa82818;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ec8428c9d971dc6c4623114d4db4f41232a2858f0eee6a4381d081e5f3998b067c0005f24ef1c3bfd621ed0bf8c2c1ac17dac6895c99d2e10e15887d2d3ae750baec4ac8f8250cb622ec7c7b8c2512cc2e22417bbc23230b76168b22ffaf4d528ab718471e1cae3fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e307cc0cb9fa4589a8efb25940fabbcb937844603f9e258c8715039817d2db26112f5bcdf410473f24ca824c4d6e5b1d9a1a349a8097638156d3b48fd40d117e6b1ed5ff7c033b82f8022537dd0dba8d7fa0233b171808442dea1481daf6a438df2e599c62b65c6c6f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9cafb8472e90ee9db666dada42008af2a4b56bc8aa55daf2c564c5eda8797d0b840b5ecf4a9c99c7854461f63b3e2daaabc4274a38a2eb5e8a1ff4d4552792e0353e94dd3655863e6ada27b062bc7a28b95c561aaa3c91d3970a235b282fd74e077d56c87c05c909b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h313e8c14a3cc14933e3d9fcd23139361ed926f0b37afa1a0d86ab454004c9f272865084397d87bd2251b11b93190c568f8ac955ff46b41369c84905963ebec6b072c049082019247421561c08ae5043af0d961fcf93616c4aa7a4c4db59c2f9f9f523a50928c21e95;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b98998fdb5718f6c9b454ac7b1685baa6fc1f1745695657ef2ce043ee9026909127cdf22245129a507a1282e706cf41ea7ec11ec1941861007542e640a462b33dd36fee9a601d8abb4d578b2c17c8cd0e3a42c83e3e33e6fb94b26ba5735034d64d1e8f3a1754a157f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h73fb90a9fe1dad3c4f90808dc64b2929bc2636da72b4c0001afafb98e84f58729f5a42cedad54b8a18cc07b78c1281c32182c9b6f11985a10f061e0242449d1cd3ebecb7799192cc4b494ecc17c808307f45afc98d60666e34929c7e0a86132a55b89b9eb7e9d64b0a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h508e79e6eff1ff60edf2009f074842f2e5807a2c7697c6ae065750cc318727ffb7e855d5aded046452d84aea434cefd4cc4e1ee42b1178cfe7bedd661f759f4db4b62d7d3cd938170cc2ba85b52dfc5b52800366a49791682164225a8c6e557ffb4d55b8083d322e96;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1441ccd0754f13b9cb2489d7f83754bd79af10bb250e02cad975a1bd7aad18de6105737e098388b04e04b5350b9f1a7373668c89bc149005c1263d3ad8ade0f1f50730dd171769eeee79dc428fe4bf0e3495559516aa6c7ec9e2cb9e3afdaae8fcd419b47148685d342;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h239cf224d1fc5f4d6133a738b7ec648546e7e4ec3c851a099f1fc6b27e0ff826bdc5050e8891fa759d2ee6d6a46b1be02a9186eeda3cb3545f3e8f802ef5022b4b1bfd298d6ebf1249d25695fd77832ab583d5154824febe85335cc1f4971bb2c32027479438f5ddf7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha71492f4071c14d33d84c47ca231061257ff7fec5175426566eb67e6a20bab693f94f05b78d13e6ea9efa4b24a6837024c0effce4064921db7a78bf25fec9515b7d4f6548f32950b401e90e36d6a2de873fb82495f1d61ebfbcaf175aef3dab5f7c434edf48bc63f41;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f11a1a8f10edb24ec9ddd22bbcbcfe6e48093ffcc64271641fb0d4db90d2739e1c7bc97f2c18a78e86237a491335872dd890bbaaf503f875d411bac1214923ba5e0cb2f4ee38123c974e21c187f21446a853d0d3332302bbff03816efe144d95ec77d29e87bbae9289;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10854fde4597654eecbb68ee504feb729c7bc0979d1a8d83ee382c038aa8eb8eba3f4162010c78a940f1491d62fc29f68c3f965d69e5b863d3f2662f4a14dcf78284f119fab8d4694e1cfee9307983bd4fb080078d1a780d9b513452d3b6127a3433051d47b4e0c33da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h82036bb02fb95f7474f8ba3a70cc9b5a4b14bbc6af56ec3e7861277a7c07445c9859e37320a550867a386c1542a2c5ae7388b1b8ef85c35c9190ffb5e003273a3a30e9d158f7a4f80d59b19b9f762f0e0a303d91d80df1103d25a60f193389d32f3a9621402e467925;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155aaaea0bb46265d15370888614e5db0c85c51d8f43c7d34096adc6d8584bc2c81ff09cb3ca99041abdb1070cb075ad2e31fca657d1620b73f48c9914d2334ef8a7d5634dfdfd445b8e6d781b0f0e1a3aa84ae027905761d483ff53298927b1ecc8945fab90cd38ba5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b2fa1c5764692889c61f97ed5b99b83b899136f00716e0995998b8e024572dc780ca87c1ac63f3f0c61df2447d5b4040164daeffdc1d205c89ab5160ec8c6f656be474dda5b4e35bd91d6f8ffb297587119b3934a7af62309977308271714b60402cc1cfc7a2c0a3d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1430986737c31958d324d00d907182d68293d94b53b7d189a83ec7fc19e6aaa9995c0ca3a0a13af23dce4264b5175defd3ff735c9545d8da0881f2764e09304e7351bf5c62c76592675d88f9d6030ac052d7ea6393767eb92c0a0e101526087a16af5e3d45cdbb68366;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144818ff68bec7115f8ce81b394dc74bde1f16bf3ee19d6f048d629fcae77bb5735ac98656fe9ed0dae11beeb5fb09e68cde66f70927fdd058469fdfea4973068ecb55bd4ed8a6a19eaf8b0969ecd207d981880cb3469f0de09004ba546913915611523185c5bc7427;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c135e9343c14322e7dce57d59a17dfde97e51500ea7de7a31a5602536e6ec999e214f731a8dbdd004874447e2f8710a547e1421cd5b9b7b0bedf779878860ebb21bc85fa4d66a6ee6740cf5d40217d5e1e61587aa34659f1d45eb842c5015e1b4321de6dc9268418d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ae25e1437ace185608faaad90350ed9388a793eaa9b0c548cbf7f7543a6887cfeb9f7b6179cbb13491bd66b56e4d3b84a7e0bd029ac8b497af281914360cfb9bdec7bd8153171c75c849e5a1214521aec06df1a367b35e3df85b4262b8135c8c8c33258af1d732d52f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfcdd897a0fb153e6ba6403c0ab49ac489726673b844898f37f98b96e78b687ed47835591ef9ed4e8caf098afcb646908adb928ccb83099602ba205d49c8957174af45006bcba2397880c36299b8636a7e484e88c1fb9b5b22944c5a8ec2e5b5502ca19fe8156b1c1f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b53b37c7628742a9481e0b624d51e03f67c43b219d1fb165b70a21e5bd02cc01d24e5ebbefd1fc4ca27827a40025bece434bd21fa7382ee548f65abb0ce64d2e4c0559920f11e26bc3c2cd78e00eef121fa83a9ebeb0c6c823074ecfd754a935c15633a5604ca9ad22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1400d5209546b2354876f2e2faa8c7c367bd0c469482141a5ae4bc0f6a5d287b6f1bf1d0799efc233d8293ab72ecd24ec226fafe19cb8eef318444132c20f32e0a700f99419edb548e5963c29c2a353eb86456e96fdb1e6fca5d45239a045eafde3b3e50ca413d1e857;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1271283edd8e7856baede592f0578b326fa09dbb20839c09f30ca498cb35e474ef83028d611e897802eaab85c83f399642f5a91b70198b6e8e8a0b19516dfa3f2163ccd5192eca798fd103b8a4ac08e6b460aed6b60e1fb764e93bd6815928378f627c9cc178f8c5da8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9bd50373215cd0caaa16225c5995069ff6c59754b1081ef5768998de39095b3bafbb1f841fbe3b53c55435ac16b4ee8daafdf64a4354061c9811fccfd5b24a34a56a7c7fd95864abd8293aa61b52afad1af1ef4e452ac7b8e0c2eb8aff3a6c3f4ea2d0fbde27cacc8f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h185fb27c329866ec4ec43c23d35196f29f04c318c589d40a20f5e7f49b26b91bd4f3a266859d77031a78bf688ed7fe76d185e91ea28db19033704adbd91c14087e71d0ef2f38ac62033cad10ecb349f260087ea5c201316a68ab6fb86a5bf26387d52bda4e2ec8303af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1894eadbb5d352200a0601d4e22ad05bcfd80b6d8e1b0fe19402acb8deffcbaa2feb34a534f9e3aa44f8ecf19e326ba77015c5a6aa7121fdcd93f4931b0c31768756ed317db753fbd712fa341a7c753e54ee0746a661e14092ea079a8e213521975aaa9ecfd878fe286;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1377cb4d7e9796129d9102378ab8d5d45a4dcbb9d5696ce3a395847567cfef72de73ae4614e5d5c63101463dd2ca309c2c6d9c7928e5e07632ca4d773a7bee0a225e6f8da801b5f47e557fcf46817d9dc1e0cf4ea1a59a81257b51b44ae832bfd676d18cb80c2d500f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db24f1dbe21305c0641b84385f92d87ba8bc87da3cd5e9d9ad3a912a11ff69e3362302087d18c59b5c8ba64a69acf8c59dfded8422c0938be89accabc66a12953af3354e3941f418113661961895e0bb3de68c43e0c54aa9b2eceb6fb50cbba8d5cb6dc1c807f92fb4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1029c19d69c51699dda9171d550929bd199c3b07f49cf853a8fddff6c0c0b0e814282972d7cc6485597376e4a6ac44b69a951e00515ca5d49028bb5c83def4bfcb2f50a3ae2300f25ba3f779f889ab499b35cf7698fdf70a1188f992a5a9e2143cbccac770493f6cae0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1162b2a9516789fa32543a327190e691498665aec4aa1fbd6d8a80361cb6d13b38998610b071804784d12b9819de9f85c9ad882e1f13393031053611aaea355339eaef7d794df03eb649be2946ce6b951b83ece5a71b84790bcba9b54db2d82163870b53ab69e0aff4e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a833f5cc64a27da6f0ef27a418ace6398b4da6f33d4d93d5625f57d52974228a4daf7d2fd0088f7d34ea44c43220577864d0da347c8066e2b5407ee98572dda459e70d00949c0f83d8aa59008b6777c5c94a183ec741a43c33b9afc258a609ea0852e4a45bd5e02df;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16518e2b8dfb314e2e23b3de784a05a6126144d758ecacf289bedbc73418f61e95db15ed8930e3c5fc56a2ee0ba699df0ba0ca7d219b70834b7eaac2b8c5e571d59735fbca49d02273237231278476c78d9370b547957da2fc4d575827697799c6d48788d1fef929e91;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd2759f83f7a825b1edf7fb0e49753fdabcc0350ff2d2be6576fe7dac4c05d4ba1d8962afb5ada519a470571de895a622d2b8c9edd8f4e0d3cd689aef4925ecf7470994567cfab035d3b56a517a6c1f0a0d886e633bf3664078ed5f83966397970ef9540fcdf85cb21;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15dc89061b798161a073742a01870c2c92662e988b3dd7a3cf84e4e0352fc48f0ae9f06a65db32309e603d542781f0269b0a6a41faf03802aef214a5f330dae06b69893c01e7178aa26497a60f5374c75a95f813a2cc8feb551209978a9fb6656b813964e20030597be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d7a2b0d4e42be63d901f8394bdf903e8b4a42f7b9ec5f8f7b29668d7d46f757e7c49d70ecd26751d8744d82fc93118f344333576707f7dbd5746048c01bf1496bc99374d91693bb38c50d197a83ff613e1cb3259e841bbb1f322b832834073da8f8ef11b694db48b2a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9f6c9d9319cead0554f1f5e7e2da67b336f0e0b4dcfc971d98ad9e95ccafce95463fdf8dcf4f51a265932abaf4ff981e3d8e347adc4fc0a4c2eb53f48fe7c90e15ef2f9371f95de335c4c52c934a1758e9335b07199b90aa4ee3ecd65e7fa949b6016e4557089bbbcd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h93e8809239ed3532673cade0c5eeaec154d3c43b66d8f467090a21d1c461448a6d2e179eb1680392fa1228d78f4ed7057e0c954e07add493f8de91c55de244d42fabcb338f2d9bfe34764aff3dd2d1e72e6acb51095f55150f0422716391a6e91b1bd346724bca2ca6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15478a573c04b9487059716d311a1f7d6dbee85cf1c0bd74e7dbdb2dca352106975a620b3ef427c83840e102c6062ad40caca2813301a2331f450261b33ea5a03baceb5ad66463cb17afff595f6d2d1eb42bc50c5ab98726527125c702392c2d4804be4f0ae862596a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bedf06fcbf7dbcbf50bc0a752b4043770e6141852ec2444daf5fc1d551be9db5fe26dd1eb2b29315655b26fd56b020ae7b4193995fd7cd4c00cc62a565dcf9029d5cd777af42ba7f6bb6cab14c7bf069f15ab8e1b7c4a8f3f25af261944435c21c13a65964b908ca91;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd17b734de5f04acdd692e4fa1580f6afb4043aab7922fbaf3d0a97d4c78cbd073f1e5828d0a38a1610525642b52918e618f68abbdc1ec1604b4d7463d146cbbb1bc76a2b078a5df167bb932a86255374a383cd76e8816ddde119aad29c9d2c429bdf730ef96c68b6a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff1f7645877f177d66b2aa6c5e5e0d823bd12582f785b0776ed3c2e7860e18015b67f23b1904be9d60a644c6b6badfffbbb2a54d4dcf82c9f8aa54c5e7a5cc545f05523cac2529b38d200a5de8581dbec3d97b257002181f876698e2af081f4383f7071dee326abede;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hda9f61c449b96fc7000e5924207c15146198b8a7c1cf129a9b9d00be33195973d7f8c444641bb3bcbc11143213b47487122c7fcdbfd776f4ef333af2320ef184e52decdf2839a16380da2a83057f0633281e0e886a1824d8d8ac1f6fc6a6c2e6ea84c6cda0f3d4fd0b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b6aaac37cf4085f46d69d1b629ce0f2910e76fab09dea9a2d864d6c996f693c5e2b0739d84966ad48359b4b7a43467c5639e62e4a4d213f42f4ce6ce5d346125fd08aba138278c17f56f2d63c93dccbc87c4f58fbad25f7d8d2233dcefbfbb9bcb079f6a2de613ac7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f6d710043db0eddfc6a549c780a5635ce7378eec97e626a351e9bece02231c20f700828df058a4bb6d9e741ca6e6bcc14a7d4ffebea849533528a2f0363186bc2dcf5a119ad03f5e00bf4456185ebf68a86a4e3033249113668e10f6c849c406dc7a8d685a7b67a16;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ca6349126fa3e5c589a287098d7a188fc551ed585f74f2ff2f8e3f3ea99eb28547e1eb5fc861ad8e0ee2241de97362f80190f69074fb3133f195674ff1f057c4dfb9970b5f3c3da51b5180fd66a3cc124fd2dc3367052c74b39e88465c49fc54a618fbabada9841f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c9a5490fada91afcdc36bc41c1dccec16a6cefd512a35b1f86407fc4f126835c15fedb96047dd0248d4ee13faa60adcf197ae2fda0777b6520c1d6a87bd4efd8f90a7e9b9f3238ee102b42701186dea7e63ab62ef8dcc6779639f356b4ceacae3cc659d27b94b0970;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf3aa951ffb93e6f3994a534a80166547e3709e98629b8e3062c55ee1f0d688e4ac1131a7446e9ba5cb3f172a08233d51c6f71e5b77a4edb830dfbde40605bdbc17e47d9f176840711e4514b2b8add4bf97603bed7fb77bb5af8969a0825b3db91daa5b0780d683fbd2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf37ca19f0619ae06a3e446294ac77b84739eb75fde966e30d7f5ae257bf18c56aa5572b6e9285d8ccbaff56a845fbf0b87e51635e014f73d684bd6420149a25a160e8891f3624e3f1cb02c74e44cf504b88f0ff95eb217eb29c0b548f470c18d1a8fad9bf04292df96;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h149fd6016fa17ffbced9db40d98f7d34742e8f218d1e52a684da76fe5d2188edef39717c16673792cbc4a6ed93624c93f30a76b284288b1cdca51ace90b1d7e1b96166e3a1e61212d6169564eacde64da1c6fff53c8811faf7dbe47625d4b5e1de99aebe0878448acf0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e823be325510cff6c43673d528a6c8502124cb63e389e7e6876540e25dcfcd1ee9963c45ae31991d3eddefb0e409ee1b28c31b61777d31908d7d70bf33cdbb45751aab87432276ba69c77581af88a9545a363126b0d8b6ebc3935a615053d4bdca178a0b20956940;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7613637e9ecbf49a123edaf84d096f3c01ea255dba2e0ebe9113489f9bfadabc19c0167569ca8c932b83cda60c6350ee3de0b4ed7956017d07575b4cd25733492f8243b673b621f3d3011c8c1ef4319b3436c5ce0997773ff94690b00103d456316a5d8f5927db2d6d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e8030ab4526ee95cdb1a8006a0152cc6c79751b198f6f0ec90b4c58270f9fa805189363a97ce6a5184774acb085591c118f643d2ceca1647ca82896ed7897b148fd92b6b5c854aa78262a0f243cbe4ffa68d76ba21854f0448ec0da2d62a4beb13270ae8af43a3f90;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1de01dbca6096e7448de10fc1b39a9fb306d90e788a2b2f3acbd4271824c12fb04ffff85d459a5f650083dbe6380de2bbd4a3a69e7d85b4d16f3f91d9b847d4bff5f479da600399c940e3479a3c97409275920ae9a12bd88e559aad959f2cc70a4e0fccb9f78fb99350;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f80daefd5a42ee62b640e9dc4a8124f6a860f5e586084729ba2ae6e2eba6f202a299b200f328be3ed705fb92ff7faffe623e022b87a31e996c5ec82de54594435cb9db2964e7bbdc4405a5046ca765f3b455d170c34f571212be635b16828fd701e5c0ac73cf38c51c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e2c4bc1b704585675fd4bfc74d3f4c2b009d7acfdaefdfd6fe33246f6e6274ec5435d3f92989cd293567ffe7805dcc86258d57d2110320eca1bd192c1e5238d9c8089a79a0d7ea52033c5d23182574084690684343138cf79965ec9725d52291c13e97160241d678d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf30ecb505a46bb940b6ac1a49a6093a34ef3ccb10b6d4dbe1b2b60c9b003525fc122592e69d5ece8aa0a660731624c74501ece443b5e7b6e3e04d0a736b654002999d7c1a4a604e2503ef9e1434813112b229396781c34a8b4d21b98a7fb32e2c4390dd85b9d1ea3c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h345d78f0a47bbf29305c7124fef31d0df7f463ff6385a081a531246db3678f77bbd7579dac1ca1c31a105c13a498ccf7cbf568bcf6ab3b885b723e0629cf5041a11387008f6061c85eb72ddabe1c52b8ef250db82b6561647472148feab54f78e6482d8f0294984010;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11193a53e0c67308210146435993a446f1ce0d705f358f597ae0fb1a936931c74a3c7917b5696129eebfbb212104acee12d38316be546952c55b16a40b064b8f251f604b159ec9ecdeb9a8a43ce9a1f81bd2fe44fd31f3157e9bc0ddd10b808db3b96ea71f5acf4eeda;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2dac1b89d6d00aaee3eddc379ceb4f01e952e6f2aa2181c6e1743116b9f99342ffd4bca67da9cf528bc993a3fec37bbadf9af722c478820acc9e79b0bcaec7cf38a10684026fa9d33ecf8cf9de5154ccf790489f9d79ceb9cd9a90ab3212e9d3e43e7ba1120be14edd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5282fae577273f22b31312db4f98b78b2f7dbd8609c7eaff2cc3bc6aba4f0f1b482731c945c20f629b56807008b01d28633afc6303646298f58f97a127a0d3db0e5633336dde3f33406e99ba7587d0201694d238dcb61763e55fc6a75d6a54c0acf1017ca86c067f60;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e27633f09907cbc681b2ae0ec7ff1fab8ec9969d51d2e4c0badcca2ea7ab162bdea7ac4aec3fcffde67bd6b9829667cad54f01530fcebc4250a77fe4c8dd8b0ac72331bbdaf97fa431144e867ee586dd942837fa909edad7a2e3c003552d72aa19bbbaa0bc24e31bc6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h198d17e145d60a4766be383583091da3a86507ecd3c7ffb57cd9dac0b995f16a87ac621d57226d0975aedc466b09734666083f75360cc0f9f1a7bba25cef500d8a92d7f0f0b98360443c39f5b72ac2712aaf632610159dbaab8f1616b45cec07f6f0699dbc43d471d26;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118ef0e6f0823d1a033310124d03884e5ac46cc74f92d30245714e04613f18262de2757ef7d227e697bfa6501449f8e7d158c2eabf499d1e2bb44d8dd913e38493719dbd113f5d2d7a13f08e87463f1e3c41ce6a3ead4a6d82ab4621990009cf94d6f4d1810e224a7c5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf17224d21a9377c9d8b0c40e4f147aaf93ca6e4ec5b12d7abc05e1db7b97adc2e6d602e2e2125ec4ca6660324be2e4ee17c7ed258808b487dab62e844abdfabe9611e6bb8d2f14d984192e50cb8e665070abf1d46be607dd9ea950b27fdb7c7e44c19836ab23a5dcb2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13b201c8c9bc43bde22f9c85df2d7802f22215304b87505faa2c028dc1168dc8aa699f4f578202fb5fc44c6f4524664d9b4aca90f3dcac125588bd83de1f9b8dd4cde05653873e2de7fd724e130828ba26a5e0a4e49f7d7f4f9eea6fd48afd7acc13c3d7fdf3ba2be1b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90bc3a40e6c04a7c5bb42368088421275d2df3304761869359d3f3a33dc07a54706062e163caf0b925b2beffeaa15495155c34d42867fd4db22610e25e8e783a7c128735a6d35d935a3d76550b760eb79cbf1e16439b6983dddc6413752571a506143f7a51871d9354;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10ae96ae9cc4c6a5f2b1e1b02853749aa1b81154477be1602bc2563ec098af427f9b109d3a4e7e2044972b1a996a379867fb7243acb475db96b977fcd04d924149b37534084c83f3b08401e88d2617b58fa6575706e6f28a1b922ac89473895b2131740abc0f3f8af09;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b5b4b21cd23b8cf7de3153d39d0f4de718f19ca3dcc53338db0583139a78bab4102e964e584ed17ce3d829794bae2f8e7e8fca708ed60dfff0a0b8a9a8df445a568b700d6ad60c0c1277350ccdf289bdc8a577c1ed02c5792e40c9a3bd45d27343c5d8343b8934180;
        #1
        $finish();
    end
endmodule
