// probclass: mul
// size:      13
// stage:     8
// cost:      21
// elapsed:   351.28018522262573
module compressor (
      input wire [0:0] src0,
      input wire [1:0] src1,
      input wire [2:0] src2,
      input wire [3:0] src3,
      input wire [4:0] src4,
      input wire [5:0] src5,
      input wire [6:0] src6,
      input wire [7:0] src7,
      input wire [8:0] src8,
      input wire [9:0] src9,
      input wire [10:0] src10,
      input wire [11:0] src11,
      input wire [12:0] src12,
      input wire [11:0] src13,
      input wire [10:0] src14,
      input wire [9:0] src15,
      input wire [8:0] src16,
      input wire [7:0] src17,
      input wire [6:0] src18,
      input wire [5:0] src19,
      input wire [4:0] src20,
      input wire [3:0] src21,
      input wire [2:0] src22,
      input wire [1:0] src23,
      input wire [0:0] src24,
      output wire [0:0] dst0,
      output wire [0:0] dst1,
      output wire [0:0] dst2,
      output wire [0:0] dst3,
      output wire [0:0] dst4,
      output wire [0:0] dst5,
      output wire [0:0] dst6,
      output wire [0:0] dst7,
      output wire [0:0] dst8,
      output wire [0:0] dst9,
      output wire [0:0] dst10,
      output wire [0:0] dst11,
      output wire [0:0] dst12,
      output wire [0:0] dst13,
      output wire [0:0] dst14,
      output wire [0:0] dst15,
      output wire [0:0] dst16,
      output wire [0:0] dst17,
      output wire [0:0] dst18,
      output wire [0:0] dst19,
      output wire [0:0] dst20,
      output wire [0:0] dst21,
      output wire [0:0] dst22,
      output wire [0:0] dst23,
      output wire [0:0] dst24,
      output wire [0:0] dst25);

   wire [0:0] stage0_0;
   wire [1:0] stage0_1;
   wire [2:0] stage0_2;
   wire [3:0] stage0_3;
   wire [4:0] stage0_4;
   wire [5:0] stage0_5;
   wire [6:0] stage0_6;
   wire [7:0] stage0_7;
   wire [8:0] stage0_8;
   wire [9:0] stage0_9;
   wire [10:0] stage0_10;
   wire [11:0] stage0_11;
   wire [12:0] stage0_12;
   wire [11:0] stage0_13;
   wire [10:0] stage0_14;
   wire [9:0] stage0_15;
   wire [8:0] stage0_16;
   wire [7:0] stage0_17;
   wire [6:0] stage0_18;
   wire [5:0] stage0_19;
   wire [4:0] stage0_20;
   wire [3:0] stage0_21;
   wire [2:0] stage0_22;
   wire [1:0] stage0_23;
   wire [0:0] stage0_24;
   wire [0:0] stage1_0;
   wire [0:0] stage1_1;
   wire [0:0] stage1_2;
   wire [0:0] stage1_3;
   wire [5:0] stage1_4;
   wire [6:0] stage1_5;
   wire [0:0] stage1_6;
   wire [2:0] stage1_7;
   wire [4:0] stage1_8;
   wire [5:0] stage1_9;
   wire [6:0] stage1_10;
   wire [3:0] stage1_11;
   wire [8:0] stage1_12;
   wire [2:0] stage1_13;
   wire [7:0] stage1_14;
   wire [6:0] stage1_15;
   wire [4:0] stage1_16;
   wire [5:0] stage1_17;
   wire [7:0] stage1_18;
   wire [6:0] stage1_19;
   wire [4:0] stage1_20;
   wire [3:0] stage1_21;
   wire [2:0] stage1_22;
   wire [1:0] stage1_23;
   wire [0:0] stage1_24;
   wire [0:0] stage2_0;
   wire [0:0] stage2_1;
   wire [0:0] stage2_2;
   wire [0:0] stage2_3;
   wire [0:0] stage2_4;
   wire [5:0] stage2_5;
   wire [0:0] stage2_6;
   wire [1:0] stage2_7;
   wire [0:0] stage2_8;
   wire [4:0] stage2_9;
   wire [6:0] stage2_10;
   wire [1:0] stage2_11;
   wire [5:0] stage2_12;
   wire [1:0] stage2_13;
   wire [7:0] stage2_14;
   wire [7:0] stage2_15;
   wire [4:0] stage2_16;
   wire [5:0] stage2_17;
   wire [7:0] stage2_18;
   wire [6:0] stage2_19;
   wire [4:0] stage2_20;
   wire [3:0] stage2_21;
   wire [2:0] stage2_22;
   wire [1:0] stage2_23;
   wire [0:0] stage2_24;
   wire [0:0] stage3_0;
   wire [0:0] stage3_1;
   wire [0:0] stage3_2;
   wire [0:0] stage3_3;
   wire [0:0] stage3_4;
   wire [0:0] stage3_5;
   wire [0:0] stage3_6;
   wire [0:0] stage3_7;
   wire [0:0] stage3_8;
   wire [5:0] stage3_9;
   wire [0:0] stage3_10;
   wire [2:0] stage3_11;
   wire [0:0] stage3_12;
   wire [2:0] stage3_13;
   wire [8:0] stage3_14;
   wire [1:0] stage3_15;
   wire [5:0] stage3_16;
   wire [0:0] stage3_17;
   wire [8:0] stage3_18;
   wire [1:0] stage3_19;
   wire [5:0] stage3_20;
   wire [0:0] stage3_21;
   wire [2:0] stage3_22;
   wire [2:0] stage3_23;
   wire [0:0] stage3_24;
   wire [0:0] stage4_0;
   wire [0:0] stage4_1;
   wire [0:0] stage4_2;
   wire [0:0] stage4_3;
   wire [0:0] stage4_4;
   wire [0:0] stage4_5;
   wire [0:0] stage4_6;
   wire [0:0] stage4_7;
   wire [0:0] stage4_8;
   wire [0:0] stage4_9;
   wire [0:0] stage4_10;
   wire [0:0] stage4_11;
   wire [0:0] stage4_12;
   wire [3:0] stage4_13;
   wire [2:0] stage4_14;
   wire [2:0] stage4_15;
   wire [0:0] stage4_16;
   wire [1:0] stage4_17;
   wire [3:0] stage4_18;
   wire [2:0] stage4_19;
   wire [0:0] stage4_20;
   wire [1:0] stage4_21;
   wire [3:0] stage4_22;
   wire [2:0] stage4_23;
   wire [0:0] stage4_24;
   wire [0:0] stage5_0;
   wire [0:0] stage5_1;
   wire [0:0] stage5_2;
   wire [0:0] stage5_3;
   wire [0:0] stage5_4;
   wire [0:0] stage5_5;
   wire [0:0] stage5_6;
   wire [0:0] stage5_7;
   wire [0:0] stage5_8;
   wire [0:0] stage5_9;
   wire [0:0] stage5_10;
   wire [0:0] stage5_11;
   wire [0:0] stage5_12;
   wire [0:0] stage5_13;
   wire [0:0] stage5_14;
   wire [0:0] stage5_15;
   wire [0:0] stage5_16;
   wire [2:0] stage5_17;
   wire [3:0] stage5_18;
   wire [2:0] stage5_19;
   wire [0:0] stage5_20;
   wire [1:0] stage5_21;
   wire [3:0] stage5_22;
   wire [2:0] stage5_23;
   wire [0:0] stage5_24;
   wire [0:0] stage6_0;
   wire [0:0] stage6_1;
   wire [0:0] stage6_2;
   wire [0:0] stage6_3;
   wire [0:0] stage6_4;
   wire [0:0] stage6_5;
   wire [0:0] stage6_6;
   wire [0:0] stage6_7;
   wire [0:0] stage6_8;
   wire [0:0] stage6_9;
   wire [0:0] stage6_10;
   wire [0:0] stage6_11;
   wire [0:0] stage6_12;
   wire [0:0] stage6_13;
   wire [0:0] stage6_14;
   wire [0:0] stage6_15;
   wire [0:0] stage6_16;
   wire [0:0] stage6_17;
   wire [0:0] stage6_18;
   wire [0:0] stage6_19;
   wire [0:0] stage6_20;
   wire [2:0] stage6_21;
   wire [3:0] stage6_22;
   wire [2:0] stage6_23;
   wire [0:0] stage6_24;
   wire [0:0] stage7_0;
   wire [0:0] stage7_1;
   wire [0:0] stage7_2;
   wire [0:0] stage7_3;
   wire [0:0] stage7_4;
   wire [0:0] stage7_5;
   wire [0:0] stage7_6;
   wire [0:0] stage7_7;
   wire [0:0] stage7_8;
   wire [0:0] stage7_9;
   wire [0:0] stage7_10;
   wire [0:0] stage7_11;
   wire [0:0] stage7_12;
   wire [0:0] stage7_13;
   wire [0:0] stage7_14;
   wire [0:0] stage7_15;
   wire [0:0] stage7_16;
   wire [0:0] stage7_17;
   wire [0:0] stage7_18;
   wire [0:0] stage7_19;
   wire [0:0] stage7_20;
   wire [0:0] stage7_21;
   wire [0:0] stage7_22;
   wire [0:0] stage7_23;
   wire [0:0] stage7_24;
   wire [0:0] stage7_25;
   wire [0:0] stage8_0;
   wire [0:0] stage8_1;
   wire [0:0] stage8_2;
   wire [0:0] stage8_3;
   wire [0:0] stage8_4;
   wire [0:0] stage8_5;
   wire [0:0] stage8_6;
   wire [0:0] stage8_7;
   wire [0:0] stage8_8;
   wire [0:0] stage8_9;
   wire [0:0] stage8_10;
   wire [0:0] stage8_11;
   wire [0:0] stage8_12;
   wire [0:0] stage8_13;
   wire [0:0] stage8_14;
   wire [0:0] stage8_15;
   wire [0:0] stage8_16;
   wire [0:0] stage8_17;
   wire [0:0] stage8_18;
   wire [0:0] stage8_19;
   wire [0:0] stage8_20;
   wire [0:0] stage8_21;
   wire [0:0] stage8_22;
   wire [0:0] stage8_23;
   wire [0:0] stage8_24;
   wire [0:0] stage8_25;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;
   assign dst25 = stage8_25;

   gpc433_5 gpc0 (
      {stage0_1[0], stage0_1[1], 1'b0},
      {stage0_2[0], stage0_2[1], stage0_2[2]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3]},
      {stage1_5[0],stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0]}
   );
   gpc607_5 gpc1 (
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[0],stage1_8[0],stage1_7[0],stage1_6[0]}
   );
   gpc607_5 gpc2 (
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[1],stage1_9[1],stage1_8[1],stage1_7[1]}
   );
   gpc607_5 gpc3 (
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[0],stage1_12[0],stage1_11[1],stage1_10[2]}
   );
   gpc607_5 gpc4 (
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[1],stage1_13[1],stage1_12[1],stage1_11[2]}
   );
   gpc615_5 gpc5 (
      {stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage0_12[6]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[2],stage1_13[2],stage1_12[2],stage1_11[3]}
   );
   gpc607_5 gpc6 (
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5], stage0_14[6]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[0],stage1_16[0],stage1_15[2],stage1_14[3]}
   );
   gpc1407_5 gpc7 (
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5], stage0_15[6]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3]},
      {stage0_18[0]},
      {stage1_19[0],stage1_18[1],stage1_17[1],stage1_16[1],stage1_15[3]}
   );
   gpc1_1 gpc8 (
      {stage0_0[0]},
      {stage1_0[0]}
   );
   gpc1_1 gpc9 (
      {stage0_4[0]},
      {stage1_4[1]}
   );
   gpc1_1 gpc10 (
      {stage0_4[1]},
      {stage1_4[2]}
   );
   gpc1_1 gpc11 (
      {stage0_4[2]},
      {stage1_4[3]}
   );
   gpc1_1 gpc12 (
      {stage0_4[3]},
      {stage1_4[4]}
   );
   gpc1_1 gpc13 (
      {stage0_4[4]},
      {stage1_4[5]}
   );
   gpc1_1 gpc14 (
      {stage0_5[0]},
      {stage1_5[1]}
   );
   gpc1_1 gpc15 (
      {stage0_5[1]},
      {stage1_5[2]}
   );
   gpc1_1 gpc16 (
      {stage0_5[2]},
      {stage1_5[3]}
   );
   gpc1_1 gpc17 (
      {stage0_5[3]},
      {stage1_5[4]}
   );
   gpc1_1 gpc18 (
      {stage0_5[4]},
      {stage1_5[5]}
   );
   gpc1_1 gpc19 (
      {stage0_5[5]},
      {stage1_5[6]}
   );
   gpc1_1 gpc20 (
      {stage0_7[7]},
      {stage1_7[2]}
   );
   gpc1_1 gpc21 (
      {stage0_8[6]},
      {stage1_8[2]}
   );
   gpc1_1 gpc22 (
      {stage0_8[7]},
      {stage1_8[3]}
   );
   gpc1_1 gpc23 (
      {stage0_8[8]},
      {stage1_8[4]}
   );
   gpc1_1 gpc24 (
      {stage0_9[6]},
      {stage1_9[2]}
   );
   gpc1_1 gpc25 (
      {stage0_9[7]},
      {stage1_9[3]}
   );
   gpc1_1 gpc26 (
      {stage0_9[8]},
      {stage1_9[4]}
   );
   gpc1_1 gpc27 (
      {stage0_9[9]},
      {stage1_9[5]}
   );
   gpc1_1 gpc28 (
      {stage0_10[7]},
      {stage1_10[3]}
   );
   gpc1_1 gpc29 (
      {stage0_10[8]},
      {stage1_10[4]}
   );
   gpc1_1 gpc30 (
      {stage0_10[9]},
      {stage1_10[5]}
   );
   gpc1_1 gpc31 (
      {stage0_10[10]},
      {stage1_10[6]}
   );
   gpc1_1 gpc32 (
      {stage0_12[7]},
      {stage1_12[3]}
   );
   gpc1_1 gpc33 (
      {stage0_12[8]},
      {stage1_12[4]}
   );
   gpc1_1 gpc34 (
      {stage0_12[9]},
      {stage1_12[5]}
   );
   gpc1_1 gpc35 (
      {stage0_12[10]},
      {stage1_12[6]}
   );
   gpc1_1 gpc36 (
      {stage0_12[11]},
      {stage1_12[7]}
   );
   gpc1_1 gpc37 (
      {stage0_12[12]},
      {stage1_12[8]}
   );
   gpc1_1 gpc38 (
      {stage0_14[7]},
      {stage1_14[4]}
   );
   gpc1_1 gpc39 (
      {stage0_14[8]},
      {stage1_14[5]}
   );
   gpc1_1 gpc40 (
      {stage0_14[9]},
      {stage1_14[6]}
   );
   gpc1_1 gpc41 (
      {stage0_14[10]},
      {stage1_14[7]}
   );
   gpc1_1 gpc42 (
      {stage0_15[7]},
      {stage1_15[4]}
   );
   gpc1_1 gpc43 (
      {stage0_15[8]},
      {stage1_15[5]}
   );
   gpc1_1 gpc44 (
      {stage0_15[9]},
      {stage1_15[6]}
   );
   gpc1_1 gpc45 (
      {stage0_16[6]},
      {stage1_16[2]}
   );
   gpc1_1 gpc46 (
      {stage0_16[7]},
      {stage1_16[3]}
   );
   gpc1_1 gpc47 (
      {stage0_16[8]},
      {stage1_16[4]}
   );
   gpc1_1 gpc48 (
      {stage0_17[4]},
      {stage1_17[2]}
   );
   gpc1_1 gpc49 (
      {stage0_17[5]},
      {stage1_17[3]}
   );
   gpc1_1 gpc50 (
      {stage0_17[6]},
      {stage1_17[4]}
   );
   gpc1_1 gpc51 (
      {stage0_17[7]},
      {stage1_17[5]}
   );
   gpc1_1 gpc52 (
      {stage0_18[1]},
      {stage1_18[2]}
   );
   gpc1_1 gpc53 (
      {stage0_18[2]},
      {stage1_18[3]}
   );
   gpc1_1 gpc54 (
      {stage0_18[3]},
      {stage1_18[4]}
   );
   gpc1_1 gpc55 (
      {stage0_18[4]},
      {stage1_18[5]}
   );
   gpc1_1 gpc56 (
      {stage0_18[5]},
      {stage1_18[6]}
   );
   gpc1_1 gpc57 (
      {stage0_18[6]},
      {stage1_18[7]}
   );
   gpc1_1 gpc58 (
      {stage0_19[0]},
      {stage1_19[1]}
   );
   gpc1_1 gpc59 (
      {stage0_19[1]},
      {stage1_19[2]}
   );
   gpc1_1 gpc60 (
      {stage0_19[2]},
      {stage1_19[3]}
   );
   gpc1_1 gpc61 (
      {stage0_19[3]},
      {stage1_19[4]}
   );
   gpc1_1 gpc62 (
      {stage0_19[4]},
      {stage1_19[5]}
   );
   gpc1_1 gpc63 (
      {stage0_19[5]},
      {stage1_19[6]}
   );
   gpc1_1 gpc64 (
      {stage0_20[0]},
      {stage1_20[0]}
   );
   gpc1_1 gpc65 (
      {stage0_20[1]},
      {stage1_20[1]}
   );
   gpc1_1 gpc66 (
      {stage0_20[2]},
      {stage1_20[2]}
   );
   gpc1_1 gpc67 (
      {stage0_20[3]},
      {stage1_20[3]}
   );
   gpc1_1 gpc68 (
      {stage0_20[4]},
      {stage1_20[4]}
   );
   gpc1_1 gpc69 (
      {stage0_21[0]},
      {stage1_21[0]}
   );
   gpc1_1 gpc70 (
      {stage0_21[1]},
      {stage1_21[1]}
   );
   gpc1_1 gpc71 (
      {stage0_21[2]},
      {stage1_21[2]}
   );
   gpc1_1 gpc72 (
      {stage0_21[3]},
      {stage1_21[3]}
   );
   gpc1_1 gpc73 (
      {stage0_22[0]},
      {stage1_22[0]}
   );
   gpc1_1 gpc74 (
      {stage0_22[1]},
      {stage1_22[1]}
   );
   gpc1_1 gpc75 (
      {stage0_22[2]},
      {stage1_22[2]}
   );
   gpc1_1 gpc76 (
      {stage0_23[0]},
      {stage1_23[0]}
   );
   gpc1_1 gpc77 (
      {stage0_23[1]},
      {stage1_23[1]}
   );
   gpc1_1 gpc78 (
      {stage0_24[0]},
      {stage1_24[0]}
   );
   gpc126_4 gpc79 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_5[0], stage1_5[1]},
      {stage1_6[0]},
      {stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[0]}
   );
   gpc1253_5 gpc80 (
      {stage1_7[0], stage1_7[1], stage1_7[2]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4]},
      {stage1_9[0], stage1_9[1]},
      {stage1_10[0]},
      {stage2_11[0],stage2_10[0],stage2_9[0],stage2_8[0],stage2_7[1]}
   );
   gpc1244_5 gpc81 (
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3]},
      {stage1_13[0], stage1_13[1]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[0],stage2_13[0],stage2_12[0],stage2_11[1]}
   );
   gpc1_1 gpc82 (
      {stage1_0[0]},
      {stage2_0[0]}
   );
   gpc1_1 gpc83 (
      {stage1_1[0]},
      {stage2_1[0]}
   );
   gpc1_1 gpc84 (
      {stage1_2[0]},
      {stage2_2[0]}
   );
   gpc1_1 gpc85 (
      {stage1_3[0]},
      {stage2_3[0]}
   );
   gpc1_1 gpc86 (
      {stage1_5[2]},
      {stage2_5[1]}
   );
   gpc1_1 gpc87 (
      {stage1_5[3]},
      {stage2_5[2]}
   );
   gpc1_1 gpc88 (
      {stage1_5[4]},
      {stage2_5[3]}
   );
   gpc1_1 gpc89 (
      {stage1_5[5]},
      {stage2_5[4]}
   );
   gpc1_1 gpc90 (
      {stage1_5[6]},
      {stage2_5[5]}
   );
   gpc1_1 gpc91 (
      {stage1_9[2]},
      {stage2_9[1]}
   );
   gpc1_1 gpc92 (
      {stage1_9[3]},
      {stage2_9[2]}
   );
   gpc1_1 gpc93 (
      {stage1_9[4]},
      {stage2_9[3]}
   );
   gpc1_1 gpc94 (
      {stage1_9[5]},
      {stage2_9[4]}
   );
   gpc1_1 gpc95 (
      {stage1_10[1]},
      {stage2_10[1]}
   );
   gpc1_1 gpc96 (
      {stage1_10[2]},
      {stage2_10[2]}
   );
   gpc1_1 gpc97 (
      {stage1_10[3]},
      {stage2_10[3]}
   );
   gpc1_1 gpc98 (
      {stage1_10[4]},
      {stage2_10[4]}
   );
   gpc1_1 gpc99 (
      {stage1_10[5]},
      {stage2_10[5]}
   );
   gpc1_1 gpc100 (
      {stage1_10[6]},
      {stage2_10[6]}
   );
   gpc1_1 gpc101 (
      {stage1_12[4]},
      {stage2_12[1]}
   );
   gpc1_1 gpc102 (
      {stage1_12[5]},
      {stage2_12[2]}
   );
   gpc1_1 gpc103 (
      {stage1_12[6]},
      {stage2_12[3]}
   );
   gpc1_1 gpc104 (
      {stage1_12[7]},
      {stage2_12[4]}
   );
   gpc1_1 gpc105 (
      {stage1_12[8]},
      {stage2_12[5]}
   );
   gpc1_1 gpc106 (
      {stage1_13[2]},
      {stage2_13[1]}
   );
   gpc1_1 gpc107 (
      {stage1_14[1]},
      {stage2_14[1]}
   );
   gpc1_1 gpc108 (
      {stage1_14[2]},
      {stage2_14[2]}
   );
   gpc1_1 gpc109 (
      {stage1_14[3]},
      {stage2_14[3]}
   );
   gpc1_1 gpc110 (
      {stage1_14[4]},
      {stage2_14[4]}
   );
   gpc1_1 gpc111 (
      {stage1_14[5]},
      {stage2_14[5]}
   );
   gpc1_1 gpc112 (
      {stage1_14[6]},
      {stage2_14[6]}
   );
   gpc1_1 gpc113 (
      {stage1_14[7]},
      {stage2_14[7]}
   );
   gpc1_1 gpc114 (
      {stage1_15[0]},
      {stage2_15[1]}
   );
   gpc1_1 gpc115 (
      {stage1_15[1]},
      {stage2_15[2]}
   );
   gpc1_1 gpc116 (
      {stage1_15[2]},
      {stage2_15[3]}
   );
   gpc1_1 gpc117 (
      {stage1_15[3]},
      {stage2_15[4]}
   );
   gpc1_1 gpc118 (
      {stage1_15[4]},
      {stage2_15[5]}
   );
   gpc1_1 gpc119 (
      {stage1_15[5]},
      {stage2_15[6]}
   );
   gpc1_1 gpc120 (
      {stage1_15[6]},
      {stage2_15[7]}
   );
   gpc1_1 gpc121 (
      {stage1_16[0]},
      {stage2_16[0]}
   );
   gpc1_1 gpc122 (
      {stage1_16[1]},
      {stage2_16[1]}
   );
   gpc1_1 gpc123 (
      {stage1_16[2]},
      {stage2_16[2]}
   );
   gpc1_1 gpc124 (
      {stage1_16[3]},
      {stage2_16[3]}
   );
   gpc1_1 gpc125 (
      {stage1_16[4]},
      {stage2_16[4]}
   );
   gpc1_1 gpc126 (
      {stage1_17[0]},
      {stage2_17[0]}
   );
   gpc1_1 gpc127 (
      {stage1_17[1]},
      {stage2_17[1]}
   );
   gpc1_1 gpc128 (
      {stage1_17[2]},
      {stage2_17[2]}
   );
   gpc1_1 gpc129 (
      {stage1_17[3]},
      {stage2_17[3]}
   );
   gpc1_1 gpc130 (
      {stage1_17[4]},
      {stage2_17[4]}
   );
   gpc1_1 gpc131 (
      {stage1_17[5]},
      {stage2_17[5]}
   );
   gpc1_1 gpc132 (
      {stage1_18[0]},
      {stage2_18[0]}
   );
   gpc1_1 gpc133 (
      {stage1_18[1]},
      {stage2_18[1]}
   );
   gpc1_1 gpc134 (
      {stage1_18[2]},
      {stage2_18[2]}
   );
   gpc1_1 gpc135 (
      {stage1_18[3]},
      {stage2_18[3]}
   );
   gpc1_1 gpc136 (
      {stage1_18[4]},
      {stage2_18[4]}
   );
   gpc1_1 gpc137 (
      {stage1_18[5]},
      {stage2_18[5]}
   );
   gpc1_1 gpc138 (
      {stage1_18[6]},
      {stage2_18[6]}
   );
   gpc1_1 gpc139 (
      {stage1_18[7]},
      {stage2_18[7]}
   );
   gpc1_1 gpc140 (
      {stage1_19[0]},
      {stage2_19[0]}
   );
   gpc1_1 gpc141 (
      {stage1_19[1]},
      {stage2_19[1]}
   );
   gpc1_1 gpc142 (
      {stage1_19[2]},
      {stage2_19[2]}
   );
   gpc1_1 gpc143 (
      {stage1_19[3]},
      {stage2_19[3]}
   );
   gpc1_1 gpc144 (
      {stage1_19[4]},
      {stage2_19[4]}
   );
   gpc1_1 gpc145 (
      {stage1_19[5]},
      {stage2_19[5]}
   );
   gpc1_1 gpc146 (
      {stage1_19[6]},
      {stage2_19[6]}
   );
   gpc1_1 gpc147 (
      {stage1_20[0]},
      {stage2_20[0]}
   );
   gpc1_1 gpc148 (
      {stage1_20[1]},
      {stage2_20[1]}
   );
   gpc1_1 gpc149 (
      {stage1_20[2]},
      {stage2_20[2]}
   );
   gpc1_1 gpc150 (
      {stage1_20[3]},
      {stage2_20[3]}
   );
   gpc1_1 gpc151 (
      {stage1_20[4]},
      {stage2_20[4]}
   );
   gpc1_1 gpc152 (
      {stage1_21[0]},
      {stage2_21[0]}
   );
   gpc1_1 gpc153 (
      {stage1_21[1]},
      {stage2_21[1]}
   );
   gpc1_1 gpc154 (
      {stage1_21[2]},
      {stage2_21[2]}
   );
   gpc1_1 gpc155 (
      {stage1_21[3]},
      {stage2_21[3]}
   );
   gpc1_1 gpc156 (
      {stage1_22[0]},
      {stage2_22[0]}
   );
   gpc1_1 gpc157 (
      {stage1_22[1]},
      {stage2_22[1]}
   );
   gpc1_1 gpc158 (
      {stage1_22[2]},
      {stage2_22[2]}
   );
   gpc1_1 gpc159 (
      {stage1_23[0]},
      {stage2_23[0]}
   );
   gpc1_1 gpc160 (
      {stage1_23[1]},
      {stage2_23[1]}
   );
   gpc1_1 gpc161 (
      {stage1_24[0]},
      {stage2_24[0]}
   );
   gpc1316_5 gpc162 (
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage2_6[0]},
      {stage2_7[0], stage2_7[1], 1'b0},
      {stage2_8[0]},
      {stage3_9[0],stage3_8[0],stage3_7[0],stage3_6[0],stage3_5[0]}
   );
   gpc607_5 gpc163 (
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5], stage2_10[6]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[0],stage3_11[0],stage3_10[0]}
   );
   gpc607_5 gpc164 (
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[0],stage3_17[0],stage3_16[0],stage3_15[0]}
   );
   gpc1407_5 gpc165 (
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5], stage2_19[6]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3]},
      {stage2_22[0]},
      {stage3_23[0],stage3_22[0],stage3_21[0],stage3_20[0],stage3_19[1]}
   );
   gpc1_1 gpc166 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc167 (
      {stage2_1[0]},
      {stage3_1[0]}
   );
   gpc1_1 gpc168 (
      {stage2_2[0]},
      {stage3_2[0]}
   );
   gpc1_1 gpc169 (
      {stage2_3[0]},
      {stage3_3[0]}
   );
   gpc1_1 gpc170 (
      {stage2_4[0]},
      {stage3_4[0]}
   );
   gpc1_1 gpc171 (
      {stage2_9[0]},
      {stage3_9[1]}
   );
   gpc1_1 gpc172 (
      {stage2_9[1]},
      {stage3_9[2]}
   );
   gpc1_1 gpc173 (
      {stage2_9[2]},
      {stage3_9[3]}
   );
   gpc1_1 gpc174 (
      {stage2_9[3]},
      {stage3_9[4]}
   );
   gpc1_1 gpc175 (
      {stage2_9[4]},
      {stage3_9[5]}
   );
   gpc1_1 gpc176 (
      {stage2_11[0]},
      {stage3_11[1]}
   );
   gpc1_1 gpc177 (
      {stage2_11[1]},
      {stage3_11[2]}
   );
   gpc1_1 gpc178 (
      {stage2_13[0]},
      {stage3_13[1]}
   );
   gpc1_1 gpc179 (
      {stage2_13[1]},
      {stage3_13[2]}
   );
   gpc1_1 gpc180 (
      {stage2_14[0]},
      {stage3_14[1]}
   );
   gpc1_1 gpc181 (
      {stage2_14[1]},
      {stage3_14[2]}
   );
   gpc1_1 gpc182 (
      {stage2_14[2]},
      {stage3_14[3]}
   );
   gpc1_1 gpc183 (
      {stage2_14[3]},
      {stage3_14[4]}
   );
   gpc1_1 gpc184 (
      {stage2_14[4]},
      {stage3_14[5]}
   );
   gpc1_1 gpc185 (
      {stage2_14[5]},
      {stage3_14[6]}
   );
   gpc1_1 gpc186 (
      {stage2_14[6]},
      {stage3_14[7]}
   );
   gpc1_1 gpc187 (
      {stage2_14[7]},
      {stage3_14[8]}
   );
   gpc1_1 gpc188 (
      {stage2_15[7]},
      {stage3_15[1]}
   );
   gpc1_1 gpc189 (
      {stage2_16[0]},
      {stage3_16[1]}
   );
   gpc1_1 gpc190 (
      {stage2_16[1]},
      {stage3_16[2]}
   );
   gpc1_1 gpc191 (
      {stage2_16[2]},
      {stage3_16[3]}
   );
   gpc1_1 gpc192 (
      {stage2_16[3]},
      {stage3_16[4]}
   );
   gpc1_1 gpc193 (
      {stage2_16[4]},
      {stage3_16[5]}
   );
   gpc1_1 gpc194 (
      {stage2_18[0]},
      {stage3_18[1]}
   );
   gpc1_1 gpc195 (
      {stage2_18[1]},
      {stage3_18[2]}
   );
   gpc1_1 gpc196 (
      {stage2_18[2]},
      {stage3_18[3]}
   );
   gpc1_1 gpc197 (
      {stage2_18[3]},
      {stage3_18[4]}
   );
   gpc1_1 gpc198 (
      {stage2_18[4]},
      {stage3_18[5]}
   );
   gpc1_1 gpc199 (
      {stage2_18[5]},
      {stage3_18[6]}
   );
   gpc1_1 gpc200 (
      {stage2_18[6]},
      {stage3_18[7]}
   );
   gpc1_1 gpc201 (
      {stage2_18[7]},
      {stage3_18[8]}
   );
   gpc1_1 gpc202 (
      {stage2_20[0]},
      {stage3_20[1]}
   );
   gpc1_1 gpc203 (
      {stage2_20[1]},
      {stage3_20[2]}
   );
   gpc1_1 gpc204 (
      {stage2_20[2]},
      {stage3_20[3]}
   );
   gpc1_1 gpc205 (
      {stage2_20[3]},
      {stage3_20[4]}
   );
   gpc1_1 gpc206 (
      {stage2_20[4]},
      {stage3_20[5]}
   );
   gpc1_1 gpc207 (
      {stage2_22[1]},
      {stage3_22[1]}
   );
   gpc1_1 gpc208 (
      {stage2_22[2]},
      {stage3_22[2]}
   );
   gpc1_1 gpc209 (
      {stage2_23[0]},
      {stage3_23[1]}
   );
   gpc1_1 gpc210 (
      {stage2_23[1]},
      {stage3_23[2]}
   );
   gpc1_1 gpc211 (
      {stage2_24[0]},
      {stage3_24[0]}
   );
   gpc1316_5 gpc212 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_10[0]},
      {stage3_11[0], stage3_11[1], stage3_11[2]},
      {stage3_12[0]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[0]}
   );
   gpc607_5 gpc213 (
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[0],stage4_16[0],stage4_15[0],stage4_14[0]}
   );
   gpc607_5 gpc214 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5], stage3_18[6]},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage4_22[0],stage4_21[0],stage4_20[0],stage4_19[0],stage4_18[1]}
   );
   gpc1_1 gpc215 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc216 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc217 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc218 (
      {stage3_3[0]},
      {stage4_3[0]}
   );
   gpc1_1 gpc219 (
      {stage3_4[0]},
      {stage4_4[0]}
   );
   gpc1_1 gpc220 (
      {stage3_5[0]},
      {stage4_5[0]}
   );
   gpc1_1 gpc221 (
      {stage3_6[0]},
      {stage4_6[0]}
   );
   gpc1_1 gpc222 (
      {stage3_7[0]},
      {stage4_7[0]}
   );
   gpc1_1 gpc223 (
      {stage3_8[0]},
      {stage4_8[0]}
   );
   gpc1_1 gpc224 (
      {stage3_13[0]},
      {stage4_13[1]}
   );
   gpc1_1 gpc225 (
      {stage3_13[1]},
      {stage4_13[2]}
   );
   gpc1_1 gpc226 (
      {stage3_13[2]},
      {stage4_13[3]}
   );
   gpc1_1 gpc227 (
      {stage3_14[7]},
      {stage4_14[1]}
   );
   gpc1_1 gpc228 (
      {stage3_14[8]},
      {stage4_14[2]}
   );
   gpc1_1 gpc229 (
      {stage3_15[0]},
      {stage4_15[1]}
   );
   gpc1_1 gpc230 (
      {stage3_15[1]},
      {stage4_15[2]}
   );
   gpc1_1 gpc231 (
      {stage3_17[0]},
      {stage4_17[1]}
   );
   gpc1_1 gpc232 (
      {stage3_18[7]},
      {stage4_18[2]}
   );
   gpc1_1 gpc233 (
      {stage3_18[8]},
      {stage4_18[3]}
   );
   gpc1_1 gpc234 (
      {stage3_19[0]},
      {stage4_19[1]}
   );
   gpc1_1 gpc235 (
      {stage3_19[1]},
      {stage4_19[2]}
   );
   gpc1_1 gpc236 (
      {stage3_21[0]},
      {stage4_21[1]}
   );
   gpc1_1 gpc237 (
      {stage3_22[0]},
      {stage4_22[1]}
   );
   gpc1_1 gpc238 (
      {stage3_22[1]},
      {stage4_22[2]}
   );
   gpc1_1 gpc239 (
      {stage3_22[2]},
      {stage4_22[3]}
   );
   gpc1_1 gpc240 (
      {stage3_23[0]},
      {stage4_23[0]}
   );
   gpc1_1 gpc241 (
      {stage3_23[1]},
      {stage4_23[1]}
   );
   gpc1_1 gpc242 (
      {stage3_23[2]},
      {stage4_23[2]}
   );
   gpc1_1 gpc243 (
      {stage3_24[0]},
      {stage4_24[0]}
   );
   gpc1334_5 gpc244 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3]},
      {stage4_14[0], stage4_14[1], stage4_14[2]},
      {stage4_15[0], stage4_15[1], stage4_15[2]},
      {stage4_16[0]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[0]}
   );
   gpc1_1 gpc245 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc246 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc247 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc248 (
      {stage4_3[0]},
      {stage5_3[0]}
   );
   gpc1_1 gpc249 (
      {stage4_4[0]},
      {stage5_4[0]}
   );
   gpc1_1 gpc250 (
      {stage4_5[0]},
      {stage5_5[0]}
   );
   gpc1_1 gpc251 (
      {stage4_6[0]},
      {stage5_6[0]}
   );
   gpc1_1 gpc252 (
      {stage4_7[0]},
      {stage5_7[0]}
   );
   gpc1_1 gpc253 (
      {stage4_8[0]},
      {stage5_8[0]}
   );
   gpc1_1 gpc254 (
      {stage4_9[0]},
      {stage5_9[0]}
   );
   gpc1_1 gpc255 (
      {stage4_10[0]},
      {stage5_10[0]}
   );
   gpc1_1 gpc256 (
      {stage4_11[0]},
      {stage5_11[0]}
   );
   gpc1_1 gpc257 (
      {stage4_12[0]},
      {stage5_12[0]}
   );
   gpc1_1 gpc258 (
      {stage4_17[0]},
      {stage5_17[1]}
   );
   gpc1_1 gpc259 (
      {stage4_17[1]},
      {stage5_17[2]}
   );
   gpc1_1 gpc260 (
      {stage4_18[0]},
      {stage5_18[0]}
   );
   gpc1_1 gpc261 (
      {stage4_18[1]},
      {stage5_18[1]}
   );
   gpc1_1 gpc262 (
      {stage4_18[2]},
      {stage5_18[2]}
   );
   gpc1_1 gpc263 (
      {stage4_18[3]},
      {stage5_18[3]}
   );
   gpc1_1 gpc264 (
      {stage4_19[0]},
      {stage5_19[0]}
   );
   gpc1_1 gpc265 (
      {stage4_19[1]},
      {stage5_19[1]}
   );
   gpc1_1 gpc266 (
      {stage4_19[2]},
      {stage5_19[2]}
   );
   gpc1_1 gpc267 (
      {stage4_20[0]},
      {stage5_20[0]}
   );
   gpc1_1 gpc268 (
      {stage4_21[0]},
      {stage5_21[0]}
   );
   gpc1_1 gpc269 (
      {stage4_21[1]},
      {stage5_21[1]}
   );
   gpc1_1 gpc270 (
      {stage4_22[0]},
      {stage5_22[0]}
   );
   gpc1_1 gpc271 (
      {stage4_22[1]},
      {stage5_22[1]}
   );
   gpc1_1 gpc272 (
      {stage4_22[2]},
      {stage5_22[2]}
   );
   gpc1_1 gpc273 (
      {stage4_22[3]},
      {stage5_22[3]}
   );
   gpc1_1 gpc274 (
      {stage4_23[0]},
      {stage5_23[0]}
   );
   gpc1_1 gpc275 (
      {stage4_23[1]},
      {stage5_23[1]}
   );
   gpc1_1 gpc276 (
      {stage4_23[2]},
      {stage5_23[2]}
   );
   gpc1_1 gpc277 (
      {stage4_24[0]},
      {stage5_24[0]}
   );
   gpc1343_5 gpc278 (
      {stage5_17[0], stage5_17[1], stage5_17[2]},
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3]},
      {stage5_19[0], stage5_19[1], stage5_19[2]},
      {stage5_20[0]},
      {stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[0]}
   );
   gpc1_1 gpc279 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc280 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc281 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc282 (
      {stage5_3[0]},
      {stage6_3[0]}
   );
   gpc1_1 gpc283 (
      {stage5_4[0]},
      {stage6_4[0]}
   );
   gpc1_1 gpc284 (
      {stage5_5[0]},
      {stage6_5[0]}
   );
   gpc1_1 gpc285 (
      {stage5_6[0]},
      {stage6_6[0]}
   );
   gpc1_1 gpc286 (
      {stage5_7[0]},
      {stage6_7[0]}
   );
   gpc1_1 gpc287 (
      {stage5_8[0]},
      {stage6_8[0]}
   );
   gpc1_1 gpc288 (
      {stage5_9[0]},
      {stage6_9[0]}
   );
   gpc1_1 gpc289 (
      {stage5_10[0]},
      {stage6_10[0]}
   );
   gpc1_1 gpc290 (
      {stage5_11[0]},
      {stage6_11[0]}
   );
   gpc1_1 gpc291 (
      {stage5_12[0]},
      {stage6_12[0]}
   );
   gpc1_1 gpc292 (
      {stage5_13[0]},
      {stage6_13[0]}
   );
   gpc1_1 gpc293 (
      {stage5_14[0]},
      {stage6_14[0]}
   );
   gpc1_1 gpc294 (
      {stage5_15[0]},
      {stage6_15[0]}
   );
   gpc1_1 gpc295 (
      {stage5_16[0]},
      {stage6_16[0]}
   );
   gpc1_1 gpc296 (
      {stage5_21[0]},
      {stage6_21[1]}
   );
   gpc1_1 gpc297 (
      {stage5_21[1]},
      {stage6_21[2]}
   );
   gpc1_1 gpc298 (
      {stage5_22[0]},
      {stage6_22[0]}
   );
   gpc1_1 gpc299 (
      {stage5_22[1]},
      {stage6_22[1]}
   );
   gpc1_1 gpc300 (
      {stage5_22[2]},
      {stage6_22[2]}
   );
   gpc1_1 gpc301 (
      {stage5_22[3]},
      {stage6_22[3]}
   );
   gpc1_1 gpc302 (
      {stage5_23[0]},
      {stage6_23[0]}
   );
   gpc1_1 gpc303 (
      {stage5_23[1]},
      {stage6_23[1]}
   );
   gpc1_1 gpc304 (
      {stage5_23[2]},
      {stage6_23[2]}
   );
   gpc1_1 gpc305 (
      {stage5_24[0]},
      {stage6_24[0]}
   );
   gpc1343_5 gpc306 (
      {stage6_21[0], stage6_21[1], stage6_21[2]},
      {stage6_22[0], stage6_22[1], stage6_22[2], stage6_22[3]},
      {stage6_23[0], stage6_23[1], stage6_23[2]},
      {stage6_24[0]},
      {stage7_25[0],stage7_24[0],stage7_23[0],stage7_22[0],stage7_21[0]}
   );
   gpc1_1 gpc307 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc308 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc309 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc310 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc311 (
      {stage6_4[0]},
      {stage7_4[0]}
   );
   gpc1_1 gpc312 (
      {stage6_5[0]},
      {stage7_5[0]}
   );
   gpc1_1 gpc313 (
      {stage6_6[0]},
      {stage7_6[0]}
   );
   gpc1_1 gpc314 (
      {stage6_7[0]},
      {stage7_7[0]}
   );
   gpc1_1 gpc315 (
      {stage6_8[0]},
      {stage7_8[0]}
   );
   gpc1_1 gpc316 (
      {stage6_9[0]},
      {stage7_9[0]}
   );
   gpc1_1 gpc317 (
      {stage6_10[0]},
      {stage7_10[0]}
   );
   gpc1_1 gpc318 (
      {stage6_11[0]},
      {stage7_11[0]}
   );
   gpc1_1 gpc319 (
      {stage6_12[0]},
      {stage7_12[0]}
   );
   gpc1_1 gpc320 (
      {stage6_13[0]},
      {stage7_13[0]}
   );
   gpc1_1 gpc321 (
      {stage6_14[0]},
      {stage7_14[0]}
   );
   gpc1_1 gpc322 (
      {stage6_15[0]},
      {stage7_15[0]}
   );
   gpc1_1 gpc323 (
      {stage6_16[0]},
      {stage7_16[0]}
   );
   gpc1_1 gpc324 (
      {stage6_17[0]},
      {stage7_17[0]}
   );
   gpc1_1 gpc325 (
      {stage6_18[0]},
      {stage7_18[0]}
   );
   gpc1_1 gpc326 (
      {stage6_19[0]},
      {stage7_19[0]}
   );
   gpc1_1 gpc327 (
      {stage6_20[0]},
      {stage7_20[0]}
   );
   gpc1_1 gpc328 (
      {stage7_0[0]},
      {stage8_0[0]}
   );
   gpc1_1 gpc329 (
      {stage7_1[0]},
      {stage8_1[0]}
   );
   gpc1_1 gpc330 (
      {stage7_2[0]},
      {stage8_2[0]}
   );
   gpc1_1 gpc331 (
      {stage7_3[0]},
      {stage8_3[0]}
   );
   gpc1_1 gpc332 (
      {stage7_4[0]},
      {stage8_4[0]}
   );
   gpc1_1 gpc333 (
      {stage7_5[0]},
      {stage8_5[0]}
   );
   gpc1_1 gpc334 (
      {stage7_6[0]},
      {stage8_6[0]}
   );
   gpc1_1 gpc335 (
      {stage7_7[0]},
      {stage8_7[0]}
   );
   gpc1_1 gpc336 (
      {stage7_8[0]},
      {stage8_8[0]}
   );
   gpc1_1 gpc337 (
      {stage7_9[0]},
      {stage8_9[0]}
   );
   gpc1_1 gpc338 (
      {stage7_10[0]},
      {stage8_10[0]}
   );
   gpc1_1 gpc339 (
      {stage7_11[0]},
      {stage8_11[0]}
   );
   gpc1_1 gpc340 (
      {stage7_12[0]},
      {stage8_12[0]}
   );
   gpc1_1 gpc341 (
      {stage7_13[0]},
      {stage8_13[0]}
   );
   gpc1_1 gpc342 (
      {stage7_14[0]},
      {stage8_14[0]}
   );
   gpc1_1 gpc343 (
      {stage7_15[0]},
      {stage8_15[0]}
   );
   gpc1_1 gpc344 (
      {stage7_16[0]},
      {stage8_16[0]}
   );
   gpc1_1 gpc345 (
      {stage7_17[0]},
      {stage8_17[0]}
   );
   gpc1_1 gpc346 (
      {stage7_18[0]},
      {stage8_18[0]}
   );
   gpc1_1 gpc347 (
      {stage7_19[0]},
      {stage8_19[0]}
   );
   gpc1_1 gpc348 (
      {stage7_20[0]},
      {stage8_20[0]}
   );
   gpc1_1 gpc349 (
      {stage7_21[0]},
      {stage8_21[0]}
   );
   gpc1_1 gpc350 (
      {stage7_22[0]},
      {stage8_22[0]}
   );
   gpc1_1 gpc351 (
      {stage7_23[0]},
      {stage8_23[0]}
   );
   gpc1_1 gpc352 (
      {stage7_24[0]},
      {stage8_24[0]}
   );
   gpc1_1 gpc353 (
      {stage7_25[0]},
      {stage8_25[0]}
   );
endmodule
