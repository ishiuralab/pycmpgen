module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [16:0] src18;
    reg [15:0] src19;
    reg [14:0] src20;
    reg [13:0] src21;
    reg [12:0] src22;
    reg [11:0] src23;
    reg [10:0] src24;
    reg [9:0] src25;
    reg [8:0] src26;
    reg [7:0] src27;
    reg [6:0] src28;
    reg [5:0] src29;
    reg [4:0] src30;
    reg [3:0] src31;
    reg [2:0] src32;
    reg [1:0] src33;
    reg [0:0] src34;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [35:0] srcsum;
    wire [35:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3])<<31) + ((src32[0] + src32[1] + src32[2])<<32) + ((src33[0] + src33[1])<<33) + ((src34[0])<<34);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98a99fc87cfd2cd2524afd18fd3d9cf83127b6313deaf8695379919b1c42169daa250c0c9bbd22037;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h676ec7ef961f25fbef26d148fba41b21464546ce9651e3ffa62b9fcef5ab4d2b88affdebb35f9a714;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc439d0103dcd7ec18b4492487375f79890ccc9d7fd0252dc1778f02e9d1211fc49dd84e0b4d0e6de6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7721ceb3c61b11254d50f22fcc59d3278fe52b4c27f2b15bd44333e8dcc40b1b01f1506ac4049217a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb6b4d8860989b117e2ccae31ecf62a4fdd4f048c8ec41124d7a568df786e13c54993fd3d11e56d5b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3890a0d29d9254b88261971140ea7f4e9407c253b75b09ab6ec3d491dbbcb339d4a390f531378b1d0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf5f5b792cfc4ade72881b52a12ceae31040f69164105ae633cd6e639c55125fa1a10686d83d59704;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfeb518a597501e5648bebc5392667472ad4cd20d8735c0a182a56804ccea70d642b0d87fbeaf6efb6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd69ee2175b7d111a2512616699819f255903a1476e3dd6250df8bf1db74d0954a212e78043189d530;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1afc2c6dd6e33746c19afdca977e202f0a7f8d4ffc0216dc4d6cde1f186058ef63d04e27d8d8b8af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f1b51d513638eb3bb939a768d4b8e29451a239934f3dc7de7ab8459b7b84eae1452d540fc2b7d01b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h437278f09791c90339c1d204e7d8fb302f7645b80f6cd77bc5b442a6b33d68010719a1a38e4ff43c3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32ab2dcbf9d5a75f96f42b6b36c50d226b0cd59612940849b84d2935224741965da56f285807477ef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a779cc4c934991ece4988d54839fb5ee00c8c6b53ebcc79915c1580b56b31642c0b79b2f857d40af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd489908ded1142a9fc856d41d61126aafc0486e8ff7386c9401604606ef753426bbcb8af2514ce41;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5d728f39c06fa2cb5c4ea3d280c5ca1d4fd136b0a7cc616599450e88108bb3f508cd70b71da02aca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c18179c137af474d4da61820c705eee9985e74b8a4895868c6210f762857f188cafbefd5aa1bd8fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he874c848dee6c35a7fade365dda7c8ed2ff0907804fe1035a2e8e98f41555eb67ba5ee25c9ea2cedd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1549762880ea9dc4fbfad059da3c045e0819d5e93bf2671995dbe790c2aea1895c81fb0a2d57a4e1a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha14ec90517df083a0bc765c49a83352988dea40f7a92056e50a98b4690ab2f80c21747062e395fc68;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83e503e1b91899707c5d57f9160f42af21b35ba8d5cab6248e73b4c7a22cc36c17be963a4e90cce0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h33415791b1eb610ba7d9b8304428569a532c298d5dc0ed20ce3c47c10c6965812ba2792fa93b2e0df;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he74956b42da55d028f13ff336f738191f66d9ce49b6375219bff5de90244c354c78b47b546b693748;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35ef3b3627d9ad84245ffea557155b92b9c509e1c8fcb0bdfccb7ff157e8bd20ac80547ee1de47728;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d38f0bb6d99ca733183d6fae4002ac9cea0f15724afa1129748956499fffe90a1b1e7ab2a43da3a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba59099b7545969d3e5a5faa0138ab0666e0ed9a0dc9b3c2ba25c1936dcb2dc285514ba2f7b2ada04;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6dfd103f3b4ae3780511410bd9b2964f19b6051d7b7b5857b77a9388dc2ce84656beb43e08f89a561;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86530314c789c278fdf33a1eef4547216097fc12f819ecfb7ca0cfcc1057769c4f60c9c520fb0b802;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha433dbf021fdeca9d55920838765623bcc4225d05fc291b58d88e55d3754419d945d96378b46f4f11;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb49ef11f78852d3f682b4661593be77f37b65184a6b13f61dc9777bfe41d958b9aff9bc12e90b1069;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf5005f5730d805249414303b7c0935b7a2a0e974db25e896c622ce74a2eebe680f0b518dcff210b0d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc342c6d3479a44d661750de493c175bc56310b5b14364a3b54b48fab2211e25f3a1d5e1db57772afa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7f728bd390392a2df7084c9a91483889269e435a0c22323df6fd349e804bbb1ea2d5160a08ea442;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc60acb6777178862521f7e85a96737c336273abd2ecc9470d694f4363f4d91181bed19c1e5bbc66ff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc82bd740e1181539291f5978f4191156dd1377fe6ab9717ef7c0df566e9d1bfcd732b2fa6514e91;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9166a4385d3f76a9fa27fc0d42999889cf0c2bbfeda1816167fcf1a252b8e8f61aec8f9ba6cd9a8c0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82d31e96a55cc46379fbcb11b77340a10d3e73e143212ab03805436a4567dede19db5b2fe2e78ed59;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b23d726cb64d7c3633d9a0b097277eec59e91f4eb7389c65d41b87ec60e84da563095d67268dce9c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf1643a0671dfa6d99c91680948be4608703824246f2fc8d1c286c3eb59bb8d6babb45dfb779c662;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7cf0896e0c4048083d29dcd9a682aa0789cdc08e4036fdae26e06ef5449231c81c16f2b092d36817d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c321c4f675f98dfd63dc951644561b067bf2f4f2ba059a7ce95542b06aebd58b5d034bd14ecbe3a1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61aad466eba25f6235bd8cdee6e73078b2561e91232e3265e9802c6e32d7f53c2d5719e25c9035eff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1c2fe465618fc75863821f4afe8c854498d5bdf5dac05f8ca1bc6042ba4aaf4697c4de3e3c2053be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8fa4e1cb6d60a7d41becc9f71bfefacf5c4d78b469eb98692f779e331b82c2f099658242a29e7dc84;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0604dd9c9aa0831691987621d198f768bd258d30f255e532681d383dbfba05c88806da358ebf2d83;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3211126a8ab986648dd85fa573b7537a35172f2aa1ba57d147a15fb204104fd704a73bc95bbd6cd0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb697adcbb64202c976175a8680850f3cbad4e66827e08183e08a40ecb78c1851a7749bfcd733ddb72;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h218df1915c68fa3d8b0b7acc3084b514bf61a35d12745f26fdd37a8e11bde7655db847b210b01556;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b2b0fae5d50a7d0cc2f5506ae3b85d6c1e8a074a69195f3ebeea8865dbf7186c5e52dadb2db32e1d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1dd00728ddb2d26f2db3bfb6311c8c718cc99992d7874a84164a4285d3a16266efe053829f9e2f242;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a73d406649c4571bfcd40c9713e8f17fb7bd4a31a9825f02dfb98e9cf5dfa6ed1bdcfec9f7d8159a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c65b88f8626bd74b194da522de2d9c54f31ce360cdc5e36f62a9a7e81748d84d208b42bc81fb5c29;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4cd23dfcaa5c6cad16bf5f27c7f1554e54578845482352b2719a438bb147e16dd13dc5e60c458b003;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95692effcd905c53cdefb57e6849bd452abe7b514dd43a40d12b0a945775a8ecf01ff26054afbd9e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54a84efd966ddfb18d1449434a7374c29e07a76de111d3736279a1d36e51f0986350d6b6faeac73e2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde85d5d5432b2e9f2930a0afefc7750e207a2e47d9e48c43f4b596a6d98c3aea1e5a9bb9523dfa0c2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc914a4c30e76ee5efd8eb8a7d68a3290ce3f6881c3eee5d1cac3732b8979495ba943a22eaa19bc7f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99047feb74e4debc19fc26b1b83965be55504de7f8ffbb95a1e6d8bfbf3c3ef6ebed28292169fa42d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbda1a21e2133307e7489707204f335676a1e57e945fca7ac26c0be50c28c97d6664cceca868c51ceb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7b5629036b87fbd9b64846a9f234a7bc5ee3b148f19f5ff7b38422211fd672013d1b172e7525a147;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c8d2e396e61bd9075ee63d0572f62de775fa33b2cacf988ac39a40e0c7474da91b628dc908e0e2d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85990b2c076ab5a68c3061a7eff27bbc6ed1dd22367b55e024d0d3129f1961b9a47527bdc7529d08c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2eee7c431be7d30e790b659f010b86c407752d591270c4b14e7ba79441e08da34e9e1222c4eb997;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3105fcd43059388c582105b54e2be7507f6e2fe6feb1a1e8ed9dc3770e5b9032a9acb5a309151b1df;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha84b0417f3d079c2e1f7ccb5d15efe80f2ca6913d637a9522d76f46047cb41e7db30904feea96eea3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa12f6095b3ec3b4d6d9a035af2919e63c5be09d6c4979e99636d54a3cfa0c8e980b6d12ff67df9a4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha029a4852a3827a03e579ea2448386501137846341ff52fa04c8d6f8e874675a0f9e02d86a7850650;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ae2fa694290ac20c1ffe8ecfd25fbe26eaa9483b4f6468d6a764db2e140ceff9c9e391efca8cd199;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h106c06f1dfb4c6507e19b8f2b563b868d13ee8a6297694a4fa37f60030740aec243017d06aa393e5d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e0f5987428d0bf6202b8261e139ba9ad2d6de19cbc2a5f9cb8016ff9e604fc596d37ef8055c24aac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4d31d55366b42a102ce6d64fc48d96f2455817b5a00a84cdb46a8d24c1ee39f0bf4d51d1717951af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf328a3fc42f0ed127c332b2d53f370ad05d4c137ac330e0481768e2fbf242f26a6e2afbe781aa75;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7591afd6d3d2b785736a424ac4a2d68be56c42d1528bc7f50dca1b90b649e9d9cfea1479e112a35f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6de5eb7c533286aa96e422adada4ee6b96fafb9fd190899277fca9aaa0c52ebdc697e8477f25b2a9b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8cf9ad1e55aee7ca234b29660f58f150362eac63fd2c58e9cfea01da4d5f4550255564769221640bf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha02c90b9d49012501ceab3defe766b33ca0395a850444090d182d0e251d1cf481c6b1c8e8ed439646;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c9780c54d90837a6cb35286cb46afbe399e7f5ab122e1b1df4b5adcb8daff72564836921e92dd255;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffe28c6bbe2eaaf4f32b0f06a7552ba57822c3b1e662758125de5d405f2029959d99a670f766c4630;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3149dc749c9ae3f24df90356103c99f68f70d9fc09f12d7df7ffd889745347607f13f0aed3411f43d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd527208b89a92ecf42dc53e3055fada789a8b8311b60ee4ea79190d6d804d37f7e05336dea359a502;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ef755b356be93ec4780714684df67ae2f4f933e9b7eaff3ce714163032524c8d9d1cca7b059f6ede;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99cd20d9d0421016ec6528dcbd1dee45328907bde583fe6737b374ef456d64e394c3bfcb09e8f3522;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h284d440c15d109cc72a1e9581e8a1462db9da2d39a3ab92f43f5893b5e98f04ff231c1490d08c3de6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12969c8e06217c290ccfc781b943ef4d0854add4c4b163ae433060a0fe5728fff9f406c61949df095;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22fa5afc07895b43a5595fa306b9ef76f26b563e57690feef1f54171d5ad09bfb643e8f0f287c5269;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb655aad6aa82992336625be51e46262046afe23576d5b72afafdbc11e642c24118f7fdbd104a7c13b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20edbe9ae8ffa1d3368ef61f13f4295d95a9773e104768ac08556a3043c42a42d0bd49f066bb01271;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ea4eef43af76937659e2aae4116ea34161931f2d8b5be3444f370ca9e562d7232cc3d0d5f007d236;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h555a33ef4a9268315fa9667f2247640c572eab1349546b6d88de35fd1c107b193a1b06cbd400bdb4f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94ba74157ba3baab79769a57565d4cf766577afa513780f57fffb889e6c8cebc6b7d2193f79d3160f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd90f7397572601f38e6d68af6f0f7467be63ef1afa63583c842a94c627806e25e9225b37456a34b79;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5bfe90bcb06d7771b69b556ddb5602f49f3b15f9b5aff8ed773dcf66458a2b9011f03eecac7600c58;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a1c5855627b1f030a806b687832baf1e65d2b888cbbef94336d70a3ea0652a220f0115638c805853;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf06fb2c60d8c106f39cd646a5c50882769380f0ee76ecaed5030404a4ca38d48f92e602f1b6fd54e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61bba6b98394ee4341ef4e5ae05aab16a573978500d8fe41d15abe53faec60608bb3d865a294c39cc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h579a781aa472e56fb08d26334584eb6984238e7f4d876c4af8934e393eba621a35de2f766355afe64;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h669563b207cd1f0229fe5ea239c793d6f2990be5a6b434fb88e3920881f88af74d3bb048207a98018;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5828c742d095da654d41e2c410a8e58675b5732830a6f3f92ca1037a50dc72505ff5a4e733318a78d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16ee01f2f22db9ba840c40e577499d1f2431f2b736cfdc12a2292144d0c56a3714686efbf211ffa64;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9616b7977b590dfa9716fc239263f10fb81a71c6c5b91b6c18caf46429b559888be17f2c49f6cd48a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hccfa6453ba37a7e6a0a09ea4a9b3eaa32ff805227e7eed1ba7855d864b841ff4c1f60d7124366a0f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he04dea033c63bea7b1da074b1ef48c5ab9f7157beb1175f91d7bd695ad4633143de82cb0a352d0f0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcb790b9fe3c68dbef230090e094a419ecee0e181e27bafe683a99aa07715220c610c9f5eb9d3d100;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h951826f33e896145447d47076d9c0eae5cafb2d9c6849186546afbd4bbdb35f42795d12086a3c1af8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63c4f28c119f7cb96920641fa3ac1eff389fe47aa568481a14faaac6ef90d006387df6818c00bea02;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h291ceef90d0fe57a3ea70459028cec0023cc9ac1024fb1674207cb760cad7404a85c224f3eb508700;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde2c826e1394d3c029da7d6fd075905f6a44b336d78aad9a15a3da6eebe5d2107e4d1242d5d9c493b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c013f5b07f3ded5ddf42edfadb2cd89cf3eb12b5c6cd3d71f5ede44fdd666d68cd4396c3d76f1a99;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f8e634dd5b5e7f037aca8bcb97048a0c7f9b658e926fd172bc3ffc0bed0d301e2db661e711a64444;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42dceff64feed43840aef39c7e58c282e7e4d78ae45c872fe35d18a8510f1a76353034f429f856dab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4735919566fc542582ed819a397838efd08db5a9c92e6d777e421850bf038760a301891b130f3b651;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he051af3bb68163ca61a466d705be448269a53b3d54bb01ae3297f400fadfea4171707835d63142e0d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7b729d7cda2d70c021e7a98a406b02f17d21325c4f4fd96ed9f133df6ac5ffe9ee29acc3052c9176;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h431f60c60ece8dd6b0bc6560c1d39766637277269193bb46b5d334df491e076a2464bd8a9a63ebe39;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51c8c69c589a9edd519cd7499eac162c08e99a4bfbc44088946c4ae6b41ee76ff79ead57190a66765;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4edf9eefc558ba828f10271587b44222ff653f0f18b8007cf17c39a8b8d57773db45a94a820b750b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf828cde526aa1dc6f193f7f9710b53f55d831f96f9e3293c743c613fdfc4206313e6cafcbd83503b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e45180e85eb576452c5e91c1cc3c52a9e1ef39876ce7e23cd2e24ed5677bb6db1f7b559482dbf841;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65e263f78564bfa586a7fb765157f47ba07a231a4d26c2da89172bb69876627421b006c2626e214e3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b48f8e30614d1f119b52bc25e53c12c5f2f5197edffb01be0bc02332b80e36431fedff97c5162a1b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a8c40bd43358bd168e1239a1e1309a9458c772dadf42bcf27c53b7d8a20f0e0c75fd88269ca3ee38;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he006a49b8af997a53e27319789dab5afcdc670bde190d3e8719e2b03861990744bf75ac74514c7ecd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafb4d6b7bf2195f04e5fe29228b8a4240a9c91d21906e4f074d340a207d12f65f3c8cceab06158992;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7564140022ab72fce32d7a70dd1287d4f57200927dc0527feb6338b9773bbe2ee5a58e5bed8e7811f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6eaf3c043b9c94abfe55e7e83cb84633f4e46cd027736095db79df17094d5487fb7d600b75f098e6a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h913e706b56abb63a3e605b398c120fdbe5306a8e595b6b39425ec6d22dd82bc7a13a97329f68a0739;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h233dabb28e6f394dae334ca317ca5d8be7e573769ca8129b3da259ed92bda4a3d8b51a13dbd93c8a8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17c166bc3eadc1cecafa8e44725e5437323058c3605474e710c21ff92731e87b148d14db5a4ca9079;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87ead7edc521bf48f4f7ba565ac0cd810e169ab0a15594ac66ba6268dbc95644e9e0b5e5bcd7c1383;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f7f47692e40af592a4931c9c254749790825b5f48ad79725d2a53a15f57d44efcf4e6b27644aab84;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e03f060961bb4844a253d07105663d1d8fea0d337af302c080b6a6fcc831585a05c63820654e905b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1575c7097545677fde8ddf468e630f7f149862817236c0a8fdfbe5d705aec4463ff27eb4b18dc7e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d7e2a59a927ee7138d357b7d0659f72a0b59f879a37aca14d52775d8a57a770639f841dc661e779a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc97ae202455596578aa1ae2a2ad2182952b9defc9074dd5e0e5f64ef46c2d2fe669b80b7d58f384bd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedf13f4df57a6b94c484d7a1b3ca2f2f280c024b73eae13be7ea4e2a70ef12a81d1773635e6155ebf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf85bf8ef6b5b9d7c65bf04fcc6c1b6f18699aa89d5d968c3335873ded2828c36e1cf5a931f46767e6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10bc80e9c8786471065075ffa4328a8c60c2437916d12226a86e3ededa67e259de02a561c163d02b5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7805e31a6b48529439ccdb8fe2e35a5f9a02f717e2cb8560b98214814ba957f92331641e9d88cfa0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e7d943d28759480c15a0604b8a75a02f02052ed4e49117ff84fb8b06981c2ee6b6bcdaf692c40839;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8df30f4f25712da78c145f6adb33da5bba4e8d6321e3a59adc82f211f619c952cae3f864cb8996bdb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde0e5b0c2189a88809217a72c711306518656d2f3b1950d14d49de839ab03f77d84da9b3ee8a2ddf7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h466bb7b93e4483900879ba2165e6fa6e0ac6882b526da21b2a1ea3188c439c1e8243def6e316db1ac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6ac7b57fca8defb1bbaf085d9db36dd6724c273df5057bac5060920fdce8fb7c44fbd636362dbe83;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd65c475c059a619d3d5dd1afe09371c3846f800f14374dff4115e82b675e43e5fd32e6fe44b69957;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h979b1376cd2ec78bc80ae41b8d44fcbed098a58da82388641ef0a28ebcaa4d9f3f6c7e7e1ecbb551a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1de31f63ce9d67da74690948e828971c777be676643c64ced873c16bcef7474d70d7eced0b3945e99;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc23a42e9b81ec7aaedb96ee10f896671e740e4fc779c4697d90d9678c70e6c76e9345221da2c84b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e5259e6070b7836db38f0b9b445f817eab95d9f0cc0a5f38fc0a9663ea998bc3d4ab5c4009a08a12;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd993244328a9c4559efe2c879d0fa7048d792dcdf0bc4848f3c7f470bb9d204f1c47d4ba42d676e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2832f158da8120a50907f045fb447a50dca1fda9460b66f78b8559f03aa88ea4cee25bfbd92af0f4a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he851935928c177c3b19716ce5970c3a72ab21b39cd3169e98cb4bf0cd50b20e24d9fb8513ddf88a36;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d3d0f28eccb42f9437274d67c76fb6d0a9c1c28b29e382b6d430e79d7cff706f64dbfd38f0774305;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24dbc48c8de32a795cff3faac272ddc1dc49e1dd2fd448d7ae362080500b39e98847b66c59fa477c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73c569c69fb2e96c4eac31c2a718a3afde572cd081a6fc297f63b485345613d850e772fba71529c48;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99cd0d2f4d18bcaf2f04e7a0f7069fc48a35a616115a08a1d1f6c9a7ea6b82781335ad2af408d8e37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd739da38b3785793e22685d663e2836c6a9041a9c81bdf7d13699f4d5cdb87410d297eebae892d524;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ef8b43f3a430d49dfb6162cb418283739325b5b8544d41b0b29c40552e6413a90319682819bc401a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9848bab5ada241486ef9cb0b7c2286a8f83667bb19683bd698a5bd313fb5a27e145d93cf6e29498ea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c4291e9919a12518b758c9199831847a2a022af8e77f52731cdd996d58f35852e9a9dfbe558817b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae606b9413a185b0f3caf987c7d900af477fc702c61c9714c827eaf166b215154516a0a6141c66814;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85696a151d53498147158e8e7e46e1d7474b67778342ce1abf95f690cdc749a8e174f901e32814151;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35d4a00a31d76b1621bd294a677f25346d09efcd26cf8da762e469206e83a1e76ec5cd65f93375287;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0ce78e6404cf02c0c285446960b655353f711491e575d8ec31c9f9d5de1baabd5c5e9d236b8af8ea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc67403b687bf68cf94fdb72ff733f3bf539b5d385f75f6ea5798d483476a0a768c5f5426bc5c03df8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31da39a000ac7e6692103534ebb831a190b6e12a493cbb2270935cd97a57a0c866b1405b65440e8f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36dacc3ccbdfd1a91b5ab19a8415e3260af211a0aa5eff577a742fff4150ceaab5783e766c5dd91af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc036a4cc3f6c834949bc6673bd00cd33399108fa1a55c96e053d300e8765088403c94046bc0736284;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60e33350f75d8d843922963197349043b354f06e60e8a7f91a41756476776a3ed1e59bae6d65d034c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4a92ca79a975abf5dbced024b90cdd0b26afbb4dda9c0a4ef3da4cc410ad76ff18ee33b852a0c5c3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h311f5df398980eaa9a50d429d7957dbe15f1dc91c3e1acf3e004f2111ef563c75fddfbf41edd7172e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3031f582e423529a5c0446c8b529eb0b6faa77a348a2d1a24adb6f939978aa7b68fb8511f76de8ca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbeb5d58ef4be87646c564f404e7fee78586594f6cb01b57851ed12cc000b89defb5741e5dcbd2fafe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76208184d80cdaac6ebee3460245dc5ed2cf824cdb98af6509200314a8a83c288e0909e442af43c3e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdefac6e0e36418b08565e0f59b5a039399f5579918bc26541c80ac6417c3c04758322fecc12b02f3e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf41e6bcb123621613c484fdc011a4c075e2caa0cc7a883154fcd07562d5a1367ea3e258436a3ab118;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf43581505fdd35b3ca3ef66c20e55618b2828cef305c8b2c3612349537a512ed6879cd9d5f3bf8134;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a8a373130e9d095ede68375755b71bb127f708fb4322f285191556f446a1a984656a65e22bc5a38c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h487994e6b6bf0a31de2c0162d45009b22f3d38d93c6cbce2db58bffa0bc687c7f9935b475902684df;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had7764a4674220c6c2a9e16b254471985aa3a79f4afc097373be903ad246e6c1f2b1c8e33ea17d9a1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1d5fd42d6b7dc1ff8aacb287a963cad59428aef9fb145496f57adc64957ed69f35d72635b780a67;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78fe28b4d7f4d76e45e9ca669d9ad82da6f0354ae38d9dce44269f2a059e7f88241f68bec95d32b96;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4294243c24c6587130895913bf1c695a4e9cbee2771801606bce1ae5f3c362e02eed15098e1536f0a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c95082a98917fd5221a100cfc2c7f37f1b0cc0b90c91d89ff2bb48670c8096bec351a5082ae13a52;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86aabefcb87ec17e48de9535507a0d44969a52ee926f3f8b606e592d82f0637ddbafbd7713949567c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h558652482f9d66b965c6ada6eac6bd5b38250e61d8e6c43d1679f3b7352e9051093c4ab05ebff9491;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce6e465a046176217132f16171b3f4d3769f8d42a650c90fc784dbd092f509323dd4465885467e094;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd623afec593a80630d8aa291ca1d657d5c9e7b5ffc1d948bd81f5bead4210ffd916dddf98eac9d33;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5bdc247cc98bc0b3204e99dcb83d997ee2868b31c1abd1a8215fa27883c4b53c8676948d6e8010d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20b3f452cb105341404a7844d8e203e5d203eb13b6b204410c01e4a68d684e4ef9c189ec3f914137b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h684e4abc1d4b8a91292c49d920d866518b1ae2604df82658690588e467fa3300174a1fc82887f231a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4503633fdf420218eb78ef1640c6393f6a20a191bf1a27f522a1cf7b9e4a1ebb2fcac6a13ae2eef59;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5dce91e77c520f410101873df88e5951c9ff518e006028389a9d758a7a7a4f7afc04cd560c6ebc27f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae1a5551d2732aa93758549df5da08129988715a2ab7dfc9c32db90061c40f36e093741188a9196bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbdae155295c959d45f72ed0be89486cbd9abcb9f11d241496cd18546446c151054cf551e570168bb6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb53aa569cffb16038d9cff631237a033cdda852f98555724d18ffa720adf5fbb2754e7fa5bbf33ba1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73563806f49ac91ac71bd061851af3c90d616e5c537e36e7bba55f4d150edf9e246714b99ecd1be0d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had96656295f6486411c11dbad11f58b676f2f3c7a846d6bbea9e387c8962ce8d2a080de3ca58feb6e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7085e328c91eb74fb4f453578b988177bb89cf1ef906f49239f4ec407a89e7c3723fc8dacb9c0e7da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5faef7ac738a21c6cdb77c40365881cbf22b41bad2f787e4de5ebd6645534788d9b0955cec2e6725f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a3985cb7cca8cc21249c75679cfaf8ceeca2b6cbe4d843ef473f0e68e8e096ef854bfab44af45164;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4e67de0150e06f342abadccea4307b7cc2736c61e2b07598e45eceda5a60f075cac37614250905db;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5a4ae300cad54179850b1556ea4b122914973faeb3ebaa8856ae04f0389296d32971be7c5b0cd8f5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb47e0e81efdfccd576263d274668c70020488f3b0cbaa1cb2b334b237fafe952c091e96c8454b26b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haaa1239d6b57d377527a4feb7fd03f85db9c566d6f18ab6b62cf7b8b313984878dd1488902aaf1416;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3562a6441aa3654a51109f418e8cd6681f8b6b29a74828a141a1f4cffdf5c485b866c182a7a47f79b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5daaf3d05a97594d535d60f96eb5ed52b9eba21939cb982561219d12b56154a054367e6f6fb15bb5b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f6305b3db909398295ac4c060b191ab73a8e02e9be1d221d298882100d07d299cf7a37512036b760;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63c2859f7cf950ba1d5e070b32e2e2302598f1a8b67e2df6158cc28b95b40355744a37613fe8a3406;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13874b52a03b5a701b2e19d8caa4114ce524ad871055bcd45debbedf753cd44b7013da3c727a5f01b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb13dd882295d99fca2c5f38e8b52245e5413a3218d7d990950a1e511894b2c68aa3dfca82f64b03d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc29a1abb82ce967f1f45e7d7780ee227bfe15dc7b1d14aecf7ac5632d63210c304533e24d41a3de83;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3efdffe05431f4e52beeb4d8c95df2b95b225222a5e48dd346cf1b49aaaeb8ce2d6b0cbf48e5dbe89;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d9a3cee8110e93ee30662f87d6a937ef5d9b31ccfb02d5372236ede1efbd62c4b4e026543b312786;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfefc4cc410e718bdee3b8613c7d48a8f81bbb437e2c42a2af1820fb8de6525745430f427f9c7d6691;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64755ed456bf553a803bb7693c487d323fcf0d40f98a4ea6fc6a3e224708107ae3ea56b0a6ea08dba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27f1ded0f91cc20d6a9b1f437312b705b340f514219b5329c846d4c88e1e295ed2afa875d328f072b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7018e4c67c95d5f1d5d398fb940f4b6d7471bc27f83265e908b0e620ec0681391ff22650293a6d41b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b9661e1cd2da3f8df5931e85885a53151683b87e2a141f4c9178c8be1c50a5de32c0c76517d5f49;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf34186cfea5c43bbc2a3dc395a2654650399fbf788016b14e945d9d3ea4b63726b41377b555b4dd08;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ec8aaa53c12256d0f6e6e811b21233abd0c0622e64a538453a940864365aa73536f42e700633b81b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h646f0597f5d9f728b2997a0ae5948120930139f5bd85f3bd2347971317f8b39a137d569c7ce2f98af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa68ee6ebca9ddc29d227f52292b6e8d2ab657e6c4501adebc65acc84d9f5ee316674abcf812c48df;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfa4988c6df979def82ff40881a2ec9bb4952306ec37b72c525654519e3a036bfbfc7eb7e28519920;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40465d4bef69d1275db07fde2cb922ab757f1c94e11006468950a054dd791e35423ae3ba7930e9b12;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a9e54e44ddf802bdff1dec02c4d8b83283437619d2cfd12cd14b13802d52ffd198e340083d85908f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbba3173e24e308fa9943aabef2e07cb0e17f66e8f3333b3d19529c4fcc73715542084cf972cefdcd2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85feb1c1776374961f5da7efdf3f7427d8e28b56d792d4f3cfecd85218b6e97770eaaa1194ffb74f8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd6fa443924d57cb234ace6d83eec6b9776b12390f78a23dd02bf197477033dea6bfe8b7ffc5d7324;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7826c5e64748d4517271b30f4ad72c5971e3a31f327af67a0a1d0925eae69706b461113a5face112b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5bfb2ab4ab783555ea2d8319a758be2b5683795f437a2450f9279b47d5855fbdd318838bb256dc973;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h823035ecb2510f292289fde49cdc94952d51163ce4ed4bebfa19f1da6628384665f25cc5aa1d92f43;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36b91d6f332745c552e8c01ea8c4fac9e51135e28d0de70352c4a786d8c5f940a382f6af5377b819d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15d3e2047a336c9bed51b2e23077458b98c83e13bfd1ff3159d8aabcb6a5e9a6aac4622ffd5a73f40;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71e1806a38e613a67368fbf9ceeecf2b738a2023bf25584b76f1caeadbc14006b068360448afba4ff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9ff6dbf490695067ba5b6f66028c92b2246f534f3e406f6a62dd05576116b61b75bd57fd4a8fe349;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha489bd0c9b49a101ec7837a9e93fe19fc68cf2ec6281c70424e0f1dfe7f65d121e2326d87535da7ed;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f32b798afb63c2564af2cf5df0fa140a40728c2baf8a45be8740ef5be87b653644c99e721ea8b73c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6259a2b883ace45b297fd270865f7c3d883dd238f7007e5ce7f83271824a30c6b893c07e44ac6606f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1feccc3c6648059c8cbf88d93e513ccf01b4f87a1ba133e8801e27465743bc30dc04b108abbf5995;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he72d361c5b857070015571b6cd0289ef687b9a7b35b87933db0b13f0477e4b82764eb3cceef5bf1ec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58cd9890dedc52411590895e5c69a1c75ec1c4a085dce4b98261d917de0692ac5609276f1f2afdcb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbd2b2b5213ef46116b34e403515a18944f638421fd06a22dc964a933e297fe96d2a593dd0ffa3590;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23a19bedbc9a57c0cc7b1338ea5db2914ddafaffbac3dff9f6c70dc67aaec4493b0074814a6397c80;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96982890963fed81b171cfabf1957f73aa323b01109064ec72bb08bdf66b53f727dd0ece981ded853;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2524fa0eb3fcbb206d4af0248077e9a5c2cfd28616130e77148705bb6ea2c61dfbb65e1eab84f9de0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7214069ad1ab89ad9a0b889c28d7b3c51bad1363ddc2a585344b74b365517c2978b908b5461cf4a1e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf6c761162cfa7c61d33ce9a7f86d4fcdee519395d87514477188abde759a64431d26a21a5a2e8a5d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68fd4bab7f60cedaf56c27d316e7ab6d5ca0331bbf2f944ad34c4b23c564ccea188ded62a6da5a7bf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3bed1310516e8e1034015fbaf71f96936c43e9d3410ea3c6a60fc915ed44430e5e2aed115398c2a34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h879be9203fcfd30bba1887d5d85a80cb3a064d0811c22e1e2e17049bf378d39c0381d39895ff81bad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd896bb56f954e3669f7c9a61ba85fe4cccb9e9f72d88f16df7e1151ac36a6ad2af0131a41ccfc418a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ac7d79743259bc3fa0b18900d7d9ea4369e2291622f79a5d98013031154a93a6901c5a2eb2f864a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7eeaa5695dea98b2c166cbd46dec2adaa30f5348ec0c3a2d0a22bd9dd162dcd0dcd26b0cb0c4519b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72259dc266857801a4c43d2dc1f8536bb3397bb70500fe93f4154beb9a87aeefc6384281db7db64c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb7d36b52bb8c61b843f35a379386ec4c61c79e597a32190a503bb957bc67fc12a85efa46f384c12a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h592d3dd5cf168c9b80371cc640405c0c4ab4b3f6d7840bd44aaeaeec77bdaafdbbc9785dde6df84f5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6fc49278ca5cec63abd03fc72d7ce3bbb32af28be14dc7106cce820c75bde390ed8b0f44fcf506e58;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h385158f40251a14fc523f63a7fe4a837f21058f57bfd747688e21e7b49e10e2423fc4219a9ed2a204;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h444e68ea9ef8023ec8c77d0968bc0e4e43fbc02fec00d40ce51779db77753c43bb11c583c91979d18;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63c71ee409b9f01594238acb08b63bd7027d9237be6f2e6ef944f02dc9f297cb32789296119d6c353;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h736a089d70470a680c9de5d4769aa03c371fef7ef3ae0515288951e4e14bccaf255c3536edd87c2e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69fe940fda97358c160f9da83ecd7014d92d7fbd2cb9e3f4fc3dfd48deaf65ad04ddb450ab297ab06;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27cde3be6f98db63e4b5c40db54b97936ab022b7fafd715df1ae96c29bad4eb8843cf59df07bf5597;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h268d6a10f86c392b84754162a59f6e22cf70afa0c05cbd9359874bd2b078419badd7c6ae8ecf95528;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d023e852070ce774d6bf98ea5e7dc0a59f63e9c1e3a2f0aa5ed135fce317a09d7f47c8aff002c99e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85a46bbb676bb1e2e3d05da9d5591dd77fdccc6a21dc56357ff0451715d4c202f0029d5abb5e07ca3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e0eb72fc236bd6384d229b7198cb0b45e6c523d27c2a55561326a92e7476a62511b1aa676e7be922;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha796e2edbeaf87dbb82f20542881d61ba42df412cbe0ba6a295800811e94e69ae801b731b927418e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a2189ee2416ee048fc842f98d5bb577d4aa6d0e35667235afdcdb319f9632cc6b499ca130495b68a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h405f92adc7fe2d6e215880c5a2f06bafebf995f5031505a4a875b957e12dc56b1a2a1d4e82657669a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89c919333b5c5626f6e449e8622d313fd94face7e2586ce477b65d301c31f47b8dec94eccd7781893;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h744b6bd84b79f90691a3eeab652678c304d307756fb9a9516de144b6404677c9af06e1b1ff379e531;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40f6e3a2b4fad631bc8d313c51b7f6c2c6ee437452d7a7b75a7384a91f360a748737475c8c72bd372;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11c3022776dff0308df3fea5d9158ee3245a67be5040d52a06b1c148be4e59c25a8db5753968ed60e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b9d2c53e8713793cd487a762c1f288e9e795101acfd6b1d8049e27d971cac3aca31f8e515fc375d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b1602506c0b20e307ccb02619df6a9d128efc3d89a830a221f608f3fa491b515d6e0a5325667c77c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4a5ce494440dc6c6ba2250e1db91f7e051326886a837e5e7a3041987a3de1ce0309719caa0869b8d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29d642a74b78851216d58704eceb2573605045b5847191643748668c107651479e0065e3b22b8ae85;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcaa5106931a8b4ce07178d286630977fd5f23c71c945d6f896534921d236a893b8343ad50f39fa674;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h176270de6e79d3a58ca873252985bf422528bad20007ec51cdb28bc7af6e578b2b36218b21f88976;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc5459514af4ceea358ec720266f1d585e9fb0665a7bcea77239a8a49dddec281b905610ea1298035;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h850419009f03667496e3050cbe2a78fc3c751d00c99e70fab562aee008090b98ba0d25eab637ac8f2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hacd87908ab3c4c05a1fa2e85569c015012b12c0f0c9d45eae217b2a1f9b7f792559f0040a47028772;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48d5fb829d7b6d1f69546d629a093a589770c17ec25df4299a882e82f0d05c8189ebbf28a05549066;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2d876f102a2d072d8a47bf91455f8be1609b44fa6958673f3423f6be938e1adaf4eb137370339247;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h418362a5437502cd972811461f6fd7386e77ec4a50a042b60d17e9ef3a218fae9c070a9d9a3f5fcac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h430cfb6e26d685752b44263e367293ed68d51516663a3c7ca2135e470d87202b1342c19976f974d9f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h463eb31fce0bd7b1179136d5f67d07d4952f77a670a796a240e0c0877014c5f38281b532cb77021d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h174774b2973aba05fb2081e9d3a471563091af5990feee5a87ebf6eb0a0bc15c05727bee23abc8b0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35c7966e3f3396c816758286a6eefaf51047dc5096fbfec76193318804341bc65ca4e3fa8bf4570a0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b48188eaf4485eed485e3c756f827769fdbb88a7eef00976e8dd43a7fb701ce5d9d8f9d508afa08d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f49721f3f1e13935cc331e3676ad06d52556fe91ea05a61099064ef9d584e4ff348b12bb1a9ea7eb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda4acb134a847b535ffca5419008906657cd1c05a4013058070ae4e646b5fff71de1b2ea5d36c5d8a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3101f877f1d2a490ef0c6c4e23313a4221d4356fd8dd30b8042844a40a5623c2b5f83a8465c45b45;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha422284424f13062d4c21092299cc6167bc6d4fd6793ddf8ff2e42b504e1718a97f4a5825c4894717;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h162ee7566056809d7847a22160a5c574e98b1002d4db4615fb21759680480ef6b8059c776f1a8d5e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5869d8612ae9545d4e10b13b7ad32ad428b8f6dd5a9cbe3b4338b5241c5f6b945104599aa9483ced7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e88af358329c738bbd96b13485d05c5e9cef1708cf8f9ec95ce5bc1a36393a8b6382c801fd12a89;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcc98e9e35a113465efe47e94a4feca74357f6db9724755489de8fc5a7a7338ae25fa1fc6b4b35706;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe22d4024df8c3c88ee355740c26b306a1c56ddc1e756df76376196fce1b68bf226ab633dbdca81fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd87c3492ed580015a87384aeca48625966df0a57a664805f229cb3ec3119031114a7fc66b04068749;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1bd3994d3b1696a414250082328e04219419a370959287dfd2200a255bd9c36acfd8c35cefd6b435b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdba0ac29d001f78c3da788d6c89fa438914c1c8460af5417dbe0bcf22c8ea53528e50285355a082c2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18634af7b072685f936ac3d1a9cf404b5ad7e62e224441b9c47d44f368cd47b41ed79c60cef8795a1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf062c54ea8fe99ed0b37926467baeffd31b5bc6af148837b6d9fed594368f68b95efba87a371c69e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h657d48ae27a9ab1c37fd7a327292a6d75115c97d9a437259948eb1d69a19ee4e84619f62cc5111a3b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h126a6fe0703afb148351e3c92d9a87552f5bceae9e6ca5d24baaefb9a8c4c5309e5db64ab8883a7d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67736d7321d34884d315dd736b715f1f9c66de29916921250d1fc50f7b02d399fd2549a834a642cb6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf73406dc73cad3ed662c6ab2584e4efb9d34e28523a2a04492c52aaa828adf017a0f7734d88b50afa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f06dd6dedac8fd7e5f92a9162cf6c9f0b7c2d59cc45afb0195643cef09b0e5773b2210a356f36b83;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7edd7ff1e209d94ea504af70719155dc65f6167474e4af6742c5323eb4c5121db1fa90ccadffe03fe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65d454c961a95444cb4830a6c312c5f4fd10bf1e80cf5c1accbdd6f43381ee2d08d112b096a7937f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b296be404b19803f48cb432f8967bc7709aec0a2138e1c7eb1403c1847c91c1795dfaaaaf8f0b59f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h116042a00ac3e6058b628d44250e9fe8c7e071e835540a8a35ce27e037ac29515521e3aa4cc8d9a16;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81df57521e2b6549572cc673e5ac8b0e287204e00ab595e82bf1cf42ec468845beda14b0c3ee94604;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h815d77bd473facdd29aebfeb9e5c3d9a6f071458255d70cf01f14a2e08d9ba451f310b4b8525efb24;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0a05b99b900366ad1d8ae02b4f06bbab2461797bae46e6d6d6ee4ac510db5c944f1c1e9346dc8c33;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8412a5c5e71d1e9b2c03d6fda7d364aa14498f5064a037c047d6454a17c0e8160a5f510ddeebc331;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62887c9cb049326c3d17bf6b151cbbe884e0bba025653e54e8f55530f30cbe5c49819f5dce83c2df5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h944df811d1d67b4ed16b2e5ebcef56cfae3742eb99e176864c859898e84c0cd938955bea5b67a63af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7a39a4260061a0099207a30bbed44c297cbbf7bd7b8de0256fa881e275fa9f575424e4361f2589c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99b97542f89f3a09d3e69e57916f109318330f6d7d6e99d0a5821d425a008de6c67cc3aa6ff47d41f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45356e045ed15ca6272e99f0650510746b1ef17de343ff1eb0ee9e05e2f0d40b8439c2ca75f4bcd58;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf13af864063a7558e3c89fb5206354c4c977bab1adc9e99d18f510c9c2566b00a9509b64c2d38844b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a76d19620869a2d65fe9b1c3273d3a00794beb901ba59a1d6329a066d127d34ade11bdea0957ec2b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ea9599b0f9276539dfe4fab32d86f345c32d768548b6dfe8f93faab2a46ba4066c1cac32396f8d23;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3696dd8f1a2901937381ac0de22325f29911c5ef7134545c1859e3c00091eae4b38cd10c45051dfb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he65aab6a67181e183d3a65a738f42c40da18758af295bc655e57b2855aab6e1732a8c3f667fc93c68;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f6d30c081815af39ec728c860a49b9f0acdda07549c528c56a8662eca83312f1abe10c597c0dd2e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d5b974077bb13d04f980ff05abc7a148ec8629227e5262f83349ffd46889a8157cdb457c870d838b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41e14032bbf4ae8ff4c2f6a12ea29eb8877613ef448a9acf683c50b87b27209e748b5a050ad4f3cc8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9c50e2d5e945527c2f62ab95eb5a09475645c4f5270bc9c74a7c12dfcaa2c71bf06c09e464cc6625;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1d52d16d4bd332b340a9ec3dfd49ac8e59303c6c8c4122d0c4da1ad574b63770aeed41ce77235590;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf41f76201fca34a9dd15ede5f806991a3c2845488e5ecd43d9938445017f425458438a4c75315cf7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h285f3eb0875ebcdf82da56fb0efcdbee221dc8db785ed3fe500e0bc439e3c5d3517b6a09bf793f3fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6da26b5be99057db1c2ce2d5e2b7ca62643a281bd879e13d077df7294819b81072b2dae68b0a1228;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffa70ed4126217f2965c58004ed9cb8771c9a1f63e80f1a2e50cdf878f1c7e4aaf5696c2761b3e8f2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3d9dd94c9af028df973353f49f4cb957f06cf382ec1215232f5c084775e8ee617e4148d808884a19;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2e0ab83ef172d293b677b9db687bed7c0ad6d6bedce8a00695dee9299046c7804f4117a224a608ef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f4bfe500c340f3b29abfd431b573fab13be91ab048e709dc4028226212618a2ea5232387cbdb86c5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h307e2ffc6e4364de93f0a8815becf00b2223698ab7832edf7929a4bb8192f424f0320a24dfb4787bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h319576261cce8d2b50e66216d391851a58725be8660103159b1eeee9d04fc4e9ac146ab695fd70a9c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb719a0d7c2acedb7ff4d779f2c616f6cd97f783eac75282556a02f4bcccbde5fdf19650f39dec0765;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f9cbe2c718fc62d51156060bf18efea851273899c8d5c20ef011b3ee7123445503808b365dd832fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80f64cb787441bfb0bbf54f39193b091dea9eab582c6860705df655bbc0ab9e0adea2a885682b7cb3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f772ca77a887867d66f7e9df45debd7d9c160b9ad976579bd6423dff6de46eb08e598807868cdb91;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha051f5e59880e22bd99c3d2604e8ab783f024f552697a6e4b21589d5d1b3815296234cc900cc54a52;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1deb12e56eb020b885d53962abdcc781b895d15357469b2b896ddf99ccee31d47d017345cc2d14044;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf42527ea333f12a619e79fbd339340efbbade7326489e6acd1aefbc3b69fcd9f8a88c9be9b7e873c9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42cc344d839e44fb681189746e0f5affff01c558eb89ff3153210e2cb097dd420c82951cd7ba25003;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53760f0cbbce2593f73f2462a40fb8fda2fcc447a3eb202063e8a8d93c1e8163119490ae07ecfa61d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hebfec0ddaebf43f94f4829c5e2c828717b5d3f55cded4456ede3b351117065f36a273c758e0bf0267;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b36005fecf927839ade2fb437d92bc7a346f27dd731fedb03ec2dfc8c45456e3df1ab0723406b013;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h880b9f1366e204f5c6d0a0fe61bf32f1c26702c6b3824bb18b54d7ad7b0282e8f4694370c8d7f40ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a5ec650aac25c69242446cfabeb0386525ad013ace464d6881c0b4ad425788e943e712f3f3c16ada;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ab116bf7419d561392508f1a34484d14dbb5758aacbfd1a83fbef245cb07eb7011fd9b500db72c29;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff84d224e1d917f526af25ecffe2fa5a48afeb12371d3f5d5143dd87ca95549a3ed1a3e467d97585;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9dd40356a0c02d8261f2578ef83a640d06c1080ed0f61774a79de4bb9f7987da1991a4f3614e9af20;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4099c2e8eaa38079554ded58c3a996e2049869cea9b0510c309fc25a9128bfcb88c5437f5ec91f4d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h330282045879b9b88f9056df45859e915d84e706dd46a4319306dac67ace4fe67ecf6c974a68d6fa8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2a427065e3a25fe89a7cb2175a0d65dcee353a4ee84a547b4f9f36bc881db9cf15359be895de38a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd23118b47937680ed482120b30b2f483385d36a1f9c783f516a6f428fc8fa05be1e4d4b7e08d476c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1b037a4ec3333489f7d4cb333769b4442d2336db8bce5692a87925bdc34d2f6f98890e73934c11f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37a2b46b19bc1a69e418f73e9464cb659b288eb26c6958fc9bd078cf96ad1885faf502daf81f6abbf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7379f5fd3f204f31431e19d60789081afd0ed592107539311970bfcfcc5b4bb1d765d1103e092e4c7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf3992da16b5158f2ae432e0f4040bf190be54ed4dfec65ec3cda1f1ff5ded37a159f10ef50d485dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8269d088836c74a2646bf833b5376203f658bd8705d0972c7b98548ab3b8d822c293fe516dd452e04;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf918b1c142ec3b147d27f855dda7ab6f69f2fb580acbe7123ad20fca5a568e1715b29b1958f29c843;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h124c69fb95f5902aac477dd568a940287c5b92e560a46b3ce26ffb3c351dc6bba6ae75cdf7d76ab48;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13182c0efc670b1573c628a42b2c5d8b5dd52f8011f8db77815fc972cae46a537a66bcd8cfa649c47;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4e36ac4f2eb5820a36d77b09de3f6b7eba890bf3815353a33d9669b7b70e9c4fe8b09f292307fe0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70e0f2cd2a46ae5e394ad1df7be0ccfd065e7dd513cfa0912fbda74fee49a874cd5dd10f27b91acef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h892f1613fbd48db663875803279f4c37932dd60d01965d917130b48223a4d4a584d81f4e9cdcf46bd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha9ff02896eb29340cf14185e03d241dbcdd63bc1bd4d8065a577c5b250746d59a078019bb979ccb0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb649f7d169f58cee722dc950ae39bab088bdbbeb1fd854c0cb4e7d4b63f1feaf0073b5d9d922fff1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7033ef286f1c164c792a5c4f043cb3cd785073661a693199cf2389916dfa2bec93995991f963b3d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9447823985f5b1848b91a8046591c3056dfb6821c0862dcdb413868c5cb24813deb316160a086510b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb86f663294329d6b0786d71ead85c472796863fa8cb723e5fc995e533326081bf43ceac6522b7e5c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7b230ac96302c80f00aebd3bcc8772d2f2bf65b537135bfff9f7d819fdece7cb2e687e2ae9e38fd2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9ed981eebb0603517e0acbbc190796e12f15578329e47520fb09c7b56ff72a279b9ec1901facb9ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5d15b504520d2b0d928816a4f71dceab536aaff22152bfaf905cd7c64fb00077d9135292ea7b715d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd09801dc142c962c78b1fc3be0aae5f4e92182e69c102f13d3670162a88c7e7f14df3c8834ee878b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19f806827ce1397fe8147f9aded39a9a099628126f9d0d31715021150cfbbc9a8446f99a13a00c67b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1fceb1dc341ff184bcf302bf84df1dc64ccb9e933f13c63a2de98bbde8eeb68c450278c618620e63a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfa61c277aea267c27237d00b25c5b3dc333a0e59a0984fef3b7bf85f0df15b5778284733040cccfc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f6546b90e843a613a989b32f3b4fa9402409d970e9b786faa4811476bc9d1e5b1a499d0ae530e4c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10c39032a8263fea17f7ffa5058a14c8b641f462dab50aac7299cef5ddf0ae9b633d86a2b5b008b88;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h284d98d8648140a100aed898bb5faf7ab28a810317bce06d2b80bb07090f720eebb0fa76f3549a0a4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ddab4714a1b90f5a376db16c14d0ce8498b1435f3c90d8a0a7d2a29fe38d03db8eebd245ed872c23;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc64c7ea2c2543904005e0711318cfa29184f8071764743813324b2b3bcd3a6b2a567a53ea7dc8c93;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1a8490612c7f827ba4c20a64921b834aad5085add869903a0c5a040ba327ee670f3446241170e938;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70689ea5f94ab7d9e529b99cba2fa54358dff1b1d378c4b71213e09fe73bd73db539f201227c494b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18d0cddf94a9ba5e128b622fe018c212aa762499d87cc13eda1ba25a1490e95632a42909a9db0077b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcabc198653ab7f86cb784ad43ca394fe39eaaa68f7911f8993fb090dc9ba756a8c0a481485b54c1e3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54883f3982b283ca68f179183831328bc0e151f4e3aca77950408e94e73881ec4d19b5b2e59a66f20;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b86659fd7b2a64d7f5e941ba7ac9f7b7fb2efc7bb5568f8dac2f54d8781cfbfce7209b18e91a314f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f738d63f9bcbad0bf37632971f9ded1503c15ef69072ac2152339207c576cdbb05b96ca807db475d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h972eb07c05e3f9d23abf3a314c8a2d1287c14ea42cdbe51aa1dcae753719868927b72b9bae96e5867;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16a6e2fd55467c301bb7bccb2e60d2fe67403cb7bc1ea7bd0ecbacf1c8626e8af36061cfef80188ec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5406c4937dac435929a30127a5067947d3c31797b4b18f881baf4ad4051fd6381d71f3a303610bdb0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c727db4bd55dfadf1445edf1d7bbf3e6959e7258ac27ba4bfcf747587653ff3f4d2baf355a7a254d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfaf1afab518be61120f1a264bf095ead0beb591a56dd679f7f2b81120cf6bc0233e27afee52b52ba3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1674b0a250bbc2475f01af96bb97aa31a6cef0c89eed26d166a729a69c1ecd7e924a3ee161211ece;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28a5f8a823ef4022fa98a4ed499d2114f8047260c710b6e9bb8536980fb24e905f8281482b41a2bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f9bf82a3711a4a372b66c35aacca40d985ce16d02118285565b57c40e66443cf45c31a40e1b5e890;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h279295354600482f386afee633160b56efc454639faaa31297ec2484f8ee66bb0ec31acf473c15c7a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9118d10478ec0adf6f38d08a3e3adddba6ec7a3a1fcda7b276a40d7cf9ff8e1403fd721c4a8ab93d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h752a2f9818287110c3c964d60e7da55c8dd5a9f5054602cfe6f64f2c1606dd22bdc968887b007f213;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h56c4a1d44e0f602dd9d1362d7504adbc734cf63582e9f718e1d22a885adfc063462a346e0ab707025;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hebf0ee599060433a564edee9ba93ba3cd989d0830b6ef8abf49bec5f5d1741274d1e87e3c0a6b6b54;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb72721bb6bc33b88729837fd99b01ab98eb2c4c2925e39f10b0100dff29cf8874674cb41dbc2ad40d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h731203a0f6b8ac600032e3007a0bfee5b8f507d9d47c57298dec820df7dd4a918d6cb2b024207beda;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5111c916dfa5940a5cd4c25a868bfb43538eff464b2d12ea086b5fbe94c44795fd85d910a81fcab2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31196025437ee71fd4926d2fda4f24c81cf4768ab3a604ecdb612ab08bbd31b77b334568759b83400;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d124a314ce1bddbfb6473d1efbbd7070ac75f799243d8bdbbdf07ef11511d8ce5eeae198cce8ac72;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf618c85c592547a180aa676dd179576b5ce90e617df353e162acc6ab5113cc04868996389001ec88;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18d7591dbba81ee09c99d8dbb4da532b998d80969f8124712345988ed1458e965566f5b556b71aded;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbca970fd32d55b74733117a5464001c08c1c864b301c084f6eda476bdb2af63bb52613a586414d009;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68a70bda7a8a77f74d6573ae64e3d72ade5864cbd32f672708e44318d3d34bef4ddb8a126869e1511;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8bc9616baffaf1830ddba37e116067ed67510a255265483af1cd44a198999692deba608ae15073a1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf33ba5fe606fb20681cf28ae4460fc509c8617ac377036a772e297270f5aec316b71836db95c39423;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2dba5a890232978f85daaca20b55b022c8f302cd93a3ddf4fab1ed2ccc35d38f465b48b9d510a8845;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12f1fa32f2c4835e95497d5089b2165329beca12d80567d73eacd38b5455b9c23773b398a7c1519ac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac987cade6ba0f5a4d68fa8298e1a8f1801204ef72aa69f14ede186626c91db094ddb2e782dd21d06;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89923cb4312e550aecb0f086f0b9a4efaa5cba60c365608a83c0c912bd26b5f96cc4d2e1994a59aae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd20257ccca36f552911d543a967072f3de6c9fa824edd68fef6ce855846241d73d573a8e6113a7bf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0874e3283ffe5fd336aa95a2b172d0f58a16030de9e23b4ca707544694954f499b709f24e2dc512;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd70d98115e3aec951a4a1097340ab1142af6065afddea6e6f2deca302802dc8221e6386445a0bd383;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h876f38e1fd2e6c77fedd9f37d45280ff88b2cce80d7d965b2f2e52394b8e91ab2723c966420aeac8f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54739baa705c0a24d16b19d44a9e0a0c235110c1138bf6137f0c40e3d08b504347afc69d75876f0cc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h606f79dd53cd0bbef541ec692586a836b2840c274d1d643c3e600e1742807b8e50405afe18831836d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65f3fff924355667d462f228c412d7dafe498af7eccc9bbc2ef6482e8a90daaf267cc9914ab9eee65;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30be440e72c24c02135a5455168869d7cec2ac600e2a17465c86775079e72286c2580d6a7b532d485;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43520eab6c6c14e4cad8560cc9679991dcc68663d51b1520e31cc2eac6cf14170d02deb4164f4523;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4831c26e6018793c11fda31fc3001ca22db991404db32c0e4729da498717d7252eefaf7fdaeeaf00d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd18f60e80579964a880e52c5243487b42cb4bfebe1dba2b3adc2dee9d4324c507c1382217101b7c65;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf01bbce567d999ca05c5e91504d972994a3f3d2093d87017b7e1c9248789f02dc4e5891009bfef00f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75e2c71864ed0f5b3b0e20f9f21a7689dc940a81c867f566c602b159269757d027864a85a1acb2699;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28e933c03e0b27581bb506b5bd0ccd47e631b6e8f5a25212a1692906eada49a302c2dbe1e7b821dc5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3abde1ae6c655b20aa1cf296a4ebe1cf3d3590f1845f017c57eb1c503f95905b28f8a3588a101214;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2cd83f92c22fdbeffc7bd6f9b5db58ed87137c8070ecccc6d4cd1a7e2bb4480d80b9f84a0431af17;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5519fb0eb12ab35d15982a03f36a6244f302da3a222fd3b1f8dbe5de714eca46ec3374cd3ce8043c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e03e4e50fb83e892f5781bf3d2d0f6f19ee455aa9b7eb45c7818ebfeb8ddd6ed04703196045d026b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0a84749f83e96e63f528663579721eae00af0e5fa300da458e5536b20a9036bfc646fcd4ad1fb4af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d3780e239798e11cf247a79d0ef0db2b4b0070365a141467d0f90908178e0371ed3d975a48539c5b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6fc931c89ccdd78ca6500fab3a75ed8bd11dc439c9c1ab2ad33c924aac39713f49ef6931a6fba9a8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79d167f51e694409531b259c306d89f9443ec706c092359564b6653f5c6155e0ebe8ef3c3988e03c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5fb1d79704eb405eb84376d7beed54b7b720c1562083d6451d15974dfffd8d89ea52234baf15e749e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc543d1a62dd7a6bd35725efac46b7b45116c8469c01db81c9198a04a54fea16d2f49309e09c76f4fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2221a678a2e0f63312191651a89ab2095f853c1e34720c426890b1b0ec86ad0bd437ab0c219995518;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf2f2f12109879320329645a17074ff2567c138afc636c9b280e4e56e2045ddde663dd185b108e616;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h686bbffed5e2b2563746d903a21b7faf801f02105db70fbe92efa52bfce9cd06f6fbbdc868d840532;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h908392e5df9ad652dec1b1e099db173c717787317850239256e5b7722623f61f1f60700c13807074a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd90db07076d4c30309d062e43b8583992ecdd3631065ecc07a0eeb7babb8574167b872c1d81c91c9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he781c3a05d967d104cec0d868e30babf1c03c6b44b29294e21e7e7e828e7001de7b118a85b2f6cdd7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf080dee34a40a5256039f8b384d6ded662038aead0cc058717500c3bf5e09aff2814c79816955abd6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53b6bd4f6982dcf20fe7bd132e30b1540d51694f78d69d87db3c37e36f738d3b2f8d26aa5cba3af53;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b50dab26a943e4f4c3c1e76fa8cb866f858f117034985147c6f143b15fe6a51bb9f7149a776b7d27;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he791844f66a9629b5043959550a3dae7ee49783cae31856eaa144c5792ef528b6a9a6018aeb2f2c6f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc53f2bf657397c34b9ae20cb3efbe255541259690373e88ddf4665c65ae6094a4cb6464149fd86c99;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc44a2908c2b5e43fd1079e4a03254220e730add38488126080707e503393c910a57feabea542f8d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ef1d01b6b40f93ebdead1efba39a2cd1475228210372680a0e6d90671e0185b824e0f121b13c68c9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbd5cc60f0bbbc0282f0815a6224840bdf638efc4b661024780a1cbeb53c1abca105b0e6735236639;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0026b7ff6e5d9effa5222bc6bf677c9c811f650682260c757115774fc26096cf71cd93d61aae8bb3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he20ef46fe5f1fdae0bc6d69d11ec59d1697a2332feb8ca30141eb157205fd4a37f90b3c68dae42959;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbff54ea80b867737558695303b49c6fd8c604b565e5ccfd27689c7e2d0fc198026232ce72c100ae76;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3253c0a020bec372170bf8e0d6eb42414c356aad24b9feb77e55ed54ef0b56a7a2c9f419984736bda;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6bfd582e0922679b7e888e610cf23777b58d7953ee8bede17bf87628867fb88caa7a93d2457e84911;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf3d6469d9fbead104162836fd67bfc7bd5c7b7e19b562b72e3d68c902b39b4396067265e72c01b13;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2992d4750367906f252dcc62e01a200185b76d0c4d5630b49c80aa0a305102af7ae9f8553f49cd8b0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8e055084ee944d1357bead4db0950036b599098c7d77306213236c659df6a93e2aedcbdec91f1f2b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdafb6b47169a8dab6f3807191c1d941e00f0608a972bbcb4ac8784f5da0921f59058c0ee2bf3c09b6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d6db172e72b21fe9510dc733fb510bd2c70794c149d070d704f287f0049d73d92c0e9e8279e835d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf91dfe84bbfe535329650f4a11fa05a056fe5977d4cb4888961c5e4138442dac7eff7ee4bd427329;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2070f76398be1e2c94897304328bb0dab537c526f96429a5fe5a61756e15ed2fdf38a6bae92e29f9d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf653c5aeef6c65a167523b069ead98e194b7d0663efa9828289dddb9549354681d78a6fc69c867365;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h986a92e5295281afb4ba7c17b327e63c85bdc02f440c71ddfea2912429dfa92eed14e14b8cd042cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8763a7b1ec1015b7410d01eb528fc7280254ef4ef4722654120bdfd2963e2ca4f0819eedd7e7be32;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f76d94029eb716eda5b0dc682484f6a94824d0dd2b989953ccd4dfda1e9a9b6994884100e12dc064;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha41ad727562f0538a1da72a111b4680ae8cb911af14361814f1d48feea51bdd3f78508bfe4788579b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f3a6b4e3d7c6c131d6b44480a0835f4be51e7239b4717df60744703baeb56d16873ed66350ea4bd1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8416e6bbd0f916fe453a87f230a60789420675218ca2f83fb64443fa7259a9cd2683812a90c474f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfeee6957ffe5650dfe78354bd11736dce5fb0cefdea21768d625c03b2827ed98c744ae2bdf8accc7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a9d84e18e0e054f3d51c4d8616d7c16b5eb65a4323276af81934d3a15e6c222483fb8a38c0b1c4d8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4124afb0233a93547a2b2dd904098e45d39a3d906ccf1c8aeddbd3a495430ff9f3663885cec58759;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd7908e34f9079b81f682faa34709519aa27cb57c47cad144e9ba1a183ad67f258899a4c990200790;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb84c890f5ac001e6151e8fcbbb9af49d78f3013495f83b34fc27924173e517551a21061bff6f803b3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94b9d0c21da200dbd2bebd190651c0b06db1d93b4355a00fa5b8ea7565506fc697b2328a4ba7f4848;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1125e960560bd035711e695c51f2bfeb44a98a5aab9b4dba2ef122af402313642a92b82036dd98685;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca8f310bef18279411327f113b065e00ca547e18ea447b05c141460c8a572b940dbfe3b8fe287e02c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b92aa6a8d3275da577ca1e48c2175ea2e402d17c0cc843cad607a33165c62ddc42008d00d6e48ec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80059d467c9de562401755a337220aaa0200770659e20507337c177698b9f9c46e047125343ad732d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h262d69c077175394764556947c38145c563957d8fc7df818a94f9e5bade8aef44b1a926c8ee9f3797;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b4bda5ae383d54c74647f0ba619d3b60a9f2c1bbf03f97f66e2bc7c9c620ca467f93b37ba2aa9625;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b766a39e45a17a3d12efb604c23d16188596bf2009fa2b4a74df6e52ed5233121bf5f5ab3fecd1e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8823732c6b8a811f6a69e98f789494563280611437b4168966c4f7e6c7ee974df16cff9228d2fadb2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3b904457b83cddf9d06842f820342732d8b213613a489dc2d0a0271b064a2f6c79817242b353253b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45bbe037bc841fa460a56d4150d6b0b69e844463e51f1c075f4926f56ed2918c7200aeda828d0b92f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3925f9096698aee2092fa6eab9d31572ad4b42113407f776717b7601f2b23b179a915dae42dc254b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7686793a33ed5659fec6dc470d39df5dd8533218b94cfcdb05be61f08faa899cdbdfb3aa8104a004;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc26ce43507e3f67eba1d5076bbbbec5f2e8913f8b377b1758210d60746f9c37a859d585c4f55594b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc75d64a9b21d84b20f19644726a4e173359b77bb33f21b81c9deb56f4014ede87b0202362e4ea2b25;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14ddb09ec80d3e54204db361f920b39cd5fae1f2d2079e5bb4e684f8ff471a6b32069bf9c0b16b202;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6a00682162c8645a45bcd0019d044cd69103b9ab4ba5bb4433eb1a1cdc5d063722837ae82c986e08;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h523860feb0c97889c626b630c5c1171a9342f0a4c4acbd380d61bda9d0b68eafcc3020ee237386949;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h532b196034730a8a121a6dfe1bb2a9bfc5ff4d42b9793290d24b00448a83fd07f45773f341c6070e2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heaf65dd6782d27f5e4cbf33ef0c4c9c2d142624bc05d39f7de871a69dd4acb84e91dec1469e5bc734;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13dbb5164ddf6e52376c0647e7b2628183e7c991672b0d3719e336cb2f35bdc5cf12820e74773d0cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17b3b76cdae266b5a17f169ad97760d3dd760b1caa7e89b8c87d00d46ee96370329a2fd5c063e0c2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h709aaa335f85d42b54c46f9aa0ac8008f533692ddd07547f7a7ce52e6701be9ec16760bac16fe1a88;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h808c825bc0e23e4daeaefa8c70b18f784606732cbf6874807612c311ed9baa8b747e220e570094731;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5230dbf976d51d28af2fa029a99331a683c5e23e5708749405a7d05da8acab7b34a2bc65b8bb45c9e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24df63b0ad73e0fd4680f77f119d9de272ebd0ae1cf026681a9bfbd8db61edf22c14e3adedcebb8ae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94bbc95a334a5178d1cd80a03bfcc8d50f7820fefe1af7f1f929576dc3e48398c26db2c915ca0dfba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50bf790c5c497e1146c2bb23fc6aa273db911cdcc4fc17b1bdb11b96c32017d58c33e70aff5a075e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd22f635fbcf24c335aee3ad8e072e7292f542d3dfbafeb983fd3e2101febeba8a8814be686348187;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf64b0bb157eafc8da9249ec1fac9cc2ff3dd48f2711b3f2edeee4d7a350af7e38f4a6def97c24465d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6bba6e43a90b0ff7736247cc48593cc71b9a30e380e2c3b8cc54a509744ccaab8a71fb3305b8a90a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72e72fd562ff29633a992a69fa701e3b1a6b9d75676b3946e030083d442c6bf0cea96f5d685640b5e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd8585d60801ba71894288ead67a6ea0a151cb1b9de8faac1f4e65b8a3c95b74cc88b07655b3e9585;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20ba1e29bf70b2f1b35d7763f0da871cc0abd47b8f4dd0f7c4c148ba26379e242dd6cdbbd8bea3b1a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he43498242bc4886bc323a6f99122d36b3499938590d323c70d84e10eb881fc9e583ad5c434582e649;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3495b1f45984b47472fa959498d183a47f43a33fd9634b0e51aef41c5d3fb90dd64b1b32126410166;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c7ea08910417fdbe4e3536a5163bc0822a20da327f77a002b9fe5f13545a2aa70b52b8e8f1e6d2eb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c29c6698724f0c22d686059326ee131d6606326a472913f27a93178f093063c6312b03825a6133e2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a5a84b13ee79bf25bdead62f7c667c5b406abf93938484ab478e6ad922da0eefba3806112b181ba7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53061df77330c7352c93d34afaca83f482296b6a0ed4439a9688e083f6359401bbe7640dd26c60de9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11d90932279dc31b792f0c350902f6e9c689a43d079908c91d8c3d45d9c1c6460d46b13aa784cbe67;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h593e4fef5c2af4610f5b8330d311d3b362c78dd7c48b6a2e507e19dbefa264cf1059bb8ef472bf228;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66276db8606e28da989b016718c51491af38e297ea333d85df70fa15c03d68c09c24860fa2a58963;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2042f14d38b46ecceaf351430e73ac1f6256c9159d3601089f081e5d5924c26f23f55886d37db8d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc51c0a2343e312cadd8d131731c745a8f5c890034f4f16a8b71b0888432530af33f41ce4a7c90d8cf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd8b51d87d2fb418e5326776d75f231fbe9fc523a3ce28a166bc0277ca0bcafa889e54d8075c42b1e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he855bbedb06ee524c5f2db93174f0594f6568433c59c242530a8790313dcc59d2dbc0c1723ac1db0d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f523c6c51109d68aff01d5a40a79247374df47dd919d6c3282759e8c88c3cea59103b0209293a809;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca47608388c4344bfafb87e4eb57e4fe76388407189c82c061b6ff0a0a3ba9617a0889501ceb17614;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47177c46ba6303cac201e56aadc5827b9d9811f9d338fc53057c719a2d164784ede09713cbbc87a0f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9163705ce6c11bfe0a60b1fc1685eab4c51a2724a325408739279ac47d9256cb6737c3a72f504551d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h804b7d7b12a18f0466e0d8e2a88db737885755b5d428194e789a8abe9af40c5ea07f3a52725d82842;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52684caba651095acc2c10a3a89f081e4dbbfc98999f450aa19298e8816fa9b1be4287c26018a3ac9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bc8f106c74532f785cc00039115c21e9eb91d45f970c5895fdfaecc7bdb121048ed3623b36962ef8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98197a19d945f77c43cd22fc96cfc1a8350a99447ca837846b0604637e43bea7da3f174ce615fd171;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4ff34b44ae126c2514bfe534fe8f74ca8daf4bd0bd19ba229b157e4b6f434bdf452219faa4875673;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf565617a01484fdd50780bcd9e69e28325475df7f4df0faa97463da04e98668cce361a5fb7ea9a8b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8caf03c492dc2d98af5a3c494716d98c1ee535f3c10cb122222eb54d5a369c72d875a4142dd264b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb935767a3d20dd2283761d94e3600ebf7e5895037fc4f9374406842c4cf7093b907509aac51e336bd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h697566e21b3ba1555cecb3338317530c18d3a9224433293df3cf7a3dd9336e407e79785ef2bb35a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68cdfd98291c702b9a45d82bc88b82b8e1cc6dbef0a258f7ecbc23f12e562e93810200d5d9733fada;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h772b0c4fc1c29550e5b45051f155bbc3cd7a362215a2636f63b5a6c0ce98101d4a7bab6c7ab864dc0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5019e1cdc87b2328ecd96442a1f7902ede5ac1b7301f4f84bcdcd46b412ed1a55ea84400cfa9ab8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffb73545f276e5bc6cc3a6c5bd7f79f16c95ae1c3d5887005632cbddeb551ea68c813308d0d2b89a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3339e82cea872f03345b57cee36695af21de0b8896a753e918745b733f4b773f7075c004e095d26ac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1336c4abc8444708c81efc4f0a363cdf404bc3358d5583dbc431da0f8b50c2dc2eef3cc028e191f1b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h111e09526b0353bf5f0959a71c66843548f0a309fd3286c4ce62f566474218f19def59c7abb9a0fe3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8b1aa53e5c1f1fb4fd0af13d9e98a9b03e163b9da0a0e1a859b0c0e58c6ac732810bc6528bed531e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6bbd37fb09ac0f47b415c95d95fd49d0e78c00bcf6f5a9be1263fe223534009e50613450eb3a124a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h330847d0002096f196028b45dfb21df4cdfc6f764c2419e859515c538446165d15583c4cedab2f315;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h245f3a7d47f404157339bfdc30593ff9907b3d764443de0fdbbf15dd2cd4ed17ac8abd3e8acf6af5d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d5ded551cd448418b15a8f629550eea01629ff7f755b2e0fd49748222ed50705d9677455b30e1a68;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha637d5dcd73c57a2fae19a97454d969379d004e2ceb634f085257ddcf69ff0093ff68f987005aaa46;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20c3758525773cd043951092cd6495bc4aa955e6f5e93c3e6ee4a9afc4504935e53931bfa939941c2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29cce5d2937b268c57e535612224c94e7a0285e811a584fd6b377f40627ed1ecf470937360a9934bd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a6fe41d04988f4df91846dd0fce170ac54ba129e790b3d0c70b2fc0b709d30a8a39ff0965e2812d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2196405cfe6d78240691ff750e5695462d3c02315c0abec381ca05f06cac8bc487f92155cc89f873;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74e4a6f9177752e60eb5f28c46bb6871786cbe70ee65790dbb9d686e517796dad6bfdf47d4e2c8c54;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef28248fc739dcb7454158af02ab703f4c7c11b145288cd69404788c13869fa0538575371b9f2b525;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78f515104cae98c3a79d251396ef9fbb2851c56e7c076ed8fcf05980c588d2c34f9e38af5fdefc3f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcbd43697dab1e42e5ea727bf1982b364dff31d95a54275692a3ad9d0933fb41d22bc5e733154bc39;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5fae0a4e2b921760aec4e2c16de2cbeb525e1913a23ad9825a66899096bd7480ed9b2eac1c06f8fd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1edafe34693906b4c1efdd8c5153d0d75785999926fe90878229461ce1b1e8cb1605f6377b8600fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h753b5a34e11ae05648ea8e7c39f5a10349501fa33dbb2cd5385e26e0a6719fadbaf99a2680951056a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ea967d2316978cf7d3aafc44ece18c93ed7c16417f17dd0b7113c16b828241f668cde386269bfdd3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee47af094d104ff9ea6d384f953b9b088e69902513b5f8e6d16d6172d92f1ede4d7f0b19fb75e47de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b62da2e4fa94c0eae2cbd92356e2865924f7429157e2532e02752398e18ecd3b46c1482a3c656e54;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1163dee8ad715e21d1494bdb1b35c3711a60a0d39b9c7fc9ad04426d9d2820a0ea906a183ece00977;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a308ea00b48ea92c2053ac1ccdb50e6c674ff4efa2e02849f1e37a0ddf223f1c8904734377785c30;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21e4e682fa95c98d802caffc003b838ffc7db4307c5dfbd6d9af3cc84e751cfbafba030d4b19e9b24;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a6d07e9491923d17b48d44e158758f75604002ab68b0a06b268df77f07605754acfb7f0efcd73c15;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb522da65812a2988b6bff9ed5ad7d69997eac1419d2759cf2b1e95cca86fa3ee6626ead120e4665d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5909f1fd84c280b1452f4e430032ce491e412ac5a9ca67b3d72a07b1e1963e94a83cd56b660cc9745;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8900e1767b2e5a31a5f010d92a5e10ef5ac440dd3535a1b35a85ea97f4f757c52ff68b7a69228aa73;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e61be98fc8bc9455cbbe59ca9e69ad7d4560229f8c3c7378a753cf5f05f16c42ff928083c853b330;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93b33cf98f601805f86972e3f45ebff3e9163adf425d66de52afd0d02456f3d2d30662eda7be0b2ef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1481f601a4dc1a7c9d4089908c7148bc930e47015afcce821270c0783dc5cd0b58ff2aeac3f0706f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec861724543556b0fbc74201158294db09be08428f656374a17044e2258b5275f16bf6c3268654f4e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h422acb8b7f151399c4111da8a0198d4bf978cf76bc9db6a3364c9b1ac3a5546693f6610e71ff9a1b5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82d06ddb3b95f40fc46ed9b32a20651a1b52cbb4fc7930144f4a8cf03225480946b05eb58103bc4e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc813d3abd3ddc83c7299f88bf04fde78d023b5bbca76a62f53eb280a9aeb806b01a442717a5b16d84;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7e2ecb2e2fd49a89a2d1b43ac105a88d2fe44ed09992487c2d7d77c8f67d768380170df80ca01af1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd395bbc1fe087970540fb6719eb53cd605a208b2e186aba76754acda66876648b627531e995c7b438;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6446a27d12d41ed85b50bb09ce331a202db467b8f80696a83d87f3a6ea980d95b63a816e89809779a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b3bfbe53f49dd765a9678cce96af4c393a02e84b7be4032cc5f7eef7d6e7020e213574866f78921b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58b1240d749156a62116711cb267ff20ecc713528313af5cd33419f3b61d0e7df4aeeb4041f4c8217;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47ebd70cff440c0d9dbe27e27f1371c367aa864cef2b20b0d6a8a70cc8d6a0775a3b287a5b06a6bfc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7b8e6a61ca9a2ab8a034b561fb429b553271b5b85aff937432bfc202ae62d7b13a3ae1c29db693e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2bd1b583258a5a166488e382c72057e5312c64e5b8735cfd23e3166212077aba535d3d9a621c1a930;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e834eaeccc671b962eff802c8f6448c4f1c1d65b92492026dbd91e9e7ece1c153a88ccdf1e0ffd08;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc048c2304d7f47aab57a952aa6616e79339944b862dced1d6a6062c350b53188504c2044dbe0afa74;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdddda4468091f718a32361dde1539207d3a02e947500317b36c46f4600a8c53de27fa51d2df1a9182;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96498096cfc3f3224a0e210b8836fd0da8a6ef0f93324ca1be56b645992338b6c90250f76b403a804;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c98a9d6052737689dc3a16ea2e8da2bcce79897997442320e6020b0f1c86608d4ea9e06c64183992;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h579787d60448ed42214764ad876bed27305b82b94c97eb6291740d33ced72474701360cec8985741d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb39928043ea49943a680aa4b54e11a6b9f14686ca0514851744fffee93b00caba8576faa14b7543d1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h938be186c45dc256ad0fff0bab6a7d69b7ad4fb6ae0b3c4506d920a628ec8441e6c83f40ff15fab1f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70f8fc50ab83dfb88050de9c2c33990556c30a6c9d7a0cd1820fc71992d62a894b8abcf1aee4db3e0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78a0d070c7e2f2fde7c502879f7e52ef92a6f641e33561fa3ad866c6b201731f4713b30900c30070d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcda165c825737c03100fb6a7355bc05a4a5bdebb9b90238ac4679871becc58e7dee55e550912a30e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4a4ce3e5412fdf3111c21354656ea8ab548c4627d75efe93df4b0996f01331ea5548353e03e09561;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5866c5791ba3b60cc87f163ccb580c838fdeae4d2459aa8d590a32e69eb56b935b8b612f5927570a4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h493f8cb05d4d7961ab6c146267a15a37030fe1aeae20ca111c50ae335f8f4f305aec1475caad598bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84d39794db2d1478f56ade2c1f771cedac9060953e61b16f4596dbe2d08ba0e425cd2e1bdfddea86a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb76bcdf18478f2c5fd0362f24743f12eb805f23c7b749199cd071fd7500b36be065c283c0ab4b24a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hade2e1408095bd19e79da664e6add7c1ba3f1552fc4bf11d42531a6f10dc962c0dd7e0c8c99d433e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h689fdb996cf0f12e3552a240ed1c55ac0eb9200f66e987de38b7743f1156b182088c80d5befbb8b66;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5209ff75973e28cbc806fa1789946ce2839d46c49fb91db0350271f872c3459175b62422c1cedcf01;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29798120e81c994c85352152aa16b68bad78746bb609e1b1e4a901b5d1899ecbb53b5050726458876;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89e80aaaa6746a5adea9709a276d7aeed1d7ab338f550be96b933b8fccd21f2339b14ac43f9586298;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b105f469ee7af3d6645934b4aacf2afced014b7d291b8d8d1b8c1844770f1c4aa3af1899f4c72910;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10b941858c1b0e4a5fc96a4e66b278330e9690d3584cc9db873f59683a5a0e696705d213ea771db19;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e793ba8b2f0f07c5a10cc307da9fbf62ec913f11a8dddc6eeb3441d609098f419232411eb16d3098;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h683dabda96e26d3f76b45b0a846fce9174276290ccd9d851d9bb5aa7d995d03f8e28cdab17ec37c18;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb04e728601867701a34ecece3dfe4e64a1d2bffb1c38cacdf463c8fcfdefd275f981438a23b9ca8d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3add8bc8a34e0eba37e6a8a31406be1a0368c4b17d783f0cbbcbb8260f5a8e6692ad5d673251e0528;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda1a9618fec24154cee2b5d633bb74b1dbfc06f81a7b83074db3afb05f2e6552f1f20eaf958e8b27e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ebe888706585de775113274e79a822de658993a72d6d3035b38afdfa3482409cde29687a1c52eaf6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h516e06053e16b62cf1fa8f8add061a958baeeb0052eb9689da1da5f2ab7bb7fe0c3256a6e615b919d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa90401a51736bd638a2b5bd247b924f4de4562d3a29de5b37f2f341739c4b4703858c4398712563e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h661b9808ec1d817f19b8621c8f4f37f59d92bfe370b1aa14c07ff5cea583e146dfd7d9e38f559627e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c94a690d2f0da5e60a5f585b76734271dc17cce80c43701ffc643353704d6b0962f55f92f6bdba35;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9195898190b2663b1338c860583ccbb925a1d2007d689c2a4612003a175fd796098a9a4717562ace4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9be566615e8ee974916a140544282ce03b2ce61b31c75eab1d4bf2b4c8260a4bace11642900139c37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6006b5d8de4b62a92b86ce9cf1e45554268cc62685648b297530fdece624f45db131dda19400ba623;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27f34868ed362269bce18daef6c460f3b1520dcb6313b760173a11746fe768287d89433edb58d737f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff38f6e71e3321bf968706b6c3da7e231d45bdecb83878593da55977ac99328fe3a8c62cc03ab1f9d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd500ef5b19bf63fa5e3918c4eb4e3a7c95f3fcbf21b91b6b5cfa2cd54b5f1afa64367ade19b67c748;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8aeef460442de7379eec23e32e64012c28bb3d91505b70d2abf45d774fa59117bcf36163176df0d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87605dde8d02c62dfaa2002a023fa31f94d190721e56e4446a3703edcedfb45379d97818cb917bc90;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff3e7ab93d6a190a5d79bb61b8bd58ab1f53795cfe1c15255a5a2ecb72e68733544352f2845f6958;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2985b9bc4c3f44d3c0b2518a625e3e82aed99a4c5586e3f7e805855147c5e37050dd64761619c1216;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1540543adc4f8827cf2d9d1495cfe4a20539d47164661e2e306c042c93cf90cb2102ef40c26875b55;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hced69e5267564c5270d81862d8e7693570da9b322fbb209ba038f0438c39554e3e770658cb30df232;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc0d1534e5b9b10bf81bef9451e3cdb31a07cb607281528ec12ac4c75963fb014a3693c19d5b667ce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h414abc0b836ca3d1f4f16f9e24ecba83ece51b2507fa1fa26b94f01f6fc80a922ba6a10b14ccb44b5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbeecef079e52213d4c93d0dee8ed7df6188b5729ca28ab39242cb2350fe90522c1e91cc4b3ca8ed44;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7087983eb2de06f077b696bfe6bfbf2df47f72f20b55a77f1399c4cf815d3ba4f37f9782f4f972111;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83764ba7a1870b8dcb75d4ac09e0851eb174c95f2d2aa58de67677d8e4c3f207e1cbe9bd071386869;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe0affa1eccabb20947aa9f8ec9d1bb87b7f2847029e28962de5d4f42bc9094dd9f0a864720821196;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha31f10df44ef3cf85998bc92424647f2d2586c7ad2985b377610252fbcb40add9c36622ad3c428bc9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had818ae64ab28bd044df8b21ce9746aae2e746f6b0cb67d64916765ca2aafffb056609591b3c550e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88239ece8197c71ceb59ff2a20168f514d329bcbd8007c601215f16d407da11f499458c064218afb4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfeb7acfd320d8cabacf78e6fc1777e830d138aa980821d88cce01c61ce701ed2ae036650ad1598eae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ab761a06ba8bf6451c62758c683411c04a919b89252695b7b99a56ff91752d91677f441406ff3ffe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd06531d7a66a374b75926b90df5cda4ba25e0215318807602727cea370a665032deba57f53d66d035;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fe9edfa395ce63fb77cf5569334060fa1ec25170a98ce52ada4b1f0e15d38c5897c4effb4d91fcfa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8088020930ea229b916fa094f5b9dc958aa11dc034765efc5bb2400b084969a5e9e4d8ba31e10589f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76cd1c571a15bef6d52c29d2b9927bb5aa6e97b389c4ffa9bfe3ead79af77a74c21e9d2c9a53bc02e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1411f3dba04bcfff7eb376853eb9fc911b880637f7e7339df24358899b9433cb699cd665be6eb0b4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7aeb555bc5bf39599a1594b4a074c661087fa527336253934429134ec64713487658624ffd64d2aa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc3b9a11baea4d14cd30dd720db3df5d22c098f56d506335fd354c8396e91087960fd2eb6fbe7d863;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f81c1ee4f5c0aa374c60c33532e89ccac24c6e67873ac37e73454de74e849a411da28d23f71899f5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc999864887e37ebb4e105aba5da33a3dd96726252f796598638b677131ff5686fc02675d3afc1e87;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h464255c5419cb7d18b4a012876775b3d301eced23c0eb22ff3a4bd8b51f602b2ebd5b9adcc9111a7e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34caf8b9b8f6ea60890447ee07c290e8f49f8b67ddc41993f9ede8a2131088b6dceab462340e8e294;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7533e69e8283b58fefd5b77d5658589faafa969a057576b7a9bc6a8d17857ada0b02710b2d89b24be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80d5dadd6ab07f8a13ab982118494b77dc39583f27c24fb28c3741be19dab7a016633821dde4894aa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55e0a8ae3689955c9d47a253b65f025700837c6f151e0cf2130ff10695d2e91ed0c780ff59df67ab8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h250294d1619683c2ba254f8b346d01a1f8a527af6013510bab5fe264a0ac3d1feea374688398b20b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59d5ec04cd17073a2f155e38c9845a91accfd1fe62f9a094824acc0bcd7e2c8698b742feaf9de83d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca865b37062436098c9c0af3be15de049e41405b6065b22e558a9e84b9a9fc18cb64ddc06bfa9dc8b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3734dfbad305b25b3aac62a4934231b66d70449fe600c06740a974f0387aef0efd5533f925095349;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc01c8c5f6a21c09409fbc731c82b05c6dfdb7982a75c1469385337190da276a7a42ae67777cacad9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2112495c749a93e06a5ab87ee34d92b0094929a2df5aa26460766f6921dc643a3f6781bd9dee8e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h880c420078a892431739c280e58e301beb2da60eb04383b7833d7acab6f26afe7022e373fb2a78e25;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha306fa20f38e2c753326815a0cfeffab02db58474d9f61532683534216066e067ac5da1790a433214;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67ebcb78e7e54baea4723acb0f07846e9dc5d521c67e6b4a266cf694dd40651b09f76b96b907165d9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16cb9fecde78464f68bb474d3e9ed7053ae6f3ec899339957a1e415173898bc039a32406f6100b364;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e8a3c8247a5fcec0d37c9a69b38180dd0015012034110f1a41a49f27b9267adeb0e9df2ac70e7e53;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf7babe6e5f4b7c6a16f0644117d38f1f200c49ba32d2a7a43504a7a2a53a56499e0bfd6806ba67cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h912775442d15af4458e5704f93d30f31a59d2ccce34c8ab5fc11b2deb943c5929aaf44f0acbb6a33e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8bb38ec30c4d92c22a5c42fc145e3fa0ee73aa152a063e63092c680e2e8d378e76743bcbf5edfa28;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h291c818aa9d1f1e49d3f4a8a6912e8809719404f474198a2021cb4841700c25ed624b2bda138a28f5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha56b440cd2e673ac15eb0baae42067611f625679f147a9d4126dc63b6fae0590024faa5a35b9b93cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7d49094a63f099be6adef297bf5775ab2fd46e490228fa6c1b6fdfdebb8598c2d8a8d5886a1854c7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h157642c618cb6711cfe200f4b2b7f701cee79ce2c226d9e3260ceef1c3c8c8ddeb6f1bf2fdefe9248;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c1dbe975b95d7e21310577889c8454fe203a793ad6c63066a70a48af4b113bd763134ff9afd40667;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f4b163c7ca9bba5af7756b9498038afe74bb4204aae5cc188d9b7c6c9cf4ebd14da305023db3fb80;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f343b4e9f22081d56031805198fcfa51eab26dc07c45b3ffba58b8411e89060bfff33944b88e6941;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd162b5edad764bf294e30e8f63807554e3243b13c60b8dbf8336ff7775692e22a1e0fddcfbfd7a80;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc90e5a0f66a2d2f6eb23f2e5b91978b6458a83d6b8a721839927dbfa5c2609af66f2f186e40fb19cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf631b67331f2a7d22cd25917ce48f5319470eef177aef83135f96ea5aef9bbb6599486f7ae848a0de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f9a43b060a8a749048787b5de6dcbeb6ea08bba94b83ca12abde9992c4c15ee8a496f02638385b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7aaf61009b99979e1c292f9fae4f5ef9f1edfd632fcb7b805f52e1227131191e9dfc2bc15d85629e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8cf382be663b90a60a46a11e3436af8a50291092091f52c6f5e4e3b0a5e28420a6f996aac5981b90;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b6bd3c2993f21da9da123d66272bee4dd02556252da677a459b1f4ff1901e7ab38486589351a7e5c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heef0d1fe1b5886fd3103ad293b7c4fea5b3dc170dc7dce9946e2da199a7e1047918a616eebf04b637;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h25d45d16226ac97e8355003f016e50ec74bb568c0e14329965e5f3f761be0b9a522b37b941f03225a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d211fc21af27d6c99e52e0e75b2dd32b8a5d5c2d38e9831b57456cad521fd68ef04cfad7033f68da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2982a1341297e73b47c9cfa09433a7abcf0c9bc26f75b9535d196a53e6093101752c5e1d0d045d4d8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h776f0a2f9a73d3b994044866006ab604f39f02c3ffae50114fe4591c9a1955f476548224ff13a14d5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3d9d747fe2dcecc4580d3036c61639b7cf44b6fdcf30dad305219b81d082fb6dee1cbf0ccd19c82b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc706bd54cb4cd9381f4f51374a24d08aa9955cfd56130fcf2836484a9f2d4206c8da17ddfb4ebd578;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73ec2d73de48d915bb118ae3d094edf9cbc3ce31e30fff3dba604a0f037f8936a1a6efc1231e23f5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h915f81741e4b76cdb6a3ad27d1fbe04baa9f181dcd38a198f18a8a3153cec2387d8709d0c38430af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae3d334baf1d88ce0781d510190b02cd87f8737073d5040dcd93d9c96eb6fcd4a289e4448c8800d32;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1d1b9f171dbbbbe5a26a9704d5ddaf1954bf595e1725f2e4adc7b2e5c37431f619a6cf320f91d073;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb4b60fe9382917d27b9e3f084c59d846b7c95d8f2067744dea81c461402f9c3cda072c23f279b914;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff2859a61689435cc0a006a5e21fe296a5c6e75e459602d0bc3cece8e4f1659d772260499cc98cbed;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc85d3606b3fc2faac84186762a486adae7cf81c77d69ea37e6f722de6544b08ce2113f1759c8f275;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h767f6d5a06db74a960801a2406fc7449e74e6e2c0470868ded7f61d51b245cc0b22b8e89e37566ad0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h112d3203574d220b5fc5f8be8e5a00994c72978c18be9ca7008f95f3aca657cbde75350085d738798;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h318bc1d36af15a584917ddb3d39c921a67f6d76defa0d726a23b98e90252d10f4e7a4fa19af5e9087;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he895fe85762a33f517a12fa532a9e665fda7907b119edd26e0659e372ebe62652c8847ef3bc221301;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h797974a499960c7b29cad9f0094ca46c0f2e4e6093b02fdb56ebae6d9843683201909b19915ed1853;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9c349c2beea0bd554313f7ef43de8b1c3f973dd52095c08f5cc3b1a9e98c1e19546cdbbbf685e971;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3956a52f53112636c751f1ba47dfb858a4ef7259d14589538d19894783060410ce74b87ef406588fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84003177325298a41b00db06231782bc9dca043394cedc34ff47d31e70b96d0d539540527b0f6d47d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ed70b6087c7deed35cf6bab3055af28f9b9e688940f514313f328b3267215e52ad116f22a6a17d1d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67153753cd1ccc36e74eb09ab321cf88fdf9dafef14071e7ccee7c98b4e50f8df51a4af515610814f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde5b5df7c83093813f82ad3c3ac0088ae7dddc48d9fb5afeef1a8760b8c0751166e838ceab42bec48;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5bffd9c0b41ef7548a83a88bf010fa2782633813762b9ca8aea4e22798e4a4c6752aec57a0163ae0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h192a504026c7a1c9488ae0b0a6f4508b422728914f3e59fa01efd96d3b181ea573962d369a916e714;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1bc73052f0a0696a0c895073928ab1a3a93abf66a180a77025e292d546c79a479b817fc1ecc4e11fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c22563c177b6085288700f36e86b4f39cade00f94311b0898986a18f18641e2acd695f9aca73dd69;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd314e7ed583368544d86656bcc81422c47e8b8b31de2d81f6ef2272c83c7992c9315100d7a24aa70;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdac8ef3eaa819e5dddfb0ed0bdad4e408c165f637b4eab43fcd818523ea950604a88837f332dd5a72;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64016c76e62407bb7e8612b0cfe6cc906fc15b59d552d3305bc0c0eeedaa2425954c33cbeebc6bc53;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e7fa92e0512bbeae3c152ddf6a3a7d375f8280b6255973e778e6b2ef7bd61949d24931f3b1972e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hadf7cf3095c1a5ef1645965a04a6a2423a78bbce33596c068b3f581c4b14e598835ff3315e59163dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8db4422b66b8f429aa5285245767067089b440d675923c3ba2989fd10ac2ad14df3b49623111ac57d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1ce2955197bd4233ba64302e8a7a5c04ffc22ce328393650716a0930fd61ccf4a0f2de407cb8fbaf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8a8a2f98a1aa4497f91e1a08997475689303b6d378ac01e6b508ebd6119c375124816718a11263f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d9b46ceeb5ae2ec76cc85a338c2dd5024a3d6c9bdcb1cbef9b7cded97b2264b70c5c5a15b56926ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf379dd89674d0d1abb2c88cbd34819947436b48b5dc0d460aa5c82ec9ee083109d4095aaa5230fce3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h968d868c440ed620cfde25ecd446cfdac8d2cb329e2e661f7460de518c0fbe774248fbb375a54ce37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73c5b85d7f1dc65ed0e823cc84c164008eb0ffe2c850749353cb2114c7d04531823e69744130c3603;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h933b075be87a499ace531fb068892fa785e9ed01385cd17702df1c24d8ffb6b169b9b8808bbeebd71;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23f10779261859b43e3c7a4a8ef9097b559b7549cc4358cc76071a48aead50f32aa669c24d29a556c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ef33c993b0d21f5cb5aa657cef2e804a69887718c417215ad9ae367a1eafc9752528b452cf645743;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h940fb458ba1dce7568f2e4e5eb31a8e9f7da5f97d828a35461e6217025f80331f680b853e880c539f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7eaa0efb85a5eb6eb09c7c9bed62fba7ebdd4ab208e56284c69ecafaf34acb65b1bdeecf2890a0f32;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bcb48c03888c2903e53699b138d156715ebcede65dac349a93c266c3626834a0b6ea9e71fc3b3215;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54d49eb45c226edd2581a7c041e7cb59d46fc57506a5e3a77c75a880398c976feab8255e270b19a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4aaec03c5506c687dbf9ba401c2544a32eb780bd3267f4085d4ed6011272155df54f2984274d0c4a2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedede5bf74dd258b26c251c33c4882fd44482fcff6181edc70b770284c50d2ee35987edbf411cf070;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8bf10df33ac8b91590e721a8118ca1a3aa2cafa128450186583967465c7360439339158756d500a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28b1f71857d4815e5a58c10175418b96e3ebc1926a5771d9f980b8d93dc2b79279b2cc845030324b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hadb961d5ff04a06bae2090192cf57a377a81b67a4b85472a915fd5644a694b0ee6d8ae3810c677a4d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd94c017eebaf3bb94a21443c94b822fd6c39e35d16a413ec2adca8e5eee2f018de0f8d6e044ee3947;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd1249efb63a5c6cc0bd38a71f744727c371af942984ef80a75dced3d4b7664aed685405997dbed15;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55a283f32c5c540cff76dc97d0921a723744bce326d5f56b1a704188f108b2d5f7c81e2bc842e5d79;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he37472c76bd54f787b88bb9a7c43eed02d4052aca3b457e8fe82ff14b1a6ea02734df0a2a69d3d02d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a4331674eb8d1a9b3638b9682bfd8db9cfc26ecb27421bd3515f0f882b7cf1fbcae4755e0a42b632;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h620df18c37c73f68571261ccb161b3f90e627e5e3a34ffd74b455c52717e91c8f9d85a886edcddebb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2bcce18f08fbdbd37149f65124bc2353160e63beca153859b3e344e9a6f2b07ea1441a285a60d5b09;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2ade6228f31057c732969ed0c09e56f1abfe86d8aa2fd2671d85af7ff0dd26d5bb0c7487cd9ebc27;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffd0ae884e96cd7ed1bd37cf779aa3292233dd29cc5d6a5b8a7256c44f88cc16ec2c49f9e649b7f0d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h343916a046f92c4ba0ffb6fb824bde4eb41cd906f1dcc82325178e5fbc049dd95d9d8a2f8e5ad5c9c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4917adec3b886d4c53ef963a2b0860cec0913fb96e87ec3fbc6d933d5614e9513e2af6f0d4061e455;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h730ad6643b356e2f611f5c7f8e00ffdeab586b73c3bbdb70bd30979d04a7e0369a3a7cef41beba433;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40b3e82364a093ce9e27bb3876542527ce54c9eef7108a5cecd6da2b0d9659fcc4c48a760c1423cc4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16449d19f3e7b0adb491f088164510c055b4557a8790648d19618e26782b5b3037fc74b8c514b94f7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he33751be278ac129b19ff769b606eab00fe3d08ece5161cb9ea69e653b9f69870eec1a94354bdb948;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81c4c6258321f5f5de763253fca270f959497c9332fd96b7e67e4365e22ed50c507486080720f6741;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb216f3c0d56e38e5a4a6c917cb178aa3fb606e5a6101afbbc165e7a85a296179d50edab9b232c9cdc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b4867db14f3e9b97726b77c56f65e2a0d3c20f6634b8beb74579251c063328fdf329dd08d6a26088;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had818913995a7abca45d6a75178cd54a79755c0c0a73f1ee0ca6cee5b9f0cbb1e02da2cef44b5235b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc3505f4323781c661e07aa90208eb1a5d28fe3fc448fdd7801aa2d9101bdd52ed7dd199f6f0cec40;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76ee6aa4ddf2cd423867e8069267d12d28496535a6d854d9bc96449eb8dfbaebc0ffad4c72247fccd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9a1757df002ac78066c8701f365a84209e5e44a7d1b0784a8e7bdb650ff1acac1bb3ff38267342de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18e5c88ad17791734d195b12e682bcd270278812c141e27f1118e57df190027c253e82c450befb466;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ee88d8b88d6a2d40d8fc045f1e8e56014ee0f53ceb12ce43c892e1be9811ee9038e9f8335d27064c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21e74d81f318ed68479695e388e714030674877b034ace1863d62727d461d424d8bdadbc45484e6ca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb689c06333fff1c340b573bf9e8e5d985dd58d2cc92965d22567a8051fcb35ebfc227910f6d402910;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h914b20be468c630612ada85404db0fe901c2b050703c1c71bd3380582342c953da9cdf2b884285780;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3dfd89724f812692ed84b52be03f36555fefa85081d94a52a656ad02c5b16ce8c0f3b29191270ba10;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea6cb42bfcbaa91f551e5b9cf6d5f45ba643494cb4d3f179c82daae1428120c7e5d00d55481a15ed8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h713cb222c0a1e9d1ae970f2f16112c5e5edfecc7b2ce950f6c459a108377cb3eb89d9a2ca35260f8e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he061faa983d27c5ef6fd4e853cec968454d08f4f26cd8ed15044d2a5d723324b3f2a05bf311191670;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9bc414f47c79a64c65f2959ad72794d1f443754c571aa15628d5acafd19f8b2c08b8ba895091c909c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76977d052fd0be77aaac5e15edbfb559f4124bd6e1fd73d1d1d03cb331db4578a3140d6fbac472403;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ca9e01d570d80c6fa67e189d0ca51c68c0d62435fd81e707dd4c3a8d020cc7762c40658598e58c60;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc37e306f222dad7bfa1d88a8a887c8d7dd6ecdbb6f14cb3f51508e413d144845f90dbe0cea2380155;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe7ccef63eb92f0a57ce3c2431ab433d891b0f20c477b6a5b815de6e53342a3b468756558cda485cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd07406d252b934f1ce8e6d74c45e16309f063da46797dbb15256a66763197246a2844e5eda86634b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h270294bf10740249c20277092fff6c03735d64f517c5b64ba8347acc91582987180fe2cb8280161e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf661f095df129e944a6b09c7ad6e2b40401cb8c995f9d1f712d83ef4286dd6c35cf059d8fc5a4173c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6c81f39f2a6fd8c50123e5c370485c7d202ac01afcc36b147c57be55d7d148c25c93ef1a1546a1da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h121597004c32254a299a661b32af6a9130773027c5e6f0e0a2bfa1720b4525db8b5b175fec227e4c9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6dbf61c5c32fbd6e5c262d079f513b928f19afd4011a401884c4a4d2926ecd9ac528dfedb3306d529;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfce76f7ccb8fcaba86df9ff566cd61bf4880caf1f8c81b83de0942620e4fdca270fb7c0ed9d822844;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19542756471199a42cbb393715b278302a201032bc3be532304870b815e1efcc578643b879faffea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ff115b39c12bd38b75c97118fdbfd6d75a2a2b0c4d1cc3de793e446f0c6a636c71375de780a27cb3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62abff62708aa64cef053acaf0a99d7d0fcde8617d4871e5596a14a1ef53897425a1e5ada037f3a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84073f5eb5a79c2d574036e70466a2f28c904a645d57109e7e27eec438f1c9f4c11e4fa55583560a7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb91571828b44c643fd0a4d5361692c4efcd17e69c1c14682c29ea26813c67355cc9117444dc55a8b3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd42fdfd80a555691aed9c34c707fd8bdbcd5176cc27352b6a03c799527e0a7ec9ca36adab44551265;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82e1eb129420e044e189813f86f0046d059b06198da5447d292df40aca4e954ecd5960535b8b74c20;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1fe89b2aeebec8eedf8e93f80141450dd12f03353a0c49e2ef44f7958c7a97ffdf46e3efafeb16793;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51af6ba0c98a17c20b54cd16ee34b1dfcbae0f2025f3ee8e6ca57190f88e571b82b81edf5f15b9e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26ccafb88e658380da345e3d95779dd0476933f5eaf02d5efd57c0cae76c715805194ae438892731f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7cd21260e56f555394fcd70e20f69c3f6ab35b8bf8955b8c49a67e745f2d45452e1c0fde2d886c7a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha03b2fa65ba3eacee1e0fcbb5d4d3418858fc303d82be50956df74549d28bcf4ca54a1bdf781db4e6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf748a99947780e6eb1d6b0c51aafc8fa9c0cbcf62f9f96954c90133b246d41e539b32f551a55b36c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafda16f90c6c4cb0264b8d957c1286d0eef2b0313249a9ac3be1b2076f28b7f94a3a229038878f90a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46f9ad4ed51828fbd6bce054406f0fe93cd3acfffb1f15966c3a5837e4a805174c3b84a25d7fb6764;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15783e5c6506cb559db13b8b5df0c37da16d91cfb87a1fafe9d5dfd2026e82b3dbd3c7fe50e4b65d0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hecbf5f024e387e57ca55ce40c6868b62d60420f29a896bd4fb9040263212cf97f8fc38b2cdea8c947;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h874fede7d8cf746bc6ce46bd36cbd27d795ba6d67a4b447b66f187602e04862fb4832a6ec06ae4cae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23f11b13ce4a51e8de2b03fd436f806909d6804fcd44fc2d8f3bd6a556c1300dc350dbb582a584ed7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h946b7a93828ded52991a549ca6bd894d4c1e7d1d49e8c5dacc61f32a724ead08e48c30f8d464efff0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4331d76f79ece0a2c804d7d1c3fe5376a71fa3c4ddd8bb281ec84caad9d5260fbf05f688f9d21e3ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf139c71052da41fd290d110300c3d8cdec6c327df806faebc12ce315220d0afb8c789d29c1a4a40ab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd44f1eaacbf9f3550b7d4773233a884a4aaea030526e615359fbc98e64a55b88a4a418798b6de068;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e6903759a34d154dbc79e0fe135d6d31e0b204cef539084b2d7e15cba505df47f9054c6426065c7b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8988aad3fa608243eb528d8777c27279af86b566fc0ede7e98e476330088a70a71f380d9760ec8d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha012b66cc022d2b31334cf18f26026d408afbacf1eda5c14bf3699e9dbcb3578bf6c1346e9b05857d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h587cfc812e4323cd1b1a0a1c172b6703bb0d6d280aec07ba55e4cdd166030d5309eb51b17eca7b14d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ded8def8cc0e07def103add1f65b2c6c6439edd9b558acdf8b73ac038103779cf019c610020c2852;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28d2874b045e26fbd42de487813d83cbf0ec7a93e4d0f8dd3364015beb84e7fbacbc4b978b09f699a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcba01ec09042b5d5a8c0e572dc4ed35d5e73070f2db2e09b3e360c6ecbd1f20c506064d9617e1c3be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb03ab7842749aef9e6106bbce8f34cebefbbd80d1c9e366ed1b1fb505753f9a902c22d184f2db03f3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8f5b1bd6febce0b02463f6b3d97852832cc4c9d60c8206db59309e577f8c7751a644833e3a5ae604;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92effa1c33114cbaaea41e8ae73ef23bcf483c0b820bd3d1d55a9b3cef955f372ad33e1b566622e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3df5c7753bb4d5c3b76a8ba96096e28ebe60f4826cd857fa9fc45cad930fcf5f69ea1617479e21da4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2bba64654938c608ff5d1393635d5c9dc3d24bae6976f738ba59db5e8e593761264d875442542759;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff9463cd44ae340dd99bf34baae1f8ad40b9b47461fa33daa025cd54b1c31456371165a4ba7ca7b60;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5411680a251569efcb44ff90438a42b466a4c60b9dee3110035d768b3ab5cfcf010d8ab67bf5253b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf3bf1a2b1ce7a0100b74c261f5334b562073c4dec0ba23e0c4f0cb35a76af40194129666c311c395;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7736739bab9d0ca0741cb4daf1e5c0655ba44114ebce13001fe4bcb9ae53e6abcaad25cb189d17563;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f209cb33abd654785bdcc4bb67248f074154d097ee4af1b9a3b469f686a8be359d22986e10819baa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h875addcae059cd14211d9b8611de575f532c16823b07247cc1bc77bdcb3d8a4332ba62286bcf7ccbc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a055d2db721c47d1fbc990a31f299a8d8a8b31dcbdd5b671579e8227e2d88248a7c7dbbfbf8d0038;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe8bd483abb06300a535e3f9916b71851ea021ef51c4d64ef9196226ec651d9432b9fcc6dc68133e2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a3a2a75e60e5cdd58bba25499bc8ee01055f0085302fd1a45ff9ea59dbd34270362ca73d677d0413;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc601bf8a3cb40cb30c0f51f352089e88ef2231c73af5e058ea582592d10a90f2840b2c15ebfa0825f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h301c9f89e487cc4ede15727133de6355cfd8805030758c5afd64225bd9c9fdeffea998ef0883b29b6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf488bd783c983c78d3e63a93f3788d524b446df57aee41198f39b9923ee1d8825628edc9dc476b555;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7bcbee7b23b3443e4243c10666f7d101d8875d01600c1c4c17e6cbabea5ecde43e6f9b176c5e99d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haea739107d94ff0b8eb2a9be1a59b6427fe334a1fe792287c66dab7a8c0c5f549ca59968668be48bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e5906a64b4ad4e535760a74b1f7fba6cf0aa1520fd813586cbdb71a637f6d269667c13ae9017fc85;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76b81b0ff80b77cac96fd60c8afc0608cde20ea6b4bfcc386d2d5b8afa9a4cfe339cc1f51c0173c46;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6473be7f94863be7216e7fb14bb4c2a33ef9c9a10a2cc9635d9715043163418d188941ae18896777;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde42c99ae883689fedd3d73c9f24052490b912515a63f9098cb2f8f6e9e2352da79d5fbc020e8457d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef73629aa959243c5b9243984e42d04aaceebd160d40f6b356a7540b1936ee27c9f4dd84334d06b5e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9cea189ab7b179a953656e148da2b02246e255012341614a6934d664ec2fdc00fbed14aa2a438f5dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h954344b18430a5d1ce3553f56908acbf1e59c6f9ac52ae7f2b927dc15596222350c71d5783486a862;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf03639771d1ef84d1a356c382c3912753c031350663e616f267bb1343953592d52bd85e4867db310d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4609623a7d3fbcef9831544db9e7cd9564b28a5c9dddb82f9bcd2d50c4bc90d677d9657ebb03b0899;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1e3041343051db2512face8b4201f30dd6e5ca0939193a90072568872ccba54a765e4687eae43d15;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34ef606ee326965302e3efdd9c01014907d6cc935f599fbd58c4da97e28e3e0489bef86bca6f6f19;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c1d132bf280818ebb90905eb3b73249626f75f12bcfb868d7473c8b0bf841158af2194becab7741a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62c6c6cfc32493cecaacd141b89847f2fb602b41bcda2c997d3c473f669cd3d8ed0a3bace80824b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90f6f14b8f739fff1201a1a0fa1c806cebf8953456f759c3fa225b371e0e92c33412a921db4612e76;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10da3bc5a8dfdae9f9fcb8796d2ab0d30276e34d19202e4631b6dc33ddb3b1ba9ada51520ac341547;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d0541e6fdb0bb03ff79428c335c2c3d66bccb8a8ddf8f5ac9610753969e9467ba6b467d81923c4e6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6c7b7bd29be6ccc8b138e10f491ad84d4f8438e14cb0296e1558cda9a4f687345ab1e2a927549ec7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ed5b7c5085f1844e60b2bb9931ba38a76f67fb7266b75faa4278e62125f60cc1ea4d389deaf77d15;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h655d9eed40d568a45ebc6a59caf9c5f8c30973816ba0cb187f74440ef8f24a63f472627a349af6fde;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3234f79ed2fbb93a410f6acd43599dab90325cbfbead4cca0c82a185f05a18cd75edc6b73353f1e89;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92ee46fcc145e072c2ba7b5f49513c4940b28f3ea7e01f6b789b2453655555976af0f8492f041905a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4e6b56a70cfd5f64e9456bb935bc4d46141eb66e0778872c1005012aaba098e4db7c03b0edf3066e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdf2bae32023ea73e3f7aaf3b36f8d568a42c8e497cb5f0226ff98961f6e220ae5503bf5fefd894e93;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34237ef45796e53edc37eb6726d80d9397050461636fbffcfa1e744d7ab74d09d85ec25a1210d9288;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1ceb256658d481e623ce9d5a4907ffbf3d415c98b189a15a59e0c3f6806eb4c0fbe734d52235f681;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f7d19ee574526dbe62ba2462d41dfc1565dbb67b308fd63a55a36b2f6a5cc2165eb00fd6de8aa93d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd279ef69ef0155d7754b2af6126b6609b4bd5eddd6ecd80bad4531335c7618696b250e527b2f8cefa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1399b80a6ad046820ea2923aafc9f3bb2c9bfd26d58f4a016c6514a0e586347148ec49fef60ca460e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdea9898ac506fd19931e9221aae1f68d56386c2aefb03986932a1e7344e3abdf69d3c2ab246c8fa53;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2366b9d1262df767e72afde2a5f0d5badc5f30c1b5e14c9ceb8cfc7a4fa05fc7d7ec42129c3e96086;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3528885d82fe219ec68dfd00d0bc015a94141860acb067668db77778d0e9eb2a355f7e7067000e9f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70d00663ff305a8a4e666fb3c1b49be5c17c9b04ad4f4877389d8e6890fc765be0007a431cb58c9e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11931513bb893f76e7abb565c6b5dbf3f0eed336e3bac44bda8de7c20708cbf422f88db36d54c9971;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c1c80975251bbb7422760ab2f2c466164214c0630cf8ae734332f75576e66719a87025b872abb6e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f565e16b08af7a07e9e5fd5558e62a40dc3bec2da4f39611f389a845d5bed7ddba76fcac385f8839;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h845aa6cae8970ee283600784f57e7d0432022171a57ce3ee740013240528b57da739538fa7fa7e3b8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66eb25729261b137e7a8cb985c012f98cad2fa973ee94535d8f652e1b38920836fca62e09177ed098;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hceaa0a9863a35cd493e40e3f7b69657dbe06e29f086a29983a32a92eceb1d366031c0df8af7ac401d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1fdfedf5e4d991ae284361aab33fb0fdb9d48e01af4cab647555cd27eee9c6c16da9a5fbac5f40f11;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55aca6b710fbba901ab58a20ac47ec3585553caf07529a2ddf34bf3c9570d0dd5d7cdadbd9283df48;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f4cf1c2a5f50684c98c6ef0f92dbe4055a36109bdd3b8548bb47ed586530ab8ca7a4a6ac61a57326;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2bee3111a154404512e4aa04e15c2416137debb757d98bd8c669f74913f7f80d87e4ebd90cdac5d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd62caf88ab27f8ef9d1ca1ef2e9340a4122395245bae5288ada8c5592e0ae644e5ce422e1cadfa2b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b01fcb6023f75b5de45b79af7e0afc3c41db106e7de699e1b489373269d87edb1b38ba4855254bf7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7438999ded5cf3e27e49718f6472301655bd38df3e0a9ef5d10a9b9bf5ce0bb015a5e3b3a197db21a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb25cef34e017b32d445ab8d9042207b7bdea01487a77ed60383bdfe314cea53f9bdb4c4d0972def34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0b754a7fa84e5d293fd5008edd1e6a58adbc7a01d20c9a2c8152e55496aee2ad5e9ed3b5cc47be35;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h221a346ac2d5b2e98f2c66c06a0559a6aa0549074dad10897c5c025bf40a30f4a77434dffd3754178;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hece76a189dc84b6d96974f24310a66543eb78c322417d260f9fdf11fc3e4c4e354cab0d8351727e14;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3cc2e3105ff505682181fbf4e4eebd4c15acfb263f46b260d39ab438881bfaad08d47edb5eb2b796;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b580ea3f8d71140d0b41a5637887e2bf5e32f58a6b1d8766c54560b5380d7b8617b83667a46e9569;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b89ffa10b3d8b50dbe85aef0c18b0f60f47fd3d82cff3b0390443ddb669a04080816f0ae94dbe8c9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf867988a553feebecc5ff96d227f78a6a7ac3c16d4a1284b137949447bac1385c7caf2c2989086eff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17818260f23ddd79e2dc550f05ba49fc9e2bb75c483a3ce7dc8e0fc7c7e03a3795775b54eea217a22;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe9d616b6e23d16c61030513594cda4e729a34418a356f6b9768e6772179b68d68aaf6b0f5db4d99a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7974c10df501fc97e09747a13c7b13d86531ca10eda39f67b54de0dc3c0ec9db933ad3fb7b039e35;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he29e7c56f51a528994a188b7b794dd365b9a8406dea303206c3fa51f331b26385b4e2fb2bf668f41b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc207e7e87f4aa07f2085a55c27ae260285cd35cefd940c22d2f0bfee84b959d4e162db8d22377bfb6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35644a27afb3dff8ff17086e1e1fe029f4dc5c6d07b09cb2ed24abdb8d85450f7a077d6aca54b0f2f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5431c702794aae24a0a90807df6703c92cd21563c0f990ea745f5e8baff4cd9b350571d68b17f69da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6989dab392de6f1b467c84674f47a50da8ba1867c1b1289481b89c5dc405e76920a35d10462b88934;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d08b2fd5143cc77c6e43539a4322a574644801e62b866495227e3c2568212322436dff4479940f59;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h25702c3492f09773ca10d6c5f412d00e9012929df83243b9c97a0d9fa4fa795d6203dc6f805862ce7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5bae72638c30a2c37925683b291b5977fa1b8df5f6dca4586494d7f9788aa8b003d43f0936afdda7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9aa698919a2196d460ad209b1de385ed9bbe1d00305a03419d9036e9bcd689a3893d2a2dee218717d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7efbb1a26a9f0ab43277acf1b68aa79423892027142d63c05c6787cd2b8c5df6fc105ef1322c2364;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3663792fb4f0208baf28cbce5b0e30bd48976ff4637c1205d53f0d4f1e415751810b271d444de7e2b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14b0a1b8301b015a4f858acf5b98c98c1d563a4ca28c0c92bda6376fc97dd2d2e5700c722eaf251af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h399e26638b42305b818e51802da81526102c8eac93aac984066ee24e4608ae464f7ad7e068bdc4650;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb238246a88dad910609529d7f012ed088650cc02fc6b3467a3e0be487894f471c04c4944acbe215df;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46c12a1a622d2dc6edcb4f75c588f88a678243b304f59a312df680bdf00516463dc0a8bd23af1cdb0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4940ae2763766017a20f6f1c0054482aa4cd72887ac636b07222b07ad07449bf6b5e5cf4f8abbdc0d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb731006edb38f077e7afb1f1dcf49de87e82f9bc24f922ccc8f41988a1ab91a37e87dffa966d853;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4117b62c473317c4c399a2a5b185c872224d584a87dc966b607ba4c960cce5de3decefde221a4043;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38e7a0be45877128d2f5d89f2ee568f2aa9ad57f0ee7e55aae3e3c07c140ba7bd56dddb51f5cb4787;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84ed0b48b451f5a5a479a1bfe640092ce758d00152119b36e1ea6347e6bc170d580dde86ed3c026e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24b853570b440d442f24300c3c2e7a74e329485309bf03d3b2a6679aa8881d4ba307139ecb6f1b4f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1cf82a39fcecf46108d41e24ab3003a940cbe60059beb2e54773f45733eba627f56cf3c9a9077f13;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f345f0e6adea54f32efc61f6214b89cd5b949fe59aeb489737fdf597d301f421e2feea2b26074654;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h756e82ae6efefeeb78209fbd3f95109d11da0864fc9b80b15e59909dff66049060e429abc3345a51;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h293fc305807bb2124ea855ebfb21f5313fdf60c47c1dae8791735bd49db5baa12f68aa2d3749a2939;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0a7e266ea2f0b4a13a9184afd55d8d99174bc19678c762ef4f733ad15aaf260fb51b5fb6fc6452a0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h25d9f0f6231f0f4295a028e8b8c2c69fed60e9ad76fe424b2bb0bffbd382d34a0305f90ad64e7afb6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ccd04cfcf2431fa68716b43add61309f0e5df8bf4450bb612b9f86e2e082b6c5c4c190a2ea54698c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h594ff3d7d0c48823d79e5400c61ed8418d59ba8a7d3ee87d859795adf9cd4a98cade8c70d826bb188;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd08355f4ce7808df16f8b9d16bc9c656c0bde54bc9ef64a69782d3ac0871a80ce7e3854641b5b7c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c425457abe2ee7bc48406903ce7f05d5ff2d4e8887b9da53f12d664d2cd270c31ce06d970903ffd7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habc966e6532178eef8f69c91c81e9bd85f24532de4b57f39ea6d579b5e6ac9093a8e7dcb6c3b913b8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6c7ca12091bfe1a64ceede192f288c93cce2822548207d5b62d51ee37f5e43d74c1ca815a96db051;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf72e2512e1266638fd5989930a8c1f838c40b9e8caf9b32afc5a160d994d62cea79effad739fda5bf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67105f38bd38ed6ee3dac0570e99ef56a9d7fd3aeb91d48ec38b32897f2ec565b12fe0c6ed51ef23a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e746cb92890645bb99a6bdb4c1c85e3c5ab8e64b320a85d31b78aec860c729ca14460ca584530f11;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6870726866cbfe9e42670a6fdcfd25b2815097249e817ee2683b17d5770bb44f521d320cfbc5c8354;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ca5bea9084d4a543c096d4166caee21ff42efba2cbbf6ba5df884f839422c74e458672304dbc68c5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93f8ed253674e51f3ad5d3ea4831a263e6a5460e40610309aeb0534f9a62ff2076bad64395b4b8e7e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e9b64d17f61a1f4aa0b58cb1225f873500b0b2f84b560e9b50589cb32ac27585dee151f1b8d75fd1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h377ba04268cbdbf399e5942f1b2786754c8b57d41c013ad8f3a4881db4ad2709949277219fb0ab85e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce76754c912706f276aa7b5ad7c3c5e45bf3f2d402ab0bc64b4b951316c34663fff639d174539ef3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9855bf8aa8217f704007d141d0782865a84058780e389520cddcb2d57afbb93fbce7c3052e370c2d3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53b3bdd35358fdc192fbbe42ba50a5876bb6a5f47ebb6001ddfba6e606d04904a0a8fc11b10df298a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30b2da3eb19cce06844db3b37e8bcb70283a7ef0759128d60850f65502d7b974ce67323146f959dd4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60b828ea4b6c2817b3344c33e5df9786536022548a9504a4ea11d715568e37f9cdca9ae032ab86d23;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c981b20139562e33f44b31cfecb4fa253ed2dd58b355964e9466c7e26a81a6a0e28507239869f598;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hccf6e49442a7910e8ad5d9e41cba1bdcd7e97e4e2f6abe890523058eb208ebc48f4af87e6a32b6514;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11b5f72f785079843b973a85805e9037d344b024e0c40cd9ac25038641280bd7933d0bc39bcf46ec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83b02ad6ad35359279385f53f0f00348f5028fba68e29d18441f7b8cba2f4d6855f499dc6ebccaa65;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd49abc5a0bddf1bb512aeda46eccc517b6d96692f81abdaa461e22ccfaa4e0546b98d8a40c33b087b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84c23532d6c8654a66453c4f82f1d6020ddee974b6045126864e61fdd1905e4f36c02d329d54068c9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5622a76bdf7f16129b911bcbbdd477037ad0bea0399d205ede7aedbb42f597c17e6494a86d4ab4098;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf71d202b48107d2a303f6ed78f16b05eb1956a419c5d94ac1a5b858c55d5969396dec96d8cf483cd5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43498ec602ff45cca0539677bd8b3dc987436eb8eb2420795967b8306a7da2a0ba926d91c10d8a81f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66cf7cb4d9419cffa242f3e49635323b769b5e10586d3f9efb1179e8145c68428a23605119e8fe458;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70bdae950fa9b17d325d9c3530a0fd345a9bf1564640e5da71fe791141f131333fdf09b399826e556;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73bdac8d32ffd2e68481ebf69d71970c345f772823a40be8b10833ece60ba9818a45ffae1c5db8bcf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h259bd09f9b0a859a357e3a6ec18abff607ad525209649f84e216e1131e8e7f357a6dda35fcf426652;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1403a303d5e3e5f85c66d35f91e2fc9c0179aad4847b1c1033e54bb46622b653446e4e81d06ca3e11;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8fca5d081dfb780b034848cee869038a90f984912b1b4238abfb22bcdac1c17f2662bfcf508ba752;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0ed3db62a41d2bc1ee41dab7780575cbd653564e01382acbbfaa78fd6136d7140654390c1ca603ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h361e21249424fe8036a5a3cc88e95250534e02284eb0f15b91da7e12e3163b27e1c04c7d917017edb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb457ac30651737fac8c69b07ed671ab4fbe2d7aabe00f65ae2998b945e23562808bff01f0d2c9b47;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2bbf6c58cc41c86cb9c294acddbd17be5e5064e690c7c3f23d266fcb76e59d53cd8e710d93caee441;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdefcdc95a1e5c01dd9ee118a081b35d14d60cc00008024afa70256343bc41f23a587fb79a1de5e863;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab05d6945098678c5937531d16a8e8fcb37c2c03e66bc369d20a1fcdb34cca012a678d2e588681f7a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2276694d36c7b3b2a29c2f16fe84d3b1bba4094ccafd34e5728fb801b9cf450756b49fbcb9fdd142;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd01100932e15709f325982b37f2c744bf1446051d9fba8c986c142c2631798bc35a28b98d0151ae8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h460eb6afed2efa6ecf81e25dc9f0f54bb09c20bb72aecbe5322bf18bb57c4ec74b1613c0e774f5088;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89b921ba2ed76f507d8eabf5b268116e5747b8810f80dc23448b465a43037b7dc4f0513a864d4e8a2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b175078e73e077c6625996ffa0b50cc16774ffb7dd791fe60020281df9042807fee90162dca6ae0c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e09237603aeba81a45e188be450bd3c436f3a2efa56f5f9c1d2b9b7926ba699e81b94fa22f09077a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f4cfa31bd754929943ba27c45b535651971fad9d9dec994e8cab3b43f6b03d083b53050c4e64dd27;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c671488a0dac3ce405dc3972a34e3f7030091e5665715a44a04e92b826d6de248ab6ed3f745593a0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h906564f4047da355dcc74de477c32ea147bec211886f056c4b7535581d3ae48d6caee06082ddba96;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha22a66393fbd790acdf8b6877eb68d4ffd46f6e93d858679442aaad82a4abd10bcc3c4cfffc585598;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0bb5f30deaf34cc75d759a4b1e4f874f689bb368d5d1a5e9486d4f3134c8277433dddfef38d1d981;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hede8d1849665df3bb6d5d2d5319f44237e6ceaa387c76ee36c67a9343122f7122c62a9c66e055de79;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h513831806b74fdc3b9f975a87c793b7ad1c96fe34e3e6f1da7356200adb28a8571092f58a8809be34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2644b2bede48085c35ea0472836f65026a8515a32bc518467336b5015004f8fdc282b865523d5674;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94fbe9c93e3dfab29b98279f478fe933ed3690832c9f00aca0445b9b5ee7b6dc2a9d90a142efa73b1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7216913c21722a2aafda944f1c08eaa7624d6cf9fe9cbad664a7609122db21284237de9c945bf6f6d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haad3cae77aca30282d8f2c4bbe74bade33e60f2795be9e13a59d1b070835efc12a21db3d3137fae65;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27889f75fa41a955a51ce27fb36809dfb66b8f072d721a3b03c899556a59a6cdc0026faddadb7ebc7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha630cb54ca38c21770216ba6a7ad1471dc129682d85a7d698720befa65da230f3cf7e5176d4617ba4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e7399fd27d1be9dd7d8cf3c8b0fa34a37a8ea1134e54dac54aa063f6a8c9b471ae81df28e2158d57;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a8484616130aec08b43cb702215c22dbe89dce0e3a87cb10a942b93ddfc21e32f7ba99e66c41d53e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h734a29eba814ec67d9adce1f45a66f9d3ac18e936c06740c9e2e831d56117d0a16d756763d474502c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ece0f4439de4474ab2798bd14579bf286e23828ad68d06714e60421181ca562ea64f80c15c5a6a10;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4828603a5d49f6e531d87987e21f178047e91f82dd6149fe667deb18a6a6bfed6a806433c8515a825;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7cc078d7e411ddf7dee0b660743260590010d43bf11b535754ce78e10b096d59def4f3c67bcf74220;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c486307482dd09e2e8e5233233be5e76208327e264a26aa31bf0bb9058c18b2810ead35929bf214b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76b16c7f4da252030e1fe0f2b2f03190c0c51e98a0fa6cab689d3d75c4afe2941ce23329075acd310;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h584e18106ade5c5b6f72b3a07d7eb42880e832a86141972c9185a8632db6eb3e225b23d21c5be71b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9cc139c3b038610a0cbdb77982922dfcb3ea7fd3888c56fc82cd3c9d0de2db9beb5e933314b7c057;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8590896fb489bdc11d2b68a077938d142c9538ccf845522b064707acdbfb96275de205aea5d0b4df;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3fc54ea67e4a9f995d714debc74d16334ecf0f51caccaebd8d3389056689cb3627c5eb4f07965183;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2880cca34e03048fd5e3d15ac63fceaee444ba1425b42d3ac7748a6c67aa1a7d3640e74da6747e424;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95997e5207e19148991e51c75a2f839cb3959429d5ed6b59c99e6fba3a20f74930ea9a063c2c11649;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5731d88c23e781e9da5dca40480d5e3276a5fc62e4c791245a18f387995f6fc60366c172786ead440;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ae7b5bb99e70583f519e7804b78657f6bc34e773a5f732464ada9e58063d39e8808df34411b04104;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4374a6f4775360d402128d431682b19d4478aa0ac30ec0e6e9b2ab9b4647ee63b39d425ddf8441935;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c0c5ec71ae13faa5845597bc01f9e8e9d92d7a1629a67834dd74eafd85dd8e866f219e099bd3c2f9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb69263d53b661cedcfad39309a70a34cc82846beb0685cb58106033450520f97e1fd304b3d9fe5ae7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h120fb256ae2dba22a589634a90c2508091d76a42d03daf7f6f049bc51914ec32ea923fbd73d2fa91a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79aff1921c2fde6771e2c8cf2bafc8ec38a96213ef7934cce9cd2d4c3d504c4514af2f853d8cb3192;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16c7fa2528c8c40e7aff0cc78b4fd64bb77c7f43f5b7d135a880cde3f74b1804582c931ad56e76274;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb89efc3bde3507ac066634e2223f9c22c92122221e3ca24858611b3e38944bdefe560faba5c7e49d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h827e372551081835220ec69646b86a8b2329108785e2c7ef1163bed6f9d82d68078d749214c470b17;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58cca850db3d27bab3e1cd6e9747b91bb47e3cd7e20a56964509ce3f6a1d7eed841638de6bced66d0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d93526567ba41b230582ab58f7c6fa80e61a62a3dfa591be5c01a24ad58b8344292d8074efc748ca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea65f8b836d156d28990ae69163dcf03c49fb56c76bf55c9ac0b59d3989a475cfb91d0c6aa32d9ee9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7865a7d5ef17070ab90e21a1964af55cf3fcaa57bfccdb138999c60d90ae307167db06c461e2fb76;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h279150b7ec531bc9d71ed789dbd5816cfc183b948242e2a2ba79f3d6801f6397b4f9f135941227753;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12e539858771242710b191e9fe8607121cec2dd97d9427c1d93c5bc0b91fe3c8ac98e87206c218929;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1203757e1fa551454492fcea8fc64f60d2e1ec296c6776ae36306210ec7fdcb6753e70e226b80c0d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h687a8025ab47c4dd8a093d860023e70be105ce80b847bbeca4f96f745218cb938b98eff4674225473;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h693f123092a0573a4259852d3752be90989e663b09a0739d821d65510e679b3ecefabd10108b850e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4eb153b7bb2c8c4bd5d91c630ac2c8400799cf1d7d7d4c259cc26dd7481f4c08c55329b16579a7d1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f4bc3768c9ae5ce4eabe80d7a022c03f3a2278b6d493a8def6901a3fcadcc47ff0bf5e487cf11385;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a06d229c1f16d0f8cbb155e90858878427337063f63f460999f44195630c99d4184bffb0cc37a37b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h969cceab128efce5b2ada0aa4ff2c09ea4362a541133f9f64caa9f1921e557f7ddcfd6aab7c894e78;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h751eac950db8007bc21e6b7806fa00da478c9ecd656c36e2eada3bb9b80564cc1f62e6f19bf735507;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbaeb98ac22746d26fc45289e7ff66b653111e06f0e6fb7b7064b5e0f238b7cbea2c48a8caf25c03f5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9ad56b02203cf00a7385c5c75c5ef5509e8185cb49725b6ef43eb100adf0f02d1f5394e90d33fceb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2269bee7a4fd5bb51f18d15ba4bb11a6090e265ff793681f3fd9b84bb41ea0a0249bafb29ed0efe45;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b36a8ce49f8aca2cc2887fccaa18c634199f74d795e5bb3c528580c7935db60667c2f11ccc696e8b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50929680809c359fc7a31b2f96ca303158d1a7433f0788c688ee41c889dfc767f723e312775073808;
        #1
        $finish();
    end
endmodule
