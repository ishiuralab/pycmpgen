module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69,
        output wire [0:0] dst70,
        output wire [0:0] dst71,
        output wire [0:0] dst72);
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    reg [485:0] src16;
    reg [485:0] src17;
    reg [485:0] src18;
    reg [485:0] src19;
    reg [485:0] src20;
    reg [485:0] src21;
    reg [485:0] src22;
    reg [485:0] src23;
    reg [485:0] src24;
    reg [485:0] src25;
    reg [485:0] src26;
    reg [485:0] src27;
    reg [485:0] src28;
    reg [485:0] src29;
    reg [485:0] src30;
    reg [485:0] src31;
    reg [485:0] src32;
    reg [485:0] src33;
    reg [485:0] src34;
    reg [485:0] src35;
    reg [485:0] src36;
    reg [485:0] src37;
    reg [485:0] src38;
    reg [485:0] src39;
    reg [485:0] src40;
    reg [485:0] src41;
    reg [485:0] src42;
    reg [485:0] src43;
    reg [485:0] src44;
    reg [485:0] src45;
    reg [485:0] src46;
    reg [485:0] src47;
    reg [485:0] src48;
    reg [485:0] src49;
    reg [485:0] src50;
    reg [485:0] src51;
    reg [485:0] src52;
    reg [485:0] src53;
    reg [485:0] src54;
    reg [485:0] src55;
    reg [485:0] src56;
    reg [485:0] src57;
    reg [485:0] src58;
    reg [485:0] src59;
    reg [485:0] src60;
    reg [485:0] src61;
    reg [485:0] src62;
    reg [485:0] src63;
    compressor_CLA486_64 compressor_CLA486_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69),
            .dst70(dst70),
            .dst71(dst71),
            .dst72(dst72));
    initial begin
        src0 <= 486'h0;
        src1 <= 486'h0;
        src2 <= 486'h0;
        src3 <= 486'h0;
        src4 <= 486'h0;
        src5 <= 486'h0;
        src6 <= 486'h0;
        src7 <= 486'h0;
        src8 <= 486'h0;
        src9 <= 486'h0;
        src10 <= 486'h0;
        src11 <= 486'h0;
        src12 <= 486'h0;
        src13 <= 486'h0;
        src14 <= 486'h0;
        src15 <= 486'h0;
        src16 <= 486'h0;
        src17 <= 486'h0;
        src18 <= 486'h0;
        src19 <= 486'h0;
        src20 <= 486'h0;
        src21 <= 486'h0;
        src22 <= 486'h0;
        src23 <= 486'h0;
        src24 <= 486'h0;
        src25 <= 486'h0;
        src26 <= 486'h0;
        src27 <= 486'h0;
        src28 <= 486'h0;
        src29 <= 486'h0;
        src30 <= 486'h0;
        src31 <= 486'h0;
        src32 <= 486'h0;
        src33 <= 486'h0;
        src34 <= 486'h0;
        src35 <= 486'h0;
        src36 <= 486'h0;
        src37 <= 486'h0;
        src38 <= 486'h0;
        src39 <= 486'h0;
        src40 <= 486'h0;
        src41 <= 486'h0;
        src42 <= 486'h0;
        src43 <= 486'h0;
        src44 <= 486'h0;
        src45 <= 486'h0;
        src46 <= 486'h0;
        src47 <= 486'h0;
        src48 <= 486'h0;
        src49 <= 486'h0;
        src50 <= 486'h0;
        src51 <= 486'h0;
        src52 <= 486'h0;
        src53 <= 486'h0;
        src54 <= 486'h0;
        src55 <= 486'h0;
        src56 <= 486'h0;
        src57 <= 486'h0;
        src58 <= 486'h0;
        src59 <= 486'h0;
        src60 <= 486'h0;
        src61 <= 486'h0;
        src62 <= 486'h0;
        src63 <= 486'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA486_64(
    input [485:0]src0,
    input [485:0]src1,
    input [485:0]src2,
    input [485:0]src3,
    input [485:0]src4,
    input [485:0]src5,
    input [485:0]src6,
    input [485:0]src7,
    input [485:0]src8,
    input [485:0]src9,
    input [485:0]src10,
    input [485:0]src11,
    input [485:0]src12,
    input [485:0]src13,
    input [485:0]src14,
    input [485:0]src15,
    input [485:0]src16,
    input [485:0]src17,
    input [485:0]src18,
    input [485:0]src19,
    input [485:0]src20,
    input [485:0]src21,
    input [485:0]src22,
    input [485:0]src23,
    input [485:0]src24,
    input [485:0]src25,
    input [485:0]src26,
    input [485:0]src27,
    input [485:0]src28,
    input [485:0]src29,
    input [485:0]src30,
    input [485:0]src31,
    input [485:0]src32,
    input [485:0]src33,
    input [485:0]src34,
    input [485:0]src35,
    input [485:0]src36,
    input [485:0]src37,
    input [485:0]src38,
    input [485:0]src39,
    input [485:0]src40,
    input [485:0]src41,
    input [485:0]src42,
    input [485:0]src43,
    input [485:0]src44,
    input [485:0]src45,
    input [485:0]src46,
    input [485:0]src47,
    input [485:0]src48,
    input [485:0]src49,
    input [485:0]src50,
    input [485:0]src51,
    input [485:0]src52,
    input [485:0]src53,
    input [485:0]src54,
    input [485:0]src55,
    input [485:0]src56,
    input [485:0]src57,
    input [485:0]src58,
    input [485:0]src59,
    input [485:0]src60,
    input [485:0]src61,
    input [485:0]src62,
    input [485:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69,
    output dst70,
    output dst71,
    output dst72);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [0:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [0:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [1:0] comp_out68;
    wire [1:0] comp_out69;
    wire [1:0] comp_out70;
    wire [1:0] comp_out71;
    wire [1:0] comp_out72;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69),
        .dst70(comp_out70),
        .dst71(comp_out71),
        .dst72(comp_out72)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out72[0], comp_out71[0], comp_out70[0], comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out72[1], comp_out71[1], comp_out70[1], comp_out69[1], comp_out68[1], comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], 1'h0, comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], 1'h0, comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], 1'h0}),
        .dst({dst72, dst71, dst70, dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [485:0] src0,
      input wire [485:0] src1,
      input wire [485:0] src2,
      input wire [485:0] src3,
      input wire [485:0] src4,
      input wire [485:0] src5,
      input wire [485:0] src6,
      input wire [485:0] src7,
      input wire [485:0] src8,
      input wire [485:0] src9,
      input wire [485:0] src10,
      input wire [485:0] src11,
      input wire [485:0] src12,
      input wire [485:0] src13,
      input wire [485:0] src14,
      input wire [485:0] src15,
      input wire [485:0] src16,
      input wire [485:0] src17,
      input wire [485:0] src18,
      input wire [485:0] src19,
      input wire [485:0] src20,
      input wire [485:0] src21,
      input wire [485:0] src22,
      input wire [485:0] src23,
      input wire [485:0] src24,
      input wire [485:0] src25,
      input wire [485:0] src26,
      input wire [485:0] src27,
      input wire [485:0] src28,
      input wire [485:0] src29,
      input wire [485:0] src30,
      input wire [485:0] src31,
      input wire [485:0] src32,
      input wire [485:0] src33,
      input wire [485:0] src34,
      input wire [485:0] src35,
      input wire [485:0] src36,
      input wire [485:0] src37,
      input wire [485:0] src38,
      input wire [485:0] src39,
      input wire [485:0] src40,
      input wire [485:0] src41,
      input wire [485:0] src42,
      input wire [485:0] src43,
      input wire [485:0] src44,
      input wire [485:0] src45,
      input wire [485:0] src46,
      input wire [485:0] src47,
      input wire [485:0] src48,
      input wire [485:0] src49,
      input wire [485:0] src50,
      input wire [485:0] src51,
      input wire [485:0] src52,
      input wire [485:0] src53,
      input wire [485:0] src54,
      input wire [485:0] src55,
      input wire [485:0] src56,
      input wire [485:0] src57,
      input wire [485:0] src58,
      input wire [485:0] src59,
      input wire [485:0] src60,
      input wire [485:0] src61,
      input wire [485:0] src62,
      input wire [485:0] src63,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [0:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [0:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [1:0] dst69,
      output wire [1:0] dst70,
      output wire [1:0] dst71,
      output wire [1:0] dst72);

   wire [485:0] stage0_0;
   wire [485:0] stage0_1;
   wire [485:0] stage0_2;
   wire [485:0] stage0_3;
   wire [485:0] stage0_4;
   wire [485:0] stage0_5;
   wire [485:0] stage0_6;
   wire [485:0] stage0_7;
   wire [485:0] stage0_8;
   wire [485:0] stage0_9;
   wire [485:0] stage0_10;
   wire [485:0] stage0_11;
   wire [485:0] stage0_12;
   wire [485:0] stage0_13;
   wire [485:0] stage0_14;
   wire [485:0] stage0_15;
   wire [485:0] stage0_16;
   wire [485:0] stage0_17;
   wire [485:0] stage0_18;
   wire [485:0] stage0_19;
   wire [485:0] stage0_20;
   wire [485:0] stage0_21;
   wire [485:0] stage0_22;
   wire [485:0] stage0_23;
   wire [485:0] stage0_24;
   wire [485:0] stage0_25;
   wire [485:0] stage0_26;
   wire [485:0] stage0_27;
   wire [485:0] stage0_28;
   wire [485:0] stage0_29;
   wire [485:0] stage0_30;
   wire [485:0] stage0_31;
   wire [485:0] stage0_32;
   wire [485:0] stage0_33;
   wire [485:0] stage0_34;
   wire [485:0] stage0_35;
   wire [485:0] stage0_36;
   wire [485:0] stage0_37;
   wire [485:0] stage0_38;
   wire [485:0] stage0_39;
   wire [485:0] stage0_40;
   wire [485:0] stage0_41;
   wire [485:0] stage0_42;
   wire [485:0] stage0_43;
   wire [485:0] stage0_44;
   wire [485:0] stage0_45;
   wire [485:0] stage0_46;
   wire [485:0] stage0_47;
   wire [485:0] stage0_48;
   wire [485:0] stage0_49;
   wire [485:0] stage0_50;
   wire [485:0] stage0_51;
   wire [485:0] stage0_52;
   wire [485:0] stage0_53;
   wire [485:0] stage0_54;
   wire [485:0] stage0_55;
   wire [485:0] stage0_56;
   wire [485:0] stage0_57;
   wire [485:0] stage0_58;
   wire [485:0] stage0_59;
   wire [485:0] stage0_60;
   wire [485:0] stage0_61;
   wire [485:0] stage0_62;
   wire [485:0] stage0_63;
   wire [124:0] stage1_0;
   wire [175:0] stage1_1;
   wire [157:0] stage1_2;
   wire [214:0] stage1_3;
   wire [227:0] stage1_4;
   wire [197:0] stage1_5;
   wire [213:0] stage1_6;
   wire [220:0] stage1_7;
   wire [205:0] stage1_8;
   wire [213:0] stage1_9;
   wire [284:0] stage1_10;
   wire [276:0] stage1_11;
   wire [188:0] stage1_12;
   wire [304:0] stage1_13;
   wire [218:0] stage1_14;
   wire [170:0] stage1_15;
   wire [221:0] stage1_16;
   wire [228:0] stage1_17;
   wire [208:0] stage1_18;
   wire [275:0] stage1_19;
   wire [267:0] stage1_20;
   wire [189:0] stage1_21;
   wire [170:0] stage1_22;
   wire [286:0] stage1_23;
   wire [213:0] stage1_24;
   wire [183:0] stage1_25;
   wire [250:0] stage1_26;
   wire [205:0] stage1_27;
   wire [223:0] stage1_28;
   wire [228:0] stage1_29;
   wire [191:0] stage1_30;
   wire [217:0] stage1_31;
   wire [216:0] stage1_32;
   wire [258:0] stage1_33;
   wire [189:0] stage1_34;
   wire [216:0] stage1_35;
   wire [201:0] stage1_36;
   wire [307:0] stage1_37;
   wire [264:0] stage1_38;
   wire [212:0] stage1_39;
   wire [303:0] stage1_40;
   wire [170:0] stage1_41;
   wire [173:0] stage1_42;
   wire [253:0] stage1_43;
   wire [255:0] stage1_44;
   wire [211:0] stage1_45;
   wire [297:0] stage1_46;
   wire [235:0] stage1_47;
   wire [197:0] stage1_48;
   wire [172:0] stage1_49;
   wire [189:0] stage1_50;
   wire [274:0] stage1_51;
   wire [198:0] stage1_52;
   wire [168:0] stage1_53;
   wire [230:0] stage1_54;
   wire [266:0] stage1_55;
   wire [186:0] stage1_56;
   wire [188:0] stage1_57;
   wire [219:0] stage1_58;
   wire [205:0] stage1_59;
   wire [214:0] stage1_60;
   wire [218:0] stage1_61;
   wire [192:0] stage1_62;
   wire [307:0] stage1_63;
   wire [123:0] stage1_64;
   wire [53:0] stage1_65;
   wire [37:0] stage2_0;
   wire [53:0] stage2_1;
   wire [62:0] stage2_2;
   wire [113:0] stage2_3;
   wire [111:0] stage2_4;
   wire [151:0] stage2_5;
   wire [91:0] stage2_6;
   wire [72:0] stage2_7;
   wire [159:0] stage2_8;
   wire [142:0] stage2_9;
   wire [163:0] stage2_10;
   wire [138:0] stage2_11;
   wire [106:0] stage2_12;
   wire [77:0] stage2_13;
   wire [107:0] stage2_14;
   wire [140:0] stage2_15;
   wire [82:0] stage2_16;
   wire [86:0] stage2_17;
   wire [118:0] stage2_18;
   wire [112:0] stage2_19;
   wire [92:0] stage2_20;
   wire [127:0] stage2_21;
   wire [107:0] stage2_22;
   wire [75:0] stage2_23;
   wire [101:0] stage2_24;
   wire [95:0] stage2_25;
   wire [84:0] stage2_26;
   wire [105:0] stage2_27;
   wire [91:0] stage2_28;
   wire [86:0] stage2_29;
   wire [116:0] stage2_30;
   wire [98:0] stage2_31;
   wire [105:0] stage2_32;
   wire [75:0] stage2_33;
   wire [131:0] stage2_34;
   wire [132:0] stage2_35;
   wire [74:0] stage2_36;
   wire [89:0] stage2_37;
   wire [139:0] stage2_38;
   wire [136:0] stage2_39;
   wire [112:0] stage2_40;
   wire [105:0] stage2_41;
   wire [85:0] stage2_42;
   wire [78:0] stage2_43;
   wire [118:0] stage2_44;
   wire [117:0] stage2_45;
   wire [87:0] stage2_46;
   wire [103:0] stage2_47;
   wire [129:0] stage2_48;
   wire [95:0] stage2_49;
   wire [85:0] stage2_50;
   wire [87:0] stage2_51;
   wire [104:0] stage2_52;
   wire [114:0] stage2_53;
   wire [99:0] stage2_54;
   wire [105:0] stage2_55;
   wire [114:0] stage2_56;
   wire [65:0] stage2_57;
   wire [85:0] stage2_58;
   wire [109:0] stage2_59;
   wire [84:0] stage2_60;
   wire [74:0] stage2_61;
   wire [104:0] stage2_62;
   wire [98:0] stage2_63;
   wire [141:0] stage2_64;
   wire [55:0] stage2_65;
   wire [41:0] stage2_66;
   wire [20:0] stage3_0;
   wire [21:0] stage3_1;
   wire [42:0] stage3_2;
   wire [28:0] stage3_3;
   wire [111:0] stage3_4;
   wire [52:0] stage3_5;
   wire [77:0] stage3_6;
   wire [50:0] stage3_7;
   wire [34:0] stage3_8;
   wire [53:0] stage3_9;
   wire [99:0] stage3_10;
   wire [57:0] stage3_11;
   wire [67:0] stage3_12;
   wire [56:0] stage3_13;
   wire [31:0] stage3_14;
   wire [47:0] stage3_15;
   wire [50:0] stage3_16;
   wire [35:0] stage3_17;
   wire [59:0] stage3_18;
   wire [47:0] stage3_19;
   wire [82:0] stage3_20;
   wire [38:0] stage3_21;
   wire [72:0] stage3_22;
   wire [42:0] stage3_23;
   wire [28:0] stage3_24;
   wire [32:0] stage3_25;
   wire [48:0] stage3_26;
   wire [48:0] stage3_27;
   wire [56:0] stage3_28;
   wire [47:0] stage3_29;
   wire [41:0] stage3_30;
   wire [37:0] stage3_31;
   wire [53:0] stage3_32;
   wire [45:0] stage3_33;
   wire [41:0] stage3_34;
   wire [56:0] stage3_35;
   wire [45:0] stage3_36;
   wire [52:0] stage3_37;
   wire [59:0] stage3_38;
   wire [57:0] stage3_39;
   wire [51:0] stage3_40;
   wire [42:0] stage3_41;
   wire [49:0] stage3_42;
   wire [45:0] stage3_43;
   wire [40:0] stage3_44;
   wire [43:0] stage3_45;
   wire [57:0] stage3_46;
   wire [43:0] stage3_47;
   wire [41:0] stage3_48;
   wire [41:0] stage3_49;
   wire [46:0] stage3_50;
   wire [62:0] stage3_51;
   wire [62:0] stage3_52;
   wire [74:0] stage3_53;
   wire [38:0] stage3_54;
   wire [66:0] stage3_55;
   wire [31:0] stage3_56;
   wire [53:0] stage3_57;
   wire [61:0] stage3_58;
   wire [49:0] stage3_59;
   wire [41:0] stage3_60;
   wire [52:0] stage3_61;
   wire [33:0] stage3_62;
   wire [47:0] stage3_63;
   wire [50:0] stage3_64;
   wire [37:0] stage3_65;
   wire [37:0] stage3_66;
   wire [13:0] stage3_67;
   wire [5:0] stage3_68;
   wire [8:0] stage4_0;
   wire [6:0] stage4_1;
   wire [10:0] stage4_2;
   wire [16:0] stage4_3;
   wire [30:0] stage4_4;
   wire [35:0] stage4_5;
   wire [23:0] stage4_6;
   wire [38:0] stage4_7;
   wire [27:0] stage4_8;
   wire [13:0] stage4_9;
   wire [41:0] stage4_10;
   wire [28:0] stage4_11;
   wire [23:0] stage4_12;
   wire [31:0] stage4_13;
   wire [29:0] stage4_14;
   wire [14:0] stage4_15;
   wire [26:0] stage4_16;
   wire [17:0] stage4_17;
   wire [20:0] stage4_18;
   wire [28:0] stage4_19;
   wire [33:0] stage4_20;
   wire [36:0] stage4_21;
   wire [17:0] stage4_22;
   wire [20:0] stage4_23;
   wire [21:0] stage4_24;
   wire [20:0] stage4_25;
   wire [18:0] stage4_26;
   wire [26:0] stage4_27;
   wire [18:0] stage4_28;
   wire [21:0] stage4_29;
   wire [32:0] stage4_30;
   wire [14:0] stage4_31;
   wire [29:0] stage4_32;
   wire [28:0] stage4_33;
   wire [18:0] stage4_34;
   wire [35:0] stage4_35;
   wire [35:0] stage4_36;
   wire [17:0] stage4_37;
   wire [19:0] stage4_38;
   wire [23:0] stage4_39;
   wire [27:0] stage4_40;
   wire [19:0] stage4_41;
   wire [37:0] stage4_42;
   wire [13:0] stage4_43;
   wire [24:0] stage4_44;
   wire [28:0] stage4_45;
   wire [16:0] stage4_46;
   wire [20:0] stage4_47;
   wire [22:0] stage4_48;
   wire [12:0] stage4_49;
   wire [21:0] stage4_50;
   wire [35:0] stage4_51;
   wire [18:0] stage4_52;
   wire [43:0] stage4_53;
   wire [25:0] stage4_54;
   wire [38:0] stage4_55;
   wire [13:0] stage4_56;
   wire [25:0] stage4_57;
   wire [23:0] stage4_58;
   wire [20:0] stage4_59;
   wire [21:0] stage4_60;
   wire [31:0] stage4_61;
   wire [16:0] stage4_62;
   wire [13:0] stage4_63;
   wire [33:0] stage4_64;
   wire [35:0] stage4_65;
   wire [10:0] stage4_66;
   wire [10:0] stage4_67;
   wire [13:0] stage4_68;
   wire [1:0] stage4_69;
   wire [4:0] stage5_0;
   wire [1:0] stage5_1;
   wire [4:0] stage5_2;
   wire [7:0] stage5_3;
   wire [10:0] stage5_4;
   wire [15:0] stage5_5;
   wire [9:0] stage5_6;
   wire [10:0] stage5_7;
   wire [18:0] stage5_8;
   wire [10:0] stage5_9;
   wire [20:0] stage5_10;
   wire [13:0] stage5_11;
   wire [10:0] stage5_12;
   wire [14:0] stage5_13;
   wire [15:0] stage5_14;
   wire [11:0] stage5_15;
   wire [7:0] stage5_16;
   wire [6:0] stage5_17;
   wire [11:0] stage5_18;
   wire [15:0] stage5_19;
   wire [13:0] stage5_20;
   wire [10:0] stage5_21;
   wire [13:0] stage5_22;
   wire [9:0] stage5_23;
   wire [8:0] stage5_24;
   wire [9:0] stage5_25;
   wire [14:0] stage5_26;
   wire [5:0] stage5_27;
   wire [9:0] stage5_28;
   wire [14:0] stage5_29;
   wire [8:0] stage5_30;
   wire [9:0] stage5_31;
   wire [19:0] stage5_32;
   wire [11:0] stage5_33;
   wire [13:0] stage5_34;
   wire [13:0] stage5_35;
   wire [12:0] stage5_36;
   wire [10:0] stage5_37;
   wire [9:0] stage5_38;
   wire [9:0] stage5_39;
   wire [10:0] stage5_40;
   wire [8:0] stage5_41;
   wire [18:0] stage5_42;
   wire [10:0] stage5_43;
   wire [12:0] stage5_44;
   wire [14:0] stage5_45;
   wire [11:0] stage5_46;
   wire [11:0] stage5_47;
   wire [13:0] stage5_48;
   wire [5:0] stage5_49;
   wire [11:0] stage5_50;
   wire [18:0] stage5_51;
   wire [9:0] stage5_52;
   wire [12:0] stage5_53;
   wire [16:0] stage5_54;
   wire [21:0] stage5_55;
   wire [8:0] stage5_56;
   wire [13:0] stage5_57;
   wire [15:0] stage5_58;
   wire [7:0] stage5_59;
   wire [14:0] stage5_60;
   wire [15:0] stage5_61;
   wire [11:0] stage5_62;
   wire [8:0] stage5_63;
   wire [14:0] stage5_64;
   wire [17:0] stage5_65;
   wire [7:0] stage5_66;
   wire [10:0] stage5_67;
   wire [13:0] stage5_68;
   wire [2:0] stage5_69;
   wire [0:0] stage5_70;
   wire [4:0] stage6_0;
   wire [1:0] stage6_1;
   wire [4:0] stage6_2;
   wire [1:0] stage6_3;
   wire [5:0] stage6_4;
   wire [3:0] stage6_5;
   wire [7:0] stage6_6;
   wire [4:0] stage6_7;
   wire [5:0] stage6_8;
   wire [9:0] stage6_9;
   wire [4:0] stage6_10;
   wire [6:0] stage6_11;
   wire [6:0] stage6_12;
   wire [9:0] stage6_13;
   wire [6:0] stage6_14;
   wire [5:0] stage6_15;
   wire [4:0] stage6_16;
   wire [4:0] stage6_17;
   wire [5:0] stage6_18;
   wire [4:0] stage6_19;
   wire [5:0] stage6_20;
   wire [5:0] stage6_21;
   wire [5:0] stage6_22;
   wire [6:0] stage6_23;
   wire [6:0] stage6_24;
   wire [2:0] stage6_25;
   wire [7:0] stage6_26;
   wire [4:0] stage6_27;
   wire [5:0] stage6_28;
   wire [5:0] stage6_29;
   wire [4:0] stage6_30;
   wire [5:0] stage6_31;
   wire [5:0] stage6_32;
   wire [5:0] stage6_33;
   wire [8:0] stage6_34;
   wire [4:0] stage6_35;
   wire [5:0] stage6_36;
   wire [5:0] stage6_37;
   wire [4:0] stage6_38;
   wire [3:0] stage6_39;
   wire [5:0] stage6_40;
   wire [7:0] stage6_41;
   wire [6:0] stage6_42;
   wire [6:0] stage6_43;
   wire [4:0] stage6_44;
   wire [8:0] stage6_45;
   wire [4:0] stage6_46;
   wire [6:0] stage6_47;
   wire [4:0] stage6_48;
   wire [5:0] stage6_49;
   wire [2:0] stage6_50;
   wire [7:0] stage6_51;
   wire [6:0] stage6_52;
   wire [4:0] stage6_53;
   wire [5:0] stage6_54;
   wire [9:0] stage6_55;
   wire [9:0] stage6_56;
   wire [6:0] stage6_57;
   wire [5:0] stage6_58;
   wire [4:0] stage6_59;
   wire [4:0] stage6_60;
   wire [8:0] stage6_61;
   wire [5:0] stage6_62;
   wire [4:0] stage6_63;
   wire [8:0] stage6_64;
   wire [4:0] stage6_65;
   wire [4:0] stage6_66;
   wire [4:0] stage6_67;
   wire [16:0] stage6_68;
   wire [4:0] stage6_69;
   wire [0:0] stage6_70;
   wire [4:0] stage7_0;
   wire [1:0] stage7_1;
   wire [4:0] stage7_2;
   wire [1:0] stage7_3;
   wire [0:0] stage7_4;
   wire [1:0] stage7_5;
   wire [2:0] stage7_6;
   wire [2:0] stage7_7;
   wire [4:0] stage7_8;
   wire [5:0] stage7_9;
   wire [1:0] stage7_10;
   wire [3:0] stage7_11;
   wire [1:0] stage7_12;
   wire [5:0] stage7_13;
   wire [2:0] stage7_14;
   wire [5:0] stage7_15;
   wire [2:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [6:0] stage7_19;
   wire [2:0] stage7_20;
   wire [5:0] stage7_21;
   wire [6:0] stage7_22;
   wire [0:0] stage7_23;
   wire [3:0] stage7_24;
   wire [1:0] stage7_25;
   wire [5:0] stage7_26;
   wire [4:0] stage7_27;
   wire [0:0] stage7_28;
   wire [4:0] stage7_29;
   wire [6:0] stage7_30;
   wire [1:0] stage7_31;
   wire [5:0] stage7_32;
   wire [0:0] stage7_33;
   wire [5:0] stage7_34;
   wire [5:0] stage7_35;
   wire [0:0] stage7_36;
   wire [1:0] stage7_37;
   wire [6:0] stage7_38;
   wire [0:0] stage7_39;
   wire [6:0] stage7_40;
   wire [4:0] stage7_41;
   wire [2:0] stage7_42;
   wire [3:0] stage7_43;
   wire [1:0] stage7_44;
   wire [4:0] stage7_45;
   wire [2:0] stage7_46;
   wire [7:0] stage7_47;
   wire [0:0] stage7_48;
   wire [1:0] stage7_49;
   wire [2:0] stage7_50;
   wire [3:0] stage7_51;
   wire [3:0] stage7_52;
   wire [5:0] stage7_53;
   wire [0:0] stage7_54;
   wire [6:0] stage7_55;
   wire [6:0] stage7_56;
   wire [1:0] stage7_57;
   wire [1:0] stage7_58;
   wire [6:0] stage7_59;
   wire [5:0] stage7_60;
   wire [1:0] stage7_61;
   wire [1:0] stage7_62;
   wire [2:0] stage7_63;
   wire [3:0] stage7_64;
   wire [2:0] stage7_65;
   wire [5:0] stage7_66;
   wire [0:0] stage7_67;
   wire [4:0] stage7_68;
   wire [4:0] stage7_69;
   wire [2:0] stage7_70;
   wire [1:0] stage7_71;
   wire [0:0] stage8_0;
   wire [1:0] stage8_1;
   wire [1:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [1:0] stage8_5;
   wire [0:0] stage8_6;
   wire [1:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [1:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [1:0] stage8_24;
   wire [1:0] stage8_25;
   wire [1:0] stage8_26;
   wire [1:0] stage8_27;
   wire [1:0] stage8_28;
   wire [1:0] stage8_29;
   wire [1:0] stage8_30;
   wire [1:0] stage8_31;
   wire [1:0] stage8_32;
   wire [1:0] stage8_33;
   wire [1:0] stage8_34;
   wire [1:0] stage8_35;
   wire [1:0] stage8_36;
   wire [1:0] stage8_37;
   wire [1:0] stage8_38;
   wire [1:0] stage8_39;
   wire [1:0] stage8_40;
   wire [1:0] stage8_41;
   wire [1:0] stage8_42;
   wire [1:0] stage8_43;
   wire [1:0] stage8_44;
   wire [1:0] stage8_45;
   wire [0:0] stage8_46;
   wire [1:0] stage8_47;
   wire [1:0] stage8_48;
   wire [1:0] stage8_49;
   wire [1:0] stage8_50;
   wire [1:0] stage8_51;
   wire [1:0] stage8_52;
   wire [1:0] stage8_53;
   wire [1:0] stage8_54;
   wire [1:0] stage8_55;
   wire [1:0] stage8_56;
   wire [1:0] stage8_57;
   wire [1:0] stage8_58;
   wire [1:0] stage8_59;
   wire [1:0] stage8_60;
   wire [1:0] stage8_61;
   wire [1:0] stage8_62;
   wire [1:0] stage8_63;
   wire [1:0] stage8_64;
   wire [1:0] stage8_65;
   wire [1:0] stage8_66;
   wire [1:0] stage8_67;
   wire [1:0] stage8_68;
   wire [1:0] stage8_69;
   wire [1:0] stage8_70;
   wire [1:0] stage8_71;
   wire [1:0] stage8_72;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;
   assign dst25 = stage8_25;
   assign dst26 = stage8_26;
   assign dst27 = stage8_27;
   assign dst28 = stage8_28;
   assign dst29 = stage8_29;
   assign dst30 = stage8_30;
   assign dst31 = stage8_31;
   assign dst32 = stage8_32;
   assign dst33 = stage8_33;
   assign dst34 = stage8_34;
   assign dst35 = stage8_35;
   assign dst36 = stage8_36;
   assign dst37 = stage8_37;
   assign dst38 = stage8_38;
   assign dst39 = stage8_39;
   assign dst40 = stage8_40;
   assign dst41 = stage8_41;
   assign dst42 = stage8_42;
   assign dst43 = stage8_43;
   assign dst44 = stage8_44;
   assign dst45 = stage8_45;
   assign dst46 = stage8_46;
   assign dst47 = stage8_47;
   assign dst48 = stage8_48;
   assign dst49 = stage8_49;
   assign dst50 = stage8_50;
   assign dst51 = stage8_51;
   assign dst52 = stage8_52;
   assign dst53 = stage8_53;
   assign dst54 = stage8_54;
   assign dst55 = stage8_55;
   assign dst56 = stage8_56;
   assign dst57 = stage8_57;
   assign dst58 = stage8_58;
   assign dst59 = stage8_59;
   assign dst60 = stage8_60;
   assign dst61 = stage8_61;
   assign dst62 = stage8_62;
   assign dst63 = stage8_63;
   assign dst64 = stage8_64;
   assign dst65 = stage8_65;
   assign dst66 = stage8_66;
   assign dst67 = stage8_67;
   assign dst68 = stage8_68;
   assign dst69 = stage8_69;
   assign dst70 = stage8_70;
   assign dst71 = stage8_71;
   assign dst72 = stage8_72;

   gpc117_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6]},
      {stage0_1[0]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[1]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[2]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27]},
      {stage0_1[3]},
      {stage0_2[3]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[4]},
      {stage0_2[4]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc117_4 gpc5 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_1[5]},
      {stage0_2[5]},
      {stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc117_4 gpc6 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_1[6]},
      {stage0_2[6]},
      {stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc117_4 gpc7 (
      {stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_1[7]},
      {stage0_2[7]},
      {stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc117_4 gpc8 (
      {stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[8]},
      {stage0_2[8]},
      {stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc117_4 gpc9 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[9]},
      {stage0_2[9]},
      {stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc117_4 gpc10 (
      {stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76]},
      {stage0_1[10]},
      {stage0_2[10]},
      {stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc117_4 gpc11 (
      {stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_1[11]},
      {stage0_2[11]},
      {stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc117_4 gpc12 (
      {stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_1[12]},
      {stage0_2[12]},
      {stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_2[13]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[94], stage0_0[95], stage0_0[96]},
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_2[14]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_2[15]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[100], stage0_0[101], stage0_0[102]},
      {stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36]},
      {stage0_2[16]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42]},
      {stage0_2[17]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48]},
      {stage0_2[18]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54]},
      {stage0_2[19]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60]},
      {stage0_2[20]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66]},
      {stage0_2[21]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72]},
      {stage0_2[22]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78]},
      {stage0_2[23]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84]},
      {stage0_2[24]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90]},
      {stage0_2[25]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96]},
      {stage0_2[26]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102]},
      {stage0_2[27]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108]},
      {stage0_2[28]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114]},
      {stage0_2[29]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120]},
      {stage0_2[30]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126]},
      {stage0_2[31]},
      {stage0_3[18]},
      {stage1_4[18],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[148], stage0_0[149], stage0_0[150]},
      {stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132]},
      {stage0_2[32]},
      {stage0_3[19]},
      {stage1_4[19],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138]},
      {stage0_2[33]},
      {stage0_3[20]},
      {stage1_4[20],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144]},
      {stage0_2[34]},
      {stage0_3[21]},
      {stage1_4[21],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150]},
      {stage0_2[35]},
      {stage0_3[22]},
      {stage1_4[22],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[160], stage0_0[161], stage0_0[162]},
      {stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156]},
      {stage0_2[36]},
      {stage0_3[23]},
      {stage1_4[23],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162]},
      {stage0_2[37]},
      {stage0_3[24]},
      {stage1_4[24],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[166], stage0_0[167], stage0_0[168]},
      {stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168]},
      {stage0_2[38]},
      {stage0_3[25]},
      {stage1_4[25],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174]},
      {stage0_2[39]},
      {stage0_3[26]},
      {stage1_4[26],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[172], stage0_0[173], stage0_0[174]},
      {stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180]},
      {stage0_2[40]},
      {stage0_3[27]},
      {stage1_4[27],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186]},
      {stage0_2[41]},
      {stage0_3[28]},
      {stage1_4[28],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[29],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[30],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195]},
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59]},
      {stage1_4[31],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201]},
      {stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65]},
      {stage1_4[32],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207]},
      {stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71]},
      {stage1_4[33],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213]},
      {stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77]},
      {stage1_4[34],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219]},
      {stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83]},
      {stage1_4[35],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225]},
      {stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89]},
      {stage1_4[36],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231]},
      {stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95]},
      {stage1_4[37],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237]},
      {stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101]},
      {stage1_4[38],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243]},
      {stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107]},
      {stage1_4[39],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249]},
      {stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113]},
      {stage1_4[40],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[250], stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255]},
      {stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119]},
      {stage1_4[41],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[256], stage0_0[257], stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261]},
      {stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125]},
      {stage1_4[42],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[262], stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267]},
      {stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131]},
      {stage1_4[43],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[268], stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272], stage0_0[273]},
      {stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137]},
      {stage1_4[44],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[274], stage0_0[275], stage0_0[276], stage0_0[277], stage0_0[278], stage0_0[279]},
      {stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143]},
      {stage1_4[45],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[280], stage0_0[281], stage0_0[282], stage0_0[283], stage0_0[284], stage0_0[285]},
      {stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149]},
      {stage1_4[46],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[286], stage0_0[287], stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291]},
      {stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155]},
      {stage1_4[47],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[292], stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297]},
      {stage0_2[156], stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161]},
      {stage1_4[48],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[298], stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302], stage0_0[303]},
      {stage0_2[162], stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167]},
      {stage1_4[49],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[304], stage0_0[305], stage0_0[306], stage0_0[307], stage0_0[308], stage0_0[309]},
      {stage0_2[168], stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173]},
      {stage1_4[50],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[310], stage0_0[311], stage0_0[312], stage0_0[313], stage0_0[314], stage0_0[315]},
      {stage0_2[174], stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179]},
      {stage1_4[51],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[316], stage0_0[317], stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321]},
      {stage0_2[180], stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185]},
      {stage1_4[52],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[322], stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327]},
      {stage0_2[186], stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191]},
      {stage1_4[53],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[328], stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332], stage0_0[333]},
      {stage0_2[192], stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197]},
      {stage1_4[54],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[334], stage0_0[335], stage0_0[336], stage0_0[337], stage0_0[338], stage0_0[339]},
      {stage0_2[198], stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203]},
      {stage1_4[55],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[340], stage0_0[341], stage0_0[342], stage0_0[343], stage0_0[344], stage0_0[345]},
      {stage0_2[204], stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209]},
      {stage1_4[56],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[346], stage0_0[347], stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351]},
      {stage0_2[210], stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215]},
      {stage1_4[57],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[352], stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357]},
      {stage0_2[216], stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221]},
      {stage1_4[58],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[358], stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362], stage0_0[363]},
      {stage0_2[222], stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227]},
      {stage1_4[59],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[364], stage0_0[365], stage0_0[366], stage0_0[367], stage0_0[368], stage0_0[369]},
      {stage0_2[228], stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233]},
      {stage1_4[60],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[370], stage0_0[371], stage0_0[372], stage0_0[373], stage0_0[374], stage0_0[375]},
      {stage0_2[234], stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239]},
      {stage1_4[61],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[376], stage0_0[377], stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381]},
      {stage0_2[240], stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245]},
      {stage1_4[62],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[382], stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387]},
      {stage0_2[246], stage0_2[247], stage0_2[248], stage0_2[249], stage0_2[250], stage0_2[251]},
      {stage1_4[63],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[388], stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392], stage0_0[393]},
      {stage0_2[252], stage0_2[253], stage0_2[254], stage0_2[255], stage0_2[256], stage0_2[257]},
      {stage1_4[64],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[394], stage0_0[395], stage0_0[396], stage0_0[397], stage0_0[398], stage0_0[399]},
      {stage0_2[258], stage0_2[259], stage0_2[260], stage0_2[261], stage0_2[262], stage0_2[263]},
      {stage1_4[65],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[400], stage0_0[401], stage0_0[402], stage0_0[403], stage0_0[404], stage0_0[405]},
      {stage0_2[264], stage0_2[265], stage0_2[266], stage0_2[267], stage0_2[268], stage0_2[269]},
      {stage1_4[66],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[406], stage0_0[407], stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411]},
      {stage0_2[270], stage0_2[271], stage0_2[272], stage0_2[273], stage0_2[274], stage0_2[275]},
      {stage1_4[67],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[412], stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417]},
      {stage0_2[276], stage0_2[277], stage0_2[278], stage0_2[279], stage0_2[280], stage0_2[281]},
      {stage1_4[68],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[418], stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422], stage0_0[423]},
      {stage0_2[282], stage0_2[283], stage0_2[284], stage0_2[285], stage0_2[286], stage0_2[287]},
      {stage1_4[69],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[424], stage0_0[425], stage0_0[426], stage0_0[427], stage0_0[428], stage0_0[429]},
      {stage0_2[288], stage0_2[289], stage0_2[290], stage0_2[291], stage0_2[292], stage0_2[293]},
      {stage1_4[70],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[430], stage0_0[431], stage0_0[432], stage0_0[433], stage0_0[434], stage0_0[435]},
      {stage0_2[294], stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299]},
      {stage1_4[71],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_0[436], stage0_0[437], stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441]},
      {stage0_2[300], stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305]},
      {stage1_4[72],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc606_5 gpc86 (
      {stage0_0[442], stage0_0[443], stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447]},
      {stage0_2[306], stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311]},
      {stage1_4[73],stage1_3[86],stage1_2[86],stage1_1[86],stage1_0[86]}
   );
   gpc606_5 gpc87 (
      {stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192]},
      {stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34]},
      {stage1_5[0],stage1_4[74],stage1_3[87],stage1_2[87],stage1_1[87]}
   );
   gpc606_5 gpc88 (
      {stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198]},
      {stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40]},
      {stage1_5[1],stage1_4[75],stage1_3[88],stage1_2[88],stage1_1[88]}
   );
   gpc606_5 gpc89 (
      {stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204]},
      {stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46]},
      {stage1_5[2],stage1_4[76],stage1_3[89],stage1_2[89],stage1_1[89]}
   );
   gpc606_5 gpc90 (
      {stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210]},
      {stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52]},
      {stage1_5[3],stage1_4[77],stage1_3[90],stage1_2[90],stage1_1[90]}
   );
   gpc606_5 gpc91 (
      {stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216]},
      {stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58]},
      {stage1_5[4],stage1_4[78],stage1_3[91],stage1_2[91],stage1_1[91]}
   );
   gpc606_5 gpc92 (
      {stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222]},
      {stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64]},
      {stage1_5[5],stage1_4[79],stage1_3[92],stage1_2[92],stage1_1[92]}
   );
   gpc606_5 gpc93 (
      {stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228]},
      {stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70]},
      {stage1_5[6],stage1_4[80],stage1_3[93],stage1_2[93],stage1_1[93]}
   );
   gpc606_5 gpc94 (
      {stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234]},
      {stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76]},
      {stage1_5[7],stage1_4[81],stage1_3[94],stage1_2[94],stage1_1[94]}
   );
   gpc606_5 gpc95 (
      {stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239], stage0_1[240]},
      {stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82]},
      {stage1_5[8],stage1_4[82],stage1_3[95],stage1_2[95],stage1_1[95]}
   );
   gpc606_5 gpc96 (
      {stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245], stage0_1[246]},
      {stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88]},
      {stage1_5[9],stage1_4[83],stage1_3[96],stage1_2[96],stage1_1[96]}
   );
   gpc606_5 gpc97 (
      {stage0_1[247], stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251], stage0_1[252]},
      {stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94]},
      {stage1_5[10],stage1_4[84],stage1_3[97],stage1_2[97],stage1_1[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[253], stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257], stage0_1[258]},
      {stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100]},
      {stage1_5[11],stage1_4[85],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[259], stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263], stage0_1[264]},
      {stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage1_5[12],stage1_4[86],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[265], stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269], stage0_1[270]},
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112]},
      {stage1_5[13],stage1_4[87],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[271], stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275], stage0_1[276]},
      {stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118]},
      {stage1_5[14],stage1_4[88],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[277], stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281], stage0_1[282]},
      {stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124]},
      {stage1_5[15],stage1_4[89],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[283], stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287], stage0_1[288]},
      {stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130]},
      {stage1_5[16],stage1_4[90],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[289], stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293], stage0_1[294]},
      {stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136]},
      {stage1_5[17],stage1_4[91],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[295], stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299], stage0_1[300]},
      {stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142]},
      {stage1_5[18],stage1_4[92],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[301], stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305], stage0_1[306]},
      {stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148]},
      {stage1_5[19],stage1_4[93],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[307], stage0_1[308], stage0_1[309], stage0_1[310], stage0_1[311], stage0_1[312]},
      {stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154]},
      {stage1_5[20],stage1_4[94],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[313], stage0_1[314], stage0_1[315], stage0_1[316], stage0_1[317], stage0_1[318]},
      {stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160]},
      {stage1_5[21],stage1_4[95],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[319], stage0_1[320], stage0_1[321], stage0_1[322], stage0_1[323], stage0_1[324]},
      {stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166]},
      {stage1_5[22],stage1_4[96],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[325], stage0_1[326], stage0_1[327], stage0_1[328], stage0_1[329], stage0_1[330]},
      {stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170], stage0_3[171], stage0_3[172]},
      {stage1_5[23],stage1_4[97],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[331], stage0_1[332], stage0_1[333], stage0_1[334], stage0_1[335], stage0_1[336]},
      {stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178]},
      {stage1_5[24],stage1_4[98],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[337], stage0_1[338], stage0_1[339], stage0_1[340], stage0_1[341], stage0_1[342]},
      {stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184]},
      {stage1_5[25],stage1_4[99],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[343], stage0_1[344], stage0_1[345], stage0_1[346], stage0_1[347], stage0_1[348]},
      {stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190]},
      {stage1_5[26],stage1_4[100],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[349], stage0_1[350], stage0_1[351], stage0_1[352], stage0_1[353], stage0_1[354]},
      {stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196]},
      {stage1_5[27],stage1_4[101],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[355], stage0_1[356], stage0_1[357], stage0_1[358], stage0_1[359], stage0_1[360]},
      {stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201], stage0_3[202]},
      {stage1_5[28],stage1_4[102],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[361], stage0_1[362], stage0_1[363], stage0_1[364], stage0_1[365], stage0_1[366]},
      {stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208]},
      {stage1_5[29],stage1_4[103],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[367], stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371], stage0_1[372]},
      {stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214]},
      {stage1_5[30],stage1_4[104],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[373], stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377], stage0_1[378]},
      {stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220]},
      {stage1_5[31],stage1_4[105],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[379], stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383], stage0_1[384]},
      {stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226]},
      {stage1_5[32],stage1_4[106],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[385], stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389], stage0_1[390]},
      {stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232]},
      {stage1_5[33],stage1_4[107],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[391], stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395], stage0_1[396]},
      {stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238]},
      {stage1_5[34],stage1_4[108],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[397], stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401], stage0_1[402]},
      {stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244]},
      {stage1_5[35],stage1_4[109],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[403], stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407], stage0_1[408]},
      {stage0_3[245], stage0_3[246], stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250]},
      {stage1_5[36],stage1_4[110],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[409], stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413], stage0_1[414]},
      {stage0_3[251], stage0_3[252], stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256]},
      {stage1_5[37],stage1_4[111],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[415], stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419], stage0_1[420]},
      {stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260], stage0_3[261], stage0_3[262]},
      {stage1_5[38],stage1_4[112],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[421], stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425], stage0_1[426]},
      {stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266], stage0_3[267], stage0_3[268]},
      {stage1_5[39],stage1_4[113],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[427], stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431], stage0_1[432]},
      {stage0_3[269], stage0_3[270], stage0_3[271], stage0_3[272], stage0_3[273], stage0_3[274]},
      {stage1_5[40],stage1_4[114],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[433], stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437], stage0_1[438]},
      {stage0_3[275], stage0_3[276], stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280]},
      {stage1_5[41],stage1_4[115],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_2[312], stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[42],stage1_4[116],stage1_3[129],stage1_2[129]}
   );
   gpc606_5 gpc130 (
      {stage0_2[318], stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[43],stage1_4[117],stage1_3[130],stage1_2[130]}
   );
   gpc606_5 gpc131 (
      {stage0_2[324], stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[44],stage1_4[118],stage1_3[131],stage1_2[131]}
   );
   gpc606_5 gpc132 (
      {stage0_2[330], stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[45],stage1_4[119],stage1_3[132],stage1_2[132]}
   );
   gpc606_5 gpc133 (
      {stage0_2[336], stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[46],stage1_4[120],stage1_3[133],stage1_2[133]}
   );
   gpc606_5 gpc134 (
      {stage0_2[342], stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[47],stage1_4[121],stage1_3[134],stage1_2[134]}
   );
   gpc606_5 gpc135 (
      {stage0_2[348], stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[48],stage1_4[122],stage1_3[135],stage1_2[135]}
   );
   gpc606_5 gpc136 (
      {stage0_2[354], stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358], stage0_2[359]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[49],stage1_4[123],stage1_3[136],stage1_2[136]}
   );
   gpc606_5 gpc137 (
      {stage0_2[360], stage0_2[361], stage0_2[362], stage0_2[363], stage0_2[364], stage0_2[365]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[50],stage1_4[124],stage1_3[137],stage1_2[137]}
   );
   gpc606_5 gpc138 (
      {stage0_2[366], stage0_2[367], stage0_2[368], stage0_2[369], stage0_2[370], stage0_2[371]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[51],stage1_4[125],stage1_3[138],stage1_2[138]}
   );
   gpc606_5 gpc139 (
      {stage0_2[372], stage0_2[373], stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[52],stage1_4[126],stage1_3[139],stage1_2[139]}
   );
   gpc606_5 gpc140 (
      {stage0_2[378], stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[53],stage1_4[127],stage1_3[140],stage1_2[140]}
   );
   gpc606_5 gpc141 (
      {stage0_2[384], stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388], stage0_2[389]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[54],stage1_4[128],stage1_3[141],stage1_2[141]}
   );
   gpc606_5 gpc142 (
      {stage0_2[390], stage0_2[391], stage0_2[392], stage0_2[393], stage0_2[394], stage0_2[395]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[55],stage1_4[129],stage1_3[142],stage1_2[142]}
   );
   gpc606_5 gpc143 (
      {stage0_2[396], stage0_2[397], stage0_2[398], stage0_2[399], stage0_2[400], stage0_2[401]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[56],stage1_4[130],stage1_3[143],stage1_2[143]}
   );
   gpc606_5 gpc144 (
      {stage0_2[402], stage0_2[403], stage0_2[404], stage0_2[405], stage0_2[406], stage0_2[407]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[57],stage1_4[131],stage1_3[144],stage1_2[144]}
   );
   gpc606_5 gpc145 (
      {stage0_2[408], stage0_2[409], stage0_2[410], stage0_2[411], stage0_2[412], stage0_2[413]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[58],stage1_4[132],stage1_3[145],stage1_2[145]}
   );
   gpc606_5 gpc146 (
      {stage0_2[414], stage0_2[415], stage0_2[416], stage0_2[417], stage0_2[418], stage0_2[419]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[59],stage1_4[133],stage1_3[146],stage1_2[146]}
   );
   gpc606_5 gpc147 (
      {stage0_2[420], stage0_2[421], stage0_2[422], stage0_2[423], stage0_2[424], stage0_2[425]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage1_6[18],stage1_5[60],stage1_4[134],stage1_3[147],stage1_2[147]}
   );
   gpc606_5 gpc148 (
      {stage0_2[426], stage0_2[427], stage0_2[428], stage0_2[429], stage0_2[430], stage0_2[431]},
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage1_6[19],stage1_5[61],stage1_4[135],stage1_3[148],stage1_2[148]}
   );
   gpc606_5 gpc149 (
      {stage0_2[432], stage0_2[433], stage0_2[434], stage0_2[435], stage0_2[436], stage0_2[437]},
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage1_6[20],stage1_5[62],stage1_4[136],stage1_3[149],stage1_2[149]}
   );
   gpc606_5 gpc150 (
      {stage0_2[438], stage0_2[439], stage0_2[440], stage0_2[441], stage0_2[442], stage0_2[443]},
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage1_6[21],stage1_5[63],stage1_4[137],stage1_3[150],stage1_2[150]}
   );
   gpc606_5 gpc151 (
      {stage0_2[444], stage0_2[445], stage0_2[446], stage0_2[447], stage0_2[448], stage0_2[449]},
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage1_6[22],stage1_5[64],stage1_4[138],stage1_3[151],stage1_2[151]}
   );
   gpc606_5 gpc152 (
      {stage0_2[450], stage0_2[451], stage0_2[452], stage0_2[453], stage0_2[454], stage0_2[455]},
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage1_6[23],stage1_5[65],stage1_4[139],stage1_3[152],stage1_2[152]}
   );
   gpc606_5 gpc153 (
      {stage0_2[456], stage0_2[457], stage0_2[458], stage0_2[459], stage0_2[460], stage0_2[461]},
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage1_6[24],stage1_5[66],stage1_4[140],stage1_3[153],stage1_2[153]}
   );
   gpc606_5 gpc154 (
      {stage0_2[462], stage0_2[463], stage0_2[464], stage0_2[465], stage0_2[466], stage0_2[467]},
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage1_6[25],stage1_5[67],stage1_4[141],stage1_3[154],stage1_2[154]}
   );
   gpc606_5 gpc155 (
      {stage0_2[468], stage0_2[469], stage0_2[470], stage0_2[471], stage0_2[472], stage0_2[473]},
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage1_6[26],stage1_5[68],stage1_4[142],stage1_3[155],stage1_2[155]}
   );
   gpc606_5 gpc156 (
      {stage0_2[474], stage0_2[475], stage0_2[476], stage0_2[477], stage0_2[478], stage0_2[479]},
      {stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167]},
      {stage1_6[27],stage1_5[69],stage1_4[143],stage1_3[156],stage1_2[156]}
   );
   gpc606_5 gpc157 (
      {stage0_2[480], stage0_2[481], stage0_2[482], stage0_2[483], stage0_2[484], stage0_2[485]},
      {stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173]},
      {stage1_6[28],stage1_5[70],stage1_4[144],stage1_3[157],stage1_2[157]}
   );
   gpc615_5 gpc158 (
      {stage0_3[281], stage0_3[282], stage0_3[283], stage0_3[284], stage0_3[285]},
      {stage0_4[174]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[29],stage1_5[71],stage1_4[145],stage1_3[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[286], stage0_3[287], stage0_3[288], stage0_3[289], stage0_3[290]},
      {stage0_4[175]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[30],stage1_5[72],stage1_4[146],stage1_3[159]}
   );
   gpc615_5 gpc160 (
      {stage0_3[291], stage0_3[292], stage0_3[293], stage0_3[294], stage0_3[295]},
      {stage0_4[176]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[31],stage1_5[73],stage1_4[147],stage1_3[160]}
   );
   gpc615_5 gpc161 (
      {stage0_3[296], stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300]},
      {stage0_4[177]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[32],stage1_5[74],stage1_4[148],stage1_3[161]}
   );
   gpc615_5 gpc162 (
      {stage0_3[301], stage0_3[302], stage0_3[303], stage0_3[304], stage0_3[305]},
      {stage0_4[178]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[33],stage1_5[75],stage1_4[149],stage1_3[162]}
   );
   gpc615_5 gpc163 (
      {stage0_3[306], stage0_3[307], stage0_3[308], stage0_3[309], stage0_3[310]},
      {stage0_4[179]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[34],stage1_5[76],stage1_4[150],stage1_3[163]}
   );
   gpc615_5 gpc164 (
      {stage0_3[311], stage0_3[312], stage0_3[313], stage0_3[314], stage0_3[315]},
      {stage0_4[180]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[35],stage1_5[77],stage1_4[151],stage1_3[164]}
   );
   gpc615_5 gpc165 (
      {stage0_3[316], stage0_3[317], stage0_3[318], stage0_3[319], stage0_3[320]},
      {stage0_4[181]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[36],stage1_5[78],stage1_4[152],stage1_3[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[321], stage0_3[322], stage0_3[323], stage0_3[324], stage0_3[325]},
      {stage0_4[182]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[37],stage1_5[79],stage1_4[153],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[326], stage0_3[327], stage0_3[328], stage0_3[329], stage0_3[330]},
      {stage0_4[183]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[38],stage1_5[80],stage1_4[154],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[331], stage0_3[332], stage0_3[333], stage0_3[334], stage0_3[335]},
      {stage0_4[184]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[39],stage1_5[81],stage1_4[155],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[336], stage0_3[337], stage0_3[338], stage0_3[339], stage0_3[340]},
      {stage0_4[185]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[40],stage1_5[82],stage1_4[156],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[341], stage0_3[342], stage0_3[343], stage0_3[344], stage0_3[345]},
      {stage0_4[186]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[41],stage1_5[83],stage1_4[157],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[346], stage0_3[347], stage0_3[348], stage0_3[349], stage0_3[350]},
      {stage0_4[187]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[42],stage1_5[84],stage1_4[158],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[351], stage0_3[352], stage0_3[353], stage0_3[354], stage0_3[355]},
      {stage0_4[188]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[43],stage1_5[85],stage1_4[159],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[356], stage0_3[357], stage0_3[358], stage0_3[359], stage0_3[360]},
      {stage0_4[189]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[44],stage1_5[86],stage1_4[160],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[361], stage0_3[362], stage0_3[363], stage0_3[364], stage0_3[365]},
      {stage0_4[190]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[45],stage1_5[87],stage1_4[161],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[366], stage0_3[367], stage0_3[368], stage0_3[369], stage0_3[370]},
      {stage0_4[191]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[46],stage1_5[88],stage1_4[162],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[371], stage0_3[372], stage0_3[373], stage0_3[374], stage0_3[375]},
      {stage0_4[192]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[47],stage1_5[89],stage1_4[163],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[376], stage0_3[377], stage0_3[378], stage0_3[379], stage0_3[380]},
      {stage0_4[193]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[48],stage1_5[90],stage1_4[164],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[381], stage0_3[382], stage0_3[383], stage0_3[384], stage0_3[385]},
      {stage0_4[194]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[49],stage1_5[91],stage1_4[165],stage1_3[178]}
   );
   gpc615_5 gpc179 (
      {stage0_3[386], stage0_3[387], stage0_3[388], stage0_3[389], stage0_3[390]},
      {stage0_4[195]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[50],stage1_5[92],stage1_4[166],stage1_3[179]}
   );
   gpc615_5 gpc180 (
      {stage0_3[391], stage0_3[392], stage0_3[393], stage0_3[394], stage0_3[395]},
      {stage0_4[196]},
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage1_7[22],stage1_6[51],stage1_5[93],stage1_4[167],stage1_3[180]}
   );
   gpc615_5 gpc181 (
      {stage0_3[396], stage0_3[397], stage0_3[398], stage0_3[399], stage0_3[400]},
      {stage0_4[197]},
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage1_7[23],stage1_6[52],stage1_5[94],stage1_4[168],stage1_3[181]}
   );
   gpc615_5 gpc182 (
      {stage0_3[401], stage0_3[402], stage0_3[403], stage0_3[404], stage0_3[405]},
      {stage0_4[198]},
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage1_7[24],stage1_6[53],stage1_5[95],stage1_4[169],stage1_3[182]}
   );
   gpc615_5 gpc183 (
      {stage0_3[406], stage0_3[407], stage0_3[408], stage0_3[409], stage0_3[410]},
      {stage0_4[199]},
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage1_7[25],stage1_6[54],stage1_5[96],stage1_4[170],stage1_3[183]}
   );
   gpc615_5 gpc184 (
      {stage0_3[411], stage0_3[412], stage0_3[413], stage0_3[414], stage0_3[415]},
      {stage0_4[200]},
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage1_7[26],stage1_6[55],stage1_5[97],stage1_4[171],stage1_3[184]}
   );
   gpc615_5 gpc185 (
      {stage0_3[416], stage0_3[417], stage0_3[418], stage0_3[419], stage0_3[420]},
      {stage0_4[201]},
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage1_7[27],stage1_6[56],stage1_5[98],stage1_4[172],stage1_3[185]}
   );
   gpc615_5 gpc186 (
      {stage0_3[421], stage0_3[422], stage0_3[423], stage0_3[424], stage0_3[425]},
      {stage0_4[202]},
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage1_7[28],stage1_6[57],stage1_5[99],stage1_4[173],stage1_3[186]}
   );
   gpc615_5 gpc187 (
      {stage0_3[426], stage0_3[427], stage0_3[428], stage0_3[429], stage0_3[430]},
      {stage0_4[203]},
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage1_7[29],stage1_6[58],stage1_5[100],stage1_4[174],stage1_3[187]}
   );
   gpc615_5 gpc188 (
      {stage0_3[431], stage0_3[432], stage0_3[433], stage0_3[434], stage0_3[435]},
      {stage0_4[204]},
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage1_7[30],stage1_6[59],stage1_5[101],stage1_4[175],stage1_3[188]}
   );
   gpc615_5 gpc189 (
      {stage0_3[436], stage0_3[437], stage0_3[438], stage0_3[439], stage0_3[440]},
      {stage0_4[205]},
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage1_7[31],stage1_6[60],stage1_5[102],stage1_4[176],stage1_3[189]}
   );
   gpc615_5 gpc190 (
      {stage0_3[441], stage0_3[442], stage0_3[443], stage0_3[444], stage0_3[445]},
      {stage0_4[206]},
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage1_7[32],stage1_6[61],stage1_5[103],stage1_4[177],stage1_3[190]}
   );
   gpc615_5 gpc191 (
      {stage0_3[446], stage0_3[447], stage0_3[448], stage0_3[449], stage0_3[450]},
      {stage0_4[207]},
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage1_7[33],stage1_6[62],stage1_5[104],stage1_4[178],stage1_3[191]}
   );
   gpc615_5 gpc192 (
      {stage0_3[451], stage0_3[452], stage0_3[453], stage0_3[454], stage0_3[455]},
      {stage0_4[208]},
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage1_7[34],stage1_6[63],stage1_5[105],stage1_4[179],stage1_3[192]}
   );
   gpc615_5 gpc193 (
      {stage0_3[456], stage0_3[457], stage0_3[458], stage0_3[459], stage0_3[460]},
      {stage0_4[209]},
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage1_7[35],stage1_6[64],stage1_5[106],stage1_4[180],stage1_3[193]}
   );
   gpc615_5 gpc194 (
      {stage0_3[461], stage0_3[462], stage0_3[463], stage0_3[464], stage0_3[465]},
      {stage0_4[210]},
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage1_7[36],stage1_6[65],stage1_5[107],stage1_4[181],stage1_3[194]}
   );
   gpc606_5 gpc195 (
      {stage0_4[211], stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[37],stage1_6[66],stage1_5[108],stage1_4[182]}
   );
   gpc606_5 gpc196 (
      {stage0_4[217], stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[38],stage1_6[67],stage1_5[109],stage1_4[183]}
   );
   gpc606_5 gpc197 (
      {stage0_4[223], stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[39],stage1_6[68],stage1_5[110],stage1_4[184]}
   );
   gpc606_5 gpc198 (
      {stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[40],stage1_6[69],stage1_5[111],stage1_4[185]}
   );
   gpc606_5 gpc199 (
      {stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[41],stage1_6[70],stage1_5[112],stage1_4[186]}
   );
   gpc606_5 gpc200 (
      {stage0_4[241], stage0_4[242], stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[42],stage1_6[71],stage1_5[113],stage1_4[187]}
   );
   gpc606_5 gpc201 (
      {stage0_4[247], stage0_4[248], stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[43],stage1_6[72],stage1_5[114],stage1_4[188]}
   );
   gpc606_5 gpc202 (
      {stage0_4[253], stage0_4[254], stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[44],stage1_6[73],stage1_5[115],stage1_4[189]}
   );
   gpc606_5 gpc203 (
      {stage0_4[259], stage0_4[260], stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[45],stage1_6[74],stage1_5[116],stage1_4[190]}
   );
   gpc606_5 gpc204 (
      {stage0_4[265], stage0_4[266], stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[46],stage1_6[75],stage1_5[117],stage1_4[191]}
   );
   gpc606_5 gpc205 (
      {stage0_4[271], stage0_4[272], stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[47],stage1_6[76],stage1_5[118],stage1_4[192]}
   );
   gpc606_5 gpc206 (
      {stage0_4[277], stage0_4[278], stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[48],stage1_6[77],stage1_5[119],stage1_4[193]}
   );
   gpc606_5 gpc207 (
      {stage0_4[283], stage0_4[284], stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[49],stage1_6[78],stage1_5[120],stage1_4[194]}
   );
   gpc606_5 gpc208 (
      {stage0_4[289], stage0_4[290], stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[50],stage1_6[79],stage1_5[121],stage1_4[195]}
   );
   gpc606_5 gpc209 (
      {stage0_4[295], stage0_4[296], stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[51],stage1_6[80],stage1_5[122],stage1_4[196]}
   );
   gpc606_5 gpc210 (
      {stage0_4[301], stage0_4[302], stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[52],stage1_6[81],stage1_5[123],stage1_4[197]}
   );
   gpc606_5 gpc211 (
      {stage0_4[307], stage0_4[308], stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[53],stage1_6[82],stage1_5[124],stage1_4[198]}
   );
   gpc606_5 gpc212 (
      {stage0_4[313], stage0_4[314], stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[54],stage1_6[83],stage1_5[125],stage1_4[199]}
   );
   gpc606_5 gpc213 (
      {stage0_4[319], stage0_4[320], stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[55],stage1_6[84],stage1_5[126],stage1_4[200]}
   );
   gpc606_5 gpc214 (
      {stage0_4[325], stage0_4[326], stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[56],stage1_6[85],stage1_5[127],stage1_4[201]}
   );
   gpc606_5 gpc215 (
      {stage0_4[331], stage0_4[332], stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[57],stage1_6[86],stage1_5[128],stage1_4[202]}
   );
   gpc606_5 gpc216 (
      {stage0_4[337], stage0_4[338], stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[58],stage1_6[87],stage1_5[129],stage1_4[203]}
   );
   gpc606_5 gpc217 (
      {stage0_4[343], stage0_4[344], stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[59],stage1_6[88],stage1_5[130],stage1_4[204]}
   );
   gpc606_5 gpc218 (
      {stage0_4[349], stage0_4[350], stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[60],stage1_6[89],stage1_5[131],stage1_4[205]}
   );
   gpc606_5 gpc219 (
      {stage0_4[355], stage0_4[356], stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[61],stage1_6[90],stage1_5[132],stage1_4[206]}
   );
   gpc606_5 gpc220 (
      {stage0_4[361], stage0_4[362], stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[62],stage1_6[91],stage1_5[133],stage1_4[207]}
   );
   gpc606_5 gpc221 (
      {stage0_4[367], stage0_4[368], stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[63],stage1_6[92],stage1_5[134],stage1_4[208]}
   );
   gpc606_5 gpc222 (
      {stage0_4[373], stage0_4[374], stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[64],stage1_6[93],stage1_5[135],stage1_4[209]}
   );
   gpc606_5 gpc223 (
      {stage0_4[379], stage0_4[380], stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[65],stage1_6[94],stage1_5[136],stage1_4[210]}
   );
   gpc606_5 gpc224 (
      {stage0_4[385], stage0_4[386], stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[66],stage1_6[95],stage1_5[137],stage1_4[211]}
   );
   gpc606_5 gpc225 (
      {stage0_4[391], stage0_4[392], stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[67],stage1_6[96],stage1_5[138],stage1_4[212]}
   );
   gpc606_5 gpc226 (
      {stage0_4[397], stage0_4[398], stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[68],stage1_6[97],stage1_5[139],stage1_4[213]}
   );
   gpc606_5 gpc227 (
      {stage0_4[403], stage0_4[404], stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[69],stage1_6[98],stage1_5[140],stage1_4[214]}
   );
   gpc606_5 gpc228 (
      {stage0_4[409], stage0_4[410], stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[70],stage1_6[99],stage1_5[141],stage1_4[215]}
   );
   gpc606_5 gpc229 (
      {stage0_4[415], stage0_4[416], stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[71],stage1_6[100],stage1_5[142],stage1_4[216]}
   );
   gpc606_5 gpc230 (
      {stage0_4[421], stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[72],stage1_6[101],stage1_5[143],stage1_4[217]}
   );
   gpc606_5 gpc231 (
      {stage0_4[427], stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431], stage0_4[432]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[73],stage1_6[102],stage1_5[144],stage1_4[218]}
   );
   gpc606_5 gpc232 (
      {stage0_4[433], stage0_4[434], stage0_4[435], stage0_4[436], stage0_4[437], stage0_4[438]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[74],stage1_6[103],stage1_5[145],stage1_4[219]}
   );
   gpc606_5 gpc233 (
      {stage0_4[439], stage0_4[440], stage0_4[441], stage0_4[442], stage0_4[443], stage0_4[444]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[75],stage1_6[104],stage1_5[146],stage1_4[220]}
   );
   gpc606_5 gpc234 (
      {stage0_4[445], stage0_4[446], stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[76],stage1_6[105],stage1_5[147],stage1_4[221]}
   );
   gpc606_5 gpc235 (
      {stage0_4[451], stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455], stage0_4[456]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[77],stage1_6[106],stage1_5[148],stage1_4[222]}
   );
   gpc606_5 gpc236 (
      {stage0_4[457], stage0_4[458], stage0_4[459], stage0_4[460], stage0_4[461], stage0_4[462]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[78],stage1_6[107],stage1_5[149],stage1_4[223]}
   );
   gpc606_5 gpc237 (
      {stage0_4[463], stage0_4[464], stage0_4[465], stage0_4[466], stage0_4[467], stage0_4[468]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[79],stage1_6[108],stage1_5[150],stage1_4[224]}
   );
   gpc606_5 gpc238 (
      {stage0_4[469], stage0_4[470], stage0_4[471], stage0_4[472], stage0_4[473], stage0_4[474]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[80],stage1_6[109],stage1_5[151],stage1_4[225]}
   );
   gpc606_5 gpc239 (
      {stage0_4[475], stage0_4[476], stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[81],stage1_6[110],stage1_5[152],stage1_4[226]}
   );
   gpc606_5 gpc240 (
      {stage0_4[481], stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485], 1'b0},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[82],stage1_6[111],stage1_5[153],stage1_4[227]}
   );
   gpc606_5 gpc241 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[46],stage1_7[83],stage1_6[112],stage1_5[154]}
   );
   gpc606_5 gpc242 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[47],stage1_7[84],stage1_6[113],stage1_5[155]}
   );
   gpc606_5 gpc243 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[48],stage1_7[85],stage1_6[114],stage1_5[156]}
   );
   gpc606_5 gpc244 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[49],stage1_7[86],stage1_6[115],stage1_5[157]}
   );
   gpc606_5 gpc245 (
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[50],stage1_7[87],stage1_6[116],stage1_5[158]}
   );
   gpc606_5 gpc246 (
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[51],stage1_7[88],stage1_6[117],stage1_5[159]}
   );
   gpc606_5 gpc247 (
      {stage0_5[258], stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[52],stage1_7[89],stage1_6[118],stage1_5[160]}
   );
   gpc606_5 gpc248 (
      {stage0_5[264], stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[53],stage1_7[90],stage1_6[119],stage1_5[161]}
   );
   gpc606_5 gpc249 (
      {stage0_5[270], stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[54],stage1_7[91],stage1_6[120],stage1_5[162]}
   );
   gpc606_5 gpc250 (
      {stage0_5[276], stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[55],stage1_7[92],stage1_6[121],stage1_5[163]}
   );
   gpc606_5 gpc251 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[56],stage1_7[93],stage1_6[122],stage1_5[164]}
   );
   gpc606_5 gpc252 (
      {stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[57],stage1_7[94],stage1_6[123],stage1_5[165]}
   );
   gpc606_5 gpc253 (
      {stage0_5[294], stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[58],stage1_7[95],stage1_6[124],stage1_5[166]}
   );
   gpc606_5 gpc254 (
      {stage0_5[300], stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[59],stage1_7[96],stage1_6[125],stage1_5[167]}
   );
   gpc606_5 gpc255 (
      {stage0_5[306], stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[60],stage1_7[97],stage1_6[126],stage1_5[168]}
   );
   gpc606_5 gpc256 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[61],stage1_7[98],stage1_6[127],stage1_5[169]}
   );
   gpc606_5 gpc257 (
      {stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[62],stage1_7[99],stage1_6[128],stage1_5[170]}
   );
   gpc606_5 gpc258 (
      {stage0_5[324], stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[63],stage1_7[100],stage1_6[129],stage1_5[171]}
   );
   gpc606_5 gpc259 (
      {stage0_5[330], stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[64],stage1_7[101],stage1_6[130],stage1_5[172]}
   );
   gpc606_5 gpc260 (
      {stage0_5[336], stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[65],stage1_7[102],stage1_6[131],stage1_5[173]}
   );
   gpc606_5 gpc261 (
      {stage0_5[342], stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[66],stage1_7[103],stage1_6[132],stage1_5[174]}
   );
   gpc606_5 gpc262 (
      {stage0_5[348], stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[67],stage1_7[104],stage1_6[133],stage1_5[175]}
   );
   gpc606_5 gpc263 (
      {stage0_5[354], stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[68],stage1_7[105],stage1_6[134],stage1_5[176]}
   );
   gpc606_5 gpc264 (
      {stage0_5[360], stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[69],stage1_7[106],stage1_6[135],stage1_5[177]}
   );
   gpc606_5 gpc265 (
      {stage0_5[366], stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[70],stage1_7[107],stage1_6[136],stage1_5[178]}
   );
   gpc606_5 gpc266 (
      {stage0_5[372], stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[71],stage1_7[108],stage1_6[137],stage1_5[179]}
   );
   gpc606_5 gpc267 (
      {stage0_5[378], stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[72],stage1_7[109],stage1_6[138],stage1_5[180]}
   );
   gpc606_5 gpc268 (
      {stage0_5[384], stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[73],stage1_7[110],stage1_6[139],stage1_5[181]}
   );
   gpc606_5 gpc269 (
      {stage0_5[390], stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[74],stage1_7[111],stage1_6[140],stage1_5[182]}
   );
   gpc606_5 gpc270 (
      {stage0_5[396], stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[75],stage1_7[112],stage1_6[141],stage1_5[183]}
   );
   gpc606_5 gpc271 (
      {stage0_5[402], stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[76],stage1_7[113],stage1_6[142],stage1_5[184]}
   );
   gpc606_5 gpc272 (
      {stage0_5[408], stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[77],stage1_7[114],stage1_6[143],stage1_5[185]}
   );
   gpc606_5 gpc273 (
      {stage0_5[414], stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[78],stage1_7[115],stage1_6[144],stage1_5[186]}
   );
   gpc606_5 gpc274 (
      {stage0_5[420], stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[79],stage1_7[116],stage1_6[145],stage1_5[187]}
   );
   gpc606_5 gpc275 (
      {stage0_5[426], stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[80],stage1_7[117],stage1_6[146],stage1_5[188]}
   );
   gpc606_5 gpc276 (
      {stage0_5[432], stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[81],stage1_7[118],stage1_6[147],stage1_5[189]}
   );
   gpc606_5 gpc277 (
      {stage0_5[438], stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[82],stage1_7[119],stage1_6[148],stage1_5[190]}
   );
   gpc606_5 gpc278 (
      {stage0_5[444], stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[83],stage1_7[120],stage1_6[149],stage1_5[191]}
   );
   gpc606_5 gpc279 (
      {stage0_5[450], stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[84],stage1_7[121],stage1_6[150],stage1_5[192]}
   );
   gpc606_5 gpc280 (
      {stage0_5[456], stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[85],stage1_7[122],stage1_6[151],stage1_5[193]}
   );
   gpc606_5 gpc281 (
      {stage0_5[462], stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[86],stage1_7[123],stage1_6[152],stage1_5[194]}
   );
   gpc606_5 gpc282 (
      {stage0_5[468], stage0_5[469], stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[87],stage1_7[124],stage1_6[153],stage1_5[195]}
   );
   gpc606_5 gpc283 (
      {stage0_5[474], stage0_5[475], stage0_5[476], stage0_5[477], stage0_5[478], stage0_5[479]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[88],stage1_7[125],stage1_6[154],stage1_5[196]}
   );
   gpc606_5 gpc284 (
      {stage0_5[480], stage0_5[481], stage0_5[482], stage0_5[483], stage0_5[484], stage0_5[485]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[89],stage1_7[126],stage1_6[155],stage1_5[197]}
   );
   gpc615_5 gpc285 (
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280]},
      {stage0_7[264]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[44],stage1_8[90],stage1_7[127],stage1_6[156]}
   );
   gpc615_5 gpc286 (
      {stage0_6[281], stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285]},
      {stage0_7[265]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[45],stage1_8[91],stage1_7[128],stage1_6[157]}
   );
   gpc615_5 gpc287 (
      {stage0_6[286], stage0_6[287], stage0_6[288], stage0_6[289], stage0_6[290]},
      {stage0_7[266]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[46],stage1_8[92],stage1_7[129],stage1_6[158]}
   );
   gpc615_5 gpc288 (
      {stage0_6[291], stage0_6[292], stage0_6[293], stage0_6[294], stage0_6[295]},
      {stage0_7[267]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[47],stage1_8[93],stage1_7[130],stage1_6[159]}
   );
   gpc615_5 gpc289 (
      {stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299], stage0_6[300]},
      {stage0_7[268]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[48],stage1_8[94],stage1_7[131],stage1_6[160]}
   );
   gpc615_5 gpc290 (
      {stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage0_7[269]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[49],stage1_8[95],stage1_7[132],stage1_6[161]}
   );
   gpc615_5 gpc291 (
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310]},
      {stage0_7[270]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[50],stage1_8[96],stage1_7[133],stage1_6[162]}
   );
   gpc615_5 gpc292 (
      {stage0_6[311], stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315]},
      {stage0_7[271]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[51],stage1_8[97],stage1_7[134],stage1_6[163]}
   );
   gpc615_5 gpc293 (
      {stage0_6[316], stage0_6[317], stage0_6[318], stage0_6[319], stage0_6[320]},
      {stage0_7[272]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[52],stage1_8[98],stage1_7[135],stage1_6[164]}
   );
   gpc615_5 gpc294 (
      {stage0_6[321], stage0_6[322], stage0_6[323], stage0_6[324], stage0_6[325]},
      {stage0_7[273]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[53],stage1_8[99],stage1_7[136],stage1_6[165]}
   );
   gpc615_5 gpc295 (
      {stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329], stage0_6[330]},
      {stage0_7[274]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[54],stage1_8[100],stage1_7[137],stage1_6[166]}
   );
   gpc615_5 gpc296 (
      {stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335]},
      {stage0_7[275]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[55],stage1_8[101],stage1_7[138],stage1_6[167]}
   );
   gpc615_5 gpc297 (
      {stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340]},
      {stage0_7[276]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[56],stage1_8[102],stage1_7[139],stage1_6[168]}
   );
   gpc615_5 gpc298 (
      {stage0_6[341], stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345]},
      {stage0_7[277]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[57],stage1_8[103],stage1_7[140],stage1_6[169]}
   );
   gpc615_5 gpc299 (
      {stage0_6[346], stage0_6[347], stage0_6[348], stage0_6[349], stage0_6[350]},
      {stage0_7[278]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[58],stage1_8[104],stage1_7[141],stage1_6[170]}
   );
   gpc615_5 gpc300 (
      {stage0_6[351], stage0_6[352], stage0_6[353], stage0_6[354], stage0_6[355]},
      {stage0_7[279]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[59],stage1_8[105],stage1_7[142],stage1_6[171]}
   );
   gpc615_5 gpc301 (
      {stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359], stage0_6[360]},
      {stage0_7[280]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[60],stage1_8[106],stage1_7[143],stage1_6[172]}
   );
   gpc615_5 gpc302 (
      {stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365]},
      {stage0_7[281]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[61],stage1_8[107],stage1_7[144],stage1_6[173]}
   );
   gpc615_5 gpc303 (
      {stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370]},
      {stage0_7[282]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[62],stage1_8[108],stage1_7[145],stage1_6[174]}
   );
   gpc615_5 gpc304 (
      {stage0_6[371], stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375]},
      {stage0_7[283]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[63],stage1_8[109],stage1_7[146],stage1_6[175]}
   );
   gpc615_5 gpc305 (
      {stage0_6[376], stage0_6[377], stage0_6[378], stage0_6[379], stage0_6[380]},
      {stage0_7[284]},
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage1_10[20],stage1_9[64],stage1_8[110],stage1_7[147],stage1_6[176]}
   );
   gpc615_5 gpc306 (
      {stage0_6[381], stage0_6[382], stage0_6[383], stage0_6[384], stage0_6[385]},
      {stage0_7[285]},
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage1_10[21],stage1_9[65],stage1_8[111],stage1_7[148],stage1_6[177]}
   );
   gpc615_5 gpc307 (
      {stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389], stage0_6[390]},
      {stage0_7[286]},
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage1_10[22],stage1_9[66],stage1_8[112],stage1_7[149],stage1_6[178]}
   );
   gpc615_5 gpc308 (
      {stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395]},
      {stage0_7[287]},
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage1_10[23],stage1_9[67],stage1_8[113],stage1_7[150],stage1_6[179]}
   );
   gpc615_5 gpc309 (
      {stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400]},
      {stage0_7[288]},
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage1_10[24],stage1_9[68],stage1_8[114],stage1_7[151],stage1_6[180]}
   );
   gpc615_5 gpc310 (
      {stage0_6[401], stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405]},
      {stage0_7[289]},
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage1_10[25],stage1_9[69],stage1_8[115],stage1_7[152],stage1_6[181]}
   );
   gpc615_5 gpc311 (
      {stage0_6[406], stage0_6[407], stage0_6[408], stage0_6[409], stage0_6[410]},
      {stage0_7[290]},
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage1_10[26],stage1_9[70],stage1_8[116],stage1_7[153],stage1_6[182]}
   );
   gpc615_5 gpc312 (
      {stage0_6[411], stage0_6[412], stage0_6[413], stage0_6[414], stage0_6[415]},
      {stage0_7[291]},
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage1_10[27],stage1_9[71],stage1_8[117],stage1_7[154],stage1_6[183]}
   );
   gpc615_5 gpc313 (
      {stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419], stage0_6[420]},
      {stage0_7[292]},
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage1_10[28],stage1_9[72],stage1_8[118],stage1_7[155],stage1_6[184]}
   );
   gpc615_5 gpc314 (
      {stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425]},
      {stage0_7[293]},
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage1_10[29],stage1_9[73],stage1_8[119],stage1_7[156],stage1_6[185]}
   );
   gpc615_5 gpc315 (
      {stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430]},
      {stage0_7[294]},
      {stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185]},
      {stage1_10[30],stage1_9[74],stage1_8[120],stage1_7[157],stage1_6[186]}
   );
   gpc615_5 gpc316 (
      {stage0_6[431], stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435]},
      {stage0_7[295]},
      {stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191]},
      {stage1_10[31],stage1_9[75],stage1_8[121],stage1_7[158],stage1_6[187]}
   );
   gpc615_5 gpc317 (
      {stage0_6[436], stage0_6[437], stage0_6[438], stage0_6[439], stage0_6[440]},
      {stage0_7[296]},
      {stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage1_10[32],stage1_9[76],stage1_8[122],stage1_7[159],stage1_6[188]}
   );
   gpc615_5 gpc318 (
      {stage0_6[441], stage0_6[442], stage0_6[443], stage0_6[444], stage0_6[445]},
      {stage0_7[297]},
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203]},
      {stage1_10[33],stage1_9[77],stage1_8[123],stage1_7[160],stage1_6[189]}
   );
   gpc615_5 gpc319 (
      {stage0_6[446], stage0_6[447], stage0_6[448], stage0_6[449], stage0_6[450]},
      {stage0_7[298]},
      {stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage1_10[34],stage1_9[78],stage1_8[124],stage1_7[161],stage1_6[190]}
   );
   gpc615_5 gpc320 (
      {stage0_6[451], stage0_6[452], stage0_6[453], stage0_6[454], stage0_6[455]},
      {stage0_7[299]},
      {stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215]},
      {stage1_10[35],stage1_9[79],stage1_8[125],stage1_7[162],stage1_6[191]}
   );
   gpc615_5 gpc321 (
      {stage0_6[456], stage0_6[457], stage0_6[458], stage0_6[459], stage0_6[460]},
      {stage0_7[300]},
      {stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221]},
      {stage1_10[36],stage1_9[80],stage1_8[126],stage1_7[163],stage1_6[192]}
   );
   gpc615_5 gpc322 (
      {stage0_6[461], stage0_6[462], stage0_6[463], stage0_6[464], stage0_6[465]},
      {stage0_7[301]},
      {stage0_8[222], stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227]},
      {stage1_10[37],stage1_9[81],stage1_8[127],stage1_7[164],stage1_6[193]}
   );
   gpc615_5 gpc323 (
      {stage0_7[302], stage0_7[303], stage0_7[304], stage0_7[305], stage0_7[306]},
      {stage0_8[228]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[38],stage1_9[82],stage1_8[128],stage1_7[165]}
   );
   gpc615_5 gpc324 (
      {stage0_7[307], stage0_7[308], stage0_7[309], stage0_7[310], stage0_7[311]},
      {stage0_8[229]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[39],stage1_9[83],stage1_8[129],stage1_7[166]}
   );
   gpc615_5 gpc325 (
      {stage0_7[312], stage0_7[313], stage0_7[314], stage0_7[315], stage0_7[316]},
      {stage0_8[230]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[40],stage1_9[84],stage1_8[130],stage1_7[167]}
   );
   gpc615_5 gpc326 (
      {stage0_7[317], stage0_7[318], stage0_7[319], stage0_7[320], stage0_7[321]},
      {stage0_8[231]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[41],stage1_9[85],stage1_8[131],stage1_7[168]}
   );
   gpc615_5 gpc327 (
      {stage0_7[322], stage0_7[323], stage0_7[324], stage0_7[325], stage0_7[326]},
      {stage0_8[232]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[42],stage1_9[86],stage1_8[132],stage1_7[169]}
   );
   gpc615_5 gpc328 (
      {stage0_7[327], stage0_7[328], stage0_7[329], stage0_7[330], stage0_7[331]},
      {stage0_8[233]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[43],stage1_9[87],stage1_8[133],stage1_7[170]}
   );
   gpc615_5 gpc329 (
      {stage0_7[332], stage0_7[333], stage0_7[334], stage0_7[335], stage0_7[336]},
      {stage0_8[234]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[44],stage1_9[88],stage1_8[134],stage1_7[171]}
   );
   gpc615_5 gpc330 (
      {stage0_7[337], stage0_7[338], stage0_7[339], stage0_7[340], stage0_7[341]},
      {stage0_8[235]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[45],stage1_9[89],stage1_8[135],stage1_7[172]}
   );
   gpc615_5 gpc331 (
      {stage0_7[342], stage0_7[343], stage0_7[344], stage0_7[345], stage0_7[346]},
      {stage0_8[236]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[46],stage1_9[90],stage1_8[136],stage1_7[173]}
   );
   gpc615_5 gpc332 (
      {stage0_7[347], stage0_7[348], stage0_7[349], stage0_7[350], stage0_7[351]},
      {stage0_8[237]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[47],stage1_9[91],stage1_8[137],stage1_7[174]}
   );
   gpc615_5 gpc333 (
      {stage0_7[352], stage0_7[353], stage0_7[354], stage0_7[355], stage0_7[356]},
      {stage0_8[238]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[48],stage1_9[92],stage1_8[138],stage1_7[175]}
   );
   gpc615_5 gpc334 (
      {stage0_7[357], stage0_7[358], stage0_7[359], stage0_7[360], stage0_7[361]},
      {stage0_8[239]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[49],stage1_9[93],stage1_8[139],stage1_7[176]}
   );
   gpc615_5 gpc335 (
      {stage0_7[362], stage0_7[363], stage0_7[364], stage0_7[365], stage0_7[366]},
      {stage0_8[240]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[50],stage1_9[94],stage1_8[140],stage1_7[177]}
   );
   gpc615_5 gpc336 (
      {stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370], stage0_7[371]},
      {stage0_8[241]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[51],stage1_9[95],stage1_8[141],stage1_7[178]}
   );
   gpc615_5 gpc337 (
      {stage0_7[372], stage0_7[373], stage0_7[374], stage0_7[375], stage0_7[376]},
      {stage0_8[242]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[52],stage1_9[96],stage1_8[142],stage1_7[179]}
   );
   gpc615_5 gpc338 (
      {stage0_7[377], stage0_7[378], stage0_7[379], stage0_7[380], stage0_7[381]},
      {stage0_8[243]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[53],stage1_9[97],stage1_8[143],stage1_7[180]}
   );
   gpc615_5 gpc339 (
      {stage0_7[382], stage0_7[383], stage0_7[384], stage0_7[385], stage0_7[386]},
      {stage0_8[244]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[54],stage1_9[98],stage1_8[144],stage1_7[181]}
   );
   gpc615_5 gpc340 (
      {stage0_7[387], stage0_7[388], stage0_7[389], stage0_7[390], stage0_7[391]},
      {stage0_8[245]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[55],stage1_9[99],stage1_8[145],stage1_7[182]}
   );
   gpc615_5 gpc341 (
      {stage0_7[392], stage0_7[393], stage0_7[394], stage0_7[395], stage0_7[396]},
      {stage0_8[246]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[56],stage1_9[100],stage1_8[146],stage1_7[183]}
   );
   gpc615_5 gpc342 (
      {stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400], stage0_7[401]},
      {stage0_8[247]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[57],stage1_9[101],stage1_8[147],stage1_7[184]}
   );
   gpc615_5 gpc343 (
      {stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405], stage0_7[406]},
      {stage0_8[248]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[58],stage1_9[102],stage1_8[148],stage1_7[185]}
   );
   gpc615_5 gpc344 (
      {stage0_7[407], stage0_7[408], stage0_7[409], stage0_7[410], stage0_7[411]},
      {stage0_8[249]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[59],stage1_9[103],stage1_8[149],stage1_7[186]}
   );
   gpc615_5 gpc345 (
      {stage0_7[412], stage0_7[413], stage0_7[414], stage0_7[415], stage0_7[416]},
      {stage0_8[250]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[60],stage1_9[104],stage1_8[150],stage1_7[187]}
   );
   gpc615_5 gpc346 (
      {stage0_7[417], stage0_7[418], stage0_7[419], stage0_7[420], stage0_7[421]},
      {stage0_8[251]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[61],stage1_9[105],stage1_8[151],stage1_7[188]}
   );
   gpc615_5 gpc347 (
      {stage0_7[422], stage0_7[423], stage0_7[424], stage0_7[425], stage0_7[426]},
      {stage0_8[252]},
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage1_11[24],stage1_10[62],stage1_9[106],stage1_8[152],stage1_7[189]}
   );
   gpc615_5 gpc348 (
      {stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430], stage0_7[431]},
      {stage0_8[253]},
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage1_11[25],stage1_10[63],stage1_9[107],stage1_8[153],stage1_7[190]}
   );
   gpc615_5 gpc349 (
      {stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435], stage0_7[436]},
      {stage0_8[254]},
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage1_11[26],stage1_10[64],stage1_9[108],stage1_8[154],stage1_7[191]}
   );
   gpc615_5 gpc350 (
      {stage0_7[437], stage0_7[438], stage0_7[439], stage0_7[440], stage0_7[441]},
      {stage0_8[255]},
      {stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167]},
      {stage1_11[27],stage1_10[65],stage1_9[109],stage1_8[155],stage1_7[192]}
   );
   gpc615_5 gpc351 (
      {stage0_7[442], stage0_7[443], stage0_7[444], stage0_7[445], stage0_7[446]},
      {stage0_8[256]},
      {stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173]},
      {stage1_11[28],stage1_10[66],stage1_9[110],stage1_8[156],stage1_7[193]}
   );
   gpc615_5 gpc352 (
      {stage0_7[447], stage0_7[448], stage0_7[449], stage0_7[450], stage0_7[451]},
      {stage0_8[257]},
      {stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179]},
      {stage1_11[29],stage1_10[67],stage1_9[111],stage1_8[157],stage1_7[194]}
   );
   gpc615_5 gpc353 (
      {stage0_7[452], stage0_7[453], stage0_7[454], stage0_7[455], stage0_7[456]},
      {stage0_8[258]},
      {stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage1_11[30],stage1_10[68],stage1_9[112],stage1_8[158],stage1_7[195]}
   );
   gpc615_5 gpc354 (
      {stage0_7[457], stage0_7[458], stage0_7[459], stage0_7[460], stage0_7[461]},
      {stage0_8[259]},
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191]},
      {stage1_11[31],stage1_10[69],stage1_9[113],stage1_8[159],stage1_7[196]}
   );
   gpc606_5 gpc355 (
      {stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264], stage0_8[265]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[32],stage1_10[70],stage1_9[114],stage1_8[160]}
   );
   gpc606_5 gpc356 (
      {stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270], stage0_8[271]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[33],stage1_10[71],stage1_9[115],stage1_8[161]}
   );
   gpc606_5 gpc357 (
      {stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276], stage0_8[277]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[34],stage1_10[72],stage1_9[116],stage1_8[162]}
   );
   gpc606_5 gpc358 (
      {stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282], stage0_8[283]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[35],stage1_10[73],stage1_9[117],stage1_8[163]}
   );
   gpc606_5 gpc359 (
      {stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288], stage0_8[289]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[36],stage1_10[74],stage1_9[118],stage1_8[164]}
   );
   gpc606_5 gpc360 (
      {stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294], stage0_8[295]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[37],stage1_10[75],stage1_9[119],stage1_8[165]}
   );
   gpc606_5 gpc361 (
      {stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300], stage0_8[301]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[38],stage1_10[76],stage1_9[120],stage1_8[166]}
   );
   gpc606_5 gpc362 (
      {stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306], stage0_8[307]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[39],stage1_10[77],stage1_9[121],stage1_8[167]}
   );
   gpc606_5 gpc363 (
      {stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312], stage0_8[313]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[40],stage1_10[78],stage1_9[122],stage1_8[168]}
   );
   gpc606_5 gpc364 (
      {stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318], stage0_8[319]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[41],stage1_10[79],stage1_9[123],stage1_8[169]}
   );
   gpc606_5 gpc365 (
      {stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324], stage0_8[325]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[42],stage1_10[80],stage1_9[124],stage1_8[170]}
   );
   gpc606_5 gpc366 (
      {stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330], stage0_8[331]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[43],stage1_10[81],stage1_9[125],stage1_8[171]}
   );
   gpc606_5 gpc367 (
      {stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336], stage0_8[337]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[44],stage1_10[82],stage1_9[126],stage1_8[172]}
   );
   gpc606_5 gpc368 (
      {stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341], stage0_8[342], stage0_8[343]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[45],stage1_10[83],stage1_9[127],stage1_8[173]}
   );
   gpc606_5 gpc369 (
      {stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347], stage0_8[348], stage0_8[349]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[46],stage1_10[84],stage1_9[128],stage1_8[174]}
   );
   gpc606_5 gpc370 (
      {stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353], stage0_8[354], stage0_8[355]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[47],stage1_10[85],stage1_9[129],stage1_8[175]}
   );
   gpc606_5 gpc371 (
      {stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360], stage0_8[361]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[48],stage1_10[86],stage1_9[130],stage1_8[176]}
   );
   gpc606_5 gpc372 (
      {stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366], stage0_8[367]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[49],stage1_10[87],stage1_9[131],stage1_8[177]}
   );
   gpc606_5 gpc373 (
      {stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371], stage0_8[372], stage0_8[373]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[50],stage1_10[88],stage1_9[132],stage1_8[178]}
   );
   gpc606_5 gpc374 (
      {stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377], stage0_8[378], stage0_8[379]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[51],stage1_10[89],stage1_9[133],stage1_8[179]}
   );
   gpc606_5 gpc375 (
      {stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383], stage0_8[384], stage0_8[385]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[52],stage1_10[90],stage1_9[134],stage1_8[180]}
   );
   gpc606_5 gpc376 (
      {stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389], stage0_8[390], stage0_8[391]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[53],stage1_10[91],stage1_9[135],stage1_8[181]}
   );
   gpc606_5 gpc377 (
      {stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395], stage0_8[396], stage0_8[397]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[54],stage1_10[92],stage1_9[136],stage1_8[182]}
   );
   gpc606_5 gpc378 (
      {stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401], stage0_8[402], stage0_8[403]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[55],stage1_10[93],stage1_9[137],stage1_8[183]}
   );
   gpc606_5 gpc379 (
      {stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407], stage0_8[408], stage0_8[409]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[56],stage1_10[94],stage1_9[138],stage1_8[184]}
   );
   gpc606_5 gpc380 (
      {stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413], stage0_8[414], stage0_8[415]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[57],stage1_10[95],stage1_9[139],stage1_8[185]}
   );
   gpc606_5 gpc381 (
      {stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419], stage0_8[420], stage0_8[421]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[58],stage1_10[96],stage1_9[140],stage1_8[186]}
   );
   gpc606_5 gpc382 (
      {stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425], stage0_8[426], stage0_8[427]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[59],stage1_10[97],stage1_9[141],stage1_8[187]}
   );
   gpc606_5 gpc383 (
      {stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431], stage0_8[432], stage0_8[433]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[60],stage1_10[98],stage1_9[142],stage1_8[188]}
   );
   gpc606_5 gpc384 (
      {stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437], stage0_8[438], stage0_8[439]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[61],stage1_10[99],stage1_9[143],stage1_8[189]}
   );
   gpc606_5 gpc385 (
      {stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443], stage0_8[444], stage0_8[445]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[62],stage1_10[100],stage1_9[144],stage1_8[190]}
   );
   gpc606_5 gpc386 (
      {stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449], stage0_8[450], stage0_8[451]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[63],stage1_10[101],stage1_9[145],stage1_8[191]}
   );
   gpc606_5 gpc387 (
      {stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455], stage0_8[456], stage0_8[457]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[64],stage1_10[102],stage1_9[146],stage1_8[192]}
   );
   gpc606_5 gpc388 (
      {stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461], stage0_8[462], stage0_8[463]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[65],stage1_10[103],stage1_9[147],stage1_8[193]}
   );
   gpc606_5 gpc389 (
      {stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467], stage0_8[468], stage0_8[469]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[66],stage1_10[104],stage1_9[148],stage1_8[194]}
   );
   gpc606_5 gpc390 (
      {stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473], stage0_8[474], stage0_8[475]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[67],stage1_10[105],stage1_9[149],stage1_8[195]}
   );
   gpc606_5 gpc391 (
      {stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[36],stage1_11[68],stage1_10[106],stage1_9[150]}
   );
   gpc606_5 gpc392 (
      {stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[37],stage1_11[69],stage1_10[107],stage1_9[151]}
   );
   gpc606_5 gpc393 (
      {stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[38],stage1_11[70],stage1_10[108],stage1_9[152]}
   );
   gpc606_5 gpc394 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[39],stage1_11[71],stage1_10[109],stage1_9[153]}
   );
   gpc606_5 gpc395 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220], stage0_9[221]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[40],stage1_11[72],stage1_10[110],stage1_9[154]}
   );
   gpc606_5 gpc396 (
      {stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225], stage0_9[226], stage0_9[227]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[41],stage1_11[73],stage1_10[111],stage1_9[155]}
   );
   gpc606_5 gpc397 (
      {stage0_9[228], stage0_9[229], stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[42],stage1_11[74],stage1_10[112],stage1_9[156]}
   );
   gpc606_5 gpc398 (
      {stage0_9[234], stage0_9[235], stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[43],stage1_11[75],stage1_10[113],stage1_9[157]}
   );
   gpc606_5 gpc399 (
      {stage0_9[240], stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[44],stage1_11[76],stage1_10[114],stage1_9[158]}
   );
   gpc606_5 gpc400 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250], stage0_9[251]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[45],stage1_11[77],stage1_10[115],stage1_9[159]}
   );
   gpc606_5 gpc401 (
      {stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255], stage0_9[256], stage0_9[257]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[46],stage1_11[78],stage1_10[116],stage1_9[160]}
   );
   gpc606_5 gpc402 (
      {stage0_9[258], stage0_9[259], stage0_9[260], stage0_9[261], stage0_9[262], stage0_9[263]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[47],stage1_11[79],stage1_10[117],stage1_9[161]}
   );
   gpc606_5 gpc403 (
      {stage0_9[264], stage0_9[265], stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[48],stage1_11[80],stage1_10[118],stage1_9[162]}
   );
   gpc606_5 gpc404 (
      {stage0_9[270], stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[49],stage1_11[81],stage1_10[119],stage1_9[163]}
   );
   gpc606_5 gpc405 (
      {stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280], stage0_9[281]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[50],stage1_11[82],stage1_10[120],stage1_9[164]}
   );
   gpc606_5 gpc406 (
      {stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285], stage0_9[286], stage0_9[287]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[51],stage1_11[83],stage1_10[121],stage1_9[165]}
   );
   gpc606_5 gpc407 (
      {stage0_9[288], stage0_9[289], stage0_9[290], stage0_9[291], stage0_9[292], stage0_9[293]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[52],stage1_11[84],stage1_10[122],stage1_9[166]}
   );
   gpc606_5 gpc408 (
      {stage0_9[294], stage0_9[295], stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[53],stage1_11[85],stage1_10[123],stage1_9[167]}
   );
   gpc606_5 gpc409 (
      {stage0_9[300], stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[54],stage1_11[86],stage1_10[124],stage1_9[168]}
   );
   gpc606_5 gpc410 (
      {stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310], stage0_9[311]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[55],stage1_11[87],stage1_10[125],stage1_9[169]}
   );
   gpc606_5 gpc411 (
      {stage0_9[312], stage0_9[313], stage0_9[314], stage0_9[315], stage0_9[316], stage0_9[317]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[56],stage1_11[88],stage1_10[126],stage1_9[170]}
   );
   gpc606_5 gpc412 (
      {stage0_9[318], stage0_9[319], stage0_9[320], stage0_9[321], stage0_9[322], stage0_9[323]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[57],stage1_11[89],stage1_10[127],stage1_9[171]}
   );
   gpc606_5 gpc413 (
      {stage0_9[324], stage0_9[325], stage0_9[326], stage0_9[327], stage0_9[328], stage0_9[329]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[58],stage1_11[90],stage1_10[128],stage1_9[172]}
   );
   gpc606_5 gpc414 (
      {stage0_9[330], stage0_9[331], stage0_9[332], stage0_9[333], stage0_9[334], stage0_9[335]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[59],stage1_11[91],stage1_10[129],stage1_9[173]}
   );
   gpc606_5 gpc415 (
      {stage0_9[336], stage0_9[337], stage0_9[338], stage0_9[339], stage0_9[340], stage0_9[341]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[60],stage1_11[92],stage1_10[130],stage1_9[174]}
   );
   gpc606_5 gpc416 (
      {stage0_9[342], stage0_9[343], stage0_9[344], stage0_9[345], stage0_9[346], stage0_9[347]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[61],stage1_11[93],stage1_10[131],stage1_9[175]}
   );
   gpc606_5 gpc417 (
      {stage0_9[348], stage0_9[349], stage0_9[350], stage0_9[351], stage0_9[352], stage0_9[353]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[62],stage1_11[94],stage1_10[132],stage1_9[176]}
   );
   gpc606_5 gpc418 (
      {stage0_9[354], stage0_9[355], stage0_9[356], stage0_9[357], stage0_9[358], stage0_9[359]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[63],stage1_11[95],stage1_10[133],stage1_9[177]}
   );
   gpc606_5 gpc419 (
      {stage0_9[360], stage0_9[361], stage0_9[362], stage0_9[363], stage0_9[364], stage0_9[365]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[64],stage1_11[96],stage1_10[134],stage1_9[178]}
   );
   gpc606_5 gpc420 (
      {stage0_9[366], stage0_9[367], stage0_9[368], stage0_9[369], stage0_9[370], stage0_9[371]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[65],stage1_11[97],stage1_10[135],stage1_9[179]}
   );
   gpc606_5 gpc421 (
      {stage0_9[372], stage0_9[373], stage0_9[374], stage0_9[375], stage0_9[376], stage0_9[377]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[66],stage1_11[98],stage1_10[136],stage1_9[180]}
   );
   gpc606_5 gpc422 (
      {stage0_9[378], stage0_9[379], stage0_9[380], stage0_9[381], stage0_9[382], stage0_9[383]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[67],stage1_11[99],stage1_10[137],stage1_9[181]}
   );
   gpc606_5 gpc423 (
      {stage0_9[384], stage0_9[385], stage0_9[386], stage0_9[387], stage0_9[388], stage0_9[389]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[68],stage1_11[100],stage1_10[138],stage1_9[182]}
   );
   gpc606_5 gpc424 (
      {stage0_9[390], stage0_9[391], stage0_9[392], stage0_9[393], stage0_9[394], stage0_9[395]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[69],stage1_11[101],stage1_10[139],stage1_9[183]}
   );
   gpc606_5 gpc425 (
      {stage0_9[396], stage0_9[397], stage0_9[398], stage0_9[399], stage0_9[400], stage0_9[401]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[70],stage1_11[102],stage1_10[140],stage1_9[184]}
   );
   gpc606_5 gpc426 (
      {stage0_9[402], stage0_9[403], stage0_9[404], stage0_9[405], stage0_9[406], stage0_9[407]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[71],stage1_11[103],stage1_10[141],stage1_9[185]}
   );
   gpc606_5 gpc427 (
      {stage0_9[408], stage0_9[409], stage0_9[410], stage0_9[411], stage0_9[412], stage0_9[413]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[72],stage1_11[104],stage1_10[142],stage1_9[186]}
   );
   gpc606_5 gpc428 (
      {stage0_9[414], stage0_9[415], stage0_9[416], stage0_9[417], stage0_9[418], stage0_9[419]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[73],stage1_11[105],stage1_10[143],stage1_9[187]}
   );
   gpc606_5 gpc429 (
      {stage0_9[420], stage0_9[421], stage0_9[422], stage0_9[423], stage0_9[424], stage0_9[425]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[74],stage1_11[106],stage1_10[144],stage1_9[188]}
   );
   gpc606_5 gpc430 (
      {stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429], stage0_9[430], stage0_9[431]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[75],stage1_11[107],stage1_10[145],stage1_9[189]}
   );
   gpc606_5 gpc431 (
      {stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435], stage0_9[436], stage0_9[437]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[76],stage1_11[108],stage1_10[146],stage1_9[190]}
   );
   gpc606_5 gpc432 (
      {stage0_9[438], stage0_9[439], stage0_9[440], stage0_9[441], stage0_9[442], stage0_9[443]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[77],stage1_11[109],stage1_10[147],stage1_9[191]}
   );
   gpc606_5 gpc433 (
      {stage0_9[444], stage0_9[445], stage0_9[446], stage0_9[447], stage0_9[448], stage0_9[449]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[78],stage1_11[110],stage1_10[148],stage1_9[192]}
   );
   gpc606_5 gpc434 (
      {stage0_9[450], stage0_9[451], stage0_9[452], stage0_9[453], stage0_9[454], stage0_9[455]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[79],stage1_11[111],stage1_10[149],stage1_9[193]}
   );
   gpc606_5 gpc435 (
      {stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459], stage0_9[460], stage0_9[461]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[80],stage1_11[112],stage1_10[150],stage1_9[194]}
   );
   gpc606_5 gpc436 (
      {stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465], stage0_9[466], stage0_9[467]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[81],stage1_11[113],stage1_10[151],stage1_9[195]}
   );
   gpc2135_5 gpc437 (
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220]},
      {stage0_11[276], stage0_11[277], stage0_11[278]},
      {stage0_12[0]},
      {stage0_13[0], stage0_13[1]},
      {stage1_14[0],stage1_13[46],stage1_12[82],stage1_11[114],stage1_10[152]}
   );
   gpc2135_5 gpc438 (
      {stage0_10[221], stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225]},
      {stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage0_12[1]},
      {stage0_13[2], stage0_13[3]},
      {stage1_14[1],stage1_13[47],stage1_12[83],stage1_11[115],stage1_10[153]}
   );
   gpc2135_5 gpc439 (
      {stage0_10[226], stage0_10[227], stage0_10[228], stage0_10[229], stage0_10[230]},
      {stage0_11[282], stage0_11[283], stage0_11[284]},
      {stage0_12[2]},
      {stage0_13[4], stage0_13[5]},
      {stage1_14[2],stage1_13[48],stage1_12[84],stage1_11[116],stage1_10[154]}
   );
   gpc2135_5 gpc440 (
      {stage0_10[231], stage0_10[232], stage0_10[233], stage0_10[234], stage0_10[235]},
      {stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage0_12[3]},
      {stage0_13[6], stage0_13[7]},
      {stage1_14[3],stage1_13[49],stage1_12[85],stage1_11[117],stage1_10[155]}
   );
   gpc606_5 gpc441 (
      {stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239], stage0_10[240], stage0_10[241]},
      {stage0_12[4], stage0_12[5], stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9]},
      {stage1_14[4],stage1_13[50],stage1_12[86],stage1_11[118],stage1_10[156]}
   );
   gpc606_5 gpc442 (
      {stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245], stage0_10[246], stage0_10[247]},
      {stage0_12[10], stage0_12[11], stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15]},
      {stage1_14[5],stage1_13[51],stage1_12[87],stage1_11[119],stage1_10[157]}
   );
   gpc606_5 gpc443 (
      {stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251], stage0_10[252], stage0_10[253]},
      {stage0_12[16], stage0_12[17], stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21]},
      {stage1_14[6],stage1_13[52],stage1_12[88],stage1_11[120],stage1_10[158]}
   );
   gpc606_5 gpc444 (
      {stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257], stage0_10[258], stage0_10[259]},
      {stage0_12[22], stage0_12[23], stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27]},
      {stage1_14[7],stage1_13[53],stage1_12[89],stage1_11[121],stage1_10[159]}
   );
   gpc606_5 gpc445 (
      {stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263], stage0_10[264], stage0_10[265]},
      {stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33]},
      {stage1_14[8],stage1_13[54],stage1_12[90],stage1_11[122],stage1_10[160]}
   );
   gpc606_5 gpc446 (
      {stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269], stage0_10[270], stage0_10[271]},
      {stage0_12[34], stage0_12[35], stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39]},
      {stage1_14[9],stage1_13[55],stage1_12[91],stage1_11[123],stage1_10[161]}
   );
   gpc606_5 gpc447 (
      {stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275], stage0_10[276], stage0_10[277]},
      {stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45]},
      {stage1_14[10],stage1_13[56],stage1_12[92],stage1_11[124],stage1_10[162]}
   );
   gpc606_5 gpc448 (
      {stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281], stage0_10[282], stage0_10[283]},
      {stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51]},
      {stage1_14[11],stage1_13[57],stage1_12[93],stage1_11[125],stage1_10[163]}
   );
   gpc606_5 gpc449 (
      {stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287], stage0_10[288], stage0_10[289]},
      {stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57]},
      {stage1_14[12],stage1_13[58],stage1_12[94],stage1_11[126],stage1_10[164]}
   );
   gpc606_5 gpc450 (
      {stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293], stage0_10[294], stage0_10[295]},
      {stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63]},
      {stage1_14[13],stage1_13[59],stage1_12[95],stage1_11[127],stage1_10[165]}
   );
   gpc606_5 gpc451 (
      {stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299], stage0_10[300], stage0_10[301]},
      {stage0_12[64], stage0_12[65], stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69]},
      {stage1_14[14],stage1_13[60],stage1_12[96],stage1_11[128],stage1_10[166]}
   );
   gpc606_5 gpc452 (
      {stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305], stage0_10[306], stage0_10[307]},
      {stage0_12[70], stage0_12[71], stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75]},
      {stage1_14[15],stage1_13[61],stage1_12[97],stage1_11[129],stage1_10[167]}
   );
   gpc606_5 gpc453 (
      {stage0_10[308], stage0_10[309], stage0_10[310], stage0_10[311], stage0_10[312], stage0_10[313]},
      {stage0_12[76], stage0_12[77], stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81]},
      {stage1_14[16],stage1_13[62],stage1_12[98],stage1_11[130],stage1_10[168]}
   );
   gpc615_5 gpc454 (
      {stage0_10[314], stage0_10[315], stage0_10[316], stage0_10[317], stage0_10[318]},
      {stage0_11[288]},
      {stage0_12[82], stage0_12[83], stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87]},
      {stage1_14[17],stage1_13[63],stage1_12[99],stage1_11[131],stage1_10[169]}
   );
   gpc615_5 gpc455 (
      {stage0_10[319], stage0_10[320], stage0_10[321], stage0_10[322], stage0_10[323]},
      {stage0_11[289]},
      {stage0_12[88], stage0_12[89], stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93]},
      {stage1_14[18],stage1_13[64],stage1_12[100],stage1_11[132],stage1_10[170]}
   );
   gpc615_5 gpc456 (
      {stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327], stage0_10[328]},
      {stage0_11[290]},
      {stage0_12[94], stage0_12[95], stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99]},
      {stage1_14[19],stage1_13[65],stage1_12[101],stage1_11[133],stage1_10[171]}
   );
   gpc615_5 gpc457 (
      {stage0_10[329], stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333]},
      {stage0_11[291]},
      {stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105]},
      {stage1_14[20],stage1_13[66],stage1_12[102],stage1_11[134],stage1_10[172]}
   );
   gpc615_5 gpc458 (
      {stage0_10[334], stage0_10[335], stage0_10[336], stage0_10[337], stage0_10[338]},
      {stage0_11[292]},
      {stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111]},
      {stage1_14[21],stage1_13[67],stage1_12[103],stage1_11[135],stage1_10[173]}
   );
   gpc615_5 gpc459 (
      {stage0_10[339], stage0_10[340], stage0_10[341], stage0_10[342], stage0_10[343]},
      {stage0_11[293]},
      {stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117]},
      {stage1_14[22],stage1_13[68],stage1_12[104],stage1_11[136],stage1_10[174]}
   );
   gpc615_5 gpc460 (
      {stage0_10[344], stage0_10[345], stage0_10[346], stage0_10[347], stage0_10[348]},
      {stage0_11[294]},
      {stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123]},
      {stage1_14[23],stage1_13[69],stage1_12[105],stage1_11[137],stage1_10[175]}
   );
   gpc615_5 gpc461 (
      {stage0_10[349], stage0_10[350], stage0_10[351], stage0_10[352], stage0_10[353]},
      {stage0_11[295]},
      {stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129]},
      {stage1_14[24],stage1_13[70],stage1_12[106],stage1_11[138],stage1_10[176]}
   );
   gpc615_5 gpc462 (
      {stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357], stage0_10[358]},
      {stage0_11[296]},
      {stage0_12[130], stage0_12[131], stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135]},
      {stage1_14[25],stage1_13[71],stage1_12[107],stage1_11[139],stage1_10[177]}
   );
   gpc615_5 gpc463 (
      {stage0_10[359], stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363]},
      {stage0_11[297]},
      {stage0_12[136], stage0_12[137], stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141]},
      {stage1_14[26],stage1_13[72],stage1_12[108],stage1_11[140],stage1_10[178]}
   );
   gpc615_5 gpc464 (
      {stage0_10[364], stage0_10[365], stage0_10[366], stage0_10[367], stage0_10[368]},
      {stage0_11[298]},
      {stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147]},
      {stage1_14[27],stage1_13[73],stage1_12[109],stage1_11[141],stage1_10[179]}
   );
   gpc615_5 gpc465 (
      {stage0_10[369], stage0_10[370], stage0_10[371], stage0_10[372], stage0_10[373]},
      {stage0_11[299]},
      {stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153]},
      {stage1_14[28],stage1_13[74],stage1_12[110],stage1_11[142],stage1_10[180]}
   );
   gpc615_5 gpc466 (
      {stage0_10[374], stage0_10[375], stage0_10[376], stage0_10[377], stage0_10[378]},
      {stage0_11[300]},
      {stage0_12[154], stage0_12[155], stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159]},
      {stage1_14[29],stage1_13[75],stage1_12[111],stage1_11[143],stage1_10[181]}
   );
   gpc615_5 gpc467 (
      {stage0_10[379], stage0_10[380], stage0_10[381], stage0_10[382], stage0_10[383]},
      {stage0_11[301]},
      {stage0_12[160], stage0_12[161], stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165]},
      {stage1_14[30],stage1_13[76],stage1_12[112],stage1_11[144],stage1_10[182]}
   );
   gpc615_5 gpc468 (
      {stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305], stage0_11[306]},
      {stage0_12[166]},
      {stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11], stage0_13[12], stage0_13[13]},
      {stage1_15[0],stage1_14[31],stage1_13[77],stage1_12[113],stage1_11[145]}
   );
   gpc615_5 gpc469 (
      {stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage0_12[167]},
      {stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17], stage0_13[18], stage0_13[19]},
      {stage1_15[1],stage1_14[32],stage1_13[78],stage1_12[114],stage1_11[146]}
   );
   gpc615_5 gpc470 (
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316]},
      {stage0_12[168]},
      {stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23], stage0_13[24], stage0_13[25]},
      {stage1_15[2],stage1_14[33],stage1_13[79],stage1_12[115],stage1_11[147]}
   );
   gpc615_5 gpc471 (
      {stage0_11[317], stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321]},
      {stage0_12[169]},
      {stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29], stage0_13[30], stage0_13[31]},
      {stage1_15[3],stage1_14[34],stage1_13[80],stage1_12[116],stage1_11[148]}
   );
   gpc615_5 gpc472 (
      {stage0_11[322], stage0_11[323], stage0_11[324], stage0_11[325], stage0_11[326]},
      {stage0_12[170]},
      {stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35], stage0_13[36], stage0_13[37]},
      {stage1_15[4],stage1_14[35],stage1_13[81],stage1_12[117],stage1_11[149]}
   );
   gpc615_5 gpc473 (
      {stage0_11[327], stage0_11[328], stage0_11[329], stage0_11[330], stage0_11[331]},
      {stage0_12[171]},
      {stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41], stage0_13[42], stage0_13[43]},
      {stage1_15[5],stage1_14[36],stage1_13[82],stage1_12[118],stage1_11[150]}
   );
   gpc615_5 gpc474 (
      {stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335], stage0_11[336]},
      {stage0_12[172]},
      {stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47], stage0_13[48], stage0_13[49]},
      {stage1_15[6],stage1_14[37],stage1_13[83],stage1_12[119],stage1_11[151]}
   );
   gpc615_5 gpc475 (
      {stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage0_12[173]},
      {stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53], stage0_13[54], stage0_13[55]},
      {stage1_15[7],stage1_14[38],stage1_13[84],stage1_12[120],stage1_11[152]}
   );
   gpc615_5 gpc476 (
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346]},
      {stage0_12[174]},
      {stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61]},
      {stage1_15[8],stage1_14[39],stage1_13[85],stage1_12[121],stage1_11[153]}
   );
   gpc615_5 gpc477 (
      {stage0_11[347], stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351]},
      {stage0_12[175]},
      {stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65], stage0_13[66], stage0_13[67]},
      {stage1_15[9],stage1_14[40],stage1_13[86],stage1_12[122],stage1_11[154]}
   );
   gpc615_5 gpc478 (
      {stage0_11[352], stage0_11[353], stage0_11[354], stage0_11[355], stage0_11[356]},
      {stage0_12[176]},
      {stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71], stage0_13[72], stage0_13[73]},
      {stage1_15[10],stage1_14[41],stage1_13[87],stage1_12[123],stage1_11[155]}
   );
   gpc615_5 gpc479 (
      {stage0_11[357], stage0_11[358], stage0_11[359], stage0_11[360], stage0_11[361]},
      {stage0_12[177]},
      {stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77], stage0_13[78], stage0_13[79]},
      {stage1_15[11],stage1_14[42],stage1_13[88],stage1_12[124],stage1_11[156]}
   );
   gpc615_5 gpc480 (
      {stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365], stage0_11[366]},
      {stage0_12[178]},
      {stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85]},
      {stage1_15[12],stage1_14[43],stage1_13[89],stage1_12[125],stage1_11[157]}
   );
   gpc615_5 gpc481 (
      {stage0_12[179], stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183]},
      {stage0_13[86]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[13],stage1_14[44],stage1_13[90],stage1_12[126]}
   );
   gpc615_5 gpc482 (
      {stage0_12[184], stage0_12[185], stage0_12[186], stage0_12[187], stage0_12[188]},
      {stage0_13[87]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[14],stage1_14[45],stage1_13[91],stage1_12[127]}
   );
   gpc615_5 gpc483 (
      {stage0_12[189], stage0_12[190], stage0_12[191], stage0_12[192], stage0_12[193]},
      {stage0_13[88]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[15],stage1_14[46],stage1_13[92],stage1_12[128]}
   );
   gpc615_5 gpc484 (
      {stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197], stage0_12[198]},
      {stage0_13[89]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[16],stage1_14[47],stage1_13[93],stage1_12[129]}
   );
   gpc615_5 gpc485 (
      {stage0_12[199], stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203]},
      {stage0_13[90]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[17],stage1_14[48],stage1_13[94],stage1_12[130]}
   );
   gpc615_5 gpc486 (
      {stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208]},
      {stage0_13[91]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[18],stage1_14[49],stage1_13[95],stage1_12[131]}
   );
   gpc615_5 gpc487 (
      {stage0_12[209], stage0_12[210], stage0_12[211], stage0_12[212], stage0_12[213]},
      {stage0_13[92]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[19],stage1_14[50],stage1_13[96],stage1_12[132]}
   );
   gpc615_5 gpc488 (
      {stage0_12[214], stage0_12[215], stage0_12[216], stage0_12[217], stage0_12[218]},
      {stage0_13[93]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[20],stage1_14[51],stage1_13[97],stage1_12[133]}
   );
   gpc615_5 gpc489 (
      {stage0_12[219], stage0_12[220], stage0_12[221], stage0_12[222], stage0_12[223]},
      {stage0_13[94]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[21],stage1_14[52],stage1_13[98],stage1_12[134]}
   );
   gpc615_5 gpc490 (
      {stage0_12[224], stage0_12[225], stage0_12[226], stage0_12[227], stage0_12[228]},
      {stage0_13[95]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[22],stage1_14[53],stage1_13[99],stage1_12[135]}
   );
   gpc615_5 gpc491 (
      {stage0_12[229], stage0_12[230], stage0_12[231], stage0_12[232], stage0_12[233]},
      {stage0_13[96]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[23],stage1_14[54],stage1_13[100],stage1_12[136]}
   );
   gpc615_5 gpc492 (
      {stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237], stage0_12[238]},
      {stage0_13[97]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[24],stage1_14[55],stage1_13[101],stage1_12[137]}
   );
   gpc615_5 gpc493 (
      {stage0_12[239], stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243]},
      {stage0_13[98]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[25],stage1_14[56],stage1_13[102],stage1_12[138]}
   );
   gpc615_5 gpc494 (
      {stage0_12[244], stage0_12[245], stage0_12[246], stage0_12[247], stage0_12[248]},
      {stage0_13[99]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[26],stage1_14[57],stage1_13[103],stage1_12[139]}
   );
   gpc615_5 gpc495 (
      {stage0_12[249], stage0_12[250], stage0_12[251], stage0_12[252], stage0_12[253]},
      {stage0_13[100]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[27],stage1_14[58],stage1_13[104],stage1_12[140]}
   );
   gpc615_5 gpc496 (
      {stage0_12[254], stage0_12[255], stage0_12[256], stage0_12[257], stage0_12[258]},
      {stage0_13[101]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[28],stage1_14[59],stage1_13[105],stage1_12[141]}
   );
   gpc615_5 gpc497 (
      {stage0_12[259], stage0_12[260], stage0_12[261], stage0_12[262], stage0_12[263]},
      {stage0_13[102]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[29],stage1_14[60],stage1_13[106],stage1_12[142]}
   );
   gpc615_5 gpc498 (
      {stage0_12[264], stage0_12[265], stage0_12[266], stage0_12[267], stage0_12[268]},
      {stage0_13[103]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[30],stage1_14[61],stage1_13[107],stage1_12[143]}
   );
   gpc615_5 gpc499 (
      {stage0_12[269], stage0_12[270], stage0_12[271], stage0_12[272], stage0_12[273]},
      {stage0_13[104]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[31],stage1_14[62],stage1_13[108],stage1_12[144]}
   );
   gpc615_5 gpc500 (
      {stage0_12[274], stage0_12[275], stage0_12[276], stage0_12[277], stage0_12[278]},
      {stage0_13[105]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[32],stage1_14[63],stage1_13[109],stage1_12[145]}
   );
   gpc615_5 gpc501 (
      {stage0_12[279], stage0_12[280], stage0_12[281], stage0_12[282], stage0_12[283]},
      {stage0_13[106]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[33],stage1_14[64],stage1_13[110],stage1_12[146]}
   );
   gpc615_5 gpc502 (
      {stage0_12[284], stage0_12[285], stage0_12[286], stage0_12[287], stage0_12[288]},
      {stage0_13[107]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[34],stage1_14[65],stage1_13[111],stage1_12[147]}
   );
   gpc615_5 gpc503 (
      {stage0_12[289], stage0_12[290], stage0_12[291], stage0_12[292], stage0_12[293]},
      {stage0_13[108]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[35],stage1_14[66],stage1_13[112],stage1_12[148]}
   );
   gpc615_5 gpc504 (
      {stage0_12[294], stage0_12[295], stage0_12[296], stage0_12[297], stage0_12[298]},
      {stage0_13[109]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[36],stage1_14[67],stage1_13[113],stage1_12[149]}
   );
   gpc615_5 gpc505 (
      {stage0_12[299], stage0_12[300], stage0_12[301], stage0_12[302], stage0_12[303]},
      {stage0_13[110]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[37],stage1_14[68],stage1_13[114],stage1_12[150]}
   );
   gpc615_5 gpc506 (
      {stage0_12[304], stage0_12[305], stage0_12[306], stage0_12[307], stage0_12[308]},
      {stage0_13[111]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[38],stage1_14[69],stage1_13[115],stage1_12[151]}
   );
   gpc615_5 gpc507 (
      {stage0_12[309], stage0_12[310], stage0_12[311], stage0_12[312], stage0_12[313]},
      {stage0_13[112]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[39],stage1_14[70],stage1_13[116],stage1_12[152]}
   );
   gpc615_5 gpc508 (
      {stage0_12[314], stage0_12[315], stage0_12[316], stage0_12[317], stage0_12[318]},
      {stage0_13[113]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[40],stage1_14[71],stage1_13[117],stage1_12[153]}
   );
   gpc615_5 gpc509 (
      {stage0_12[319], stage0_12[320], stage0_12[321], stage0_12[322], stage0_12[323]},
      {stage0_13[114]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[41],stage1_14[72],stage1_13[118],stage1_12[154]}
   );
   gpc615_5 gpc510 (
      {stage0_12[324], stage0_12[325], stage0_12[326], stage0_12[327], stage0_12[328]},
      {stage0_13[115]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[42],stage1_14[73],stage1_13[119],stage1_12[155]}
   );
   gpc615_5 gpc511 (
      {stage0_12[329], stage0_12[330], stage0_12[331], stage0_12[332], stage0_12[333]},
      {stage0_13[116]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[43],stage1_14[74],stage1_13[120],stage1_12[156]}
   );
   gpc615_5 gpc512 (
      {stage0_12[334], stage0_12[335], stage0_12[336], stage0_12[337], stage0_12[338]},
      {stage0_13[117]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[44],stage1_14[75],stage1_13[121],stage1_12[157]}
   );
   gpc615_5 gpc513 (
      {stage0_12[339], stage0_12[340], stage0_12[341], stage0_12[342], stage0_12[343]},
      {stage0_13[118]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[45],stage1_14[76],stage1_13[122],stage1_12[158]}
   );
   gpc615_5 gpc514 (
      {stage0_12[344], stage0_12[345], stage0_12[346], stage0_12[347], stage0_12[348]},
      {stage0_13[119]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[46],stage1_14[77],stage1_13[123],stage1_12[159]}
   );
   gpc615_5 gpc515 (
      {stage0_12[349], stage0_12[350], stage0_12[351], stage0_12[352], stage0_12[353]},
      {stage0_13[120]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[47],stage1_14[78],stage1_13[124],stage1_12[160]}
   );
   gpc615_5 gpc516 (
      {stage0_12[354], stage0_12[355], stage0_12[356], stage0_12[357], stage0_12[358]},
      {stage0_13[121]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[48],stage1_14[79],stage1_13[125],stage1_12[161]}
   );
   gpc615_5 gpc517 (
      {stage0_12[359], stage0_12[360], stage0_12[361], stage0_12[362], stage0_12[363]},
      {stage0_13[122]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[49],stage1_14[80],stage1_13[126],stage1_12[162]}
   );
   gpc615_5 gpc518 (
      {stage0_12[364], stage0_12[365], stage0_12[366], stage0_12[367], stage0_12[368]},
      {stage0_13[123]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[50],stage1_14[81],stage1_13[127],stage1_12[163]}
   );
   gpc615_5 gpc519 (
      {stage0_12[369], stage0_12[370], stage0_12[371], stage0_12[372], stage0_12[373]},
      {stage0_13[124]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[51],stage1_14[82],stage1_13[128],stage1_12[164]}
   );
   gpc615_5 gpc520 (
      {stage0_12[374], stage0_12[375], stage0_12[376], stage0_12[377], stage0_12[378]},
      {stage0_13[125]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[52],stage1_14[83],stage1_13[129],stage1_12[165]}
   );
   gpc615_5 gpc521 (
      {stage0_12[379], stage0_12[380], stage0_12[381], stage0_12[382], stage0_12[383]},
      {stage0_13[126]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[53],stage1_14[84],stage1_13[130],stage1_12[166]}
   );
   gpc615_5 gpc522 (
      {stage0_12[384], stage0_12[385], stage0_12[386], stage0_12[387], stage0_12[388]},
      {stage0_13[127]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[54],stage1_14[85],stage1_13[131],stage1_12[167]}
   );
   gpc615_5 gpc523 (
      {stage0_12[389], stage0_12[390], stage0_12[391], stage0_12[392], stage0_12[393]},
      {stage0_13[128]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[55],stage1_14[86],stage1_13[132],stage1_12[168]}
   );
   gpc615_5 gpc524 (
      {stage0_12[394], stage0_12[395], stage0_12[396], stage0_12[397], stage0_12[398]},
      {stage0_13[129]},
      {stage0_14[258], stage0_14[259], stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263]},
      {stage1_16[43],stage1_15[56],stage1_14[87],stage1_13[133],stage1_12[169]}
   );
   gpc615_5 gpc525 (
      {stage0_12[399], stage0_12[400], stage0_12[401], stage0_12[402], stage0_12[403]},
      {stage0_13[130]},
      {stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269]},
      {stage1_16[44],stage1_15[57],stage1_14[88],stage1_13[134],stage1_12[170]}
   );
   gpc615_5 gpc526 (
      {stage0_12[404], stage0_12[405], stage0_12[406], stage0_12[407], stage0_12[408]},
      {stage0_13[131]},
      {stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275]},
      {stage1_16[45],stage1_15[58],stage1_14[89],stage1_13[135],stage1_12[171]}
   );
   gpc615_5 gpc527 (
      {stage0_12[409], stage0_12[410], stage0_12[411], stage0_12[412], stage0_12[413]},
      {stage0_13[132]},
      {stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281]},
      {stage1_16[46],stage1_15[59],stage1_14[90],stage1_13[136],stage1_12[172]}
   );
   gpc615_5 gpc528 (
      {stage0_12[414], stage0_12[415], stage0_12[416], stage0_12[417], stage0_12[418]},
      {stage0_13[133]},
      {stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287]},
      {stage1_16[47],stage1_15[60],stage1_14[91],stage1_13[137],stage1_12[173]}
   );
   gpc615_5 gpc529 (
      {stage0_12[419], stage0_12[420], stage0_12[421], stage0_12[422], stage0_12[423]},
      {stage0_13[134]},
      {stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293]},
      {stage1_16[48],stage1_15[61],stage1_14[92],stage1_13[138],stage1_12[174]}
   );
   gpc615_5 gpc530 (
      {stage0_12[424], stage0_12[425], stage0_12[426], stage0_12[427], stage0_12[428]},
      {stage0_13[135]},
      {stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299]},
      {stage1_16[49],stage1_15[62],stage1_14[93],stage1_13[139],stage1_12[175]}
   );
   gpc615_5 gpc531 (
      {stage0_12[429], stage0_12[430], stage0_12[431], stage0_12[432], stage0_12[433]},
      {stage0_13[136]},
      {stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305]},
      {stage1_16[50],stage1_15[63],stage1_14[94],stage1_13[140],stage1_12[176]}
   );
   gpc615_5 gpc532 (
      {stage0_12[434], stage0_12[435], stage0_12[436], stage0_12[437], stage0_12[438]},
      {stage0_13[137]},
      {stage0_14[306], stage0_14[307], stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311]},
      {stage1_16[51],stage1_15[64],stage1_14[95],stage1_13[141],stage1_12[177]}
   );
   gpc615_5 gpc533 (
      {stage0_12[439], stage0_12[440], stage0_12[441], stage0_12[442], stage0_12[443]},
      {stage0_13[138]},
      {stage0_14[312], stage0_14[313], stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317]},
      {stage1_16[52],stage1_15[65],stage1_14[96],stage1_13[142],stage1_12[178]}
   );
   gpc615_5 gpc534 (
      {stage0_12[444], stage0_12[445], stage0_12[446], stage0_12[447], stage0_12[448]},
      {stage0_13[139]},
      {stage0_14[318], stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage1_16[53],stage1_15[66],stage1_14[97],stage1_13[143],stage1_12[179]}
   );
   gpc615_5 gpc535 (
      {stage0_12[449], stage0_12[450], stage0_12[451], stage0_12[452], stage0_12[453]},
      {stage0_13[140]},
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329]},
      {stage1_16[54],stage1_15[67],stage1_14[98],stage1_13[144],stage1_12[180]}
   );
   gpc615_5 gpc536 (
      {stage0_12[454], stage0_12[455], stage0_12[456], stage0_12[457], stage0_12[458]},
      {stage0_13[141]},
      {stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335]},
      {stage1_16[55],stage1_15[68],stage1_14[99],stage1_13[145],stage1_12[181]}
   );
   gpc615_5 gpc537 (
      {stage0_12[459], stage0_12[460], stage0_12[461], stage0_12[462], stage0_12[463]},
      {stage0_13[142]},
      {stage0_14[336], stage0_14[337], stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341]},
      {stage1_16[56],stage1_15[69],stage1_14[100],stage1_13[146],stage1_12[182]}
   );
   gpc615_5 gpc538 (
      {stage0_12[464], stage0_12[465], stage0_12[466], stage0_12[467], stage0_12[468]},
      {stage0_13[143]},
      {stage0_14[342], stage0_14[343], stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347]},
      {stage1_16[57],stage1_15[70],stage1_14[101],stage1_13[147],stage1_12[183]}
   );
   gpc615_5 gpc539 (
      {stage0_12[469], stage0_12[470], stage0_12[471], stage0_12[472], stage0_12[473]},
      {stage0_13[144]},
      {stage0_14[348], stage0_14[349], stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353]},
      {stage1_16[58],stage1_15[71],stage1_14[102],stage1_13[148],stage1_12[184]}
   );
   gpc615_5 gpc540 (
      {stage0_12[474], stage0_12[475], stage0_12[476], stage0_12[477], stage0_12[478]},
      {stage0_13[145]},
      {stage0_14[354], stage0_14[355], stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359]},
      {stage1_16[59],stage1_15[72],stage1_14[103],stage1_13[149],stage1_12[185]}
   );
   gpc615_5 gpc541 (
      {stage0_12[479], stage0_12[480], stage0_12[481], stage0_12[482], stage0_12[483]},
      {stage0_13[146]},
      {stage0_14[360], stage0_14[361], stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365]},
      {stage1_16[60],stage1_15[73],stage1_14[104],stage1_13[150],stage1_12[186]}
   );
   gpc606_5 gpc542 (
      {stage0_13[147], stage0_13[148], stage0_13[149], stage0_13[150], stage0_13[151], stage0_13[152]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[61],stage1_15[74],stage1_14[105],stage1_13[151]}
   );
   gpc606_5 gpc543 (
      {stage0_13[153], stage0_13[154], stage0_13[155], stage0_13[156], stage0_13[157], stage0_13[158]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[62],stage1_15[75],stage1_14[106],stage1_13[152]}
   );
   gpc606_5 gpc544 (
      {stage0_13[159], stage0_13[160], stage0_13[161], stage0_13[162], stage0_13[163], stage0_13[164]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[63],stage1_15[76],stage1_14[107],stage1_13[153]}
   );
   gpc606_5 gpc545 (
      {stage0_13[165], stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169], stage0_13[170]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[64],stage1_15[77],stage1_14[108],stage1_13[154]}
   );
   gpc606_5 gpc546 (
      {stage0_13[171], stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175], stage0_13[176]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[65],stage1_15[78],stage1_14[109],stage1_13[155]}
   );
   gpc606_5 gpc547 (
      {stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181], stage0_13[182]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[66],stage1_15[79],stage1_14[110],stage1_13[156]}
   );
   gpc606_5 gpc548 (
      {stage0_13[183], stage0_13[184], stage0_13[185], stage0_13[186], stage0_13[187], stage0_13[188]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[67],stage1_15[80],stage1_14[111],stage1_13[157]}
   );
   gpc606_5 gpc549 (
      {stage0_13[189], stage0_13[190], stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[68],stage1_15[81],stage1_14[112],stage1_13[158]}
   );
   gpc606_5 gpc550 (
      {stage0_13[195], stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[69],stage1_15[82],stage1_14[113],stage1_13[159]}
   );
   gpc615_5 gpc551 (
      {stage0_13[201], stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205]},
      {stage0_14[366]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[70],stage1_15[83],stage1_14[114],stage1_13[160]}
   );
   gpc615_5 gpc552 (
      {stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210]},
      {stage0_14[367]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[71],stage1_15[84],stage1_14[115],stage1_13[161]}
   );
   gpc615_5 gpc553 (
      {stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215]},
      {stage0_14[368]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[72],stage1_15[85],stage1_14[116],stage1_13[162]}
   );
   gpc615_5 gpc554 (
      {stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220]},
      {stage0_14[369]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[73],stage1_15[86],stage1_14[117],stage1_13[163]}
   );
   gpc615_5 gpc555 (
      {stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225]},
      {stage0_14[370]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[74],stage1_15[87],stage1_14[118],stage1_13[164]}
   );
   gpc615_5 gpc556 (
      {stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230]},
      {stage0_14[371]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[75],stage1_15[88],stage1_14[119],stage1_13[165]}
   );
   gpc615_5 gpc557 (
      {stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235]},
      {stage0_14[372]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[76],stage1_15[89],stage1_14[120],stage1_13[166]}
   );
   gpc615_5 gpc558 (
      {stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240]},
      {stage0_14[373]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[77],stage1_15[90],stage1_14[121],stage1_13[167]}
   );
   gpc615_5 gpc559 (
      {stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage0_14[374]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[78],stage1_15[91],stage1_14[122],stage1_13[168]}
   );
   gpc615_5 gpc560 (
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250]},
      {stage0_14[375]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[79],stage1_15[92],stage1_14[123],stage1_13[169]}
   );
   gpc615_5 gpc561 (
      {stage0_13[251], stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255]},
      {stage0_14[376]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[80],stage1_15[93],stage1_14[124],stage1_13[170]}
   );
   gpc615_5 gpc562 (
      {stage0_13[256], stage0_13[257], stage0_13[258], stage0_13[259], stage0_13[260]},
      {stage0_14[377]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[81],stage1_15[94],stage1_14[125],stage1_13[171]}
   );
   gpc615_5 gpc563 (
      {stage0_13[261], stage0_13[262], stage0_13[263], stage0_13[264], stage0_13[265]},
      {stage0_14[378]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[82],stage1_15[95],stage1_14[126],stage1_13[172]}
   );
   gpc615_5 gpc564 (
      {stage0_13[266], stage0_13[267], stage0_13[268], stage0_13[269], stage0_13[270]},
      {stage0_14[379]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[83],stage1_15[96],stage1_14[127],stage1_13[173]}
   );
   gpc615_5 gpc565 (
      {stage0_13[271], stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275]},
      {stage0_14[380]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[84],stage1_15[97],stage1_14[128],stage1_13[174]}
   );
   gpc615_5 gpc566 (
      {stage0_13[276], stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280]},
      {stage0_14[381]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[85],stage1_15[98],stage1_14[129],stage1_13[175]}
   );
   gpc615_5 gpc567 (
      {stage0_13[281], stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285]},
      {stage0_14[382]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[86],stage1_15[99],stage1_14[130],stage1_13[176]}
   );
   gpc615_5 gpc568 (
      {stage0_13[286], stage0_13[287], stage0_13[288], stage0_13[289], stage0_13[290]},
      {stage0_14[383]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[87],stage1_15[100],stage1_14[131],stage1_13[177]}
   );
   gpc615_5 gpc569 (
      {stage0_13[291], stage0_13[292], stage0_13[293], stage0_13[294], stage0_13[295]},
      {stage0_14[384]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[88],stage1_15[101],stage1_14[132],stage1_13[178]}
   );
   gpc615_5 gpc570 (
      {stage0_13[296], stage0_13[297], stage0_13[298], stage0_13[299], stage0_13[300]},
      {stage0_14[385]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[89],stage1_15[102],stage1_14[133],stage1_13[179]}
   );
   gpc615_5 gpc571 (
      {stage0_13[301], stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305]},
      {stage0_14[386]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[90],stage1_15[103],stage1_14[134],stage1_13[180]}
   );
   gpc615_5 gpc572 (
      {stage0_13[306], stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310]},
      {stage0_14[387]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[91],stage1_15[104],stage1_14[135],stage1_13[181]}
   );
   gpc615_5 gpc573 (
      {stage0_13[311], stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315]},
      {stage0_14[388]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[92],stage1_15[105],stage1_14[136],stage1_13[182]}
   );
   gpc615_5 gpc574 (
      {stage0_13[316], stage0_13[317], stage0_13[318], stage0_13[319], stage0_13[320]},
      {stage0_14[389]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[93],stage1_15[106],stage1_14[137],stage1_13[183]}
   );
   gpc615_5 gpc575 (
      {stage0_13[321], stage0_13[322], stage0_13[323], stage0_13[324], stage0_13[325]},
      {stage0_14[390]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[94],stage1_15[107],stage1_14[138],stage1_13[184]}
   );
   gpc615_5 gpc576 (
      {stage0_13[326], stage0_13[327], stage0_13[328], stage0_13[329], stage0_13[330]},
      {stage0_14[391]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[95],stage1_15[108],stage1_14[139],stage1_13[185]}
   );
   gpc615_5 gpc577 (
      {stage0_13[331], stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335]},
      {stage0_14[392]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[96],stage1_15[109],stage1_14[140],stage1_13[186]}
   );
   gpc615_5 gpc578 (
      {stage0_13[336], stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340]},
      {stage0_14[393]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[97],stage1_15[110],stage1_14[141],stage1_13[187]}
   );
   gpc615_5 gpc579 (
      {stage0_13[341], stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345]},
      {stage0_14[394]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[98],stage1_15[111],stage1_14[142],stage1_13[188]}
   );
   gpc615_5 gpc580 (
      {stage0_13[346], stage0_13[347], stage0_13[348], stage0_13[349], stage0_13[350]},
      {stage0_14[395]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[99],stage1_15[112],stage1_14[143],stage1_13[189]}
   );
   gpc615_5 gpc581 (
      {stage0_13[351], stage0_13[352], stage0_13[353], stage0_13[354], stage0_13[355]},
      {stage0_14[396]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[100],stage1_15[113],stage1_14[144],stage1_13[190]}
   );
   gpc615_5 gpc582 (
      {stage0_13[356], stage0_13[357], stage0_13[358], stage0_13[359], stage0_13[360]},
      {stage0_14[397]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[101],stage1_15[114],stage1_14[145],stage1_13[191]}
   );
   gpc615_5 gpc583 (
      {stage0_13[361], stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365]},
      {stage0_14[398]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[102],stage1_15[115],stage1_14[146],stage1_13[192]}
   );
   gpc615_5 gpc584 (
      {stage0_13[366], stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370]},
      {stage0_14[399]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[103],stage1_15[116],stage1_14[147],stage1_13[193]}
   );
   gpc615_5 gpc585 (
      {stage0_13[371], stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375]},
      {stage0_14[400]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[104],stage1_15[117],stage1_14[148],stage1_13[194]}
   );
   gpc606_5 gpc586 (
      {stage0_14[401], stage0_14[402], stage0_14[403], stage0_14[404], stage0_14[405], stage0_14[406]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[44],stage1_16[105],stage1_15[118],stage1_14[149]}
   );
   gpc606_5 gpc587 (
      {stage0_14[407], stage0_14[408], stage0_14[409], stage0_14[410], stage0_14[411], stage0_14[412]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[45],stage1_16[106],stage1_15[119],stage1_14[150]}
   );
   gpc606_5 gpc588 (
      {stage0_14[413], stage0_14[414], stage0_14[415], stage0_14[416], stage0_14[417], stage0_14[418]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[46],stage1_16[107],stage1_15[120],stage1_14[151]}
   );
   gpc615_5 gpc589 (
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268]},
      {stage0_16[18]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[3],stage1_17[47],stage1_16[108],stage1_15[121]}
   );
   gpc615_5 gpc590 (
      {stage0_15[269], stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273]},
      {stage0_16[19]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[4],stage1_17[48],stage1_16[109],stage1_15[122]}
   );
   gpc615_5 gpc591 (
      {stage0_15[274], stage0_15[275], stage0_15[276], stage0_15[277], stage0_15[278]},
      {stage0_16[20]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[5],stage1_17[49],stage1_16[110],stage1_15[123]}
   );
   gpc615_5 gpc592 (
      {stage0_15[279], stage0_15[280], stage0_15[281], stage0_15[282], stage0_15[283]},
      {stage0_16[21]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[6],stage1_17[50],stage1_16[111],stage1_15[124]}
   );
   gpc615_5 gpc593 (
      {stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287], stage0_15[288]},
      {stage0_16[22]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[7],stage1_17[51],stage1_16[112],stage1_15[125]}
   );
   gpc615_5 gpc594 (
      {stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage0_16[23]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[8],stage1_17[52],stage1_16[113],stage1_15[126]}
   );
   gpc615_5 gpc595 (
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298]},
      {stage0_16[24]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[9],stage1_17[53],stage1_16[114],stage1_15[127]}
   );
   gpc615_5 gpc596 (
      {stage0_15[299], stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303]},
      {stage0_16[25]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[10],stage1_17[54],stage1_16[115],stage1_15[128]}
   );
   gpc615_5 gpc597 (
      {stage0_15[304], stage0_15[305], stage0_15[306], stage0_15[307], stage0_15[308]},
      {stage0_16[26]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[11],stage1_17[55],stage1_16[116],stage1_15[129]}
   );
   gpc615_5 gpc598 (
      {stage0_15[309], stage0_15[310], stage0_15[311], stage0_15[312], stage0_15[313]},
      {stage0_16[27]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[12],stage1_17[56],stage1_16[117],stage1_15[130]}
   );
   gpc615_5 gpc599 (
      {stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317], stage0_15[318]},
      {stage0_16[28]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[13],stage1_17[57],stage1_16[118],stage1_15[131]}
   );
   gpc615_5 gpc600 (
      {stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage0_16[29]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[14],stage1_17[58],stage1_16[119],stage1_15[132]}
   );
   gpc615_5 gpc601 (
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328]},
      {stage0_16[30]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[15],stage1_17[59],stage1_16[120],stage1_15[133]}
   );
   gpc615_5 gpc602 (
      {stage0_15[329], stage0_15[330], stage0_15[331], stage0_15[332], stage0_15[333]},
      {stage0_16[31]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[16],stage1_17[60],stage1_16[121],stage1_15[134]}
   );
   gpc615_5 gpc603 (
      {stage0_15[334], stage0_15[335], stage0_15[336], stage0_15[337], stage0_15[338]},
      {stage0_16[32]},
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage1_19[14],stage1_18[17],stage1_17[61],stage1_16[122],stage1_15[135]}
   );
   gpc615_5 gpc604 (
      {stage0_15[339], stage0_15[340], stage0_15[341], stage0_15[342], stage0_15[343]},
      {stage0_16[33]},
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage1_19[15],stage1_18[18],stage1_17[62],stage1_16[123],stage1_15[136]}
   );
   gpc615_5 gpc605 (
      {stage0_15[344], stage0_15[345], stage0_15[346], stage0_15[347], stage0_15[348]},
      {stage0_16[34]},
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage1_19[16],stage1_18[19],stage1_17[63],stage1_16[124],stage1_15[137]}
   );
   gpc615_5 gpc606 (
      {stage0_15[349], stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353]},
      {stage0_16[35]},
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage1_19[17],stage1_18[20],stage1_17[64],stage1_16[125],stage1_15[138]}
   );
   gpc615_5 gpc607 (
      {stage0_15[354], stage0_15[355], stage0_15[356], stage0_15[357], stage0_15[358]},
      {stage0_16[36]},
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage1_19[18],stage1_18[21],stage1_17[65],stage1_16[126],stage1_15[139]}
   );
   gpc615_5 gpc608 (
      {stage0_15[359], stage0_15[360], stage0_15[361], stage0_15[362], stage0_15[363]},
      {stage0_16[37]},
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage1_19[19],stage1_18[22],stage1_17[66],stage1_16[127],stage1_15[140]}
   );
   gpc615_5 gpc609 (
      {stage0_15[364], stage0_15[365], stage0_15[366], stage0_15[367], stage0_15[368]},
      {stage0_16[38]},
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage1_19[20],stage1_18[23],stage1_17[67],stage1_16[128],stage1_15[141]}
   );
   gpc615_5 gpc610 (
      {stage0_15[369], stage0_15[370], stage0_15[371], stage0_15[372], stage0_15[373]},
      {stage0_16[39]},
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage1_19[21],stage1_18[24],stage1_17[68],stage1_16[129],stage1_15[142]}
   );
   gpc615_5 gpc611 (
      {stage0_15[374], stage0_15[375], stage0_15[376], stage0_15[377], stage0_15[378]},
      {stage0_16[40]},
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage1_19[22],stage1_18[25],stage1_17[69],stage1_16[130],stage1_15[143]}
   );
   gpc615_5 gpc612 (
      {stage0_15[379], stage0_15[380], stage0_15[381], stage0_15[382], stage0_15[383]},
      {stage0_16[41]},
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage1_19[23],stage1_18[26],stage1_17[70],stage1_16[131],stage1_15[144]}
   );
   gpc615_5 gpc613 (
      {stage0_15[384], stage0_15[385], stage0_15[386], stage0_15[387], stage0_15[388]},
      {stage0_16[42]},
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage1_19[24],stage1_18[27],stage1_17[71],stage1_16[132],stage1_15[145]}
   );
   gpc615_5 gpc614 (
      {stage0_15[389], stage0_15[390], stage0_15[391], stage0_15[392], stage0_15[393]},
      {stage0_16[43]},
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage1_19[25],stage1_18[28],stage1_17[72],stage1_16[133],stage1_15[146]}
   );
   gpc615_5 gpc615 (
      {stage0_15[394], stage0_15[395], stage0_15[396], stage0_15[397], stage0_15[398]},
      {stage0_16[44]},
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage1_19[26],stage1_18[29],stage1_17[73],stage1_16[134],stage1_15[147]}
   );
   gpc615_5 gpc616 (
      {stage0_15[399], stage0_15[400], stage0_15[401], stage0_15[402], stage0_15[403]},
      {stage0_16[45]},
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166], stage0_17[167]},
      {stage1_19[27],stage1_18[30],stage1_17[74],stage1_16[135],stage1_15[148]}
   );
   gpc615_5 gpc617 (
      {stage0_15[404], stage0_15[405], stage0_15[406], stage0_15[407], stage0_15[408]},
      {stage0_16[46]},
      {stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172], stage0_17[173]},
      {stage1_19[28],stage1_18[31],stage1_17[75],stage1_16[136],stage1_15[149]}
   );
   gpc615_5 gpc618 (
      {stage0_15[409], stage0_15[410], stage0_15[411], stage0_15[412], stage0_15[413]},
      {stage0_16[47]},
      {stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178], stage0_17[179]},
      {stage1_19[29],stage1_18[32],stage1_17[76],stage1_16[137],stage1_15[150]}
   );
   gpc615_5 gpc619 (
      {stage0_15[414], stage0_15[415], stage0_15[416], stage0_15[417], stage0_15[418]},
      {stage0_16[48]},
      {stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185]},
      {stage1_19[30],stage1_18[33],stage1_17[77],stage1_16[138],stage1_15[151]}
   );
   gpc615_5 gpc620 (
      {stage0_15[419], stage0_15[420], stage0_15[421], stage0_15[422], stage0_15[423]},
      {stage0_16[49]},
      {stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage1_19[31],stage1_18[34],stage1_17[78],stage1_16[139],stage1_15[152]}
   );
   gpc615_5 gpc621 (
      {stage0_15[424], stage0_15[425], stage0_15[426], stage0_15[427], stage0_15[428]},
      {stage0_16[50]},
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196], stage0_17[197]},
      {stage1_19[32],stage1_18[35],stage1_17[79],stage1_16[140],stage1_15[153]}
   );
   gpc615_5 gpc622 (
      {stage0_15[429], stage0_15[430], stage0_15[431], stage0_15[432], stage0_15[433]},
      {stage0_16[51]},
      {stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202], stage0_17[203]},
      {stage1_19[33],stage1_18[36],stage1_17[80],stage1_16[141],stage1_15[154]}
   );
   gpc615_5 gpc623 (
      {stage0_15[434], stage0_15[435], stage0_15[436], stage0_15[437], stage0_15[438]},
      {stage0_16[52]},
      {stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208], stage0_17[209]},
      {stage1_19[34],stage1_18[37],stage1_17[81],stage1_16[142],stage1_15[155]}
   );
   gpc615_5 gpc624 (
      {stage0_15[439], stage0_15[440], stage0_15[441], stage0_15[442], stage0_15[443]},
      {stage0_16[53]},
      {stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215]},
      {stage1_19[35],stage1_18[38],stage1_17[82],stage1_16[143],stage1_15[156]}
   );
   gpc615_5 gpc625 (
      {stage0_15[444], stage0_15[445], stage0_15[446], stage0_15[447], stage0_15[448]},
      {stage0_16[54]},
      {stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage1_19[36],stage1_18[39],stage1_17[83],stage1_16[144],stage1_15[157]}
   );
   gpc615_5 gpc626 (
      {stage0_15[449], stage0_15[450], stage0_15[451], stage0_15[452], stage0_15[453]},
      {stage0_16[55]},
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226], stage0_17[227]},
      {stage1_19[37],stage1_18[40],stage1_17[84],stage1_16[145],stage1_15[158]}
   );
   gpc615_5 gpc627 (
      {stage0_15[454], stage0_15[455], stage0_15[456], stage0_15[457], stage0_15[458]},
      {stage0_16[56]},
      {stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232], stage0_17[233]},
      {stage1_19[38],stage1_18[41],stage1_17[85],stage1_16[146],stage1_15[159]}
   );
   gpc615_5 gpc628 (
      {stage0_15[459], stage0_15[460], stage0_15[461], stage0_15[462], stage0_15[463]},
      {stage0_16[57]},
      {stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238], stage0_17[239]},
      {stage1_19[39],stage1_18[42],stage1_17[86],stage1_16[147],stage1_15[160]}
   );
   gpc615_5 gpc629 (
      {stage0_15[464], stage0_15[465], stage0_15[466], stage0_15[467], stage0_15[468]},
      {stage0_16[58]},
      {stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245]},
      {stage1_19[40],stage1_18[43],stage1_17[87],stage1_16[148],stage1_15[161]}
   );
   gpc615_5 gpc630 (
      {stage0_15[469], stage0_15[470], stage0_15[471], stage0_15[472], stage0_15[473]},
      {stage0_16[59]},
      {stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage1_19[41],stage1_18[44],stage1_17[88],stage1_16[149],stage1_15[162]}
   );
   gpc615_5 gpc631 (
      {stage0_15[474], stage0_15[475], stage0_15[476], stage0_15[477], stage0_15[478]},
      {stage0_16[60]},
      {stage0_17[252], stage0_17[253], stage0_17[254], stage0_17[255], stage0_17[256], stage0_17[257]},
      {stage1_19[42],stage1_18[45],stage1_17[89],stage1_16[150],stage1_15[163]}
   );
   gpc606_5 gpc632 (
      {stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65], stage0_16[66]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[43],stage1_18[46],stage1_17[90],stage1_16[151]}
   );
   gpc606_5 gpc633 (
      {stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71], stage0_16[72]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[44],stage1_18[47],stage1_17[91],stage1_16[152]}
   );
   gpc606_5 gpc634 (
      {stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77], stage0_16[78]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[45],stage1_18[48],stage1_17[92],stage1_16[153]}
   );
   gpc606_5 gpc635 (
      {stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83], stage0_16[84]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[46],stage1_18[49],stage1_17[93],stage1_16[154]}
   );
   gpc606_5 gpc636 (
      {stage0_16[85], stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89], stage0_16[90]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[47],stage1_18[50],stage1_17[94],stage1_16[155]}
   );
   gpc606_5 gpc637 (
      {stage0_16[91], stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95], stage0_16[96]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[48],stage1_18[51],stage1_17[95],stage1_16[156]}
   );
   gpc606_5 gpc638 (
      {stage0_16[97], stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[49],stage1_18[52],stage1_17[96],stage1_16[157]}
   );
   gpc606_5 gpc639 (
      {stage0_16[103], stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[50],stage1_18[53],stage1_17[97],stage1_16[158]}
   );
   gpc606_5 gpc640 (
      {stage0_16[109], stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113], stage0_16[114]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[51],stage1_18[54],stage1_17[98],stage1_16[159]}
   );
   gpc606_5 gpc641 (
      {stage0_16[115], stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119], stage0_16[120]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[52],stage1_18[55],stage1_17[99],stage1_16[160]}
   );
   gpc606_5 gpc642 (
      {stage0_16[121], stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[53],stage1_18[56],stage1_17[100],stage1_16[161]}
   );
   gpc606_5 gpc643 (
      {stage0_16[127], stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[54],stage1_18[57],stage1_17[101],stage1_16[162]}
   );
   gpc606_5 gpc644 (
      {stage0_16[133], stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[55],stage1_18[58],stage1_17[102],stage1_16[163]}
   );
   gpc606_5 gpc645 (
      {stage0_16[139], stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[56],stage1_18[59],stage1_17[103],stage1_16[164]}
   );
   gpc606_5 gpc646 (
      {stage0_16[145], stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[57],stage1_18[60],stage1_17[104],stage1_16[165]}
   );
   gpc606_5 gpc647 (
      {stage0_16[151], stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[58],stage1_18[61],stage1_17[105],stage1_16[166]}
   );
   gpc606_5 gpc648 (
      {stage0_16[157], stage0_16[158], stage0_16[159], stage0_16[160], stage0_16[161], stage0_16[162]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[59],stage1_18[62],stage1_17[106],stage1_16[167]}
   );
   gpc606_5 gpc649 (
      {stage0_16[163], stage0_16[164], stage0_16[165], stage0_16[166], stage0_16[167], stage0_16[168]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[60],stage1_18[63],stage1_17[107],stage1_16[168]}
   );
   gpc606_5 gpc650 (
      {stage0_16[169], stage0_16[170], stage0_16[171], stage0_16[172], stage0_16[173], stage0_16[174]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[61],stage1_18[64],stage1_17[108],stage1_16[169]}
   );
   gpc606_5 gpc651 (
      {stage0_16[175], stage0_16[176], stage0_16[177], stage0_16[178], stage0_16[179], stage0_16[180]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[62],stage1_18[65],stage1_17[109],stage1_16[170]}
   );
   gpc606_5 gpc652 (
      {stage0_16[181], stage0_16[182], stage0_16[183], stage0_16[184], stage0_16[185], stage0_16[186]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[63],stage1_18[66],stage1_17[110],stage1_16[171]}
   );
   gpc606_5 gpc653 (
      {stage0_16[187], stage0_16[188], stage0_16[189], stage0_16[190], stage0_16[191], stage0_16[192]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[64],stage1_18[67],stage1_17[111],stage1_16[172]}
   );
   gpc606_5 gpc654 (
      {stage0_16[193], stage0_16[194], stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[65],stage1_18[68],stage1_17[112],stage1_16[173]}
   );
   gpc606_5 gpc655 (
      {stage0_16[199], stage0_16[200], stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[66],stage1_18[69],stage1_17[113],stage1_16[174]}
   );
   gpc606_5 gpc656 (
      {stage0_16[205], stage0_16[206], stage0_16[207], stage0_16[208], stage0_16[209], stage0_16[210]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[67],stage1_18[70],stage1_17[114],stage1_16[175]}
   );
   gpc606_5 gpc657 (
      {stage0_16[211], stage0_16[212], stage0_16[213], stage0_16[214], stage0_16[215], stage0_16[216]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[68],stage1_18[71],stage1_17[115],stage1_16[176]}
   );
   gpc606_5 gpc658 (
      {stage0_16[217], stage0_16[218], stage0_16[219], stage0_16[220], stage0_16[221], stage0_16[222]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[69],stage1_18[72],stage1_17[116],stage1_16[177]}
   );
   gpc606_5 gpc659 (
      {stage0_16[223], stage0_16[224], stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[70],stage1_18[73],stage1_17[117],stage1_16[178]}
   );
   gpc606_5 gpc660 (
      {stage0_16[229], stage0_16[230], stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[71],stage1_18[74],stage1_17[118],stage1_16[179]}
   );
   gpc606_5 gpc661 (
      {stage0_16[235], stage0_16[236], stage0_16[237], stage0_16[238], stage0_16[239], stage0_16[240]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[72],stage1_18[75],stage1_17[119],stage1_16[180]}
   );
   gpc606_5 gpc662 (
      {stage0_16[241], stage0_16[242], stage0_16[243], stage0_16[244], stage0_16[245], stage0_16[246]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[73],stage1_18[76],stage1_17[120],stage1_16[181]}
   );
   gpc606_5 gpc663 (
      {stage0_16[247], stage0_16[248], stage0_16[249], stage0_16[250], stage0_16[251], stage0_16[252]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[74],stage1_18[77],stage1_17[121],stage1_16[182]}
   );
   gpc606_5 gpc664 (
      {stage0_16[253], stage0_16[254], stage0_16[255], stage0_16[256], stage0_16[257], stage0_16[258]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[75],stage1_18[78],stage1_17[122],stage1_16[183]}
   );
   gpc606_5 gpc665 (
      {stage0_16[259], stage0_16[260], stage0_16[261], stage0_16[262], stage0_16[263], stage0_16[264]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[76],stage1_18[79],stage1_17[123],stage1_16[184]}
   );
   gpc606_5 gpc666 (
      {stage0_16[265], stage0_16[266], stage0_16[267], stage0_16[268], stage0_16[269], stage0_16[270]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[77],stage1_18[80],stage1_17[124],stage1_16[185]}
   );
   gpc606_5 gpc667 (
      {stage0_16[271], stage0_16[272], stage0_16[273], stage0_16[274], stage0_16[275], stage0_16[276]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[78],stage1_18[81],stage1_17[125],stage1_16[186]}
   );
   gpc606_5 gpc668 (
      {stage0_16[277], stage0_16[278], stage0_16[279], stage0_16[280], stage0_16[281], stage0_16[282]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[79],stage1_18[82],stage1_17[126],stage1_16[187]}
   );
   gpc606_5 gpc669 (
      {stage0_16[283], stage0_16[284], stage0_16[285], stage0_16[286], stage0_16[287], stage0_16[288]},
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226], stage0_18[227]},
      {stage1_20[37],stage1_19[80],stage1_18[83],stage1_17[127],stage1_16[188]}
   );
   gpc606_5 gpc670 (
      {stage0_16[289], stage0_16[290], stage0_16[291], stage0_16[292], stage0_16[293], stage0_16[294]},
      {stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231], stage0_18[232], stage0_18[233]},
      {stage1_20[38],stage1_19[81],stage1_18[84],stage1_17[128],stage1_16[189]}
   );
   gpc606_5 gpc671 (
      {stage0_16[295], stage0_16[296], stage0_16[297], stage0_16[298], stage0_16[299], stage0_16[300]},
      {stage0_18[234], stage0_18[235], stage0_18[236], stage0_18[237], stage0_18[238], stage0_18[239]},
      {stage1_20[39],stage1_19[82],stage1_18[85],stage1_17[129],stage1_16[190]}
   );
   gpc606_5 gpc672 (
      {stage0_16[301], stage0_16[302], stage0_16[303], stage0_16[304], stage0_16[305], stage0_16[306]},
      {stage0_18[240], stage0_18[241], stage0_18[242], stage0_18[243], stage0_18[244], stage0_18[245]},
      {stage1_20[40],stage1_19[83],stage1_18[86],stage1_17[130],stage1_16[191]}
   );
   gpc606_5 gpc673 (
      {stage0_16[307], stage0_16[308], stage0_16[309], stage0_16[310], stage0_16[311], stage0_16[312]},
      {stage0_18[246], stage0_18[247], stage0_18[248], stage0_18[249], stage0_18[250], stage0_18[251]},
      {stage1_20[41],stage1_19[84],stage1_18[87],stage1_17[131],stage1_16[192]}
   );
   gpc606_5 gpc674 (
      {stage0_16[313], stage0_16[314], stage0_16[315], stage0_16[316], stage0_16[317], stage0_16[318]},
      {stage0_18[252], stage0_18[253], stage0_18[254], stage0_18[255], stage0_18[256], stage0_18[257]},
      {stage1_20[42],stage1_19[85],stage1_18[88],stage1_17[132],stage1_16[193]}
   );
   gpc606_5 gpc675 (
      {stage0_16[319], stage0_16[320], stage0_16[321], stage0_16[322], stage0_16[323], stage0_16[324]},
      {stage0_18[258], stage0_18[259], stage0_18[260], stage0_18[261], stage0_18[262], stage0_18[263]},
      {stage1_20[43],stage1_19[86],stage1_18[89],stage1_17[133],stage1_16[194]}
   );
   gpc606_5 gpc676 (
      {stage0_16[325], stage0_16[326], stage0_16[327], stage0_16[328], stage0_16[329], stage0_16[330]},
      {stage0_18[264], stage0_18[265], stage0_18[266], stage0_18[267], stage0_18[268], stage0_18[269]},
      {stage1_20[44],stage1_19[87],stage1_18[90],stage1_17[134],stage1_16[195]}
   );
   gpc606_5 gpc677 (
      {stage0_16[331], stage0_16[332], stage0_16[333], stage0_16[334], stage0_16[335], stage0_16[336]},
      {stage0_18[270], stage0_18[271], stage0_18[272], stage0_18[273], stage0_18[274], stage0_18[275]},
      {stage1_20[45],stage1_19[88],stage1_18[91],stage1_17[135],stage1_16[196]}
   );
   gpc606_5 gpc678 (
      {stage0_16[337], stage0_16[338], stage0_16[339], stage0_16[340], stage0_16[341], stage0_16[342]},
      {stage0_18[276], stage0_18[277], stage0_18[278], stage0_18[279], stage0_18[280], stage0_18[281]},
      {stage1_20[46],stage1_19[89],stage1_18[92],stage1_17[136],stage1_16[197]}
   );
   gpc606_5 gpc679 (
      {stage0_16[343], stage0_16[344], stage0_16[345], stage0_16[346], stage0_16[347], stage0_16[348]},
      {stage0_18[282], stage0_18[283], stage0_18[284], stage0_18[285], stage0_18[286], stage0_18[287]},
      {stage1_20[47],stage1_19[90],stage1_18[93],stage1_17[137],stage1_16[198]}
   );
   gpc606_5 gpc680 (
      {stage0_16[349], stage0_16[350], stage0_16[351], stage0_16[352], stage0_16[353], stage0_16[354]},
      {stage0_18[288], stage0_18[289], stage0_18[290], stage0_18[291], stage0_18[292], stage0_18[293]},
      {stage1_20[48],stage1_19[91],stage1_18[94],stage1_17[138],stage1_16[199]}
   );
   gpc606_5 gpc681 (
      {stage0_16[355], stage0_16[356], stage0_16[357], stage0_16[358], stage0_16[359], stage0_16[360]},
      {stage0_18[294], stage0_18[295], stage0_18[296], stage0_18[297], stage0_18[298], stage0_18[299]},
      {stage1_20[49],stage1_19[92],stage1_18[95],stage1_17[139],stage1_16[200]}
   );
   gpc606_5 gpc682 (
      {stage0_16[361], stage0_16[362], stage0_16[363], stage0_16[364], stage0_16[365], stage0_16[366]},
      {stage0_18[300], stage0_18[301], stage0_18[302], stage0_18[303], stage0_18[304], stage0_18[305]},
      {stage1_20[50],stage1_19[93],stage1_18[96],stage1_17[140],stage1_16[201]}
   );
   gpc606_5 gpc683 (
      {stage0_16[367], stage0_16[368], stage0_16[369], stage0_16[370], stage0_16[371], stage0_16[372]},
      {stage0_18[306], stage0_18[307], stage0_18[308], stage0_18[309], stage0_18[310], stage0_18[311]},
      {stage1_20[51],stage1_19[94],stage1_18[97],stage1_17[141],stage1_16[202]}
   );
   gpc606_5 gpc684 (
      {stage0_16[373], stage0_16[374], stage0_16[375], stage0_16[376], stage0_16[377], stage0_16[378]},
      {stage0_18[312], stage0_18[313], stage0_18[314], stage0_18[315], stage0_18[316], stage0_18[317]},
      {stage1_20[52],stage1_19[95],stage1_18[98],stage1_17[142],stage1_16[203]}
   );
   gpc606_5 gpc685 (
      {stage0_16[379], stage0_16[380], stage0_16[381], stage0_16[382], stage0_16[383], stage0_16[384]},
      {stage0_18[318], stage0_18[319], stage0_18[320], stage0_18[321], stage0_18[322], stage0_18[323]},
      {stage1_20[53],stage1_19[96],stage1_18[99],stage1_17[143],stage1_16[204]}
   );
   gpc606_5 gpc686 (
      {stage0_16[385], stage0_16[386], stage0_16[387], stage0_16[388], stage0_16[389], stage0_16[390]},
      {stage0_18[324], stage0_18[325], stage0_18[326], stage0_18[327], stage0_18[328], stage0_18[329]},
      {stage1_20[54],stage1_19[97],stage1_18[100],stage1_17[144],stage1_16[205]}
   );
   gpc606_5 gpc687 (
      {stage0_16[391], stage0_16[392], stage0_16[393], stage0_16[394], stage0_16[395], stage0_16[396]},
      {stage0_18[330], stage0_18[331], stage0_18[332], stage0_18[333], stage0_18[334], stage0_18[335]},
      {stage1_20[55],stage1_19[98],stage1_18[101],stage1_17[145],stage1_16[206]}
   );
   gpc606_5 gpc688 (
      {stage0_16[397], stage0_16[398], stage0_16[399], stage0_16[400], stage0_16[401], stage0_16[402]},
      {stage0_18[336], stage0_18[337], stage0_18[338], stage0_18[339], stage0_18[340], stage0_18[341]},
      {stage1_20[56],stage1_19[99],stage1_18[102],stage1_17[146],stage1_16[207]}
   );
   gpc606_5 gpc689 (
      {stage0_16[403], stage0_16[404], stage0_16[405], stage0_16[406], stage0_16[407], stage0_16[408]},
      {stage0_18[342], stage0_18[343], stage0_18[344], stage0_18[345], stage0_18[346], stage0_18[347]},
      {stage1_20[57],stage1_19[100],stage1_18[103],stage1_17[147],stage1_16[208]}
   );
   gpc606_5 gpc690 (
      {stage0_16[409], stage0_16[410], stage0_16[411], stage0_16[412], stage0_16[413], stage0_16[414]},
      {stage0_18[348], stage0_18[349], stage0_18[350], stage0_18[351], stage0_18[352], stage0_18[353]},
      {stage1_20[58],stage1_19[101],stage1_18[104],stage1_17[148],stage1_16[209]}
   );
   gpc606_5 gpc691 (
      {stage0_16[415], stage0_16[416], stage0_16[417], stage0_16[418], stage0_16[419], stage0_16[420]},
      {stage0_18[354], stage0_18[355], stage0_18[356], stage0_18[357], stage0_18[358], stage0_18[359]},
      {stage1_20[59],stage1_19[102],stage1_18[105],stage1_17[149],stage1_16[210]}
   );
   gpc606_5 gpc692 (
      {stage0_16[421], stage0_16[422], stage0_16[423], stage0_16[424], stage0_16[425], stage0_16[426]},
      {stage0_18[360], stage0_18[361], stage0_18[362], stage0_18[363], stage0_18[364], stage0_18[365]},
      {stage1_20[60],stage1_19[103],stage1_18[106],stage1_17[150],stage1_16[211]}
   );
   gpc606_5 gpc693 (
      {stage0_16[427], stage0_16[428], stage0_16[429], stage0_16[430], stage0_16[431], stage0_16[432]},
      {stage0_18[366], stage0_18[367], stage0_18[368], stage0_18[369], stage0_18[370], stage0_18[371]},
      {stage1_20[61],stage1_19[104],stage1_18[107],stage1_17[151],stage1_16[212]}
   );
   gpc606_5 gpc694 (
      {stage0_16[433], stage0_16[434], stage0_16[435], stage0_16[436], stage0_16[437], stage0_16[438]},
      {stage0_18[372], stage0_18[373], stage0_18[374], stage0_18[375], stage0_18[376], stage0_18[377]},
      {stage1_20[62],stage1_19[105],stage1_18[108],stage1_17[152],stage1_16[213]}
   );
   gpc606_5 gpc695 (
      {stage0_16[439], stage0_16[440], stage0_16[441], stage0_16[442], stage0_16[443], stage0_16[444]},
      {stage0_18[378], stage0_18[379], stage0_18[380], stage0_18[381], stage0_18[382], stage0_18[383]},
      {stage1_20[63],stage1_19[106],stage1_18[109],stage1_17[153],stage1_16[214]}
   );
   gpc606_5 gpc696 (
      {stage0_16[445], stage0_16[446], stage0_16[447], stage0_16[448], stage0_16[449], stage0_16[450]},
      {stage0_18[384], stage0_18[385], stage0_18[386], stage0_18[387], stage0_18[388], stage0_18[389]},
      {stage1_20[64],stage1_19[107],stage1_18[110],stage1_17[154],stage1_16[215]}
   );
   gpc606_5 gpc697 (
      {stage0_16[451], stage0_16[452], stage0_16[453], stage0_16[454], stage0_16[455], stage0_16[456]},
      {stage0_18[390], stage0_18[391], stage0_18[392], stage0_18[393], stage0_18[394], stage0_18[395]},
      {stage1_20[65],stage1_19[108],stage1_18[111],stage1_17[155],stage1_16[216]}
   );
   gpc606_5 gpc698 (
      {stage0_16[457], stage0_16[458], stage0_16[459], stage0_16[460], stage0_16[461], stage0_16[462]},
      {stage0_18[396], stage0_18[397], stage0_18[398], stage0_18[399], stage0_18[400], stage0_18[401]},
      {stage1_20[66],stage1_19[109],stage1_18[112],stage1_17[156],stage1_16[217]}
   );
   gpc606_5 gpc699 (
      {stage0_16[463], stage0_16[464], stage0_16[465], stage0_16[466], stage0_16[467], stage0_16[468]},
      {stage0_18[402], stage0_18[403], stage0_18[404], stage0_18[405], stage0_18[406], stage0_18[407]},
      {stage1_20[67],stage1_19[110],stage1_18[113],stage1_17[157],stage1_16[218]}
   );
   gpc606_5 gpc700 (
      {stage0_16[469], stage0_16[470], stage0_16[471], stage0_16[472], stage0_16[473], stage0_16[474]},
      {stage0_18[408], stage0_18[409], stage0_18[410], stage0_18[411], stage0_18[412], stage0_18[413]},
      {stage1_20[68],stage1_19[111],stage1_18[114],stage1_17[158],stage1_16[219]}
   );
   gpc606_5 gpc701 (
      {stage0_16[475], stage0_16[476], stage0_16[477], stage0_16[478], stage0_16[479], stage0_16[480]},
      {stage0_18[414], stage0_18[415], stage0_18[416], stage0_18[417], stage0_18[418], stage0_18[419]},
      {stage1_20[69],stage1_19[112],stage1_18[115],stage1_17[159],stage1_16[220]}
   );
   gpc606_5 gpc702 (
      {stage0_16[481], stage0_16[482], stage0_16[483], stage0_16[484], stage0_16[485], 1'b0},
      {stage0_18[420], stage0_18[421], stage0_18[422], stage0_18[423], stage0_18[424], stage0_18[425]},
      {stage1_20[70],stage1_19[113],stage1_18[116],stage1_17[160],stage1_16[221]}
   );
   gpc606_5 gpc703 (
      {stage0_17[258], stage0_17[259], stage0_17[260], stage0_17[261], stage0_17[262], stage0_17[263]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[71],stage1_19[114],stage1_18[117],stage1_17[161]}
   );
   gpc606_5 gpc704 (
      {stage0_17[264], stage0_17[265], stage0_17[266], stage0_17[267], stage0_17[268], stage0_17[269]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[72],stage1_19[115],stage1_18[118],stage1_17[162]}
   );
   gpc606_5 gpc705 (
      {stage0_17[270], stage0_17[271], stage0_17[272], stage0_17[273], stage0_17[274], stage0_17[275]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[73],stage1_19[116],stage1_18[119],stage1_17[163]}
   );
   gpc606_5 gpc706 (
      {stage0_17[276], stage0_17[277], stage0_17[278], stage0_17[279], stage0_17[280], stage0_17[281]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[74],stage1_19[117],stage1_18[120],stage1_17[164]}
   );
   gpc606_5 gpc707 (
      {stage0_17[282], stage0_17[283], stage0_17[284], stage0_17[285], stage0_17[286], stage0_17[287]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[75],stage1_19[118],stage1_18[121],stage1_17[165]}
   );
   gpc606_5 gpc708 (
      {stage0_17[288], stage0_17[289], stage0_17[290], stage0_17[291], stage0_17[292], stage0_17[293]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[76],stage1_19[119],stage1_18[122],stage1_17[166]}
   );
   gpc606_5 gpc709 (
      {stage0_17[294], stage0_17[295], stage0_17[296], stage0_17[297], stage0_17[298], stage0_17[299]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[77],stage1_19[120],stage1_18[123],stage1_17[167]}
   );
   gpc606_5 gpc710 (
      {stage0_17[300], stage0_17[301], stage0_17[302], stage0_17[303], stage0_17[304], stage0_17[305]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[78],stage1_19[121],stage1_18[124],stage1_17[168]}
   );
   gpc606_5 gpc711 (
      {stage0_17[306], stage0_17[307], stage0_17[308], stage0_17[309], stage0_17[310], stage0_17[311]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[79],stage1_19[122],stage1_18[125],stage1_17[169]}
   );
   gpc606_5 gpc712 (
      {stage0_17[312], stage0_17[313], stage0_17[314], stage0_17[315], stage0_17[316], stage0_17[317]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[80],stage1_19[123],stage1_18[126],stage1_17[170]}
   );
   gpc606_5 gpc713 (
      {stage0_17[318], stage0_17[319], stage0_17[320], stage0_17[321], stage0_17[322], stage0_17[323]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[81],stage1_19[124],stage1_18[127],stage1_17[171]}
   );
   gpc606_5 gpc714 (
      {stage0_17[324], stage0_17[325], stage0_17[326], stage0_17[327], stage0_17[328], stage0_17[329]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[82],stage1_19[125],stage1_18[128],stage1_17[172]}
   );
   gpc606_5 gpc715 (
      {stage0_17[330], stage0_17[331], stage0_17[332], stage0_17[333], stage0_17[334], stage0_17[335]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[83],stage1_19[126],stage1_18[129],stage1_17[173]}
   );
   gpc606_5 gpc716 (
      {stage0_17[336], stage0_17[337], stage0_17[338], stage0_17[339], stage0_17[340], stage0_17[341]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[84],stage1_19[127],stage1_18[130],stage1_17[174]}
   );
   gpc606_5 gpc717 (
      {stage0_17[342], stage0_17[343], stage0_17[344], stage0_17[345], stage0_17[346], stage0_17[347]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[85],stage1_19[128],stage1_18[131],stage1_17[175]}
   );
   gpc606_5 gpc718 (
      {stage0_17[348], stage0_17[349], stage0_17[350], stage0_17[351], stage0_17[352], stage0_17[353]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[86],stage1_19[129],stage1_18[132],stage1_17[176]}
   );
   gpc606_5 gpc719 (
      {stage0_17[354], stage0_17[355], stage0_17[356], stage0_17[357], stage0_17[358], stage0_17[359]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[87],stage1_19[130],stage1_18[133],stage1_17[177]}
   );
   gpc606_5 gpc720 (
      {stage0_17[360], stage0_17[361], stage0_17[362], stage0_17[363], stage0_17[364], stage0_17[365]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[88],stage1_19[131],stage1_18[134],stage1_17[178]}
   );
   gpc606_5 gpc721 (
      {stage0_17[366], stage0_17[367], stage0_17[368], stage0_17[369], stage0_17[370], stage0_17[371]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[89],stage1_19[132],stage1_18[135],stage1_17[179]}
   );
   gpc606_5 gpc722 (
      {stage0_17[372], stage0_17[373], stage0_17[374], stage0_17[375], stage0_17[376], stage0_17[377]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[90],stage1_19[133],stage1_18[136],stage1_17[180]}
   );
   gpc606_5 gpc723 (
      {stage0_17[378], stage0_17[379], stage0_17[380], stage0_17[381], stage0_17[382], stage0_17[383]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[91],stage1_19[134],stage1_18[137],stage1_17[181]}
   );
   gpc606_5 gpc724 (
      {stage0_17[384], stage0_17[385], stage0_17[386], stage0_17[387], stage0_17[388], stage0_17[389]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[92],stage1_19[135],stage1_18[138],stage1_17[182]}
   );
   gpc606_5 gpc725 (
      {stage0_17[390], stage0_17[391], stage0_17[392], stage0_17[393], stage0_17[394], stage0_17[395]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[93],stage1_19[136],stage1_18[139],stage1_17[183]}
   );
   gpc606_5 gpc726 (
      {stage0_17[396], stage0_17[397], stage0_17[398], stage0_17[399], stage0_17[400], stage0_17[401]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[94],stage1_19[137],stage1_18[140],stage1_17[184]}
   );
   gpc606_5 gpc727 (
      {stage0_17[402], stage0_17[403], stage0_17[404], stage0_17[405], stage0_17[406], stage0_17[407]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[95],stage1_19[138],stage1_18[141],stage1_17[185]}
   );
   gpc606_5 gpc728 (
      {stage0_17[408], stage0_17[409], stage0_17[410], stage0_17[411], stage0_17[412], stage0_17[413]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[96],stage1_19[139],stage1_18[142],stage1_17[186]}
   );
   gpc606_5 gpc729 (
      {stage0_17[414], stage0_17[415], stage0_17[416], stage0_17[417], stage0_17[418], stage0_17[419]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[97],stage1_19[140],stage1_18[143],stage1_17[187]}
   );
   gpc606_5 gpc730 (
      {stage0_17[420], stage0_17[421], stage0_17[422], stage0_17[423], stage0_17[424], stage0_17[425]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[98],stage1_19[141],stage1_18[144],stage1_17[188]}
   );
   gpc606_5 gpc731 (
      {stage0_17[426], stage0_17[427], stage0_17[428], stage0_17[429], stage0_17[430], stage0_17[431]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[99],stage1_19[142],stage1_18[145],stage1_17[189]}
   );
   gpc606_5 gpc732 (
      {stage0_17[432], stage0_17[433], stage0_17[434], stage0_17[435], stage0_17[436], stage0_17[437]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[100],stage1_19[143],stage1_18[146],stage1_17[190]}
   );
   gpc606_5 gpc733 (
      {stage0_17[438], stage0_17[439], stage0_17[440], stage0_17[441], stage0_17[442], stage0_17[443]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[101],stage1_19[144],stage1_18[147],stage1_17[191]}
   );
   gpc606_5 gpc734 (
      {stage0_17[444], stage0_17[445], stage0_17[446], stage0_17[447], stage0_17[448], stage0_17[449]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[102],stage1_19[145],stage1_18[148],stage1_17[192]}
   );
   gpc615_5 gpc735 (
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196]},
      {stage0_20[0]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[0],stage1_21[32],stage1_20[103],stage1_19[146]}
   );
   gpc615_5 gpc736 (
      {stage0_19[197], stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201]},
      {stage0_20[1]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[1],stage1_21[33],stage1_20[104],stage1_19[147]}
   );
   gpc615_5 gpc737 (
      {stage0_19[202], stage0_19[203], stage0_19[204], stage0_19[205], stage0_19[206]},
      {stage0_20[2]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[2],stage1_21[34],stage1_20[105],stage1_19[148]}
   );
   gpc615_5 gpc738 (
      {stage0_19[207], stage0_19[208], stage0_19[209], stage0_19[210], stage0_19[211]},
      {stage0_20[3]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[3],stage1_21[35],stage1_20[106],stage1_19[149]}
   );
   gpc615_5 gpc739 (
      {stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215], stage0_19[216]},
      {stage0_20[4]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[4],stage1_21[36],stage1_20[107],stage1_19[150]}
   );
   gpc615_5 gpc740 (
      {stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage0_20[5]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[5],stage1_21[37],stage1_20[108],stage1_19[151]}
   );
   gpc615_5 gpc741 (
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226]},
      {stage0_20[6]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[6],stage1_21[38],stage1_20[109],stage1_19[152]}
   );
   gpc615_5 gpc742 (
      {stage0_19[227], stage0_19[228], stage0_19[229], stage0_19[230], stage0_19[231]},
      {stage0_20[7]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[7],stage1_21[39],stage1_20[110],stage1_19[153]}
   );
   gpc615_5 gpc743 (
      {stage0_19[232], stage0_19[233], stage0_19[234], stage0_19[235], stage0_19[236]},
      {stage0_20[8]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[8],stage1_21[40],stage1_20[111],stage1_19[154]}
   );
   gpc615_5 gpc744 (
      {stage0_19[237], stage0_19[238], stage0_19[239], stage0_19[240], stage0_19[241]},
      {stage0_20[9]},
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage1_23[9],stage1_22[9],stage1_21[41],stage1_20[112],stage1_19[155]}
   );
   gpc615_5 gpc745 (
      {stage0_19[242], stage0_19[243], stage0_19[244], stage0_19[245], stage0_19[246]},
      {stage0_20[10]},
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage1_23[10],stage1_22[10],stage1_21[42],stage1_20[113],stage1_19[156]}
   );
   gpc615_5 gpc746 (
      {stage0_19[247], stage0_19[248], stage0_19[249], stage0_19[250], stage0_19[251]},
      {stage0_20[11]},
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage1_23[11],stage1_22[11],stage1_21[43],stage1_20[114],stage1_19[157]}
   );
   gpc615_5 gpc747 (
      {stage0_19[252], stage0_19[253], stage0_19[254], stage0_19[255], stage0_19[256]},
      {stage0_20[12]},
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage1_23[12],stage1_22[12],stage1_21[44],stage1_20[115],stage1_19[158]}
   );
   gpc615_5 gpc748 (
      {stage0_19[257], stage0_19[258], stage0_19[259], stage0_19[260], stage0_19[261]},
      {stage0_20[13]},
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage1_23[13],stage1_22[13],stage1_21[45],stage1_20[116],stage1_19[159]}
   );
   gpc615_5 gpc749 (
      {stage0_19[262], stage0_19[263], stage0_19[264], stage0_19[265], stage0_19[266]},
      {stage0_20[14]},
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage1_23[14],stage1_22[14],stage1_21[46],stage1_20[117],stage1_19[160]}
   );
   gpc615_5 gpc750 (
      {stage0_19[267], stage0_19[268], stage0_19[269], stage0_19[270], stage0_19[271]},
      {stage0_20[15]},
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage1_23[15],stage1_22[15],stage1_21[47],stage1_20[118],stage1_19[161]}
   );
   gpc615_5 gpc751 (
      {stage0_19[272], stage0_19[273], stage0_19[274], stage0_19[275], stage0_19[276]},
      {stage0_20[16]},
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage1_23[16],stage1_22[16],stage1_21[48],stage1_20[119],stage1_19[162]}
   );
   gpc615_5 gpc752 (
      {stage0_19[277], stage0_19[278], stage0_19[279], stage0_19[280], stage0_19[281]},
      {stage0_20[17]},
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage1_23[17],stage1_22[17],stage1_21[49],stage1_20[120],stage1_19[163]}
   );
   gpc615_5 gpc753 (
      {stage0_19[282], stage0_19[283], stage0_19[284], stage0_19[285], stage0_19[286]},
      {stage0_20[18]},
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage1_23[18],stage1_22[18],stage1_21[50],stage1_20[121],stage1_19[164]}
   );
   gpc615_5 gpc754 (
      {stage0_19[287], stage0_19[288], stage0_19[289], stage0_19[290], stage0_19[291]},
      {stage0_20[19]},
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage1_23[19],stage1_22[19],stage1_21[51],stage1_20[122],stage1_19[165]}
   );
   gpc615_5 gpc755 (
      {stage0_19[292], stage0_19[293], stage0_19[294], stage0_19[295], stage0_19[296]},
      {stage0_20[20]},
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage1_23[20],stage1_22[20],stage1_21[52],stage1_20[123],stage1_19[166]}
   );
   gpc615_5 gpc756 (
      {stage0_19[297], stage0_19[298], stage0_19[299], stage0_19[300], stage0_19[301]},
      {stage0_20[21]},
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage1_23[21],stage1_22[21],stage1_21[53],stage1_20[124],stage1_19[167]}
   );
   gpc615_5 gpc757 (
      {stage0_19[302], stage0_19[303], stage0_19[304], stage0_19[305], stage0_19[306]},
      {stage0_20[22]},
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage1_23[22],stage1_22[22],stage1_21[54],stage1_20[125],stage1_19[168]}
   );
   gpc615_5 gpc758 (
      {stage0_19[307], stage0_19[308], stage0_19[309], stage0_19[310], stage0_19[311]},
      {stage0_20[23]},
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage1_23[23],stage1_22[23],stage1_21[55],stage1_20[126],stage1_19[169]}
   );
   gpc615_5 gpc759 (
      {stage0_19[312], stage0_19[313], stage0_19[314], stage0_19[315], stage0_19[316]},
      {stage0_20[24]},
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage1_23[24],stage1_22[24],stage1_21[56],stage1_20[127],stage1_19[170]}
   );
   gpc615_5 gpc760 (
      {stage0_19[317], stage0_19[318], stage0_19[319], stage0_19[320], stage0_19[321]},
      {stage0_20[25]},
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage1_23[25],stage1_22[25],stage1_21[57],stage1_20[128],stage1_19[171]}
   );
   gpc615_5 gpc761 (
      {stage0_19[322], stage0_19[323], stage0_19[324], stage0_19[325], stage0_19[326]},
      {stage0_20[26]},
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage1_23[26],stage1_22[26],stage1_21[58],stage1_20[129],stage1_19[172]}
   );
   gpc615_5 gpc762 (
      {stage0_19[327], stage0_19[328], stage0_19[329], stage0_19[330], stage0_19[331]},
      {stage0_20[27]},
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage1_23[27],stage1_22[27],stage1_21[59],stage1_20[130],stage1_19[173]}
   );
   gpc615_5 gpc763 (
      {stage0_19[332], stage0_19[333], stage0_19[334], stage0_19[335], stage0_19[336]},
      {stage0_20[28]},
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage1_23[28],stage1_22[28],stage1_21[60],stage1_20[131],stage1_19[174]}
   );
   gpc615_5 gpc764 (
      {stage0_19[337], stage0_19[338], stage0_19[339], stage0_19[340], stage0_19[341]},
      {stage0_20[29]},
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage1_23[29],stage1_22[29],stage1_21[61],stage1_20[132],stage1_19[175]}
   );
   gpc615_5 gpc765 (
      {stage0_19[342], stage0_19[343], stage0_19[344], stage0_19[345], stage0_19[346]},
      {stage0_20[30]},
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage1_23[30],stage1_22[30],stage1_21[62],stage1_20[133],stage1_19[176]}
   );
   gpc615_5 gpc766 (
      {stage0_19[347], stage0_19[348], stage0_19[349], stage0_19[350], stage0_19[351]},
      {stage0_20[31]},
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage1_23[31],stage1_22[31],stage1_21[63],stage1_20[134],stage1_19[177]}
   );
   gpc615_5 gpc767 (
      {stage0_19[352], stage0_19[353], stage0_19[354], stage0_19[355], stage0_19[356]},
      {stage0_20[32]},
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage1_23[32],stage1_22[32],stage1_21[64],stage1_20[135],stage1_19[178]}
   );
   gpc615_5 gpc768 (
      {stage0_19[357], stage0_19[358], stage0_19[359], stage0_19[360], stage0_19[361]},
      {stage0_20[33]},
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage1_23[33],stage1_22[33],stage1_21[65],stage1_20[136],stage1_19[179]}
   );
   gpc615_5 gpc769 (
      {stage0_19[362], stage0_19[363], stage0_19[364], stage0_19[365], stage0_19[366]},
      {stage0_20[34]},
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage1_23[34],stage1_22[34],stage1_21[66],stage1_20[137],stage1_19[180]}
   );
   gpc615_5 gpc770 (
      {stage0_19[367], stage0_19[368], stage0_19[369], stage0_19[370], stage0_19[371]},
      {stage0_20[35]},
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage1_23[35],stage1_22[35],stage1_21[67],stage1_20[138],stage1_19[181]}
   );
   gpc615_5 gpc771 (
      {stage0_19[372], stage0_19[373], stage0_19[374], stage0_19[375], stage0_19[376]},
      {stage0_20[36]},
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage1_23[36],stage1_22[36],stage1_21[68],stage1_20[139],stage1_19[182]}
   );
   gpc615_5 gpc772 (
      {stage0_19[377], stage0_19[378], stage0_19[379], stage0_19[380], stage0_19[381]},
      {stage0_20[37]},
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage1_23[37],stage1_22[37],stage1_21[69],stage1_20[140],stage1_19[183]}
   );
   gpc615_5 gpc773 (
      {stage0_19[382], stage0_19[383], stage0_19[384], stage0_19[385], stage0_19[386]},
      {stage0_20[38]},
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage1_23[38],stage1_22[38],stage1_21[70],stage1_20[141],stage1_19[184]}
   );
   gpc615_5 gpc774 (
      {stage0_19[387], stage0_19[388], stage0_19[389], stage0_19[390], stage0_19[391]},
      {stage0_20[39]},
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage1_23[39],stage1_22[39],stage1_21[71],stage1_20[142],stage1_19[185]}
   );
   gpc615_5 gpc775 (
      {stage0_19[392], stage0_19[393], stage0_19[394], stage0_19[395], stage0_19[396]},
      {stage0_20[40]},
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage1_23[40],stage1_22[40],stage1_21[72],stage1_20[143],stage1_19[186]}
   );
   gpc1343_5 gpc776 (
      {stage0_20[41], stage0_20[42], stage0_20[43]},
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249]},
      {stage0_22[0], stage0_22[1], stage0_22[2]},
      {stage0_23[0]},
      {stage1_24[0],stage1_23[41],stage1_22[41],stage1_21[73],stage1_20[144]}
   );
   gpc1163_5 gpc777 (
      {stage0_20[44], stage0_20[45], stage0_20[46]},
      {stage0_21[250], stage0_21[251], stage0_21[252], stage0_21[253], stage0_21[254], stage0_21[255]},
      {stage0_22[3]},
      {stage0_23[1]},
      {stage1_24[1],stage1_23[42],stage1_22[42],stage1_21[74],stage1_20[145]}
   );
   gpc1163_5 gpc778 (
      {stage0_20[47], stage0_20[48], stage0_20[49]},
      {stage0_21[256], stage0_21[257], stage0_21[258], stage0_21[259], stage0_21[260], stage0_21[261]},
      {stage0_22[4]},
      {stage0_23[2]},
      {stage1_24[2],stage1_23[43],stage1_22[43],stage1_21[75],stage1_20[146]}
   );
   gpc1163_5 gpc779 (
      {stage0_20[50], stage0_20[51], stage0_20[52]},
      {stage0_21[262], stage0_21[263], stage0_21[264], stage0_21[265], stage0_21[266], stage0_21[267]},
      {stage0_22[5]},
      {stage0_23[3]},
      {stage1_24[3],stage1_23[44],stage1_22[44],stage1_21[76],stage1_20[147]}
   );
   gpc1163_5 gpc780 (
      {stage0_20[53], stage0_20[54], stage0_20[55]},
      {stage0_21[268], stage0_21[269], stage0_21[270], stage0_21[271], stage0_21[272], stage0_21[273]},
      {stage0_22[6]},
      {stage0_23[4]},
      {stage1_24[4],stage1_23[45],stage1_22[45],stage1_21[77],stage1_20[148]}
   );
   gpc1163_5 gpc781 (
      {stage0_20[56], stage0_20[57], stage0_20[58]},
      {stage0_21[274], stage0_21[275], stage0_21[276], stage0_21[277], stage0_21[278], stage0_21[279]},
      {stage0_22[7]},
      {stage0_23[5]},
      {stage1_24[5],stage1_23[46],stage1_22[46],stage1_21[78],stage1_20[149]}
   );
   gpc1163_5 gpc782 (
      {stage0_20[59], stage0_20[60], stage0_20[61]},
      {stage0_21[280], stage0_21[281], stage0_21[282], stage0_21[283], stage0_21[284], stage0_21[285]},
      {stage0_22[8]},
      {stage0_23[6]},
      {stage1_24[6],stage1_23[47],stage1_22[47],stage1_21[79],stage1_20[150]}
   );
   gpc606_5 gpc783 (
      {stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65], stage0_20[66], stage0_20[67]},
      {stage0_22[9], stage0_22[10], stage0_22[11], stage0_22[12], stage0_22[13], stage0_22[14]},
      {stage1_24[7],stage1_23[48],stage1_22[48],stage1_21[80],stage1_20[151]}
   );
   gpc606_5 gpc784 (
      {stage0_20[68], stage0_20[69], stage0_20[70], stage0_20[71], stage0_20[72], stage0_20[73]},
      {stage0_22[15], stage0_22[16], stage0_22[17], stage0_22[18], stage0_22[19], stage0_22[20]},
      {stage1_24[8],stage1_23[49],stage1_22[49],stage1_21[81],stage1_20[152]}
   );
   gpc606_5 gpc785 (
      {stage0_20[74], stage0_20[75], stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79]},
      {stage0_22[21], stage0_22[22], stage0_22[23], stage0_22[24], stage0_22[25], stage0_22[26]},
      {stage1_24[9],stage1_23[50],stage1_22[50],stage1_21[82],stage1_20[153]}
   );
   gpc606_5 gpc786 (
      {stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83], stage0_20[84], stage0_20[85]},
      {stage0_22[27], stage0_22[28], stage0_22[29], stage0_22[30], stage0_22[31], stage0_22[32]},
      {stage1_24[10],stage1_23[51],stage1_22[51],stage1_21[83],stage1_20[154]}
   );
   gpc606_5 gpc787 (
      {stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89], stage0_20[90], stage0_20[91]},
      {stage0_22[33], stage0_22[34], stage0_22[35], stage0_22[36], stage0_22[37], stage0_22[38]},
      {stage1_24[11],stage1_23[52],stage1_22[52],stage1_21[84],stage1_20[155]}
   );
   gpc606_5 gpc788 (
      {stage0_20[92], stage0_20[93], stage0_20[94], stage0_20[95], stage0_20[96], stage0_20[97]},
      {stage0_22[39], stage0_22[40], stage0_22[41], stage0_22[42], stage0_22[43], stage0_22[44]},
      {stage1_24[12],stage1_23[53],stage1_22[53],stage1_21[85],stage1_20[156]}
   );
   gpc606_5 gpc789 (
      {stage0_20[98], stage0_20[99], stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103]},
      {stage0_22[45], stage0_22[46], stage0_22[47], stage0_22[48], stage0_22[49], stage0_22[50]},
      {stage1_24[13],stage1_23[54],stage1_22[54],stage1_21[86],stage1_20[157]}
   );
   gpc606_5 gpc790 (
      {stage0_20[104], stage0_20[105], stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109]},
      {stage0_22[51], stage0_22[52], stage0_22[53], stage0_22[54], stage0_22[55], stage0_22[56]},
      {stage1_24[14],stage1_23[55],stage1_22[55],stage1_21[87],stage1_20[158]}
   );
   gpc606_5 gpc791 (
      {stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113], stage0_20[114], stage0_20[115]},
      {stage0_22[57], stage0_22[58], stage0_22[59], stage0_22[60], stage0_22[61], stage0_22[62]},
      {stage1_24[15],stage1_23[56],stage1_22[56],stage1_21[88],stage1_20[159]}
   );
   gpc606_5 gpc792 (
      {stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119], stage0_20[120], stage0_20[121]},
      {stage0_22[63], stage0_22[64], stage0_22[65], stage0_22[66], stage0_22[67], stage0_22[68]},
      {stage1_24[16],stage1_23[57],stage1_22[57],stage1_21[89],stage1_20[160]}
   );
   gpc606_5 gpc793 (
      {stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125], stage0_20[126], stage0_20[127]},
      {stage0_22[69], stage0_22[70], stage0_22[71], stage0_22[72], stage0_22[73], stage0_22[74]},
      {stage1_24[17],stage1_23[58],stage1_22[58],stage1_21[90],stage1_20[161]}
   );
   gpc606_5 gpc794 (
      {stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131], stage0_20[132], stage0_20[133]},
      {stage0_22[75], stage0_22[76], stage0_22[77], stage0_22[78], stage0_22[79], stage0_22[80]},
      {stage1_24[18],stage1_23[59],stage1_22[59],stage1_21[91],stage1_20[162]}
   );
   gpc606_5 gpc795 (
      {stage0_20[134], stage0_20[135], stage0_20[136], stage0_20[137], stage0_20[138], stage0_20[139]},
      {stage0_22[81], stage0_22[82], stage0_22[83], stage0_22[84], stage0_22[85], stage0_22[86]},
      {stage1_24[19],stage1_23[60],stage1_22[60],stage1_21[92],stage1_20[163]}
   );
   gpc606_5 gpc796 (
      {stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143], stage0_20[144], stage0_20[145]},
      {stage0_22[87], stage0_22[88], stage0_22[89], stage0_22[90], stage0_22[91], stage0_22[92]},
      {stage1_24[20],stage1_23[61],stage1_22[61],stage1_21[93],stage1_20[164]}
   );
   gpc606_5 gpc797 (
      {stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149], stage0_20[150], stage0_20[151]},
      {stage0_22[93], stage0_22[94], stage0_22[95], stage0_22[96], stage0_22[97], stage0_22[98]},
      {stage1_24[21],stage1_23[62],stage1_22[62],stage1_21[94],stage1_20[165]}
   );
   gpc606_5 gpc798 (
      {stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155], stage0_20[156], stage0_20[157]},
      {stage0_22[99], stage0_22[100], stage0_22[101], stage0_22[102], stage0_22[103], stage0_22[104]},
      {stage1_24[22],stage1_23[63],stage1_22[63],stage1_21[95],stage1_20[166]}
   );
   gpc606_5 gpc799 (
      {stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161], stage0_20[162], stage0_20[163]},
      {stage0_22[105], stage0_22[106], stage0_22[107], stage0_22[108], stage0_22[109], stage0_22[110]},
      {stage1_24[23],stage1_23[64],stage1_22[64],stage1_21[96],stage1_20[167]}
   );
   gpc606_5 gpc800 (
      {stage0_20[164], stage0_20[165], stage0_20[166], stage0_20[167], stage0_20[168], stage0_20[169]},
      {stage0_22[111], stage0_22[112], stage0_22[113], stage0_22[114], stage0_22[115], stage0_22[116]},
      {stage1_24[24],stage1_23[65],stage1_22[65],stage1_21[97],stage1_20[168]}
   );
   gpc606_5 gpc801 (
      {stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173], stage0_20[174], stage0_20[175]},
      {stage0_22[117], stage0_22[118], stage0_22[119], stage0_22[120], stage0_22[121], stage0_22[122]},
      {stage1_24[25],stage1_23[66],stage1_22[66],stage1_21[98],stage1_20[169]}
   );
   gpc606_5 gpc802 (
      {stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179], stage0_20[180], stage0_20[181]},
      {stage0_22[123], stage0_22[124], stage0_22[125], stage0_22[126], stage0_22[127], stage0_22[128]},
      {stage1_24[26],stage1_23[67],stage1_22[67],stage1_21[99],stage1_20[170]}
   );
   gpc606_5 gpc803 (
      {stage0_20[182], stage0_20[183], stage0_20[184], stage0_20[185], stage0_20[186], stage0_20[187]},
      {stage0_22[129], stage0_22[130], stage0_22[131], stage0_22[132], stage0_22[133], stage0_22[134]},
      {stage1_24[27],stage1_23[68],stage1_22[68],stage1_21[100],stage1_20[171]}
   );
   gpc606_5 gpc804 (
      {stage0_20[188], stage0_20[189], stage0_20[190], stage0_20[191], stage0_20[192], stage0_20[193]},
      {stage0_22[135], stage0_22[136], stage0_22[137], stage0_22[138], stage0_22[139], stage0_22[140]},
      {stage1_24[28],stage1_23[69],stage1_22[69],stage1_21[101],stage1_20[172]}
   );
   gpc606_5 gpc805 (
      {stage0_20[194], stage0_20[195], stage0_20[196], stage0_20[197], stage0_20[198], stage0_20[199]},
      {stage0_22[141], stage0_22[142], stage0_22[143], stage0_22[144], stage0_22[145], stage0_22[146]},
      {stage1_24[29],stage1_23[70],stage1_22[70],stage1_21[102],stage1_20[173]}
   );
   gpc606_5 gpc806 (
      {stage0_20[200], stage0_20[201], stage0_20[202], stage0_20[203], stage0_20[204], stage0_20[205]},
      {stage0_22[147], stage0_22[148], stage0_22[149], stage0_22[150], stage0_22[151], stage0_22[152]},
      {stage1_24[30],stage1_23[71],stage1_22[71],stage1_21[103],stage1_20[174]}
   );
   gpc606_5 gpc807 (
      {stage0_20[206], stage0_20[207], stage0_20[208], stage0_20[209], stage0_20[210], stage0_20[211]},
      {stage0_22[153], stage0_22[154], stage0_22[155], stage0_22[156], stage0_22[157], stage0_22[158]},
      {stage1_24[31],stage1_23[72],stage1_22[72],stage1_21[104],stage1_20[175]}
   );
   gpc606_5 gpc808 (
      {stage0_20[212], stage0_20[213], stage0_20[214], stage0_20[215], stage0_20[216], stage0_20[217]},
      {stage0_22[159], stage0_22[160], stage0_22[161], stage0_22[162], stage0_22[163], stage0_22[164]},
      {stage1_24[32],stage1_23[73],stage1_22[73],stage1_21[105],stage1_20[176]}
   );
   gpc606_5 gpc809 (
      {stage0_20[218], stage0_20[219], stage0_20[220], stage0_20[221], stage0_20[222], stage0_20[223]},
      {stage0_22[165], stage0_22[166], stage0_22[167], stage0_22[168], stage0_22[169], stage0_22[170]},
      {stage1_24[33],stage1_23[74],stage1_22[74],stage1_21[106],stage1_20[177]}
   );
   gpc606_5 gpc810 (
      {stage0_20[224], stage0_20[225], stage0_20[226], stage0_20[227], stage0_20[228], stage0_20[229]},
      {stage0_22[171], stage0_22[172], stage0_22[173], stage0_22[174], stage0_22[175], stage0_22[176]},
      {stage1_24[34],stage1_23[75],stage1_22[75],stage1_21[107],stage1_20[178]}
   );
   gpc606_5 gpc811 (
      {stage0_20[230], stage0_20[231], stage0_20[232], stage0_20[233], stage0_20[234], stage0_20[235]},
      {stage0_22[177], stage0_22[178], stage0_22[179], stage0_22[180], stage0_22[181], stage0_22[182]},
      {stage1_24[35],stage1_23[76],stage1_22[76],stage1_21[108],stage1_20[179]}
   );
   gpc606_5 gpc812 (
      {stage0_20[236], stage0_20[237], stage0_20[238], stage0_20[239], stage0_20[240], stage0_20[241]},
      {stage0_22[183], stage0_22[184], stage0_22[185], stage0_22[186], stage0_22[187], stage0_22[188]},
      {stage1_24[36],stage1_23[77],stage1_22[77],stage1_21[109],stage1_20[180]}
   );
   gpc606_5 gpc813 (
      {stage0_20[242], stage0_20[243], stage0_20[244], stage0_20[245], stage0_20[246], stage0_20[247]},
      {stage0_22[189], stage0_22[190], stage0_22[191], stage0_22[192], stage0_22[193], stage0_22[194]},
      {stage1_24[37],stage1_23[78],stage1_22[78],stage1_21[110],stage1_20[181]}
   );
   gpc606_5 gpc814 (
      {stage0_20[248], stage0_20[249], stage0_20[250], stage0_20[251], stage0_20[252], stage0_20[253]},
      {stage0_22[195], stage0_22[196], stage0_22[197], stage0_22[198], stage0_22[199], stage0_22[200]},
      {stage1_24[38],stage1_23[79],stage1_22[79],stage1_21[111],stage1_20[182]}
   );
   gpc606_5 gpc815 (
      {stage0_20[254], stage0_20[255], stage0_20[256], stage0_20[257], stage0_20[258], stage0_20[259]},
      {stage0_22[201], stage0_22[202], stage0_22[203], stage0_22[204], stage0_22[205], stage0_22[206]},
      {stage1_24[39],stage1_23[80],stage1_22[80],stage1_21[112],stage1_20[183]}
   );
   gpc606_5 gpc816 (
      {stage0_20[260], stage0_20[261], stage0_20[262], stage0_20[263], stage0_20[264], stage0_20[265]},
      {stage0_22[207], stage0_22[208], stage0_22[209], stage0_22[210], stage0_22[211], stage0_22[212]},
      {stage1_24[40],stage1_23[81],stage1_22[81],stage1_21[113],stage1_20[184]}
   );
   gpc606_5 gpc817 (
      {stage0_20[266], stage0_20[267], stage0_20[268], stage0_20[269], stage0_20[270], stage0_20[271]},
      {stage0_22[213], stage0_22[214], stage0_22[215], stage0_22[216], stage0_22[217], stage0_22[218]},
      {stage1_24[41],stage1_23[82],stage1_22[82],stage1_21[114],stage1_20[185]}
   );
   gpc606_5 gpc818 (
      {stage0_20[272], stage0_20[273], stage0_20[274], stage0_20[275], stage0_20[276], stage0_20[277]},
      {stage0_22[219], stage0_22[220], stage0_22[221], stage0_22[222], stage0_22[223], stage0_22[224]},
      {stage1_24[42],stage1_23[83],stage1_22[83],stage1_21[115],stage1_20[186]}
   );
   gpc606_5 gpc819 (
      {stage0_20[278], stage0_20[279], stage0_20[280], stage0_20[281], stage0_20[282], stage0_20[283]},
      {stage0_22[225], stage0_22[226], stage0_22[227], stage0_22[228], stage0_22[229], stage0_22[230]},
      {stage1_24[43],stage1_23[84],stage1_22[84],stage1_21[116],stage1_20[187]}
   );
   gpc606_5 gpc820 (
      {stage0_20[284], stage0_20[285], stage0_20[286], stage0_20[287], stage0_20[288], stage0_20[289]},
      {stage0_22[231], stage0_22[232], stage0_22[233], stage0_22[234], stage0_22[235], stage0_22[236]},
      {stage1_24[44],stage1_23[85],stage1_22[85],stage1_21[117],stage1_20[188]}
   );
   gpc606_5 gpc821 (
      {stage0_20[290], stage0_20[291], stage0_20[292], stage0_20[293], stage0_20[294], stage0_20[295]},
      {stage0_22[237], stage0_22[238], stage0_22[239], stage0_22[240], stage0_22[241], stage0_22[242]},
      {stage1_24[45],stage1_23[86],stage1_22[86],stage1_21[118],stage1_20[189]}
   );
   gpc606_5 gpc822 (
      {stage0_20[296], stage0_20[297], stage0_20[298], stage0_20[299], stage0_20[300], stage0_20[301]},
      {stage0_22[243], stage0_22[244], stage0_22[245], stage0_22[246], stage0_22[247], stage0_22[248]},
      {stage1_24[46],stage1_23[87],stage1_22[87],stage1_21[119],stage1_20[190]}
   );
   gpc606_5 gpc823 (
      {stage0_20[302], stage0_20[303], stage0_20[304], stage0_20[305], stage0_20[306], stage0_20[307]},
      {stage0_22[249], stage0_22[250], stage0_22[251], stage0_22[252], stage0_22[253], stage0_22[254]},
      {stage1_24[47],stage1_23[88],stage1_22[88],stage1_21[120],stage1_20[191]}
   );
   gpc606_5 gpc824 (
      {stage0_20[308], stage0_20[309], stage0_20[310], stage0_20[311], stage0_20[312], stage0_20[313]},
      {stage0_22[255], stage0_22[256], stage0_22[257], stage0_22[258], stage0_22[259], stage0_22[260]},
      {stage1_24[48],stage1_23[89],stage1_22[89],stage1_21[121],stage1_20[192]}
   );
   gpc606_5 gpc825 (
      {stage0_20[314], stage0_20[315], stage0_20[316], stage0_20[317], stage0_20[318], stage0_20[319]},
      {stage0_22[261], stage0_22[262], stage0_22[263], stage0_22[264], stage0_22[265], stage0_22[266]},
      {stage1_24[49],stage1_23[90],stage1_22[90],stage1_21[122],stage1_20[193]}
   );
   gpc606_5 gpc826 (
      {stage0_20[320], stage0_20[321], stage0_20[322], stage0_20[323], stage0_20[324], stage0_20[325]},
      {stage0_22[267], stage0_22[268], stage0_22[269], stage0_22[270], stage0_22[271], stage0_22[272]},
      {stage1_24[50],stage1_23[91],stage1_22[91],stage1_21[123],stage1_20[194]}
   );
   gpc606_5 gpc827 (
      {stage0_20[326], stage0_20[327], stage0_20[328], stage0_20[329], stage0_20[330], stage0_20[331]},
      {stage0_22[273], stage0_22[274], stage0_22[275], stage0_22[276], stage0_22[277], stage0_22[278]},
      {stage1_24[51],stage1_23[92],stage1_22[92],stage1_21[124],stage1_20[195]}
   );
   gpc606_5 gpc828 (
      {stage0_20[332], stage0_20[333], stage0_20[334], stage0_20[335], stage0_20[336], stage0_20[337]},
      {stage0_22[279], stage0_22[280], stage0_22[281], stage0_22[282], stage0_22[283], stage0_22[284]},
      {stage1_24[52],stage1_23[93],stage1_22[93],stage1_21[125],stage1_20[196]}
   );
   gpc606_5 gpc829 (
      {stage0_20[338], stage0_20[339], stage0_20[340], stage0_20[341], stage0_20[342], stage0_20[343]},
      {stage0_22[285], stage0_22[286], stage0_22[287], stage0_22[288], stage0_22[289], stage0_22[290]},
      {stage1_24[53],stage1_23[94],stage1_22[94],stage1_21[126],stage1_20[197]}
   );
   gpc606_5 gpc830 (
      {stage0_20[344], stage0_20[345], stage0_20[346], stage0_20[347], stage0_20[348], stage0_20[349]},
      {stage0_22[291], stage0_22[292], stage0_22[293], stage0_22[294], stage0_22[295], stage0_22[296]},
      {stage1_24[54],stage1_23[95],stage1_22[95],stage1_21[127],stage1_20[198]}
   );
   gpc606_5 gpc831 (
      {stage0_20[350], stage0_20[351], stage0_20[352], stage0_20[353], stage0_20[354], stage0_20[355]},
      {stage0_22[297], stage0_22[298], stage0_22[299], stage0_22[300], stage0_22[301], stage0_22[302]},
      {stage1_24[55],stage1_23[96],stage1_22[96],stage1_21[128],stage1_20[199]}
   );
   gpc606_5 gpc832 (
      {stage0_20[356], stage0_20[357], stage0_20[358], stage0_20[359], stage0_20[360], stage0_20[361]},
      {stage0_22[303], stage0_22[304], stage0_22[305], stage0_22[306], stage0_22[307], stage0_22[308]},
      {stage1_24[56],stage1_23[97],stage1_22[97],stage1_21[129],stage1_20[200]}
   );
   gpc606_5 gpc833 (
      {stage0_20[362], stage0_20[363], stage0_20[364], stage0_20[365], stage0_20[366], stage0_20[367]},
      {stage0_22[309], stage0_22[310], stage0_22[311], stage0_22[312], stage0_22[313], stage0_22[314]},
      {stage1_24[57],stage1_23[98],stage1_22[98],stage1_21[130],stage1_20[201]}
   );
   gpc606_5 gpc834 (
      {stage0_20[368], stage0_20[369], stage0_20[370], stage0_20[371], stage0_20[372], stage0_20[373]},
      {stage0_22[315], stage0_22[316], stage0_22[317], stage0_22[318], stage0_22[319], stage0_22[320]},
      {stage1_24[58],stage1_23[99],stage1_22[99],stage1_21[131],stage1_20[202]}
   );
   gpc606_5 gpc835 (
      {stage0_20[374], stage0_20[375], stage0_20[376], stage0_20[377], stage0_20[378], stage0_20[379]},
      {stage0_22[321], stage0_22[322], stage0_22[323], stage0_22[324], stage0_22[325], stage0_22[326]},
      {stage1_24[59],stage1_23[100],stage1_22[100],stage1_21[132],stage1_20[203]}
   );
   gpc606_5 gpc836 (
      {stage0_20[380], stage0_20[381], stage0_20[382], stage0_20[383], stage0_20[384], stage0_20[385]},
      {stage0_22[327], stage0_22[328], stage0_22[329], stage0_22[330], stage0_22[331], stage0_22[332]},
      {stage1_24[60],stage1_23[101],stage1_22[101],stage1_21[133],stage1_20[204]}
   );
   gpc606_5 gpc837 (
      {stage0_20[386], stage0_20[387], stage0_20[388], stage0_20[389], stage0_20[390], stage0_20[391]},
      {stage0_22[333], stage0_22[334], stage0_22[335], stage0_22[336], stage0_22[337], stage0_22[338]},
      {stage1_24[61],stage1_23[102],stage1_22[102],stage1_21[134],stage1_20[205]}
   );
   gpc615_5 gpc838 (
      {stage0_20[392], stage0_20[393], stage0_20[394], stage0_20[395], stage0_20[396]},
      {stage0_21[286]},
      {stage0_22[339], stage0_22[340], stage0_22[341], stage0_22[342], stage0_22[343], stage0_22[344]},
      {stage1_24[62],stage1_23[103],stage1_22[103],stage1_21[135],stage1_20[206]}
   );
   gpc615_5 gpc839 (
      {stage0_20[397], stage0_20[398], stage0_20[399], stage0_20[400], stage0_20[401]},
      {stage0_21[287]},
      {stage0_22[345], stage0_22[346], stage0_22[347], stage0_22[348], stage0_22[349], stage0_22[350]},
      {stage1_24[63],stage1_23[104],stage1_22[104],stage1_21[136],stage1_20[207]}
   );
   gpc615_5 gpc840 (
      {stage0_20[402], stage0_20[403], stage0_20[404], stage0_20[405], stage0_20[406]},
      {stage0_21[288]},
      {stage0_22[351], stage0_22[352], stage0_22[353], stage0_22[354], stage0_22[355], stage0_22[356]},
      {stage1_24[64],stage1_23[105],stage1_22[105],stage1_21[137],stage1_20[208]}
   );
   gpc615_5 gpc841 (
      {stage0_20[407], stage0_20[408], stage0_20[409], stage0_20[410], stage0_20[411]},
      {stage0_21[289]},
      {stage0_22[357], stage0_22[358], stage0_22[359], stage0_22[360], stage0_22[361], stage0_22[362]},
      {stage1_24[65],stage1_23[106],stage1_22[106],stage1_21[138],stage1_20[209]}
   );
   gpc615_5 gpc842 (
      {stage0_20[412], stage0_20[413], stage0_20[414], stage0_20[415], stage0_20[416]},
      {stage0_21[290]},
      {stage0_22[363], stage0_22[364], stage0_22[365], stage0_22[366], stage0_22[367], stage0_22[368]},
      {stage1_24[66],stage1_23[107],stage1_22[107],stage1_21[139],stage1_20[210]}
   );
   gpc615_5 gpc843 (
      {stage0_20[417], stage0_20[418], stage0_20[419], stage0_20[420], stage0_20[421]},
      {stage0_21[291]},
      {stage0_22[369], stage0_22[370], stage0_22[371], stage0_22[372], stage0_22[373], stage0_22[374]},
      {stage1_24[67],stage1_23[108],stage1_22[108],stage1_21[140],stage1_20[211]}
   );
   gpc615_5 gpc844 (
      {stage0_20[422], stage0_20[423], stage0_20[424], stage0_20[425], stage0_20[426]},
      {stage0_21[292]},
      {stage0_22[375], stage0_22[376], stage0_22[377], stage0_22[378], stage0_22[379], stage0_22[380]},
      {stage1_24[68],stage1_23[109],stage1_22[109],stage1_21[141],stage1_20[212]}
   );
   gpc615_5 gpc845 (
      {stage0_20[427], stage0_20[428], stage0_20[429], stage0_20[430], stage0_20[431]},
      {stage0_21[293]},
      {stage0_22[381], stage0_22[382], stage0_22[383], stage0_22[384], stage0_22[385], stage0_22[386]},
      {stage1_24[69],stage1_23[110],stage1_22[110],stage1_21[142],stage1_20[213]}
   );
   gpc606_5 gpc846 (
      {stage0_21[294], stage0_21[295], stage0_21[296], stage0_21[297], stage0_21[298], stage0_21[299]},
      {stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11], stage0_23[12]},
      {stage1_25[0],stage1_24[70],stage1_23[111],stage1_22[111],stage1_21[143]}
   );
   gpc606_5 gpc847 (
      {stage0_21[300], stage0_21[301], stage0_21[302], stage0_21[303], stage0_21[304], stage0_21[305]},
      {stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17], stage0_23[18]},
      {stage1_25[1],stage1_24[71],stage1_23[112],stage1_22[112],stage1_21[144]}
   );
   gpc606_5 gpc848 (
      {stage0_21[306], stage0_21[307], stage0_21[308], stage0_21[309], stage0_21[310], stage0_21[311]},
      {stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23], stage0_23[24]},
      {stage1_25[2],stage1_24[72],stage1_23[113],stage1_22[113],stage1_21[145]}
   );
   gpc606_5 gpc849 (
      {stage0_21[312], stage0_21[313], stage0_21[314], stage0_21[315], stage0_21[316], stage0_21[317]},
      {stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29], stage0_23[30]},
      {stage1_25[3],stage1_24[73],stage1_23[114],stage1_22[114],stage1_21[146]}
   );
   gpc606_5 gpc850 (
      {stage0_21[318], stage0_21[319], stage0_21[320], stage0_21[321], stage0_21[322], stage0_21[323]},
      {stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35], stage0_23[36]},
      {stage1_25[4],stage1_24[74],stage1_23[115],stage1_22[115],stage1_21[147]}
   );
   gpc606_5 gpc851 (
      {stage0_21[324], stage0_21[325], stage0_21[326], stage0_21[327], stage0_21[328], stage0_21[329]},
      {stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41], stage0_23[42]},
      {stage1_25[5],stage1_24[75],stage1_23[116],stage1_22[116],stage1_21[148]}
   );
   gpc606_5 gpc852 (
      {stage0_21[330], stage0_21[331], stage0_21[332], stage0_21[333], stage0_21[334], stage0_21[335]},
      {stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47], stage0_23[48]},
      {stage1_25[6],stage1_24[76],stage1_23[117],stage1_22[117],stage1_21[149]}
   );
   gpc606_5 gpc853 (
      {stage0_21[336], stage0_21[337], stage0_21[338], stage0_21[339], stage0_21[340], stage0_21[341]},
      {stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53], stage0_23[54]},
      {stage1_25[7],stage1_24[77],stage1_23[118],stage1_22[118],stage1_21[150]}
   );
   gpc606_5 gpc854 (
      {stage0_21[342], stage0_21[343], stage0_21[344], stage0_21[345], stage0_21[346], stage0_21[347]},
      {stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59], stage0_23[60]},
      {stage1_25[8],stage1_24[78],stage1_23[119],stage1_22[119],stage1_21[151]}
   );
   gpc606_5 gpc855 (
      {stage0_21[348], stage0_21[349], stage0_21[350], stage0_21[351], stage0_21[352], stage0_21[353]},
      {stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65], stage0_23[66]},
      {stage1_25[9],stage1_24[79],stage1_23[120],stage1_22[120],stage1_21[152]}
   );
   gpc606_5 gpc856 (
      {stage0_21[354], stage0_21[355], stage0_21[356], stage0_21[357], stage0_21[358], stage0_21[359]},
      {stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71], stage0_23[72]},
      {stage1_25[10],stage1_24[80],stage1_23[121],stage1_22[121],stage1_21[153]}
   );
   gpc606_5 gpc857 (
      {stage0_21[360], stage0_21[361], stage0_21[362], stage0_21[363], stage0_21[364], stage0_21[365]},
      {stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77], stage0_23[78]},
      {stage1_25[11],stage1_24[81],stage1_23[122],stage1_22[122],stage1_21[154]}
   );
   gpc606_5 gpc858 (
      {stage0_21[366], stage0_21[367], stage0_21[368], stage0_21[369], stage0_21[370], stage0_21[371]},
      {stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83], stage0_23[84]},
      {stage1_25[12],stage1_24[82],stage1_23[123],stage1_22[123],stage1_21[155]}
   );
   gpc606_5 gpc859 (
      {stage0_21[372], stage0_21[373], stage0_21[374], stage0_21[375], stage0_21[376], stage0_21[377]},
      {stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89], stage0_23[90]},
      {stage1_25[13],stage1_24[83],stage1_23[124],stage1_22[124],stage1_21[156]}
   );
   gpc606_5 gpc860 (
      {stage0_21[378], stage0_21[379], stage0_21[380], stage0_21[381], stage0_21[382], stage0_21[383]},
      {stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95], stage0_23[96]},
      {stage1_25[14],stage1_24[84],stage1_23[125],stage1_22[125],stage1_21[157]}
   );
   gpc606_5 gpc861 (
      {stage0_21[384], stage0_21[385], stage0_21[386], stage0_21[387], stage0_21[388], stage0_21[389]},
      {stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101], stage0_23[102]},
      {stage1_25[15],stage1_24[85],stage1_23[126],stage1_22[126],stage1_21[158]}
   );
   gpc606_5 gpc862 (
      {stage0_21[390], stage0_21[391], stage0_21[392], stage0_21[393], stage0_21[394], stage0_21[395]},
      {stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107], stage0_23[108]},
      {stage1_25[16],stage1_24[86],stage1_23[127],stage1_22[127],stage1_21[159]}
   );
   gpc606_5 gpc863 (
      {stage0_21[396], stage0_21[397], stage0_21[398], stage0_21[399], stage0_21[400], stage0_21[401]},
      {stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113], stage0_23[114]},
      {stage1_25[17],stage1_24[87],stage1_23[128],stage1_22[128],stage1_21[160]}
   );
   gpc606_5 gpc864 (
      {stage0_21[402], stage0_21[403], stage0_21[404], stage0_21[405], stage0_21[406], stage0_21[407]},
      {stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119], stage0_23[120]},
      {stage1_25[18],stage1_24[88],stage1_23[129],stage1_22[129],stage1_21[161]}
   );
   gpc606_5 gpc865 (
      {stage0_21[408], stage0_21[409], stage0_21[410], stage0_21[411], stage0_21[412], stage0_21[413]},
      {stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125], stage0_23[126]},
      {stage1_25[19],stage1_24[89],stage1_23[130],stage1_22[130],stage1_21[162]}
   );
   gpc606_5 gpc866 (
      {stage0_21[414], stage0_21[415], stage0_21[416], stage0_21[417], stage0_21[418], stage0_21[419]},
      {stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131], stage0_23[132]},
      {stage1_25[20],stage1_24[90],stage1_23[131],stage1_22[131],stage1_21[163]}
   );
   gpc606_5 gpc867 (
      {stage0_21[420], stage0_21[421], stage0_21[422], stage0_21[423], stage0_21[424], stage0_21[425]},
      {stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137], stage0_23[138]},
      {stage1_25[21],stage1_24[91],stage1_23[132],stage1_22[132],stage1_21[164]}
   );
   gpc606_5 gpc868 (
      {stage0_21[426], stage0_21[427], stage0_21[428], stage0_21[429], stage0_21[430], stage0_21[431]},
      {stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143], stage0_23[144]},
      {stage1_25[22],stage1_24[92],stage1_23[133],stage1_22[133],stage1_21[165]}
   );
   gpc606_5 gpc869 (
      {stage0_21[432], stage0_21[433], stage0_21[434], stage0_21[435], stage0_21[436], stage0_21[437]},
      {stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149], stage0_23[150]},
      {stage1_25[23],stage1_24[93],stage1_23[134],stage1_22[134],stage1_21[166]}
   );
   gpc606_5 gpc870 (
      {stage0_21[438], stage0_21[439], stage0_21[440], stage0_21[441], stage0_21[442], stage0_21[443]},
      {stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155], stage0_23[156]},
      {stage1_25[24],stage1_24[94],stage1_23[135],stage1_22[135],stage1_21[167]}
   );
   gpc606_5 gpc871 (
      {stage0_21[444], stage0_21[445], stage0_21[446], stage0_21[447], stage0_21[448], stage0_21[449]},
      {stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161], stage0_23[162]},
      {stage1_25[25],stage1_24[95],stage1_23[136],stage1_22[136],stage1_21[168]}
   );
   gpc606_5 gpc872 (
      {stage0_21[450], stage0_21[451], stage0_21[452], stage0_21[453], stage0_21[454], stage0_21[455]},
      {stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167], stage0_23[168]},
      {stage1_25[26],stage1_24[96],stage1_23[137],stage1_22[137],stage1_21[169]}
   );
   gpc606_5 gpc873 (
      {stage0_21[456], stage0_21[457], stage0_21[458], stage0_21[459], stage0_21[460], stage0_21[461]},
      {stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173], stage0_23[174]},
      {stage1_25[27],stage1_24[97],stage1_23[138],stage1_22[138],stage1_21[170]}
   );
   gpc606_5 gpc874 (
      {stage0_21[462], stage0_21[463], stage0_21[464], stage0_21[465], stage0_21[466], stage0_21[467]},
      {stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179], stage0_23[180]},
      {stage1_25[28],stage1_24[98],stage1_23[139],stage1_22[139],stage1_21[171]}
   );
   gpc615_5 gpc875 (
      {stage0_22[387], stage0_22[388], stage0_22[389], stage0_22[390], stage0_22[391]},
      {stage0_23[181]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[29],stage1_24[99],stage1_23[140],stage1_22[140]}
   );
   gpc615_5 gpc876 (
      {stage0_22[392], stage0_22[393], stage0_22[394], stage0_22[395], stage0_22[396]},
      {stage0_23[182]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[30],stage1_24[100],stage1_23[141],stage1_22[141]}
   );
   gpc615_5 gpc877 (
      {stage0_22[397], stage0_22[398], stage0_22[399], stage0_22[400], stage0_22[401]},
      {stage0_23[183]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[31],stage1_24[101],stage1_23[142],stage1_22[142]}
   );
   gpc615_5 gpc878 (
      {stage0_22[402], stage0_22[403], stage0_22[404], stage0_22[405], stage0_22[406]},
      {stage0_23[184]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[32],stage1_24[102],stage1_23[143],stage1_22[143]}
   );
   gpc615_5 gpc879 (
      {stage0_22[407], stage0_22[408], stage0_22[409], stage0_22[410], stage0_22[411]},
      {stage0_23[185]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[33],stage1_24[103],stage1_23[144],stage1_22[144]}
   );
   gpc615_5 gpc880 (
      {stage0_22[412], stage0_22[413], stage0_22[414], stage0_22[415], stage0_22[416]},
      {stage0_23[186]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[34],stage1_24[104],stage1_23[145],stage1_22[145]}
   );
   gpc615_5 gpc881 (
      {stage0_22[417], stage0_22[418], stage0_22[419], stage0_22[420], stage0_22[421]},
      {stage0_23[187]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[35],stage1_24[105],stage1_23[146],stage1_22[146]}
   );
   gpc615_5 gpc882 (
      {stage0_22[422], stage0_22[423], stage0_22[424], stage0_22[425], stage0_22[426]},
      {stage0_23[188]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[36],stage1_24[106],stage1_23[147],stage1_22[147]}
   );
   gpc615_5 gpc883 (
      {stage0_22[427], stage0_22[428], stage0_22[429], stage0_22[430], stage0_22[431]},
      {stage0_23[189]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[37],stage1_24[107],stage1_23[148],stage1_22[148]}
   );
   gpc615_5 gpc884 (
      {stage0_22[432], stage0_22[433], stage0_22[434], stage0_22[435], stage0_22[436]},
      {stage0_23[190]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[38],stage1_24[108],stage1_23[149],stage1_22[149]}
   );
   gpc615_5 gpc885 (
      {stage0_22[437], stage0_22[438], stage0_22[439], stage0_22[440], stage0_22[441]},
      {stage0_23[191]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[39],stage1_24[109],stage1_23[150],stage1_22[150]}
   );
   gpc615_5 gpc886 (
      {stage0_22[442], stage0_22[443], stage0_22[444], stage0_22[445], stage0_22[446]},
      {stage0_23[192]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[40],stage1_24[110],stage1_23[151],stage1_22[151]}
   );
   gpc615_5 gpc887 (
      {stage0_22[447], stage0_22[448], stage0_22[449], stage0_22[450], stage0_22[451]},
      {stage0_23[193]},
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage1_26[12],stage1_25[41],stage1_24[111],stage1_23[152],stage1_22[152]}
   );
   gpc615_5 gpc888 (
      {stage0_22[452], stage0_22[453], stage0_22[454], stage0_22[455], stage0_22[456]},
      {stage0_23[194]},
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage1_26[13],stage1_25[42],stage1_24[112],stage1_23[153],stage1_22[153]}
   );
   gpc615_5 gpc889 (
      {stage0_22[457], stage0_22[458], stage0_22[459], stage0_22[460], stage0_22[461]},
      {stage0_23[195]},
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage1_26[14],stage1_25[43],stage1_24[113],stage1_23[154],stage1_22[154]}
   );
   gpc615_5 gpc890 (
      {stage0_22[462], stage0_22[463], stage0_22[464], stage0_22[465], stage0_22[466]},
      {stage0_23[196]},
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage1_26[15],stage1_25[44],stage1_24[114],stage1_23[155],stage1_22[155]}
   );
   gpc615_5 gpc891 (
      {stage0_22[467], stage0_22[468], stage0_22[469], stage0_22[470], stage0_22[471]},
      {stage0_23[197]},
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage1_26[16],stage1_25[45],stage1_24[115],stage1_23[156],stage1_22[156]}
   );
   gpc615_5 gpc892 (
      {stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202]},
      {stage0_24[102]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[17],stage1_25[46],stage1_24[116],stage1_23[157]}
   );
   gpc615_5 gpc893 (
      {stage0_23[203], stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207]},
      {stage0_24[103]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[18],stage1_25[47],stage1_24[117],stage1_23[158]}
   );
   gpc615_5 gpc894 (
      {stage0_23[208], stage0_23[209], stage0_23[210], stage0_23[211], stage0_23[212]},
      {stage0_24[104]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[19],stage1_25[48],stage1_24[118],stage1_23[159]}
   );
   gpc615_5 gpc895 (
      {stage0_23[213], stage0_23[214], stage0_23[215], stage0_23[216], stage0_23[217]},
      {stage0_24[105]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[20],stage1_25[49],stage1_24[119],stage1_23[160]}
   );
   gpc615_5 gpc896 (
      {stage0_23[218], stage0_23[219], stage0_23[220], stage0_23[221], stage0_23[222]},
      {stage0_24[106]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[21],stage1_25[50],stage1_24[120],stage1_23[161]}
   );
   gpc615_5 gpc897 (
      {stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226], stage0_23[227]},
      {stage0_24[107]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[22],stage1_25[51],stage1_24[121],stage1_23[162]}
   );
   gpc615_5 gpc898 (
      {stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232]},
      {stage0_24[108]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[23],stage1_25[52],stage1_24[122],stage1_23[163]}
   );
   gpc615_5 gpc899 (
      {stage0_23[233], stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237]},
      {stage0_24[109]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[24],stage1_25[53],stage1_24[123],stage1_23[164]}
   );
   gpc615_5 gpc900 (
      {stage0_23[238], stage0_23[239], stage0_23[240], stage0_23[241], stage0_23[242]},
      {stage0_24[110]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[25],stage1_25[54],stage1_24[124],stage1_23[165]}
   );
   gpc615_5 gpc901 (
      {stage0_23[243], stage0_23[244], stage0_23[245], stage0_23[246], stage0_23[247]},
      {stage0_24[111]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[26],stage1_25[55],stage1_24[125],stage1_23[166]}
   );
   gpc615_5 gpc902 (
      {stage0_23[248], stage0_23[249], stage0_23[250], stage0_23[251], stage0_23[252]},
      {stage0_24[112]},
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage1_27[10],stage1_26[27],stage1_25[56],stage1_24[126],stage1_23[167]}
   );
   gpc615_5 gpc903 (
      {stage0_23[253], stage0_23[254], stage0_23[255], stage0_23[256], stage0_23[257]},
      {stage0_24[113]},
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage1_27[11],stage1_26[28],stage1_25[57],stage1_24[127],stage1_23[168]}
   );
   gpc615_5 gpc904 (
      {stage0_23[258], stage0_23[259], stage0_23[260], stage0_23[261], stage0_23[262]},
      {stage0_24[114]},
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage1_27[12],stage1_26[29],stage1_25[58],stage1_24[128],stage1_23[169]}
   );
   gpc615_5 gpc905 (
      {stage0_23[263], stage0_23[264], stage0_23[265], stage0_23[266], stage0_23[267]},
      {stage0_24[115]},
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage1_27[13],stage1_26[30],stage1_25[59],stage1_24[129],stage1_23[170]}
   );
   gpc615_5 gpc906 (
      {stage0_23[268], stage0_23[269], stage0_23[270], stage0_23[271], stage0_23[272]},
      {stage0_24[116]},
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage1_27[14],stage1_26[31],stage1_25[60],stage1_24[130],stage1_23[171]}
   );
   gpc615_5 gpc907 (
      {stage0_23[273], stage0_23[274], stage0_23[275], stage0_23[276], stage0_23[277]},
      {stage0_24[117]},
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage1_27[15],stage1_26[32],stage1_25[61],stage1_24[131],stage1_23[172]}
   );
   gpc615_5 gpc908 (
      {stage0_23[278], stage0_23[279], stage0_23[280], stage0_23[281], stage0_23[282]},
      {stage0_24[118]},
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage1_27[16],stage1_26[33],stage1_25[62],stage1_24[132],stage1_23[173]}
   );
   gpc615_5 gpc909 (
      {stage0_23[283], stage0_23[284], stage0_23[285], stage0_23[286], stage0_23[287]},
      {stage0_24[119]},
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage1_27[17],stage1_26[34],stage1_25[63],stage1_24[133],stage1_23[174]}
   );
   gpc615_5 gpc910 (
      {stage0_23[288], stage0_23[289], stage0_23[290], stage0_23[291], stage0_23[292]},
      {stage0_24[120]},
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113]},
      {stage1_27[18],stage1_26[35],stage1_25[64],stage1_24[134],stage1_23[175]}
   );
   gpc615_5 gpc911 (
      {stage0_23[293], stage0_23[294], stage0_23[295], stage0_23[296], stage0_23[297]},
      {stage0_24[121]},
      {stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117], stage0_25[118], stage0_25[119]},
      {stage1_27[19],stage1_26[36],stage1_25[65],stage1_24[135],stage1_23[176]}
   );
   gpc615_5 gpc912 (
      {stage0_23[298], stage0_23[299], stage0_23[300], stage0_23[301], stage0_23[302]},
      {stage0_24[122]},
      {stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125]},
      {stage1_27[20],stage1_26[37],stage1_25[66],stage1_24[136],stage1_23[177]}
   );
   gpc615_5 gpc913 (
      {stage0_23[303], stage0_23[304], stage0_23[305], stage0_23[306], stage0_23[307]},
      {stage0_24[123]},
      {stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131]},
      {stage1_27[21],stage1_26[38],stage1_25[67],stage1_24[137],stage1_23[178]}
   );
   gpc615_5 gpc914 (
      {stage0_23[308], stage0_23[309], stage0_23[310], stage0_23[311], stage0_23[312]},
      {stage0_24[124]},
      {stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137]},
      {stage1_27[22],stage1_26[39],stage1_25[68],stage1_24[138],stage1_23[179]}
   );
   gpc615_5 gpc915 (
      {stage0_23[313], stage0_23[314], stage0_23[315], stage0_23[316], stage0_23[317]},
      {stage0_24[125]},
      {stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142], stage0_25[143]},
      {stage1_27[23],stage1_26[40],stage1_25[69],stage1_24[139],stage1_23[180]}
   );
   gpc615_5 gpc916 (
      {stage0_23[318], stage0_23[319], stage0_23[320], stage0_23[321], stage0_23[322]},
      {stage0_24[126]},
      {stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147], stage0_25[148], stage0_25[149]},
      {stage1_27[24],stage1_26[41],stage1_25[70],stage1_24[140],stage1_23[181]}
   );
   gpc615_5 gpc917 (
      {stage0_23[323], stage0_23[324], stage0_23[325], stage0_23[326], stage0_23[327]},
      {stage0_24[127]},
      {stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153], stage0_25[154], stage0_25[155]},
      {stage1_27[25],stage1_26[42],stage1_25[71],stage1_24[141],stage1_23[182]}
   );
   gpc615_5 gpc918 (
      {stage0_23[328], stage0_23[329], stage0_23[330], stage0_23[331], stage0_23[332]},
      {stage0_24[128]},
      {stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159], stage0_25[160], stage0_25[161]},
      {stage1_27[26],stage1_26[43],stage1_25[72],stage1_24[142],stage1_23[183]}
   );
   gpc615_5 gpc919 (
      {stage0_23[333], stage0_23[334], stage0_23[335], stage0_23[336], stage0_23[337]},
      {stage0_24[129]},
      {stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165], stage0_25[166], stage0_25[167]},
      {stage1_27[27],stage1_26[44],stage1_25[73],stage1_24[143],stage1_23[184]}
   );
   gpc615_5 gpc920 (
      {stage0_23[338], stage0_23[339], stage0_23[340], stage0_23[341], stage0_23[342]},
      {stage0_24[130]},
      {stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171], stage0_25[172], stage0_25[173]},
      {stage1_27[28],stage1_26[45],stage1_25[74],stage1_24[144],stage1_23[185]}
   );
   gpc615_5 gpc921 (
      {stage0_23[343], stage0_23[344], stage0_23[345], stage0_23[346], stage0_23[347]},
      {stage0_24[131]},
      {stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177], stage0_25[178], stage0_25[179]},
      {stage1_27[29],stage1_26[46],stage1_25[75],stage1_24[145],stage1_23[186]}
   );
   gpc615_5 gpc922 (
      {stage0_23[348], stage0_23[349], stage0_23[350], stage0_23[351], stage0_23[352]},
      {stage0_24[132]},
      {stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183], stage0_25[184], stage0_25[185]},
      {stage1_27[30],stage1_26[47],stage1_25[76],stage1_24[146],stage1_23[187]}
   );
   gpc615_5 gpc923 (
      {stage0_23[353], stage0_23[354], stage0_23[355], stage0_23[356], stage0_23[357]},
      {stage0_24[133]},
      {stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189], stage0_25[190], stage0_25[191]},
      {stage1_27[31],stage1_26[48],stage1_25[77],stage1_24[147],stage1_23[188]}
   );
   gpc615_5 gpc924 (
      {stage0_23[358], stage0_23[359], stage0_23[360], stage0_23[361], stage0_23[362]},
      {stage0_24[134]},
      {stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195], stage0_25[196], stage0_25[197]},
      {stage1_27[32],stage1_26[49],stage1_25[78],stage1_24[148],stage1_23[189]}
   );
   gpc615_5 gpc925 (
      {stage0_23[363], stage0_23[364], stage0_23[365], stage0_23[366], stage0_23[367]},
      {stage0_24[135]},
      {stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201], stage0_25[202], stage0_25[203]},
      {stage1_27[33],stage1_26[50],stage1_25[79],stage1_24[149],stage1_23[190]}
   );
   gpc615_5 gpc926 (
      {stage0_23[368], stage0_23[369], stage0_23[370], stage0_23[371], stage0_23[372]},
      {stage0_24[136]},
      {stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207], stage0_25[208], stage0_25[209]},
      {stage1_27[34],stage1_26[51],stage1_25[80],stage1_24[150],stage1_23[191]}
   );
   gpc615_5 gpc927 (
      {stage0_23[373], stage0_23[374], stage0_23[375], stage0_23[376], stage0_23[377]},
      {stage0_24[137]},
      {stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213], stage0_25[214], stage0_25[215]},
      {stage1_27[35],stage1_26[52],stage1_25[81],stage1_24[151],stage1_23[192]}
   );
   gpc615_5 gpc928 (
      {stage0_23[378], stage0_23[379], stage0_23[380], stage0_23[381], stage0_23[382]},
      {stage0_24[138]},
      {stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219], stage0_25[220], stage0_25[221]},
      {stage1_27[36],stage1_26[53],stage1_25[82],stage1_24[152],stage1_23[193]}
   );
   gpc615_5 gpc929 (
      {stage0_23[383], stage0_23[384], stage0_23[385], stage0_23[386], stage0_23[387]},
      {stage0_24[139]},
      {stage0_25[222], stage0_25[223], stage0_25[224], stage0_25[225], stage0_25[226], stage0_25[227]},
      {stage1_27[37],stage1_26[54],stage1_25[83],stage1_24[153],stage1_23[194]}
   );
   gpc615_5 gpc930 (
      {stage0_23[388], stage0_23[389], stage0_23[390], stage0_23[391], stage0_23[392]},
      {stage0_24[140]},
      {stage0_25[228], stage0_25[229], stage0_25[230], stage0_25[231], stage0_25[232], stage0_25[233]},
      {stage1_27[38],stage1_26[55],stage1_25[84],stage1_24[154],stage1_23[195]}
   );
   gpc623_5 gpc931 (
      {stage0_23[393], stage0_23[394], stage0_23[395]},
      {stage0_24[141], stage0_24[142]},
      {stage0_25[234], stage0_25[235], stage0_25[236], stage0_25[237], stage0_25[238], stage0_25[239]},
      {stage1_27[39],stage1_26[56],stage1_25[85],stage1_24[155],stage1_23[196]}
   );
   gpc606_5 gpc932 (
      {stage0_24[143], stage0_24[144], stage0_24[145], stage0_24[146], stage0_24[147], stage0_24[148]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[40],stage1_26[57],stage1_25[86],stage1_24[156]}
   );
   gpc606_5 gpc933 (
      {stage0_24[149], stage0_24[150], stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[41],stage1_26[58],stage1_25[87],stage1_24[157]}
   );
   gpc606_5 gpc934 (
      {stage0_24[155], stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[42],stage1_26[59],stage1_25[88],stage1_24[158]}
   );
   gpc606_5 gpc935 (
      {stage0_24[161], stage0_24[162], stage0_24[163], stage0_24[164], stage0_24[165], stage0_24[166]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[43],stage1_26[60],stage1_25[89],stage1_24[159]}
   );
   gpc606_5 gpc936 (
      {stage0_24[167], stage0_24[168], stage0_24[169], stage0_24[170], stage0_24[171], stage0_24[172]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[44],stage1_26[61],stage1_25[90],stage1_24[160]}
   );
   gpc606_5 gpc937 (
      {stage0_24[173], stage0_24[174], stage0_24[175], stage0_24[176], stage0_24[177], stage0_24[178]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[45],stage1_26[62],stage1_25[91],stage1_24[161]}
   );
   gpc606_5 gpc938 (
      {stage0_24[179], stage0_24[180], stage0_24[181], stage0_24[182], stage0_24[183], stage0_24[184]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[46],stage1_26[63],stage1_25[92],stage1_24[162]}
   );
   gpc606_5 gpc939 (
      {stage0_24[185], stage0_24[186], stage0_24[187], stage0_24[188], stage0_24[189], stage0_24[190]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[47],stage1_26[64],stage1_25[93],stage1_24[163]}
   );
   gpc606_5 gpc940 (
      {stage0_24[191], stage0_24[192], stage0_24[193], stage0_24[194], stage0_24[195], stage0_24[196]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[48],stage1_26[65],stage1_25[94],stage1_24[164]}
   );
   gpc606_5 gpc941 (
      {stage0_24[197], stage0_24[198], stage0_24[199], stage0_24[200], stage0_24[201], stage0_24[202]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[49],stage1_26[66],stage1_25[95],stage1_24[165]}
   );
   gpc606_5 gpc942 (
      {stage0_24[203], stage0_24[204], stage0_24[205], stage0_24[206], stage0_24[207], stage0_24[208]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[50],stage1_26[67],stage1_25[96],stage1_24[166]}
   );
   gpc606_5 gpc943 (
      {stage0_24[209], stage0_24[210], stage0_24[211], stage0_24[212], stage0_24[213], stage0_24[214]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[51],stage1_26[68],stage1_25[97],stage1_24[167]}
   );
   gpc606_5 gpc944 (
      {stage0_24[215], stage0_24[216], stage0_24[217], stage0_24[218], stage0_24[219], stage0_24[220]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[52],stage1_26[69],stage1_25[98],stage1_24[168]}
   );
   gpc606_5 gpc945 (
      {stage0_24[221], stage0_24[222], stage0_24[223], stage0_24[224], stage0_24[225], stage0_24[226]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[53],stage1_26[70],stage1_25[99],stage1_24[169]}
   );
   gpc606_5 gpc946 (
      {stage0_24[227], stage0_24[228], stage0_24[229], stage0_24[230], stage0_24[231], stage0_24[232]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[54],stage1_26[71],stage1_25[100],stage1_24[170]}
   );
   gpc606_5 gpc947 (
      {stage0_24[233], stage0_24[234], stage0_24[235], stage0_24[236], stage0_24[237], stage0_24[238]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[55],stage1_26[72],stage1_25[101],stage1_24[171]}
   );
   gpc606_5 gpc948 (
      {stage0_24[239], stage0_24[240], stage0_24[241], stage0_24[242], stage0_24[243], stage0_24[244]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[56],stage1_26[73],stage1_25[102],stage1_24[172]}
   );
   gpc606_5 gpc949 (
      {stage0_24[245], stage0_24[246], stage0_24[247], stage0_24[248], stage0_24[249], stage0_24[250]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[57],stage1_26[74],stage1_25[103],stage1_24[173]}
   );
   gpc606_5 gpc950 (
      {stage0_24[251], stage0_24[252], stage0_24[253], stage0_24[254], stage0_24[255], stage0_24[256]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[58],stage1_26[75],stage1_25[104],stage1_24[174]}
   );
   gpc606_5 gpc951 (
      {stage0_24[257], stage0_24[258], stage0_24[259], stage0_24[260], stage0_24[261], stage0_24[262]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[59],stage1_26[76],stage1_25[105],stage1_24[175]}
   );
   gpc606_5 gpc952 (
      {stage0_24[263], stage0_24[264], stage0_24[265], stage0_24[266], stage0_24[267], stage0_24[268]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[60],stage1_26[77],stage1_25[106],stage1_24[176]}
   );
   gpc606_5 gpc953 (
      {stage0_24[269], stage0_24[270], stage0_24[271], stage0_24[272], stage0_24[273], stage0_24[274]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[61],stage1_26[78],stage1_25[107],stage1_24[177]}
   );
   gpc606_5 gpc954 (
      {stage0_24[275], stage0_24[276], stage0_24[277], stage0_24[278], stage0_24[279], stage0_24[280]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[62],stage1_26[79],stage1_25[108],stage1_24[178]}
   );
   gpc606_5 gpc955 (
      {stage0_24[281], stage0_24[282], stage0_24[283], stage0_24[284], stage0_24[285], stage0_24[286]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[63],stage1_26[80],stage1_25[109],stage1_24[179]}
   );
   gpc606_5 gpc956 (
      {stage0_24[287], stage0_24[288], stage0_24[289], stage0_24[290], stage0_24[291], stage0_24[292]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[64],stage1_26[81],stage1_25[110],stage1_24[180]}
   );
   gpc606_5 gpc957 (
      {stage0_24[293], stage0_24[294], stage0_24[295], stage0_24[296], stage0_24[297], stage0_24[298]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[65],stage1_26[82],stage1_25[111],stage1_24[181]}
   );
   gpc606_5 gpc958 (
      {stage0_24[299], stage0_24[300], stage0_24[301], stage0_24[302], stage0_24[303], stage0_24[304]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[66],stage1_26[83],stage1_25[112],stage1_24[182]}
   );
   gpc606_5 gpc959 (
      {stage0_24[305], stage0_24[306], stage0_24[307], stage0_24[308], stage0_24[309], stage0_24[310]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[67],stage1_26[84],stage1_25[113],stage1_24[183]}
   );
   gpc606_5 gpc960 (
      {stage0_24[311], stage0_24[312], stage0_24[313], stage0_24[314], stage0_24[315], stage0_24[316]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[68],stage1_26[85],stage1_25[114],stage1_24[184]}
   );
   gpc606_5 gpc961 (
      {stage0_24[317], stage0_24[318], stage0_24[319], stage0_24[320], stage0_24[321], stage0_24[322]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[69],stage1_26[86],stage1_25[115],stage1_24[185]}
   );
   gpc606_5 gpc962 (
      {stage0_24[323], stage0_24[324], stage0_24[325], stage0_24[326], stage0_24[327], stage0_24[328]},
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184], stage0_26[185]},
      {stage1_28[30],stage1_27[70],stage1_26[87],stage1_25[116],stage1_24[186]}
   );
   gpc606_5 gpc963 (
      {stage0_24[329], stage0_24[330], stage0_24[331], stage0_24[332], stage0_24[333], stage0_24[334]},
      {stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189], stage0_26[190], stage0_26[191]},
      {stage1_28[31],stage1_27[71],stage1_26[88],stage1_25[117],stage1_24[187]}
   );
   gpc606_5 gpc964 (
      {stage0_24[335], stage0_24[336], stage0_24[337], stage0_24[338], stage0_24[339], stage0_24[340]},
      {stage0_26[192], stage0_26[193], stage0_26[194], stage0_26[195], stage0_26[196], stage0_26[197]},
      {stage1_28[32],stage1_27[72],stage1_26[89],stage1_25[118],stage1_24[188]}
   );
   gpc606_5 gpc965 (
      {stage0_24[341], stage0_24[342], stage0_24[343], stage0_24[344], stage0_24[345], stage0_24[346]},
      {stage0_26[198], stage0_26[199], stage0_26[200], stage0_26[201], stage0_26[202], stage0_26[203]},
      {stage1_28[33],stage1_27[73],stage1_26[90],stage1_25[119],stage1_24[189]}
   );
   gpc606_5 gpc966 (
      {stage0_24[347], stage0_24[348], stage0_24[349], stage0_24[350], stage0_24[351], stage0_24[352]},
      {stage0_26[204], stage0_26[205], stage0_26[206], stage0_26[207], stage0_26[208], stage0_26[209]},
      {stage1_28[34],stage1_27[74],stage1_26[91],stage1_25[120],stage1_24[190]}
   );
   gpc606_5 gpc967 (
      {stage0_24[353], stage0_24[354], stage0_24[355], stage0_24[356], stage0_24[357], stage0_24[358]},
      {stage0_26[210], stage0_26[211], stage0_26[212], stage0_26[213], stage0_26[214], stage0_26[215]},
      {stage1_28[35],stage1_27[75],stage1_26[92],stage1_25[121],stage1_24[191]}
   );
   gpc606_5 gpc968 (
      {stage0_24[359], stage0_24[360], stage0_24[361], stage0_24[362], stage0_24[363], stage0_24[364]},
      {stage0_26[216], stage0_26[217], stage0_26[218], stage0_26[219], stage0_26[220], stage0_26[221]},
      {stage1_28[36],stage1_27[76],stage1_26[93],stage1_25[122],stage1_24[192]}
   );
   gpc606_5 gpc969 (
      {stage0_24[365], stage0_24[366], stage0_24[367], stage0_24[368], stage0_24[369], stage0_24[370]},
      {stage0_26[222], stage0_26[223], stage0_26[224], stage0_26[225], stage0_26[226], stage0_26[227]},
      {stage1_28[37],stage1_27[77],stage1_26[94],stage1_25[123],stage1_24[193]}
   );
   gpc606_5 gpc970 (
      {stage0_24[371], stage0_24[372], stage0_24[373], stage0_24[374], stage0_24[375], stage0_24[376]},
      {stage0_26[228], stage0_26[229], stage0_26[230], stage0_26[231], stage0_26[232], stage0_26[233]},
      {stage1_28[38],stage1_27[78],stage1_26[95],stage1_25[124],stage1_24[194]}
   );
   gpc606_5 gpc971 (
      {stage0_24[377], stage0_24[378], stage0_24[379], stage0_24[380], stage0_24[381], stage0_24[382]},
      {stage0_26[234], stage0_26[235], stage0_26[236], stage0_26[237], stage0_26[238], stage0_26[239]},
      {stage1_28[39],stage1_27[79],stage1_26[96],stage1_25[125],stage1_24[195]}
   );
   gpc606_5 gpc972 (
      {stage0_24[383], stage0_24[384], stage0_24[385], stage0_24[386], stage0_24[387], stage0_24[388]},
      {stage0_26[240], stage0_26[241], stage0_26[242], stage0_26[243], stage0_26[244], stage0_26[245]},
      {stage1_28[40],stage1_27[80],stage1_26[97],stage1_25[126],stage1_24[196]}
   );
   gpc606_5 gpc973 (
      {stage0_24[389], stage0_24[390], stage0_24[391], stage0_24[392], stage0_24[393], stage0_24[394]},
      {stage0_26[246], stage0_26[247], stage0_26[248], stage0_26[249], stage0_26[250], stage0_26[251]},
      {stage1_28[41],stage1_27[81],stage1_26[98],stage1_25[127],stage1_24[197]}
   );
   gpc606_5 gpc974 (
      {stage0_24[395], stage0_24[396], stage0_24[397], stage0_24[398], stage0_24[399], stage0_24[400]},
      {stage0_26[252], stage0_26[253], stage0_26[254], stage0_26[255], stage0_26[256], stage0_26[257]},
      {stage1_28[42],stage1_27[82],stage1_26[99],stage1_25[128],stage1_24[198]}
   );
   gpc606_5 gpc975 (
      {stage0_24[401], stage0_24[402], stage0_24[403], stage0_24[404], stage0_24[405], stage0_24[406]},
      {stage0_26[258], stage0_26[259], stage0_26[260], stage0_26[261], stage0_26[262], stage0_26[263]},
      {stage1_28[43],stage1_27[83],stage1_26[100],stage1_25[129],stage1_24[199]}
   );
   gpc606_5 gpc976 (
      {stage0_24[407], stage0_24[408], stage0_24[409], stage0_24[410], stage0_24[411], stage0_24[412]},
      {stage0_26[264], stage0_26[265], stage0_26[266], stage0_26[267], stage0_26[268], stage0_26[269]},
      {stage1_28[44],stage1_27[84],stage1_26[101],stage1_25[130],stage1_24[200]}
   );
   gpc606_5 gpc977 (
      {stage0_24[413], stage0_24[414], stage0_24[415], stage0_24[416], stage0_24[417], stage0_24[418]},
      {stage0_26[270], stage0_26[271], stage0_26[272], stage0_26[273], stage0_26[274], stage0_26[275]},
      {stage1_28[45],stage1_27[85],stage1_26[102],stage1_25[131],stage1_24[201]}
   );
   gpc606_5 gpc978 (
      {stage0_24[419], stage0_24[420], stage0_24[421], stage0_24[422], stage0_24[423], stage0_24[424]},
      {stage0_26[276], stage0_26[277], stage0_26[278], stage0_26[279], stage0_26[280], stage0_26[281]},
      {stage1_28[46],stage1_27[86],stage1_26[103],stage1_25[132],stage1_24[202]}
   );
   gpc606_5 gpc979 (
      {stage0_24[425], stage0_24[426], stage0_24[427], stage0_24[428], stage0_24[429], stage0_24[430]},
      {stage0_26[282], stage0_26[283], stage0_26[284], stage0_26[285], stage0_26[286], stage0_26[287]},
      {stage1_28[47],stage1_27[87],stage1_26[104],stage1_25[133],stage1_24[203]}
   );
   gpc606_5 gpc980 (
      {stage0_24[431], stage0_24[432], stage0_24[433], stage0_24[434], stage0_24[435], stage0_24[436]},
      {stage0_26[288], stage0_26[289], stage0_26[290], stage0_26[291], stage0_26[292], stage0_26[293]},
      {stage1_28[48],stage1_27[88],stage1_26[105],stage1_25[134],stage1_24[204]}
   );
   gpc606_5 gpc981 (
      {stage0_24[437], stage0_24[438], stage0_24[439], stage0_24[440], stage0_24[441], stage0_24[442]},
      {stage0_26[294], stage0_26[295], stage0_26[296], stage0_26[297], stage0_26[298], stage0_26[299]},
      {stage1_28[49],stage1_27[89],stage1_26[106],stage1_25[135],stage1_24[205]}
   );
   gpc606_5 gpc982 (
      {stage0_24[443], stage0_24[444], stage0_24[445], stage0_24[446], stage0_24[447], stage0_24[448]},
      {stage0_26[300], stage0_26[301], stage0_26[302], stage0_26[303], stage0_26[304], stage0_26[305]},
      {stage1_28[50],stage1_27[90],stage1_26[107],stage1_25[136],stage1_24[206]}
   );
   gpc606_5 gpc983 (
      {stage0_24[449], stage0_24[450], stage0_24[451], stage0_24[452], stage0_24[453], stage0_24[454]},
      {stage0_26[306], stage0_26[307], stage0_26[308], stage0_26[309], stage0_26[310], stage0_26[311]},
      {stage1_28[51],stage1_27[91],stage1_26[108],stage1_25[137],stage1_24[207]}
   );
   gpc606_5 gpc984 (
      {stage0_24[455], stage0_24[456], stage0_24[457], stage0_24[458], stage0_24[459], stage0_24[460]},
      {stage0_26[312], stage0_26[313], stage0_26[314], stage0_26[315], stage0_26[316], stage0_26[317]},
      {stage1_28[52],stage1_27[92],stage1_26[109],stage1_25[138],stage1_24[208]}
   );
   gpc606_5 gpc985 (
      {stage0_24[461], stage0_24[462], stage0_24[463], stage0_24[464], stage0_24[465], stage0_24[466]},
      {stage0_26[318], stage0_26[319], stage0_26[320], stage0_26[321], stage0_26[322], stage0_26[323]},
      {stage1_28[53],stage1_27[93],stage1_26[110],stage1_25[139],stage1_24[209]}
   );
   gpc606_5 gpc986 (
      {stage0_24[467], stage0_24[468], stage0_24[469], stage0_24[470], stage0_24[471], stage0_24[472]},
      {stage0_26[324], stage0_26[325], stage0_26[326], stage0_26[327], stage0_26[328], stage0_26[329]},
      {stage1_28[54],stage1_27[94],stage1_26[111],stage1_25[140],stage1_24[210]}
   );
   gpc606_5 gpc987 (
      {stage0_24[473], stage0_24[474], stage0_24[475], stage0_24[476], stage0_24[477], stage0_24[478]},
      {stage0_26[330], stage0_26[331], stage0_26[332], stage0_26[333], stage0_26[334], stage0_26[335]},
      {stage1_28[55],stage1_27[95],stage1_26[112],stage1_25[141],stage1_24[211]}
   );
   gpc606_5 gpc988 (
      {stage0_24[479], stage0_24[480], stage0_24[481], stage0_24[482], stage0_24[483], stage0_24[484]},
      {stage0_26[336], stage0_26[337], stage0_26[338], stage0_26[339], stage0_26[340], stage0_26[341]},
      {stage1_28[56],stage1_27[96],stage1_26[113],stage1_25[142],stage1_24[212]}
   );
   gpc606_5 gpc989 (
      {stage0_25[240], stage0_25[241], stage0_25[242], stage0_25[243], stage0_25[244], stage0_25[245]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[57],stage1_27[97],stage1_26[114],stage1_25[143]}
   );
   gpc606_5 gpc990 (
      {stage0_25[246], stage0_25[247], stage0_25[248], stage0_25[249], stage0_25[250], stage0_25[251]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[58],stage1_27[98],stage1_26[115],stage1_25[144]}
   );
   gpc606_5 gpc991 (
      {stage0_25[252], stage0_25[253], stage0_25[254], stage0_25[255], stage0_25[256], stage0_25[257]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[59],stage1_27[99],stage1_26[116],stage1_25[145]}
   );
   gpc606_5 gpc992 (
      {stage0_25[258], stage0_25[259], stage0_25[260], stage0_25[261], stage0_25[262], stage0_25[263]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[60],stage1_27[100],stage1_26[117],stage1_25[146]}
   );
   gpc606_5 gpc993 (
      {stage0_25[264], stage0_25[265], stage0_25[266], stage0_25[267], stage0_25[268], stage0_25[269]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[61],stage1_27[101],stage1_26[118],stage1_25[147]}
   );
   gpc606_5 gpc994 (
      {stage0_25[270], stage0_25[271], stage0_25[272], stage0_25[273], stage0_25[274], stage0_25[275]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[62],stage1_27[102],stage1_26[119],stage1_25[148]}
   );
   gpc606_5 gpc995 (
      {stage0_25[276], stage0_25[277], stage0_25[278], stage0_25[279], stage0_25[280], stage0_25[281]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[63],stage1_27[103],stage1_26[120],stage1_25[149]}
   );
   gpc606_5 gpc996 (
      {stage0_25[282], stage0_25[283], stage0_25[284], stage0_25[285], stage0_25[286], stage0_25[287]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[64],stage1_27[104],stage1_26[121],stage1_25[150]}
   );
   gpc606_5 gpc997 (
      {stage0_25[288], stage0_25[289], stage0_25[290], stage0_25[291], stage0_25[292], stage0_25[293]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[65],stage1_27[105],stage1_26[122],stage1_25[151]}
   );
   gpc606_5 gpc998 (
      {stage0_25[294], stage0_25[295], stage0_25[296], stage0_25[297], stage0_25[298], stage0_25[299]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[66],stage1_27[106],stage1_26[123],stage1_25[152]}
   );
   gpc606_5 gpc999 (
      {stage0_25[300], stage0_25[301], stage0_25[302], stage0_25[303], stage0_25[304], stage0_25[305]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[67],stage1_27[107],stage1_26[124],stage1_25[153]}
   );
   gpc606_5 gpc1000 (
      {stage0_25[306], stage0_25[307], stage0_25[308], stage0_25[309], stage0_25[310], stage0_25[311]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[68],stage1_27[108],stage1_26[125],stage1_25[154]}
   );
   gpc606_5 gpc1001 (
      {stage0_25[312], stage0_25[313], stage0_25[314], stage0_25[315], stage0_25[316], stage0_25[317]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[69],stage1_27[109],stage1_26[126],stage1_25[155]}
   );
   gpc606_5 gpc1002 (
      {stage0_25[318], stage0_25[319], stage0_25[320], stage0_25[321], stage0_25[322], stage0_25[323]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[70],stage1_27[110],stage1_26[127],stage1_25[156]}
   );
   gpc606_5 gpc1003 (
      {stage0_25[324], stage0_25[325], stage0_25[326], stage0_25[327], stage0_25[328], stage0_25[329]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[71],stage1_27[111],stage1_26[128],stage1_25[157]}
   );
   gpc606_5 gpc1004 (
      {stage0_25[330], stage0_25[331], stage0_25[332], stage0_25[333], stage0_25[334], stage0_25[335]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[72],stage1_27[112],stage1_26[129],stage1_25[158]}
   );
   gpc606_5 gpc1005 (
      {stage0_25[336], stage0_25[337], stage0_25[338], stage0_25[339], stage0_25[340], stage0_25[341]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[73],stage1_27[113],stage1_26[130],stage1_25[159]}
   );
   gpc606_5 gpc1006 (
      {stage0_25[342], stage0_25[343], stage0_25[344], stage0_25[345], stage0_25[346], stage0_25[347]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[74],stage1_27[114],stage1_26[131],stage1_25[160]}
   );
   gpc606_5 gpc1007 (
      {stage0_25[348], stage0_25[349], stage0_25[350], stage0_25[351], stage0_25[352], stage0_25[353]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[75],stage1_27[115],stage1_26[132],stage1_25[161]}
   );
   gpc606_5 gpc1008 (
      {stage0_25[354], stage0_25[355], stage0_25[356], stage0_25[357], stage0_25[358], stage0_25[359]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[76],stage1_27[116],stage1_26[133],stage1_25[162]}
   );
   gpc606_5 gpc1009 (
      {stage0_25[360], stage0_25[361], stage0_25[362], stage0_25[363], stage0_25[364], stage0_25[365]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[77],stage1_27[117],stage1_26[134],stage1_25[163]}
   );
   gpc606_5 gpc1010 (
      {stage0_25[366], stage0_25[367], stage0_25[368], stage0_25[369], stage0_25[370], stage0_25[371]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[78],stage1_27[118],stage1_26[135],stage1_25[164]}
   );
   gpc606_5 gpc1011 (
      {stage0_25[372], stage0_25[373], stage0_25[374], stage0_25[375], stage0_25[376], stage0_25[377]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[79],stage1_27[119],stage1_26[136],stage1_25[165]}
   );
   gpc606_5 gpc1012 (
      {stage0_25[378], stage0_25[379], stage0_25[380], stage0_25[381], stage0_25[382], stage0_25[383]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[80],stage1_27[120],stage1_26[137],stage1_25[166]}
   );
   gpc606_5 gpc1013 (
      {stage0_25[384], stage0_25[385], stage0_25[386], stage0_25[387], stage0_25[388], stage0_25[389]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[81],stage1_27[121],stage1_26[138],stage1_25[167]}
   );
   gpc606_5 gpc1014 (
      {stage0_25[390], stage0_25[391], stage0_25[392], stage0_25[393], stage0_25[394], stage0_25[395]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[82],stage1_27[122],stage1_26[139],stage1_25[168]}
   );
   gpc606_5 gpc1015 (
      {stage0_25[396], stage0_25[397], stage0_25[398], stage0_25[399], stage0_25[400], stage0_25[401]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[83],stage1_27[123],stage1_26[140],stage1_25[169]}
   );
   gpc606_5 gpc1016 (
      {stage0_25[402], stage0_25[403], stage0_25[404], stage0_25[405], stage0_25[406], stage0_25[407]},
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage1_29[27],stage1_28[84],stage1_27[124],stage1_26[141],stage1_25[170]}
   );
   gpc606_5 gpc1017 (
      {stage0_25[408], stage0_25[409], stage0_25[410], stage0_25[411], stage0_25[412], stage0_25[413]},
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage1_29[28],stage1_28[85],stage1_27[125],stage1_26[142],stage1_25[171]}
   );
   gpc606_5 gpc1018 (
      {stage0_25[414], stage0_25[415], stage0_25[416], stage0_25[417], stage0_25[418], stage0_25[419]},
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage1_29[29],stage1_28[86],stage1_27[126],stage1_26[143],stage1_25[172]}
   );
   gpc606_5 gpc1019 (
      {stage0_25[420], stage0_25[421], stage0_25[422], stage0_25[423], stage0_25[424], stage0_25[425]},
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage1_29[30],stage1_28[87],stage1_27[127],stage1_26[144],stage1_25[173]}
   );
   gpc606_5 gpc1020 (
      {stage0_25[426], stage0_25[427], stage0_25[428], stage0_25[429], stage0_25[430], stage0_25[431]},
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage1_29[31],stage1_28[88],stage1_27[128],stage1_26[145],stage1_25[174]}
   );
   gpc606_5 gpc1021 (
      {stage0_25[432], stage0_25[433], stage0_25[434], stage0_25[435], stage0_25[436], stage0_25[437]},
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage1_29[32],stage1_28[89],stage1_27[129],stage1_26[146],stage1_25[175]}
   );
   gpc606_5 gpc1022 (
      {stage0_25[438], stage0_25[439], stage0_25[440], stage0_25[441], stage0_25[442], stage0_25[443]},
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage1_29[33],stage1_28[90],stage1_27[130],stage1_26[147],stage1_25[176]}
   );
   gpc606_5 gpc1023 (
      {stage0_25[444], stage0_25[445], stage0_25[446], stage0_25[447], stage0_25[448], stage0_25[449]},
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208], stage0_27[209]},
      {stage1_29[34],stage1_28[91],stage1_27[131],stage1_26[148],stage1_25[177]}
   );
   gpc606_5 gpc1024 (
      {stage0_25[450], stage0_25[451], stage0_25[452], stage0_25[453], stage0_25[454], stage0_25[455]},
      {stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213], stage0_27[214], stage0_27[215]},
      {stage1_29[35],stage1_28[92],stage1_27[132],stage1_26[149],stage1_25[178]}
   );
   gpc606_5 gpc1025 (
      {stage0_25[456], stage0_25[457], stage0_25[458], stage0_25[459], stage0_25[460], stage0_25[461]},
      {stage0_27[216], stage0_27[217], stage0_27[218], stage0_27[219], stage0_27[220], stage0_27[221]},
      {stage1_29[36],stage1_28[93],stage1_27[133],stage1_26[150],stage1_25[179]}
   );
   gpc606_5 gpc1026 (
      {stage0_25[462], stage0_25[463], stage0_25[464], stage0_25[465], stage0_25[466], stage0_25[467]},
      {stage0_27[222], stage0_27[223], stage0_27[224], stage0_27[225], stage0_27[226], stage0_27[227]},
      {stage1_29[37],stage1_28[94],stage1_27[134],stage1_26[151],stage1_25[180]}
   );
   gpc606_5 gpc1027 (
      {stage0_25[468], stage0_25[469], stage0_25[470], stage0_25[471], stage0_25[472], stage0_25[473]},
      {stage0_27[228], stage0_27[229], stage0_27[230], stage0_27[231], stage0_27[232], stage0_27[233]},
      {stage1_29[38],stage1_28[95],stage1_27[135],stage1_26[152],stage1_25[181]}
   );
   gpc606_5 gpc1028 (
      {stage0_25[474], stage0_25[475], stage0_25[476], stage0_25[477], stage0_25[478], stage0_25[479]},
      {stage0_27[234], stage0_27[235], stage0_27[236], stage0_27[237], stage0_27[238], stage0_27[239]},
      {stage1_29[39],stage1_28[96],stage1_27[136],stage1_26[153],stage1_25[182]}
   );
   gpc606_5 gpc1029 (
      {stage0_25[480], stage0_25[481], stage0_25[482], stage0_25[483], stage0_25[484], stage0_25[485]},
      {stage0_27[240], stage0_27[241], stage0_27[242], stage0_27[243], stage0_27[244], stage0_27[245]},
      {stage1_29[40],stage1_28[97],stage1_27[137],stage1_26[154],stage1_25[183]}
   );
   gpc615_5 gpc1030 (
      {stage0_26[342], stage0_26[343], stage0_26[344], stage0_26[345], stage0_26[346]},
      {stage0_27[246]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[41],stage1_28[98],stage1_27[138],stage1_26[155]}
   );
   gpc615_5 gpc1031 (
      {stage0_26[347], stage0_26[348], stage0_26[349], stage0_26[350], stage0_26[351]},
      {stage0_27[247]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[42],stage1_28[99],stage1_27[139],stage1_26[156]}
   );
   gpc615_5 gpc1032 (
      {stage0_26[352], stage0_26[353], stage0_26[354], stage0_26[355], stage0_26[356]},
      {stage0_27[248]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[43],stage1_28[100],stage1_27[140],stage1_26[157]}
   );
   gpc615_5 gpc1033 (
      {stage0_26[357], stage0_26[358], stage0_26[359], stage0_26[360], stage0_26[361]},
      {stage0_27[249]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[44],stage1_28[101],stage1_27[141],stage1_26[158]}
   );
   gpc615_5 gpc1034 (
      {stage0_26[362], stage0_26[363], stage0_26[364], stage0_26[365], stage0_26[366]},
      {stage0_27[250]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[45],stage1_28[102],stage1_27[142],stage1_26[159]}
   );
   gpc615_5 gpc1035 (
      {stage0_26[367], stage0_26[368], stage0_26[369], stage0_26[370], stage0_26[371]},
      {stage0_27[251]},
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage1_30[5],stage1_29[46],stage1_28[103],stage1_27[143],stage1_26[160]}
   );
   gpc615_5 gpc1036 (
      {stage0_26[372], stage0_26[373], stage0_26[374], stage0_26[375], stage0_26[376]},
      {stage0_27[252]},
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage1_30[6],stage1_29[47],stage1_28[104],stage1_27[144],stage1_26[161]}
   );
   gpc615_5 gpc1037 (
      {stage0_26[377], stage0_26[378], stage0_26[379], stage0_26[380], stage0_26[381]},
      {stage0_27[253]},
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage1_30[7],stage1_29[48],stage1_28[105],stage1_27[145],stage1_26[162]}
   );
   gpc615_5 gpc1038 (
      {stage0_26[382], stage0_26[383], stage0_26[384], stage0_26[385], stage0_26[386]},
      {stage0_27[254]},
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage1_30[8],stage1_29[49],stage1_28[106],stage1_27[146],stage1_26[163]}
   );
   gpc615_5 gpc1039 (
      {stage0_26[387], stage0_26[388], stage0_26[389], stage0_26[390], stage0_26[391]},
      {stage0_27[255]},
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage1_30[9],stage1_29[50],stage1_28[107],stage1_27[147],stage1_26[164]}
   );
   gpc615_5 gpc1040 (
      {stage0_26[392], stage0_26[393], stage0_26[394], stage0_26[395], stage0_26[396]},
      {stage0_27[256]},
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage1_30[10],stage1_29[51],stage1_28[108],stage1_27[148],stage1_26[165]}
   );
   gpc615_5 gpc1041 (
      {stage0_26[397], stage0_26[398], stage0_26[399], stage0_26[400], stage0_26[401]},
      {stage0_27[257]},
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage1_30[11],stage1_29[52],stage1_28[109],stage1_27[149],stage1_26[166]}
   );
   gpc615_5 gpc1042 (
      {stage0_27[258], stage0_27[259], stage0_27[260], stage0_27[261], stage0_27[262]},
      {stage0_28[72]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[12],stage1_29[53],stage1_28[110],stage1_27[150]}
   );
   gpc615_5 gpc1043 (
      {stage0_27[263], stage0_27[264], stage0_27[265], stage0_27[266], stage0_27[267]},
      {stage0_28[73]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[13],stage1_29[54],stage1_28[111],stage1_27[151]}
   );
   gpc615_5 gpc1044 (
      {stage0_27[268], stage0_27[269], stage0_27[270], stage0_27[271], stage0_27[272]},
      {stage0_28[74]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[14],stage1_29[55],stage1_28[112],stage1_27[152]}
   );
   gpc615_5 gpc1045 (
      {stage0_27[273], stage0_27[274], stage0_27[275], stage0_27[276], stage0_27[277]},
      {stage0_28[75]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[15],stage1_29[56],stage1_28[113],stage1_27[153]}
   );
   gpc615_5 gpc1046 (
      {stage0_27[278], stage0_27[279], stage0_27[280], stage0_27[281], stage0_27[282]},
      {stage0_28[76]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[16],stage1_29[57],stage1_28[114],stage1_27[154]}
   );
   gpc615_5 gpc1047 (
      {stage0_27[283], stage0_27[284], stage0_27[285], stage0_27[286], stage0_27[287]},
      {stage0_28[77]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[17],stage1_29[58],stage1_28[115],stage1_27[155]}
   );
   gpc615_5 gpc1048 (
      {stage0_27[288], stage0_27[289], stage0_27[290], stage0_27[291], stage0_27[292]},
      {stage0_28[78]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[18],stage1_29[59],stage1_28[116],stage1_27[156]}
   );
   gpc615_5 gpc1049 (
      {stage0_27[293], stage0_27[294], stage0_27[295], stage0_27[296], stage0_27[297]},
      {stage0_28[79]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[19],stage1_29[60],stage1_28[117],stage1_27[157]}
   );
   gpc615_5 gpc1050 (
      {stage0_27[298], stage0_27[299], stage0_27[300], stage0_27[301], stage0_27[302]},
      {stage0_28[80]},
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage1_31[8],stage1_30[20],stage1_29[61],stage1_28[118],stage1_27[158]}
   );
   gpc615_5 gpc1051 (
      {stage0_27[303], stage0_27[304], stage0_27[305], stage0_27[306], stage0_27[307]},
      {stage0_28[81]},
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage1_31[9],stage1_30[21],stage1_29[62],stage1_28[119],stage1_27[159]}
   );
   gpc615_5 gpc1052 (
      {stage0_27[308], stage0_27[309], stage0_27[310], stage0_27[311], stage0_27[312]},
      {stage0_28[82]},
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage1_31[10],stage1_30[22],stage1_29[63],stage1_28[120],stage1_27[160]}
   );
   gpc615_5 gpc1053 (
      {stage0_27[313], stage0_27[314], stage0_27[315], stage0_27[316], stage0_27[317]},
      {stage0_28[83]},
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage1_31[11],stage1_30[23],stage1_29[64],stage1_28[121],stage1_27[161]}
   );
   gpc615_5 gpc1054 (
      {stage0_27[318], stage0_27[319], stage0_27[320], stage0_27[321], stage0_27[322]},
      {stage0_28[84]},
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage1_31[12],stage1_30[24],stage1_29[65],stage1_28[122],stage1_27[162]}
   );
   gpc615_5 gpc1055 (
      {stage0_27[323], stage0_27[324], stage0_27[325], stage0_27[326], stage0_27[327]},
      {stage0_28[85]},
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage1_31[13],stage1_30[25],stage1_29[66],stage1_28[123],stage1_27[163]}
   );
   gpc615_5 gpc1056 (
      {stage0_27[328], stage0_27[329], stage0_27[330], stage0_27[331], stage0_27[332]},
      {stage0_28[86]},
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage1_31[14],stage1_30[26],stage1_29[67],stage1_28[124],stage1_27[164]}
   );
   gpc615_5 gpc1057 (
      {stage0_27[333], stage0_27[334], stage0_27[335], stage0_27[336], stage0_27[337]},
      {stage0_28[87]},
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage1_31[15],stage1_30[27],stage1_29[68],stage1_28[125],stage1_27[165]}
   );
   gpc615_5 gpc1058 (
      {stage0_27[338], stage0_27[339], stage0_27[340], stage0_27[341], stage0_27[342]},
      {stage0_28[88]},
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage1_31[16],stage1_30[28],stage1_29[69],stage1_28[126],stage1_27[166]}
   );
   gpc615_5 gpc1059 (
      {stage0_27[343], stage0_27[344], stage0_27[345], stage0_27[346], stage0_27[347]},
      {stage0_28[89]},
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage1_31[17],stage1_30[29],stage1_29[70],stage1_28[127],stage1_27[167]}
   );
   gpc615_5 gpc1060 (
      {stage0_27[348], stage0_27[349], stage0_27[350], stage0_27[351], stage0_27[352]},
      {stage0_28[90]},
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage1_31[18],stage1_30[30],stage1_29[71],stage1_28[128],stage1_27[168]}
   );
   gpc615_5 gpc1061 (
      {stage0_27[353], stage0_27[354], stage0_27[355], stage0_27[356], stage0_27[357]},
      {stage0_28[91]},
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage1_31[19],stage1_30[31],stage1_29[72],stage1_28[129],stage1_27[169]}
   );
   gpc615_5 gpc1062 (
      {stage0_27[358], stage0_27[359], stage0_27[360], stage0_27[361], stage0_27[362]},
      {stage0_28[92]},
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage1_31[20],stage1_30[32],stage1_29[73],stage1_28[130],stage1_27[170]}
   );
   gpc615_5 gpc1063 (
      {stage0_27[363], stage0_27[364], stage0_27[365], stage0_27[366], stage0_27[367]},
      {stage0_28[93]},
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage1_31[21],stage1_30[33],stage1_29[74],stage1_28[131],stage1_27[171]}
   );
   gpc615_5 gpc1064 (
      {stage0_27[368], stage0_27[369], stage0_27[370], stage0_27[371], stage0_27[372]},
      {stage0_28[94]},
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage1_31[22],stage1_30[34],stage1_29[75],stage1_28[132],stage1_27[172]}
   );
   gpc615_5 gpc1065 (
      {stage0_27[373], stage0_27[374], stage0_27[375], stage0_27[376], stage0_27[377]},
      {stage0_28[95]},
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage1_31[23],stage1_30[35],stage1_29[76],stage1_28[133],stage1_27[173]}
   );
   gpc615_5 gpc1066 (
      {stage0_27[378], stage0_27[379], stage0_27[380], stage0_27[381], stage0_27[382]},
      {stage0_28[96]},
      {stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149]},
      {stage1_31[24],stage1_30[36],stage1_29[77],stage1_28[134],stage1_27[174]}
   );
   gpc615_5 gpc1067 (
      {stage0_27[383], stage0_27[384], stage0_27[385], stage0_27[386], stage0_27[387]},
      {stage0_28[97]},
      {stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155]},
      {stage1_31[25],stage1_30[37],stage1_29[78],stage1_28[135],stage1_27[175]}
   );
   gpc615_5 gpc1068 (
      {stage0_27[388], stage0_27[389], stage0_27[390], stage0_27[391], stage0_27[392]},
      {stage0_28[98]},
      {stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161]},
      {stage1_31[26],stage1_30[38],stage1_29[79],stage1_28[136],stage1_27[176]}
   );
   gpc615_5 gpc1069 (
      {stage0_27[393], stage0_27[394], stage0_27[395], stage0_27[396], stage0_27[397]},
      {stage0_28[99]},
      {stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167]},
      {stage1_31[27],stage1_30[39],stage1_29[80],stage1_28[137],stage1_27[177]}
   );
   gpc615_5 gpc1070 (
      {stage0_27[398], stage0_27[399], stage0_27[400], stage0_27[401], stage0_27[402]},
      {stage0_28[100]},
      {stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173]},
      {stage1_31[28],stage1_30[40],stage1_29[81],stage1_28[138],stage1_27[178]}
   );
   gpc615_5 gpc1071 (
      {stage0_27[403], stage0_27[404], stage0_27[405], stage0_27[406], stage0_27[407]},
      {stage0_28[101]},
      {stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179]},
      {stage1_31[29],stage1_30[41],stage1_29[82],stage1_28[139],stage1_27[179]}
   );
   gpc615_5 gpc1072 (
      {stage0_27[408], stage0_27[409], stage0_27[410], stage0_27[411], stage0_27[412]},
      {stage0_28[102]},
      {stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185]},
      {stage1_31[30],stage1_30[42],stage1_29[83],stage1_28[140],stage1_27[180]}
   );
   gpc615_5 gpc1073 (
      {stage0_27[413], stage0_27[414], stage0_27[415], stage0_27[416], stage0_27[417]},
      {stage0_28[103]},
      {stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190], stage0_29[191]},
      {stage1_31[31],stage1_30[43],stage1_29[84],stage1_28[141],stage1_27[181]}
   );
   gpc615_5 gpc1074 (
      {stage0_27[418], stage0_27[419], stage0_27[420], stage0_27[421], stage0_27[422]},
      {stage0_28[104]},
      {stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196], stage0_29[197]},
      {stage1_31[32],stage1_30[44],stage1_29[85],stage1_28[142],stage1_27[182]}
   );
   gpc615_5 gpc1075 (
      {stage0_27[423], stage0_27[424], stage0_27[425], stage0_27[426], stage0_27[427]},
      {stage0_28[105]},
      {stage0_29[198], stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202], stage0_29[203]},
      {stage1_31[33],stage1_30[45],stage1_29[86],stage1_28[143],stage1_27[183]}
   );
   gpc615_5 gpc1076 (
      {stage0_27[428], stage0_27[429], stage0_27[430], stage0_27[431], stage0_27[432]},
      {stage0_28[106]},
      {stage0_29[204], stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209]},
      {stage1_31[34],stage1_30[46],stage1_29[87],stage1_28[144],stage1_27[184]}
   );
   gpc615_5 gpc1077 (
      {stage0_27[433], stage0_27[434], stage0_27[435], stage0_27[436], stage0_27[437]},
      {stage0_28[107]},
      {stage0_29[210], stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215]},
      {stage1_31[35],stage1_30[47],stage1_29[88],stage1_28[145],stage1_27[185]}
   );
   gpc615_5 gpc1078 (
      {stage0_27[438], stage0_27[439], stage0_27[440], stage0_27[441], stage0_27[442]},
      {stage0_28[108]},
      {stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220], stage0_29[221]},
      {stage1_31[36],stage1_30[48],stage1_29[89],stage1_28[146],stage1_27[186]}
   );
   gpc615_5 gpc1079 (
      {stage0_27[443], stage0_27[444], stage0_27[445], stage0_27[446], stage0_27[447]},
      {stage0_28[109]},
      {stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226], stage0_29[227]},
      {stage1_31[37],stage1_30[49],stage1_29[90],stage1_28[147],stage1_27[187]}
   );
   gpc615_5 gpc1080 (
      {stage0_27[448], stage0_27[449], stage0_27[450], stage0_27[451], stage0_27[452]},
      {stage0_28[110]},
      {stage0_29[228], stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232], stage0_29[233]},
      {stage1_31[38],stage1_30[50],stage1_29[91],stage1_28[148],stage1_27[188]}
   );
   gpc615_5 gpc1081 (
      {stage0_27[453], stage0_27[454], stage0_27[455], stage0_27[456], stage0_27[457]},
      {stage0_28[111]},
      {stage0_29[234], stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239]},
      {stage1_31[39],stage1_30[51],stage1_29[92],stage1_28[149],stage1_27[189]}
   );
   gpc615_5 gpc1082 (
      {stage0_27[458], stage0_27[459], stage0_27[460], stage0_27[461], stage0_27[462]},
      {stage0_28[112]},
      {stage0_29[240], stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245]},
      {stage1_31[40],stage1_30[52],stage1_29[93],stage1_28[150],stage1_27[190]}
   );
   gpc615_5 gpc1083 (
      {stage0_27[463], stage0_27[464], stage0_27[465], stage0_27[466], stage0_27[467]},
      {stage0_28[113]},
      {stage0_29[246], stage0_29[247], stage0_29[248], stage0_29[249], stage0_29[250], stage0_29[251]},
      {stage1_31[41],stage1_30[53],stage1_29[94],stage1_28[151],stage1_27[191]}
   );
   gpc615_5 gpc1084 (
      {stage0_27[468], stage0_27[469], stage0_27[470], stage0_27[471], stage0_27[472]},
      {stage0_28[114]},
      {stage0_29[252], stage0_29[253], stage0_29[254], stage0_29[255], stage0_29[256], stage0_29[257]},
      {stage1_31[42],stage1_30[54],stage1_29[95],stage1_28[152],stage1_27[192]}
   );
   gpc606_5 gpc1085 (
      {stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[43],stage1_30[55],stage1_29[96],stage1_28[153]}
   );
   gpc606_5 gpc1086 (
      {stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[44],stage1_30[56],stage1_29[97],stage1_28[154]}
   );
   gpc606_5 gpc1087 (
      {stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[45],stage1_30[57],stage1_29[98],stage1_28[155]}
   );
   gpc606_5 gpc1088 (
      {stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[46],stage1_30[58],stage1_29[99],stage1_28[156]}
   );
   gpc606_5 gpc1089 (
      {stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143], stage0_28[144]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[47],stage1_30[59],stage1_29[100],stage1_28[157]}
   );
   gpc606_5 gpc1090 (
      {stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149], stage0_28[150]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[48],stage1_30[60],stage1_29[101],stage1_28[158]}
   );
   gpc606_5 gpc1091 (
      {stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155], stage0_28[156]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[49],stage1_30[61],stage1_29[102],stage1_28[159]}
   );
   gpc606_5 gpc1092 (
      {stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161], stage0_28[162]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[50],stage1_30[62],stage1_29[103],stage1_28[160]}
   );
   gpc606_5 gpc1093 (
      {stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167], stage0_28[168]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[51],stage1_30[63],stage1_29[104],stage1_28[161]}
   );
   gpc606_5 gpc1094 (
      {stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173], stage0_28[174]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[52],stage1_30[64],stage1_29[105],stage1_28[162]}
   );
   gpc606_5 gpc1095 (
      {stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179], stage0_28[180]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[53],stage1_30[65],stage1_29[106],stage1_28[163]}
   );
   gpc606_5 gpc1096 (
      {stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185], stage0_28[186]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[54],stage1_30[66],stage1_29[107],stage1_28[164]}
   );
   gpc606_5 gpc1097 (
      {stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191], stage0_28[192]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[55],stage1_30[67],stage1_29[108],stage1_28[165]}
   );
   gpc606_5 gpc1098 (
      {stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197], stage0_28[198]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[56],stage1_30[68],stage1_29[109],stage1_28[166]}
   );
   gpc606_5 gpc1099 (
      {stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203], stage0_28[204]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[57],stage1_30[69],stage1_29[110],stage1_28[167]}
   );
   gpc606_5 gpc1100 (
      {stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209], stage0_28[210]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[58],stage1_30[70],stage1_29[111],stage1_28[168]}
   );
   gpc606_5 gpc1101 (
      {stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215], stage0_28[216]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[59],stage1_30[71],stage1_29[112],stage1_28[169]}
   );
   gpc606_5 gpc1102 (
      {stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221], stage0_28[222]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[60],stage1_30[72],stage1_29[113],stage1_28[170]}
   );
   gpc606_5 gpc1103 (
      {stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227], stage0_28[228]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[61],stage1_30[73],stage1_29[114],stage1_28[171]}
   );
   gpc606_5 gpc1104 (
      {stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233], stage0_28[234]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[62],stage1_30[74],stage1_29[115],stage1_28[172]}
   );
   gpc606_5 gpc1105 (
      {stage0_28[235], stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239], stage0_28[240]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[63],stage1_30[75],stage1_29[116],stage1_28[173]}
   );
   gpc606_5 gpc1106 (
      {stage0_28[241], stage0_28[242], stage0_28[243], stage0_28[244], stage0_28[245], stage0_28[246]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[64],stage1_30[76],stage1_29[117],stage1_28[174]}
   );
   gpc606_5 gpc1107 (
      {stage0_28[247], stage0_28[248], stage0_28[249], stage0_28[250], stage0_28[251], stage0_28[252]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[65],stage1_30[77],stage1_29[118],stage1_28[175]}
   );
   gpc606_5 gpc1108 (
      {stage0_28[253], stage0_28[254], stage0_28[255], stage0_28[256], stage0_28[257], stage0_28[258]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[66],stage1_30[78],stage1_29[119],stage1_28[176]}
   );
   gpc606_5 gpc1109 (
      {stage0_28[259], stage0_28[260], stage0_28[261], stage0_28[262], stage0_28[263], stage0_28[264]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[67],stage1_30[79],stage1_29[120],stage1_28[177]}
   );
   gpc606_5 gpc1110 (
      {stage0_28[265], stage0_28[266], stage0_28[267], stage0_28[268], stage0_28[269], stage0_28[270]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[68],stage1_30[80],stage1_29[121],stage1_28[178]}
   );
   gpc606_5 gpc1111 (
      {stage0_28[271], stage0_28[272], stage0_28[273], stage0_28[274], stage0_28[275], stage0_28[276]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[69],stage1_30[81],stage1_29[122],stage1_28[179]}
   );
   gpc606_5 gpc1112 (
      {stage0_28[277], stage0_28[278], stage0_28[279], stage0_28[280], stage0_28[281], stage0_28[282]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[70],stage1_30[82],stage1_29[123],stage1_28[180]}
   );
   gpc606_5 gpc1113 (
      {stage0_28[283], stage0_28[284], stage0_28[285], stage0_28[286], stage0_28[287], stage0_28[288]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[71],stage1_30[83],stage1_29[124],stage1_28[181]}
   );
   gpc606_5 gpc1114 (
      {stage0_28[289], stage0_28[290], stage0_28[291], stage0_28[292], stage0_28[293], stage0_28[294]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[72],stage1_30[84],stage1_29[125],stage1_28[182]}
   );
   gpc606_5 gpc1115 (
      {stage0_28[295], stage0_28[296], stage0_28[297], stage0_28[298], stage0_28[299], stage0_28[300]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[73],stage1_30[85],stage1_29[126],stage1_28[183]}
   );
   gpc606_5 gpc1116 (
      {stage0_28[301], stage0_28[302], stage0_28[303], stage0_28[304], stage0_28[305], stage0_28[306]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[74],stage1_30[86],stage1_29[127],stage1_28[184]}
   );
   gpc606_5 gpc1117 (
      {stage0_28[307], stage0_28[308], stage0_28[309], stage0_28[310], stage0_28[311], stage0_28[312]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[75],stage1_30[87],stage1_29[128],stage1_28[185]}
   );
   gpc606_5 gpc1118 (
      {stage0_28[313], stage0_28[314], stage0_28[315], stage0_28[316], stage0_28[317], stage0_28[318]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[76],stage1_30[88],stage1_29[129],stage1_28[186]}
   );
   gpc606_5 gpc1119 (
      {stage0_28[319], stage0_28[320], stage0_28[321], stage0_28[322], stage0_28[323], stage0_28[324]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[77],stage1_30[89],stage1_29[130],stage1_28[187]}
   );
   gpc606_5 gpc1120 (
      {stage0_28[325], stage0_28[326], stage0_28[327], stage0_28[328], stage0_28[329], stage0_28[330]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[78],stage1_30[90],stage1_29[131],stage1_28[188]}
   );
   gpc606_5 gpc1121 (
      {stage0_28[331], stage0_28[332], stage0_28[333], stage0_28[334], stage0_28[335], stage0_28[336]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[79],stage1_30[91],stage1_29[132],stage1_28[189]}
   );
   gpc606_5 gpc1122 (
      {stage0_28[337], stage0_28[338], stage0_28[339], stage0_28[340], stage0_28[341], stage0_28[342]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[80],stage1_30[92],stage1_29[133],stage1_28[190]}
   );
   gpc606_5 gpc1123 (
      {stage0_28[343], stage0_28[344], stage0_28[345], stage0_28[346], stage0_28[347], stage0_28[348]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[81],stage1_30[93],stage1_29[134],stage1_28[191]}
   );
   gpc606_5 gpc1124 (
      {stage0_28[349], stage0_28[350], stage0_28[351], stage0_28[352], stage0_28[353], stage0_28[354]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[82],stage1_30[94],stage1_29[135],stage1_28[192]}
   );
   gpc606_5 gpc1125 (
      {stage0_28[355], stage0_28[356], stage0_28[357], stage0_28[358], stage0_28[359], stage0_28[360]},
      {stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243], stage0_30[244], stage0_30[245]},
      {stage1_32[40],stage1_31[83],stage1_30[95],stage1_29[136],stage1_28[193]}
   );
   gpc606_5 gpc1126 (
      {stage0_28[361], stage0_28[362], stage0_28[363], stage0_28[364], stage0_28[365], stage0_28[366]},
      {stage0_30[246], stage0_30[247], stage0_30[248], stage0_30[249], stage0_30[250], stage0_30[251]},
      {stage1_32[41],stage1_31[84],stage1_30[96],stage1_29[137],stage1_28[194]}
   );
   gpc606_5 gpc1127 (
      {stage0_28[367], stage0_28[368], stage0_28[369], stage0_28[370], stage0_28[371], stage0_28[372]},
      {stage0_30[252], stage0_30[253], stage0_30[254], stage0_30[255], stage0_30[256], stage0_30[257]},
      {stage1_32[42],stage1_31[85],stage1_30[97],stage1_29[138],stage1_28[195]}
   );
   gpc606_5 gpc1128 (
      {stage0_28[373], stage0_28[374], stage0_28[375], stage0_28[376], stage0_28[377], stage0_28[378]},
      {stage0_30[258], stage0_30[259], stage0_30[260], stage0_30[261], stage0_30[262], stage0_30[263]},
      {stage1_32[43],stage1_31[86],stage1_30[98],stage1_29[139],stage1_28[196]}
   );
   gpc606_5 gpc1129 (
      {stage0_28[379], stage0_28[380], stage0_28[381], stage0_28[382], stage0_28[383], stage0_28[384]},
      {stage0_30[264], stage0_30[265], stage0_30[266], stage0_30[267], stage0_30[268], stage0_30[269]},
      {stage1_32[44],stage1_31[87],stage1_30[99],stage1_29[140],stage1_28[197]}
   );
   gpc606_5 gpc1130 (
      {stage0_28[385], stage0_28[386], stage0_28[387], stage0_28[388], stage0_28[389], stage0_28[390]},
      {stage0_30[270], stage0_30[271], stage0_30[272], stage0_30[273], stage0_30[274], stage0_30[275]},
      {stage1_32[45],stage1_31[88],stage1_30[100],stage1_29[141],stage1_28[198]}
   );
   gpc606_5 gpc1131 (
      {stage0_28[391], stage0_28[392], stage0_28[393], stage0_28[394], stage0_28[395], stage0_28[396]},
      {stage0_30[276], stage0_30[277], stage0_30[278], stage0_30[279], stage0_30[280], stage0_30[281]},
      {stage1_32[46],stage1_31[89],stage1_30[101],stage1_29[142],stage1_28[199]}
   );
   gpc606_5 gpc1132 (
      {stage0_28[397], stage0_28[398], stage0_28[399], stage0_28[400], stage0_28[401], stage0_28[402]},
      {stage0_30[282], stage0_30[283], stage0_30[284], stage0_30[285], stage0_30[286], stage0_30[287]},
      {stage1_32[47],stage1_31[90],stage1_30[102],stage1_29[143],stage1_28[200]}
   );
   gpc606_5 gpc1133 (
      {stage0_28[403], stage0_28[404], stage0_28[405], stage0_28[406], stage0_28[407], stage0_28[408]},
      {stage0_30[288], stage0_30[289], stage0_30[290], stage0_30[291], stage0_30[292], stage0_30[293]},
      {stage1_32[48],stage1_31[91],stage1_30[103],stage1_29[144],stage1_28[201]}
   );
   gpc606_5 gpc1134 (
      {stage0_28[409], stage0_28[410], stage0_28[411], stage0_28[412], stage0_28[413], stage0_28[414]},
      {stage0_30[294], stage0_30[295], stage0_30[296], stage0_30[297], stage0_30[298], stage0_30[299]},
      {stage1_32[49],stage1_31[92],stage1_30[104],stage1_29[145],stage1_28[202]}
   );
   gpc606_5 gpc1135 (
      {stage0_28[415], stage0_28[416], stage0_28[417], stage0_28[418], stage0_28[419], stage0_28[420]},
      {stage0_30[300], stage0_30[301], stage0_30[302], stage0_30[303], stage0_30[304], stage0_30[305]},
      {stage1_32[50],stage1_31[93],stage1_30[105],stage1_29[146],stage1_28[203]}
   );
   gpc606_5 gpc1136 (
      {stage0_28[421], stage0_28[422], stage0_28[423], stage0_28[424], stage0_28[425], stage0_28[426]},
      {stage0_30[306], stage0_30[307], stage0_30[308], stage0_30[309], stage0_30[310], stage0_30[311]},
      {stage1_32[51],stage1_31[94],stage1_30[106],stage1_29[147],stage1_28[204]}
   );
   gpc606_5 gpc1137 (
      {stage0_28[427], stage0_28[428], stage0_28[429], stage0_28[430], stage0_28[431], stage0_28[432]},
      {stage0_30[312], stage0_30[313], stage0_30[314], stage0_30[315], stage0_30[316], stage0_30[317]},
      {stage1_32[52],stage1_31[95],stage1_30[107],stage1_29[148],stage1_28[205]}
   );
   gpc606_5 gpc1138 (
      {stage0_28[433], stage0_28[434], stage0_28[435], stage0_28[436], stage0_28[437], stage0_28[438]},
      {stage0_30[318], stage0_30[319], stage0_30[320], stage0_30[321], stage0_30[322], stage0_30[323]},
      {stage1_32[53],stage1_31[96],stage1_30[108],stage1_29[149],stage1_28[206]}
   );
   gpc606_5 gpc1139 (
      {stage0_28[439], stage0_28[440], stage0_28[441], stage0_28[442], stage0_28[443], stage0_28[444]},
      {stage0_30[324], stage0_30[325], stage0_30[326], stage0_30[327], stage0_30[328], stage0_30[329]},
      {stage1_32[54],stage1_31[97],stage1_30[109],stage1_29[150],stage1_28[207]}
   );
   gpc606_5 gpc1140 (
      {stage0_28[445], stage0_28[446], stage0_28[447], stage0_28[448], stage0_28[449], stage0_28[450]},
      {stage0_30[330], stage0_30[331], stage0_30[332], stage0_30[333], stage0_30[334], stage0_30[335]},
      {stage1_32[55],stage1_31[98],stage1_30[110],stage1_29[151],stage1_28[208]}
   );
   gpc606_5 gpc1141 (
      {stage0_28[451], stage0_28[452], stage0_28[453], stage0_28[454], stage0_28[455], stage0_28[456]},
      {stage0_30[336], stage0_30[337], stage0_30[338], stage0_30[339], stage0_30[340], stage0_30[341]},
      {stage1_32[56],stage1_31[99],stage1_30[111],stage1_29[152],stage1_28[209]}
   );
   gpc606_5 gpc1142 (
      {stage0_28[457], stage0_28[458], stage0_28[459], stage0_28[460], stage0_28[461], stage0_28[462]},
      {stage0_30[342], stage0_30[343], stage0_30[344], stage0_30[345], stage0_30[346], stage0_30[347]},
      {stage1_32[57],stage1_31[100],stage1_30[112],stage1_29[153],stage1_28[210]}
   );
   gpc606_5 gpc1143 (
      {stage0_28[463], stage0_28[464], stage0_28[465], stage0_28[466], stage0_28[467], stage0_28[468]},
      {stage0_30[348], stage0_30[349], stage0_30[350], stage0_30[351], stage0_30[352], stage0_30[353]},
      {stage1_32[58],stage1_31[101],stage1_30[113],stage1_29[154],stage1_28[211]}
   );
   gpc606_5 gpc1144 (
      {stage0_28[469], stage0_28[470], stage0_28[471], stage0_28[472], stage0_28[473], stage0_28[474]},
      {stage0_30[354], stage0_30[355], stage0_30[356], stage0_30[357], stage0_30[358], stage0_30[359]},
      {stage1_32[59],stage1_31[102],stage1_30[114],stage1_29[155],stage1_28[212]}
   );
   gpc606_5 gpc1145 (
      {stage0_29[258], stage0_29[259], stage0_29[260], stage0_29[261], stage0_29[262], stage0_29[263]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[60],stage1_31[103],stage1_30[115],stage1_29[156]}
   );
   gpc606_5 gpc1146 (
      {stage0_29[264], stage0_29[265], stage0_29[266], stage0_29[267], stage0_29[268], stage0_29[269]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[61],stage1_31[104],stage1_30[116],stage1_29[157]}
   );
   gpc606_5 gpc1147 (
      {stage0_29[270], stage0_29[271], stage0_29[272], stage0_29[273], stage0_29[274], stage0_29[275]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[62],stage1_31[105],stage1_30[117],stage1_29[158]}
   );
   gpc606_5 gpc1148 (
      {stage0_29[276], stage0_29[277], stage0_29[278], stage0_29[279], stage0_29[280], stage0_29[281]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[63],stage1_31[106],stage1_30[118],stage1_29[159]}
   );
   gpc606_5 gpc1149 (
      {stage0_29[282], stage0_29[283], stage0_29[284], stage0_29[285], stage0_29[286], stage0_29[287]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[64],stage1_31[107],stage1_30[119],stage1_29[160]}
   );
   gpc606_5 gpc1150 (
      {stage0_29[288], stage0_29[289], stage0_29[290], stage0_29[291], stage0_29[292], stage0_29[293]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[65],stage1_31[108],stage1_30[120],stage1_29[161]}
   );
   gpc606_5 gpc1151 (
      {stage0_29[294], stage0_29[295], stage0_29[296], stage0_29[297], stage0_29[298], stage0_29[299]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[66],stage1_31[109],stage1_30[121],stage1_29[162]}
   );
   gpc606_5 gpc1152 (
      {stage0_29[300], stage0_29[301], stage0_29[302], stage0_29[303], stage0_29[304], stage0_29[305]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[67],stage1_31[110],stage1_30[122],stage1_29[163]}
   );
   gpc606_5 gpc1153 (
      {stage0_29[306], stage0_29[307], stage0_29[308], stage0_29[309], stage0_29[310], stage0_29[311]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[68],stage1_31[111],stage1_30[123],stage1_29[164]}
   );
   gpc606_5 gpc1154 (
      {stage0_29[312], stage0_29[313], stage0_29[314], stage0_29[315], stage0_29[316], stage0_29[317]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[69],stage1_31[112],stage1_30[124],stage1_29[165]}
   );
   gpc606_5 gpc1155 (
      {stage0_29[318], stage0_29[319], stage0_29[320], stage0_29[321], stage0_29[322], stage0_29[323]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[70],stage1_31[113],stage1_30[125],stage1_29[166]}
   );
   gpc606_5 gpc1156 (
      {stage0_29[324], stage0_29[325], stage0_29[326], stage0_29[327], stage0_29[328], stage0_29[329]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[71],stage1_31[114],stage1_30[126],stage1_29[167]}
   );
   gpc606_5 gpc1157 (
      {stage0_29[330], stage0_29[331], stage0_29[332], stage0_29[333], stage0_29[334], stage0_29[335]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[72],stage1_31[115],stage1_30[127],stage1_29[168]}
   );
   gpc606_5 gpc1158 (
      {stage0_29[336], stage0_29[337], stage0_29[338], stage0_29[339], stage0_29[340], stage0_29[341]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[73],stage1_31[116],stage1_30[128],stage1_29[169]}
   );
   gpc606_5 gpc1159 (
      {stage0_29[342], stage0_29[343], stage0_29[344], stage0_29[345], stage0_29[346], stage0_29[347]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[74],stage1_31[117],stage1_30[129],stage1_29[170]}
   );
   gpc606_5 gpc1160 (
      {stage0_29[348], stage0_29[349], stage0_29[350], stage0_29[351], stage0_29[352], stage0_29[353]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[75],stage1_31[118],stage1_30[130],stage1_29[171]}
   );
   gpc606_5 gpc1161 (
      {stage0_29[354], stage0_29[355], stage0_29[356], stage0_29[357], stage0_29[358], stage0_29[359]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[76],stage1_31[119],stage1_30[131],stage1_29[172]}
   );
   gpc606_5 gpc1162 (
      {stage0_29[360], stage0_29[361], stage0_29[362], stage0_29[363], stage0_29[364], stage0_29[365]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[77],stage1_31[120],stage1_30[132],stage1_29[173]}
   );
   gpc606_5 gpc1163 (
      {stage0_29[366], stage0_29[367], stage0_29[368], stage0_29[369], stage0_29[370], stage0_29[371]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[78],stage1_31[121],stage1_30[133],stage1_29[174]}
   );
   gpc606_5 gpc1164 (
      {stage0_29[372], stage0_29[373], stage0_29[374], stage0_29[375], stage0_29[376], stage0_29[377]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[79],stage1_31[122],stage1_30[134],stage1_29[175]}
   );
   gpc606_5 gpc1165 (
      {stage0_29[378], stage0_29[379], stage0_29[380], stage0_29[381], stage0_29[382], stage0_29[383]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[80],stage1_31[123],stage1_30[135],stage1_29[176]}
   );
   gpc606_5 gpc1166 (
      {stage0_29[384], stage0_29[385], stage0_29[386], stage0_29[387], stage0_29[388], stage0_29[389]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[81],stage1_31[124],stage1_30[136],stage1_29[177]}
   );
   gpc606_5 gpc1167 (
      {stage0_29[390], stage0_29[391], stage0_29[392], stage0_29[393], stage0_29[394], stage0_29[395]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[82],stage1_31[125],stage1_30[137],stage1_29[178]}
   );
   gpc606_5 gpc1168 (
      {stage0_29[396], stage0_29[397], stage0_29[398], stage0_29[399], stage0_29[400], stage0_29[401]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[83],stage1_31[126],stage1_30[138],stage1_29[179]}
   );
   gpc606_5 gpc1169 (
      {stage0_29[402], stage0_29[403], stage0_29[404], stage0_29[405], stage0_29[406], stage0_29[407]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[84],stage1_31[127],stage1_30[139],stage1_29[180]}
   );
   gpc606_5 gpc1170 (
      {stage0_29[408], stage0_29[409], stage0_29[410], stage0_29[411], stage0_29[412], stage0_29[413]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[85],stage1_31[128],stage1_30[140],stage1_29[181]}
   );
   gpc606_5 gpc1171 (
      {stage0_29[414], stage0_29[415], stage0_29[416], stage0_29[417], stage0_29[418], stage0_29[419]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[86],stage1_31[129],stage1_30[141],stage1_29[182]}
   );
   gpc606_5 gpc1172 (
      {stage0_29[420], stage0_29[421], stage0_29[422], stage0_29[423], stage0_29[424], stage0_29[425]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[87],stage1_31[130],stage1_30[142],stage1_29[183]}
   );
   gpc606_5 gpc1173 (
      {stage0_29[426], stage0_29[427], stage0_29[428], stage0_29[429], stage0_29[430], stage0_29[431]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[88],stage1_31[131],stage1_30[143],stage1_29[184]}
   );
   gpc606_5 gpc1174 (
      {stage0_29[432], stage0_29[433], stage0_29[434], stage0_29[435], stage0_29[436], stage0_29[437]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[89],stage1_31[132],stage1_30[144],stage1_29[185]}
   );
   gpc606_5 gpc1175 (
      {stage0_29[438], stage0_29[439], stage0_29[440], stage0_29[441], stage0_29[442], stage0_29[443]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[90],stage1_31[133],stage1_30[145],stage1_29[186]}
   );
   gpc615_5 gpc1176 (
      {stage0_30[360], stage0_30[361], stage0_30[362], stage0_30[363], stage0_30[364]},
      {stage0_31[186]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[31],stage1_32[91],stage1_31[134],stage1_30[146]}
   );
   gpc615_5 gpc1177 (
      {stage0_30[365], stage0_30[366], stage0_30[367], stage0_30[368], stage0_30[369]},
      {stage0_31[187]},
      {stage0_32[6], stage0_32[7], stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11]},
      {stage1_34[1],stage1_33[32],stage1_32[92],stage1_31[135],stage1_30[147]}
   );
   gpc615_5 gpc1178 (
      {stage0_30[370], stage0_30[371], stage0_30[372], stage0_30[373], stage0_30[374]},
      {stage0_31[188]},
      {stage0_32[12], stage0_32[13], stage0_32[14], stage0_32[15], stage0_32[16], stage0_32[17]},
      {stage1_34[2],stage1_33[33],stage1_32[93],stage1_31[136],stage1_30[148]}
   );
   gpc615_5 gpc1179 (
      {stage0_30[375], stage0_30[376], stage0_30[377], stage0_30[378], stage0_30[379]},
      {stage0_31[189]},
      {stage0_32[18], stage0_32[19], stage0_32[20], stage0_32[21], stage0_32[22], stage0_32[23]},
      {stage1_34[3],stage1_33[34],stage1_32[94],stage1_31[137],stage1_30[149]}
   );
   gpc615_5 gpc1180 (
      {stage0_30[380], stage0_30[381], stage0_30[382], stage0_30[383], stage0_30[384]},
      {stage0_31[190]},
      {stage0_32[24], stage0_32[25], stage0_32[26], stage0_32[27], stage0_32[28], stage0_32[29]},
      {stage1_34[4],stage1_33[35],stage1_32[95],stage1_31[138],stage1_30[150]}
   );
   gpc615_5 gpc1181 (
      {stage0_30[385], stage0_30[386], stage0_30[387], stage0_30[388], stage0_30[389]},
      {stage0_31[191]},
      {stage0_32[30], stage0_32[31], stage0_32[32], stage0_32[33], stage0_32[34], stage0_32[35]},
      {stage1_34[5],stage1_33[36],stage1_32[96],stage1_31[139],stage1_30[151]}
   );
   gpc615_5 gpc1182 (
      {stage0_30[390], stage0_30[391], stage0_30[392], stage0_30[393], stage0_30[394]},
      {stage0_31[192]},
      {stage0_32[36], stage0_32[37], stage0_32[38], stage0_32[39], stage0_32[40], stage0_32[41]},
      {stage1_34[6],stage1_33[37],stage1_32[97],stage1_31[140],stage1_30[152]}
   );
   gpc615_5 gpc1183 (
      {stage0_30[395], stage0_30[396], stage0_30[397], stage0_30[398], stage0_30[399]},
      {stage0_31[193]},
      {stage0_32[42], stage0_32[43], stage0_32[44], stage0_32[45], stage0_32[46], stage0_32[47]},
      {stage1_34[7],stage1_33[38],stage1_32[98],stage1_31[141],stage1_30[153]}
   );
   gpc615_5 gpc1184 (
      {stage0_30[400], stage0_30[401], stage0_30[402], stage0_30[403], stage0_30[404]},
      {stage0_31[194]},
      {stage0_32[48], stage0_32[49], stage0_32[50], stage0_32[51], stage0_32[52], stage0_32[53]},
      {stage1_34[8],stage1_33[39],stage1_32[99],stage1_31[142],stage1_30[154]}
   );
   gpc615_5 gpc1185 (
      {stage0_30[405], stage0_30[406], stage0_30[407], stage0_30[408], stage0_30[409]},
      {stage0_31[195]},
      {stage0_32[54], stage0_32[55], stage0_32[56], stage0_32[57], stage0_32[58], stage0_32[59]},
      {stage1_34[9],stage1_33[40],stage1_32[100],stage1_31[143],stage1_30[155]}
   );
   gpc615_5 gpc1186 (
      {stage0_30[410], stage0_30[411], stage0_30[412], stage0_30[413], stage0_30[414]},
      {stage0_31[196]},
      {stage0_32[60], stage0_32[61], stage0_32[62], stage0_32[63], stage0_32[64], stage0_32[65]},
      {stage1_34[10],stage1_33[41],stage1_32[101],stage1_31[144],stage1_30[156]}
   );
   gpc615_5 gpc1187 (
      {stage0_30[415], stage0_30[416], stage0_30[417], stage0_30[418], stage0_30[419]},
      {stage0_31[197]},
      {stage0_32[66], stage0_32[67], stage0_32[68], stage0_32[69], stage0_32[70], stage0_32[71]},
      {stage1_34[11],stage1_33[42],stage1_32[102],stage1_31[145],stage1_30[157]}
   );
   gpc615_5 gpc1188 (
      {stage0_30[420], stage0_30[421], stage0_30[422], stage0_30[423], stage0_30[424]},
      {stage0_31[198]},
      {stage0_32[72], stage0_32[73], stage0_32[74], stage0_32[75], stage0_32[76], stage0_32[77]},
      {stage1_34[12],stage1_33[43],stage1_32[103],stage1_31[146],stage1_30[158]}
   );
   gpc615_5 gpc1189 (
      {stage0_30[425], stage0_30[426], stage0_30[427], stage0_30[428], stage0_30[429]},
      {stage0_31[199]},
      {stage0_32[78], stage0_32[79], stage0_32[80], stage0_32[81], stage0_32[82], stage0_32[83]},
      {stage1_34[13],stage1_33[44],stage1_32[104],stage1_31[147],stage1_30[159]}
   );
   gpc615_5 gpc1190 (
      {stage0_30[430], stage0_30[431], stage0_30[432], stage0_30[433], stage0_30[434]},
      {stage0_31[200]},
      {stage0_32[84], stage0_32[85], stage0_32[86], stage0_32[87], stage0_32[88], stage0_32[89]},
      {stage1_34[14],stage1_33[45],stage1_32[105],stage1_31[148],stage1_30[160]}
   );
   gpc615_5 gpc1191 (
      {stage0_30[435], stage0_30[436], stage0_30[437], stage0_30[438], stage0_30[439]},
      {stage0_31[201]},
      {stage0_32[90], stage0_32[91], stage0_32[92], stage0_32[93], stage0_32[94], stage0_32[95]},
      {stage1_34[15],stage1_33[46],stage1_32[106],stage1_31[149],stage1_30[161]}
   );
   gpc615_5 gpc1192 (
      {stage0_30[440], stage0_30[441], stage0_30[442], stage0_30[443], stage0_30[444]},
      {stage0_31[202]},
      {stage0_32[96], stage0_32[97], stage0_32[98], stage0_32[99], stage0_32[100], stage0_32[101]},
      {stage1_34[16],stage1_33[47],stage1_32[107],stage1_31[150],stage1_30[162]}
   );
   gpc615_5 gpc1193 (
      {stage0_30[445], stage0_30[446], stage0_30[447], stage0_30[448], stage0_30[449]},
      {stage0_31[203]},
      {stage0_32[102], stage0_32[103], stage0_32[104], stage0_32[105], stage0_32[106], stage0_32[107]},
      {stage1_34[17],stage1_33[48],stage1_32[108],stage1_31[151],stage1_30[163]}
   );
   gpc615_5 gpc1194 (
      {stage0_30[450], stage0_30[451], stage0_30[452], stage0_30[453], stage0_30[454]},
      {stage0_31[204]},
      {stage0_32[108], stage0_32[109], stage0_32[110], stage0_32[111], stage0_32[112], stage0_32[113]},
      {stage1_34[18],stage1_33[49],stage1_32[109],stage1_31[152],stage1_30[164]}
   );
   gpc615_5 gpc1195 (
      {stage0_30[455], stage0_30[456], stage0_30[457], stage0_30[458], stage0_30[459]},
      {stage0_31[205]},
      {stage0_32[114], stage0_32[115], stage0_32[116], stage0_32[117], stage0_32[118], stage0_32[119]},
      {stage1_34[19],stage1_33[50],stage1_32[110],stage1_31[153],stage1_30[165]}
   );
   gpc615_5 gpc1196 (
      {stage0_31[206], stage0_31[207], stage0_31[208], stage0_31[209], stage0_31[210]},
      {stage0_32[120]},
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage1_35[0],stage1_34[20],stage1_33[51],stage1_32[111],stage1_31[154]}
   );
   gpc615_5 gpc1197 (
      {stage0_31[211], stage0_31[212], stage0_31[213], stage0_31[214], stage0_31[215]},
      {stage0_32[121]},
      {stage0_33[6], stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11]},
      {stage1_35[1],stage1_34[21],stage1_33[52],stage1_32[112],stage1_31[155]}
   );
   gpc615_5 gpc1198 (
      {stage0_31[216], stage0_31[217], stage0_31[218], stage0_31[219], stage0_31[220]},
      {stage0_32[122]},
      {stage0_33[12], stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17]},
      {stage1_35[2],stage1_34[22],stage1_33[53],stage1_32[113],stage1_31[156]}
   );
   gpc615_5 gpc1199 (
      {stage0_31[221], stage0_31[222], stage0_31[223], stage0_31[224], stage0_31[225]},
      {stage0_32[123]},
      {stage0_33[18], stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23]},
      {stage1_35[3],stage1_34[23],stage1_33[54],stage1_32[114],stage1_31[157]}
   );
   gpc615_5 gpc1200 (
      {stage0_31[226], stage0_31[227], stage0_31[228], stage0_31[229], stage0_31[230]},
      {stage0_32[124]},
      {stage0_33[24], stage0_33[25], stage0_33[26], stage0_33[27], stage0_33[28], stage0_33[29]},
      {stage1_35[4],stage1_34[24],stage1_33[55],stage1_32[115],stage1_31[158]}
   );
   gpc615_5 gpc1201 (
      {stage0_31[231], stage0_31[232], stage0_31[233], stage0_31[234], stage0_31[235]},
      {stage0_32[125]},
      {stage0_33[30], stage0_33[31], stage0_33[32], stage0_33[33], stage0_33[34], stage0_33[35]},
      {stage1_35[5],stage1_34[25],stage1_33[56],stage1_32[116],stage1_31[159]}
   );
   gpc615_5 gpc1202 (
      {stage0_31[236], stage0_31[237], stage0_31[238], stage0_31[239], stage0_31[240]},
      {stage0_32[126]},
      {stage0_33[36], stage0_33[37], stage0_33[38], stage0_33[39], stage0_33[40], stage0_33[41]},
      {stage1_35[6],stage1_34[26],stage1_33[57],stage1_32[117],stage1_31[160]}
   );
   gpc615_5 gpc1203 (
      {stage0_31[241], stage0_31[242], stage0_31[243], stage0_31[244], stage0_31[245]},
      {stage0_32[127]},
      {stage0_33[42], stage0_33[43], stage0_33[44], stage0_33[45], stage0_33[46], stage0_33[47]},
      {stage1_35[7],stage1_34[27],stage1_33[58],stage1_32[118],stage1_31[161]}
   );
   gpc615_5 gpc1204 (
      {stage0_31[246], stage0_31[247], stage0_31[248], stage0_31[249], stage0_31[250]},
      {stage0_32[128]},
      {stage0_33[48], stage0_33[49], stage0_33[50], stage0_33[51], stage0_33[52], stage0_33[53]},
      {stage1_35[8],stage1_34[28],stage1_33[59],stage1_32[119],stage1_31[162]}
   );
   gpc615_5 gpc1205 (
      {stage0_31[251], stage0_31[252], stage0_31[253], stage0_31[254], stage0_31[255]},
      {stage0_32[129]},
      {stage0_33[54], stage0_33[55], stage0_33[56], stage0_33[57], stage0_33[58], stage0_33[59]},
      {stage1_35[9],stage1_34[29],stage1_33[60],stage1_32[120],stage1_31[163]}
   );
   gpc615_5 gpc1206 (
      {stage0_31[256], stage0_31[257], stage0_31[258], stage0_31[259], stage0_31[260]},
      {stage0_32[130]},
      {stage0_33[60], stage0_33[61], stage0_33[62], stage0_33[63], stage0_33[64], stage0_33[65]},
      {stage1_35[10],stage1_34[30],stage1_33[61],stage1_32[121],stage1_31[164]}
   );
   gpc615_5 gpc1207 (
      {stage0_31[261], stage0_31[262], stage0_31[263], stage0_31[264], stage0_31[265]},
      {stage0_32[131]},
      {stage0_33[66], stage0_33[67], stage0_33[68], stage0_33[69], stage0_33[70], stage0_33[71]},
      {stage1_35[11],stage1_34[31],stage1_33[62],stage1_32[122],stage1_31[165]}
   );
   gpc615_5 gpc1208 (
      {stage0_31[266], stage0_31[267], stage0_31[268], stage0_31[269], stage0_31[270]},
      {stage0_32[132]},
      {stage0_33[72], stage0_33[73], stage0_33[74], stage0_33[75], stage0_33[76], stage0_33[77]},
      {stage1_35[12],stage1_34[32],stage1_33[63],stage1_32[123],stage1_31[166]}
   );
   gpc615_5 gpc1209 (
      {stage0_31[271], stage0_31[272], stage0_31[273], stage0_31[274], stage0_31[275]},
      {stage0_32[133]},
      {stage0_33[78], stage0_33[79], stage0_33[80], stage0_33[81], stage0_33[82], stage0_33[83]},
      {stage1_35[13],stage1_34[33],stage1_33[64],stage1_32[124],stage1_31[167]}
   );
   gpc615_5 gpc1210 (
      {stage0_31[276], stage0_31[277], stage0_31[278], stage0_31[279], stage0_31[280]},
      {stage0_32[134]},
      {stage0_33[84], stage0_33[85], stage0_33[86], stage0_33[87], stage0_33[88], stage0_33[89]},
      {stage1_35[14],stage1_34[34],stage1_33[65],stage1_32[125],stage1_31[168]}
   );
   gpc615_5 gpc1211 (
      {stage0_31[281], stage0_31[282], stage0_31[283], stage0_31[284], stage0_31[285]},
      {stage0_32[135]},
      {stage0_33[90], stage0_33[91], stage0_33[92], stage0_33[93], stage0_33[94], stage0_33[95]},
      {stage1_35[15],stage1_34[35],stage1_33[66],stage1_32[126],stage1_31[169]}
   );
   gpc615_5 gpc1212 (
      {stage0_31[286], stage0_31[287], stage0_31[288], stage0_31[289], stage0_31[290]},
      {stage0_32[136]},
      {stage0_33[96], stage0_33[97], stage0_33[98], stage0_33[99], stage0_33[100], stage0_33[101]},
      {stage1_35[16],stage1_34[36],stage1_33[67],stage1_32[127],stage1_31[170]}
   );
   gpc615_5 gpc1213 (
      {stage0_31[291], stage0_31[292], stage0_31[293], stage0_31[294], stage0_31[295]},
      {stage0_32[137]},
      {stage0_33[102], stage0_33[103], stage0_33[104], stage0_33[105], stage0_33[106], stage0_33[107]},
      {stage1_35[17],stage1_34[37],stage1_33[68],stage1_32[128],stage1_31[171]}
   );
   gpc615_5 gpc1214 (
      {stage0_31[296], stage0_31[297], stage0_31[298], stage0_31[299], stage0_31[300]},
      {stage0_32[138]},
      {stage0_33[108], stage0_33[109], stage0_33[110], stage0_33[111], stage0_33[112], stage0_33[113]},
      {stage1_35[18],stage1_34[38],stage1_33[69],stage1_32[129],stage1_31[172]}
   );
   gpc615_5 gpc1215 (
      {stage0_31[301], stage0_31[302], stage0_31[303], stage0_31[304], stage0_31[305]},
      {stage0_32[139]},
      {stage0_33[114], stage0_33[115], stage0_33[116], stage0_33[117], stage0_33[118], stage0_33[119]},
      {stage1_35[19],stage1_34[39],stage1_33[70],stage1_32[130],stage1_31[173]}
   );
   gpc615_5 gpc1216 (
      {stage0_31[306], stage0_31[307], stage0_31[308], stage0_31[309], stage0_31[310]},
      {stage0_32[140]},
      {stage0_33[120], stage0_33[121], stage0_33[122], stage0_33[123], stage0_33[124], stage0_33[125]},
      {stage1_35[20],stage1_34[40],stage1_33[71],stage1_32[131],stage1_31[174]}
   );
   gpc615_5 gpc1217 (
      {stage0_31[311], stage0_31[312], stage0_31[313], stage0_31[314], stage0_31[315]},
      {stage0_32[141]},
      {stage0_33[126], stage0_33[127], stage0_33[128], stage0_33[129], stage0_33[130], stage0_33[131]},
      {stage1_35[21],stage1_34[41],stage1_33[72],stage1_32[132],stage1_31[175]}
   );
   gpc615_5 gpc1218 (
      {stage0_31[316], stage0_31[317], stage0_31[318], stage0_31[319], stage0_31[320]},
      {stage0_32[142]},
      {stage0_33[132], stage0_33[133], stage0_33[134], stage0_33[135], stage0_33[136], stage0_33[137]},
      {stage1_35[22],stage1_34[42],stage1_33[73],stage1_32[133],stage1_31[176]}
   );
   gpc615_5 gpc1219 (
      {stage0_31[321], stage0_31[322], stage0_31[323], stage0_31[324], stage0_31[325]},
      {stage0_32[143]},
      {stage0_33[138], stage0_33[139], stage0_33[140], stage0_33[141], stage0_33[142], stage0_33[143]},
      {stage1_35[23],stage1_34[43],stage1_33[74],stage1_32[134],stage1_31[177]}
   );
   gpc615_5 gpc1220 (
      {stage0_31[326], stage0_31[327], stage0_31[328], stage0_31[329], stage0_31[330]},
      {stage0_32[144]},
      {stage0_33[144], stage0_33[145], stage0_33[146], stage0_33[147], stage0_33[148], stage0_33[149]},
      {stage1_35[24],stage1_34[44],stage1_33[75],stage1_32[135],stage1_31[178]}
   );
   gpc615_5 gpc1221 (
      {stage0_31[331], stage0_31[332], stage0_31[333], stage0_31[334], stage0_31[335]},
      {stage0_32[145]},
      {stage0_33[150], stage0_33[151], stage0_33[152], stage0_33[153], stage0_33[154], stage0_33[155]},
      {stage1_35[25],stage1_34[45],stage1_33[76],stage1_32[136],stage1_31[179]}
   );
   gpc615_5 gpc1222 (
      {stage0_31[336], stage0_31[337], stage0_31[338], stage0_31[339], stage0_31[340]},
      {stage0_32[146]},
      {stage0_33[156], stage0_33[157], stage0_33[158], stage0_33[159], stage0_33[160], stage0_33[161]},
      {stage1_35[26],stage1_34[46],stage1_33[77],stage1_32[137],stage1_31[180]}
   );
   gpc615_5 gpc1223 (
      {stage0_31[341], stage0_31[342], stage0_31[343], stage0_31[344], stage0_31[345]},
      {stage0_32[147]},
      {stage0_33[162], stage0_33[163], stage0_33[164], stage0_33[165], stage0_33[166], stage0_33[167]},
      {stage1_35[27],stage1_34[47],stage1_33[78],stage1_32[138],stage1_31[181]}
   );
   gpc615_5 gpc1224 (
      {stage0_31[346], stage0_31[347], stage0_31[348], stage0_31[349], stage0_31[350]},
      {stage0_32[148]},
      {stage0_33[168], stage0_33[169], stage0_33[170], stage0_33[171], stage0_33[172], stage0_33[173]},
      {stage1_35[28],stage1_34[48],stage1_33[79],stage1_32[139],stage1_31[182]}
   );
   gpc615_5 gpc1225 (
      {stage0_31[351], stage0_31[352], stage0_31[353], stage0_31[354], stage0_31[355]},
      {stage0_32[149]},
      {stage0_33[174], stage0_33[175], stage0_33[176], stage0_33[177], stage0_33[178], stage0_33[179]},
      {stage1_35[29],stage1_34[49],stage1_33[80],stage1_32[140],stage1_31[183]}
   );
   gpc615_5 gpc1226 (
      {stage0_31[356], stage0_31[357], stage0_31[358], stage0_31[359], stage0_31[360]},
      {stage0_32[150]},
      {stage0_33[180], stage0_33[181], stage0_33[182], stage0_33[183], stage0_33[184], stage0_33[185]},
      {stage1_35[30],stage1_34[50],stage1_33[81],stage1_32[141],stage1_31[184]}
   );
   gpc615_5 gpc1227 (
      {stage0_31[361], stage0_31[362], stage0_31[363], stage0_31[364], stage0_31[365]},
      {stage0_32[151]},
      {stage0_33[186], stage0_33[187], stage0_33[188], stage0_33[189], stage0_33[190], stage0_33[191]},
      {stage1_35[31],stage1_34[51],stage1_33[82],stage1_32[142],stage1_31[185]}
   );
   gpc615_5 gpc1228 (
      {stage0_31[366], stage0_31[367], stage0_31[368], stage0_31[369], stage0_31[370]},
      {stage0_32[152]},
      {stage0_33[192], stage0_33[193], stage0_33[194], stage0_33[195], stage0_33[196], stage0_33[197]},
      {stage1_35[32],stage1_34[52],stage1_33[83],stage1_32[143],stage1_31[186]}
   );
   gpc615_5 gpc1229 (
      {stage0_31[371], stage0_31[372], stage0_31[373], stage0_31[374], stage0_31[375]},
      {stage0_32[153]},
      {stage0_33[198], stage0_33[199], stage0_33[200], stage0_33[201], stage0_33[202], stage0_33[203]},
      {stage1_35[33],stage1_34[53],stage1_33[84],stage1_32[144],stage1_31[187]}
   );
   gpc615_5 gpc1230 (
      {stage0_31[376], stage0_31[377], stage0_31[378], stage0_31[379], stage0_31[380]},
      {stage0_32[154]},
      {stage0_33[204], stage0_33[205], stage0_33[206], stage0_33[207], stage0_33[208], stage0_33[209]},
      {stage1_35[34],stage1_34[54],stage1_33[85],stage1_32[145],stage1_31[188]}
   );
   gpc615_5 gpc1231 (
      {stage0_31[381], stage0_31[382], stage0_31[383], stage0_31[384], stage0_31[385]},
      {stage0_32[155]},
      {stage0_33[210], stage0_33[211], stage0_33[212], stage0_33[213], stage0_33[214], stage0_33[215]},
      {stage1_35[35],stage1_34[55],stage1_33[86],stage1_32[146],stage1_31[189]}
   );
   gpc615_5 gpc1232 (
      {stage0_31[386], stage0_31[387], stage0_31[388], stage0_31[389], stage0_31[390]},
      {stage0_32[156]},
      {stage0_33[216], stage0_33[217], stage0_33[218], stage0_33[219], stage0_33[220], stage0_33[221]},
      {stage1_35[36],stage1_34[56],stage1_33[87],stage1_32[147],stage1_31[190]}
   );
   gpc615_5 gpc1233 (
      {stage0_31[391], stage0_31[392], stage0_31[393], stage0_31[394], stage0_31[395]},
      {stage0_32[157]},
      {stage0_33[222], stage0_33[223], stage0_33[224], stage0_33[225], stage0_33[226], stage0_33[227]},
      {stage1_35[37],stage1_34[57],stage1_33[88],stage1_32[148],stage1_31[191]}
   );
   gpc615_5 gpc1234 (
      {stage0_31[396], stage0_31[397], stage0_31[398], stage0_31[399], stage0_31[400]},
      {stage0_32[158]},
      {stage0_33[228], stage0_33[229], stage0_33[230], stage0_33[231], stage0_33[232], stage0_33[233]},
      {stage1_35[38],stage1_34[58],stage1_33[89],stage1_32[149],stage1_31[192]}
   );
   gpc615_5 gpc1235 (
      {stage0_31[401], stage0_31[402], stage0_31[403], stage0_31[404], stage0_31[405]},
      {stage0_32[159]},
      {stage0_33[234], stage0_33[235], stage0_33[236], stage0_33[237], stage0_33[238], stage0_33[239]},
      {stage1_35[39],stage1_34[59],stage1_33[90],stage1_32[150],stage1_31[193]}
   );
   gpc615_5 gpc1236 (
      {stage0_31[406], stage0_31[407], stage0_31[408], stage0_31[409], stage0_31[410]},
      {stage0_32[160]},
      {stage0_33[240], stage0_33[241], stage0_33[242], stage0_33[243], stage0_33[244], stage0_33[245]},
      {stage1_35[40],stage1_34[60],stage1_33[91],stage1_32[151],stage1_31[194]}
   );
   gpc615_5 gpc1237 (
      {stage0_31[411], stage0_31[412], stage0_31[413], stage0_31[414], stage0_31[415]},
      {stage0_32[161]},
      {stage0_33[246], stage0_33[247], stage0_33[248], stage0_33[249], stage0_33[250], stage0_33[251]},
      {stage1_35[41],stage1_34[61],stage1_33[92],stage1_32[152],stage1_31[195]}
   );
   gpc615_5 gpc1238 (
      {stage0_31[416], stage0_31[417], stage0_31[418], stage0_31[419], stage0_31[420]},
      {stage0_32[162]},
      {stage0_33[252], stage0_33[253], stage0_33[254], stage0_33[255], stage0_33[256], stage0_33[257]},
      {stage1_35[42],stage1_34[62],stage1_33[93],stage1_32[153],stage1_31[196]}
   );
   gpc615_5 gpc1239 (
      {stage0_31[421], stage0_31[422], stage0_31[423], stage0_31[424], stage0_31[425]},
      {stage0_32[163]},
      {stage0_33[258], stage0_33[259], stage0_33[260], stage0_33[261], stage0_33[262], stage0_33[263]},
      {stage1_35[43],stage1_34[63],stage1_33[94],stage1_32[154],stage1_31[197]}
   );
   gpc615_5 gpc1240 (
      {stage0_31[426], stage0_31[427], stage0_31[428], stage0_31[429], stage0_31[430]},
      {stage0_32[164]},
      {stage0_33[264], stage0_33[265], stage0_33[266], stage0_33[267], stage0_33[268], stage0_33[269]},
      {stage1_35[44],stage1_34[64],stage1_33[95],stage1_32[155],stage1_31[198]}
   );
   gpc615_5 gpc1241 (
      {stage0_31[431], stage0_31[432], stage0_31[433], stage0_31[434], stage0_31[435]},
      {stage0_32[165]},
      {stage0_33[270], stage0_33[271], stage0_33[272], stage0_33[273], stage0_33[274], stage0_33[275]},
      {stage1_35[45],stage1_34[65],stage1_33[96],stage1_32[156],stage1_31[199]}
   );
   gpc615_5 gpc1242 (
      {stage0_31[436], stage0_31[437], stage0_31[438], stage0_31[439], stage0_31[440]},
      {stage0_32[166]},
      {stage0_33[276], stage0_33[277], stage0_33[278], stage0_33[279], stage0_33[280], stage0_33[281]},
      {stage1_35[46],stage1_34[66],stage1_33[97],stage1_32[157],stage1_31[200]}
   );
   gpc615_5 gpc1243 (
      {stage0_31[441], stage0_31[442], stage0_31[443], stage0_31[444], stage0_31[445]},
      {stage0_32[167]},
      {stage0_33[282], stage0_33[283], stage0_33[284], stage0_33[285], stage0_33[286], stage0_33[287]},
      {stage1_35[47],stage1_34[67],stage1_33[98],stage1_32[158],stage1_31[201]}
   );
   gpc615_5 gpc1244 (
      {stage0_31[446], stage0_31[447], stage0_31[448], stage0_31[449], stage0_31[450]},
      {stage0_32[168]},
      {stage0_33[288], stage0_33[289], stage0_33[290], stage0_33[291], stage0_33[292], stage0_33[293]},
      {stage1_35[48],stage1_34[68],stage1_33[99],stage1_32[159],stage1_31[202]}
   );
   gpc615_5 gpc1245 (
      {stage0_31[451], stage0_31[452], stage0_31[453], stage0_31[454], stage0_31[455]},
      {stage0_32[169]},
      {stage0_33[294], stage0_33[295], stage0_33[296], stage0_33[297], stage0_33[298], stage0_33[299]},
      {stage1_35[49],stage1_34[69],stage1_33[100],stage1_32[160],stage1_31[203]}
   );
   gpc615_5 gpc1246 (
      {stage0_31[456], stage0_31[457], stage0_31[458], stage0_31[459], stage0_31[460]},
      {stage0_32[170]},
      {stage0_33[300], stage0_33[301], stage0_33[302], stage0_33[303], stage0_33[304], stage0_33[305]},
      {stage1_35[50],stage1_34[70],stage1_33[101],stage1_32[161],stage1_31[204]}
   );
   gpc615_5 gpc1247 (
      {stage0_31[461], stage0_31[462], stage0_31[463], stage0_31[464], stage0_31[465]},
      {stage0_32[171]},
      {stage0_33[306], stage0_33[307], stage0_33[308], stage0_33[309], stage0_33[310], stage0_33[311]},
      {stage1_35[51],stage1_34[71],stage1_33[102],stage1_32[162],stage1_31[205]}
   );
   gpc615_5 gpc1248 (
      {stage0_31[466], stage0_31[467], stage0_31[468], stage0_31[469], stage0_31[470]},
      {stage0_32[172]},
      {stage0_33[312], stage0_33[313], stage0_33[314], stage0_33[315], stage0_33[316], stage0_33[317]},
      {stage1_35[52],stage1_34[72],stage1_33[103],stage1_32[163],stage1_31[206]}
   );
   gpc615_5 gpc1249 (
      {stage0_31[471], stage0_31[472], stage0_31[473], stage0_31[474], stage0_31[475]},
      {stage0_32[173]},
      {stage0_33[318], stage0_33[319], stage0_33[320], stage0_33[321], stage0_33[322], stage0_33[323]},
      {stage1_35[53],stage1_34[73],stage1_33[104],stage1_32[164],stage1_31[207]}
   );
   gpc606_5 gpc1250 (
      {stage0_32[174], stage0_32[175], stage0_32[176], stage0_32[177], stage0_32[178], stage0_32[179]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[54],stage1_34[74],stage1_33[105],stage1_32[165]}
   );
   gpc606_5 gpc1251 (
      {stage0_32[180], stage0_32[181], stage0_32[182], stage0_32[183], stage0_32[184], stage0_32[185]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[55],stage1_34[75],stage1_33[106],stage1_32[166]}
   );
   gpc606_5 gpc1252 (
      {stage0_32[186], stage0_32[187], stage0_32[188], stage0_32[189], stage0_32[190], stage0_32[191]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[56],stage1_34[76],stage1_33[107],stage1_32[167]}
   );
   gpc606_5 gpc1253 (
      {stage0_32[192], stage0_32[193], stage0_32[194], stage0_32[195], stage0_32[196], stage0_32[197]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[57],stage1_34[77],stage1_33[108],stage1_32[168]}
   );
   gpc606_5 gpc1254 (
      {stage0_32[198], stage0_32[199], stage0_32[200], stage0_32[201], stage0_32[202], stage0_32[203]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[58],stage1_34[78],stage1_33[109],stage1_32[169]}
   );
   gpc606_5 gpc1255 (
      {stage0_32[204], stage0_32[205], stage0_32[206], stage0_32[207], stage0_32[208], stage0_32[209]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[59],stage1_34[79],stage1_33[110],stage1_32[170]}
   );
   gpc606_5 gpc1256 (
      {stage0_32[210], stage0_32[211], stage0_32[212], stage0_32[213], stage0_32[214], stage0_32[215]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[60],stage1_34[80],stage1_33[111],stage1_32[171]}
   );
   gpc606_5 gpc1257 (
      {stage0_32[216], stage0_32[217], stage0_32[218], stage0_32[219], stage0_32[220], stage0_32[221]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[61],stage1_34[81],stage1_33[112],stage1_32[172]}
   );
   gpc606_5 gpc1258 (
      {stage0_32[222], stage0_32[223], stage0_32[224], stage0_32[225], stage0_32[226], stage0_32[227]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[62],stage1_34[82],stage1_33[113],stage1_32[173]}
   );
   gpc606_5 gpc1259 (
      {stage0_32[228], stage0_32[229], stage0_32[230], stage0_32[231], stage0_32[232], stage0_32[233]},
      {stage0_34[54], stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage1_36[9],stage1_35[63],stage1_34[83],stage1_33[114],stage1_32[174]}
   );
   gpc606_5 gpc1260 (
      {stage0_32[234], stage0_32[235], stage0_32[236], stage0_32[237], stage0_32[238], stage0_32[239]},
      {stage0_34[60], stage0_34[61], stage0_34[62], stage0_34[63], stage0_34[64], stage0_34[65]},
      {stage1_36[10],stage1_35[64],stage1_34[84],stage1_33[115],stage1_32[175]}
   );
   gpc606_5 gpc1261 (
      {stage0_32[240], stage0_32[241], stage0_32[242], stage0_32[243], stage0_32[244], stage0_32[245]},
      {stage0_34[66], stage0_34[67], stage0_34[68], stage0_34[69], stage0_34[70], stage0_34[71]},
      {stage1_36[11],stage1_35[65],stage1_34[85],stage1_33[116],stage1_32[176]}
   );
   gpc606_5 gpc1262 (
      {stage0_32[246], stage0_32[247], stage0_32[248], stage0_32[249], stage0_32[250], stage0_32[251]},
      {stage0_34[72], stage0_34[73], stage0_34[74], stage0_34[75], stage0_34[76], stage0_34[77]},
      {stage1_36[12],stage1_35[66],stage1_34[86],stage1_33[117],stage1_32[177]}
   );
   gpc606_5 gpc1263 (
      {stage0_32[252], stage0_32[253], stage0_32[254], stage0_32[255], stage0_32[256], stage0_32[257]},
      {stage0_34[78], stage0_34[79], stage0_34[80], stage0_34[81], stage0_34[82], stage0_34[83]},
      {stage1_36[13],stage1_35[67],stage1_34[87],stage1_33[118],stage1_32[178]}
   );
   gpc606_5 gpc1264 (
      {stage0_32[258], stage0_32[259], stage0_32[260], stage0_32[261], stage0_32[262], stage0_32[263]},
      {stage0_34[84], stage0_34[85], stage0_34[86], stage0_34[87], stage0_34[88], stage0_34[89]},
      {stage1_36[14],stage1_35[68],stage1_34[88],stage1_33[119],stage1_32[179]}
   );
   gpc606_5 gpc1265 (
      {stage0_32[264], stage0_32[265], stage0_32[266], stage0_32[267], stage0_32[268], stage0_32[269]},
      {stage0_34[90], stage0_34[91], stage0_34[92], stage0_34[93], stage0_34[94], stage0_34[95]},
      {stage1_36[15],stage1_35[69],stage1_34[89],stage1_33[120],stage1_32[180]}
   );
   gpc606_5 gpc1266 (
      {stage0_32[270], stage0_32[271], stage0_32[272], stage0_32[273], stage0_32[274], stage0_32[275]},
      {stage0_34[96], stage0_34[97], stage0_34[98], stage0_34[99], stage0_34[100], stage0_34[101]},
      {stage1_36[16],stage1_35[70],stage1_34[90],stage1_33[121],stage1_32[181]}
   );
   gpc606_5 gpc1267 (
      {stage0_32[276], stage0_32[277], stage0_32[278], stage0_32[279], stage0_32[280], stage0_32[281]},
      {stage0_34[102], stage0_34[103], stage0_34[104], stage0_34[105], stage0_34[106], stage0_34[107]},
      {stage1_36[17],stage1_35[71],stage1_34[91],stage1_33[122],stage1_32[182]}
   );
   gpc606_5 gpc1268 (
      {stage0_32[282], stage0_32[283], stage0_32[284], stage0_32[285], stage0_32[286], stage0_32[287]},
      {stage0_34[108], stage0_34[109], stage0_34[110], stage0_34[111], stage0_34[112], stage0_34[113]},
      {stage1_36[18],stage1_35[72],stage1_34[92],stage1_33[123],stage1_32[183]}
   );
   gpc606_5 gpc1269 (
      {stage0_32[288], stage0_32[289], stage0_32[290], stage0_32[291], stage0_32[292], stage0_32[293]},
      {stage0_34[114], stage0_34[115], stage0_34[116], stage0_34[117], stage0_34[118], stage0_34[119]},
      {stage1_36[19],stage1_35[73],stage1_34[93],stage1_33[124],stage1_32[184]}
   );
   gpc606_5 gpc1270 (
      {stage0_32[294], stage0_32[295], stage0_32[296], stage0_32[297], stage0_32[298], stage0_32[299]},
      {stage0_34[120], stage0_34[121], stage0_34[122], stage0_34[123], stage0_34[124], stage0_34[125]},
      {stage1_36[20],stage1_35[74],stage1_34[94],stage1_33[125],stage1_32[185]}
   );
   gpc606_5 gpc1271 (
      {stage0_32[300], stage0_32[301], stage0_32[302], stage0_32[303], stage0_32[304], stage0_32[305]},
      {stage0_34[126], stage0_34[127], stage0_34[128], stage0_34[129], stage0_34[130], stage0_34[131]},
      {stage1_36[21],stage1_35[75],stage1_34[95],stage1_33[126],stage1_32[186]}
   );
   gpc606_5 gpc1272 (
      {stage0_32[306], stage0_32[307], stage0_32[308], stage0_32[309], stage0_32[310], stage0_32[311]},
      {stage0_34[132], stage0_34[133], stage0_34[134], stage0_34[135], stage0_34[136], stage0_34[137]},
      {stage1_36[22],stage1_35[76],stage1_34[96],stage1_33[127],stage1_32[187]}
   );
   gpc606_5 gpc1273 (
      {stage0_32[312], stage0_32[313], stage0_32[314], stage0_32[315], stage0_32[316], stage0_32[317]},
      {stage0_34[138], stage0_34[139], stage0_34[140], stage0_34[141], stage0_34[142], stage0_34[143]},
      {stage1_36[23],stage1_35[77],stage1_34[97],stage1_33[128],stage1_32[188]}
   );
   gpc606_5 gpc1274 (
      {stage0_32[318], stage0_32[319], stage0_32[320], stage0_32[321], stage0_32[322], stage0_32[323]},
      {stage0_34[144], stage0_34[145], stage0_34[146], stage0_34[147], stage0_34[148], stage0_34[149]},
      {stage1_36[24],stage1_35[78],stage1_34[98],stage1_33[129],stage1_32[189]}
   );
   gpc606_5 gpc1275 (
      {stage0_32[324], stage0_32[325], stage0_32[326], stage0_32[327], stage0_32[328], stage0_32[329]},
      {stage0_34[150], stage0_34[151], stage0_34[152], stage0_34[153], stage0_34[154], stage0_34[155]},
      {stage1_36[25],stage1_35[79],stage1_34[99],stage1_33[130],stage1_32[190]}
   );
   gpc606_5 gpc1276 (
      {stage0_32[330], stage0_32[331], stage0_32[332], stage0_32[333], stage0_32[334], stage0_32[335]},
      {stage0_34[156], stage0_34[157], stage0_34[158], stage0_34[159], stage0_34[160], stage0_34[161]},
      {stage1_36[26],stage1_35[80],stage1_34[100],stage1_33[131],stage1_32[191]}
   );
   gpc606_5 gpc1277 (
      {stage0_32[336], stage0_32[337], stage0_32[338], stage0_32[339], stage0_32[340], stage0_32[341]},
      {stage0_34[162], stage0_34[163], stage0_34[164], stage0_34[165], stage0_34[166], stage0_34[167]},
      {stage1_36[27],stage1_35[81],stage1_34[101],stage1_33[132],stage1_32[192]}
   );
   gpc606_5 gpc1278 (
      {stage0_32[342], stage0_32[343], stage0_32[344], stage0_32[345], stage0_32[346], stage0_32[347]},
      {stage0_34[168], stage0_34[169], stage0_34[170], stage0_34[171], stage0_34[172], stage0_34[173]},
      {stage1_36[28],stage1_35[82],stage1_34[102],stage1_33[133],stage1_32[193]}
   );
   gpc606_5 gpc1279 (
      {stage0_32[348], stage0_32[349], stage0_32[350], stage0_32[351], stage0_32[352], stage0_32[353]},
      {stage0_34[174], stage0_34[175], stage0_34[176], stage0_34[177], stage0_34[178], stage0_34[179]},
      {stage1_36[29],stage1_35[83],stage1_34[103],stage1_33[134],stage1_32[194]}
   );
   gpc606_5 gpc1280 (
      {stage0_32[354], stage0_32[355], stage0_32[356], stage0_32[357], stage0_32[358], stage0_32[359]},
      {stage0_34[180], stage0_34[181], stage0_34[182], stage0_34[183], stage0_34[184], stage0_34[185]},
      {stage1_36[30],stage1_35[84],stage1_34[104],stage1_33[135],stage1_32[195]}
   );
   gpc606_5 gpc1281 (
      {stage0_32[360], stage0_32[361], stage0_32[362], stage0_32[363], stage0_32[364], stage0_32[365]},
      {stage0_34[186], stage0_34[187], stage0_34[188], stage0_34[189], stage0_34[190], stage0_34[191]},
      {stage1_36[31],stage1_35[85],stage1_34[105],stage1_33[136],stage1_32[196]}
   );
   gpc606_5 gpc1282 (
      {stage0_32[366], stage0_32[367], stage0_32[368], stage0_32[369], stage0_32[370], stage0_32[371]},
      {stage0_34[192], stage0_34[193], stage0_34[194], stage0_34[195], stage0_34[196], stage0_34[197]},
      {stage1_36[32],stage1_35[86],stage1_34[106],stage1_33[137],stage1_32[197]}
   );
   gpc606_5 gpc1283 (
      {stage0_32[372], stage0_32[373], stage0_32[374], stage0_32[375], stage0_32[376], stage0_32[377]},
      {stage0_34[198], stage0_34[199], stage0_34[200], stage0_34[201], stage0_34[202], stage0_34[203]},
      {stage1_36[33],stage1_35[87],stage1_34[107],stage1_33[138],stage1_32[198]}
   );
   gpc606_5 gpc1284 (
      {stage0_32[378], stage0_32[379], stage0_32[380], stage0_32[381], stage0_32[382], stage0_32[383]},
      {stage0_34[204], stage0_34[205], stage0_34[206], stage0_34[207], stage0_34[208], stage0_34[209]},
      {stage1_36[34],stage1_35[88],stage1_34[108],stage1_33[139],stage1_32[199]}
   );
   gpc606_5 gpc1285 (
      {stage0_32[384], stage0_32[385], stage0_32[386], stage0_32[387], stage0_32[388], stage0_32[389]},
      {stage0_34[210], stage0_34[211], stage0_34[212], stage0_34[213], stage0_34[214], stage0_34[215]},
      {stage1_36[35],stage1_35[89],stage1_34[109],stage1_33[140],stage1_32[200]}
   );
   gpc606_5 gpc1286 (
      {stage0_32[390], stage0_32[391], stage0_32[392], stage0_32[393], stage0_32[394], stage0_32[395]},
      {stage0_34[216], stage0_34[217], stage0_34[218], stage0_34[219], stage0_34[220], stage0_34[221]},
      {stage1_36[36],stage1_35[90],stage1_34[110],stage1_33[141],stage1_32[201]}
   );
   gpc606_5 gpc1287 (
      {stage0_32[396], stage0_32[397], stage0_32[398], stage0_32[399], stage0_32[400], stage0_32[401]},
      {stage0_34[222], stage0_34[223], stage0_34[224], stage0_34[225], stage0_34[226], stage0_34[227]},
      {stage1_36[37],stage1_35[91],stage1_34[111],stage1_33[142],stage1_32[202]}
   );
   gpc606_5 gpc1288 (
      {stage0_32[402], stage0_32[403], stage0_32[404], stage0_32[405], stage0_32[406], stage0_32[407]},
      {stage0_34[228], stage0_34[229], stage0_34[230], stage0_34[231], stage0_34[232], stage0_34[233]},
      {stage1_36[38],stage1_35[92],stage1_34[112],stage1_33[143],stage1_32[203]}
   );
   gpc606_5 gpc1289 (
      {stage0_32[408], stage0_32[409], stage0_32[410], stage0_32[411], stage0_32[412], stage0_32[413]},
      {stage0_34[234], stage0_34[235], stage0_34[236], stage0_34[237], stage0_34[238], stage0_34[239]},
      {stage1_36[39],stage1_35[93],stage1_34[113],stage1_33[144],stage1_32[204]}
   );
   gpc606_5 gpc1290 (
      {stage0_32[414], stage0_32[415], stage0_32[416], stage0_32[417], stage0_32[418], stage0_32[419]},
      {stage0_34[240], stage0_34[241], stage0_34[242], stage0_34[243], stage0_34[244], stage0_34[245]},
      {stage1_36[40],stage1_35[94],stage1_34[114],stage1_33[145],stage1_32[205]}
   );
   gpc606_5 gpc1291 (
      {stage0_32[420], stage0_32[421], stage0_32[422], stage0_32[423], stage0_32[424], stage0_32[425]},
      {stage0_34[246], stage0_34[247], stage0_34[248], stage0_34[249], stage0_34[250], stage0_34[251]},
      {stage1_36[41],stage1_35[95],stage1_34[115],stage1_33[146],stage1_32[206]}
   );
   gpc606_5 gpc1292 (
      {stage0_32[426], stage0_32[427], stage0_32[428], stage0_32[429], stage0_32[430], stage0_32[431]},
      {stage0_34[252], stage0_34[253], stage0_34[254], stage0_34[255], stage0_34[256], stage0_34[257]},
      {stage1_36[42],stage1_35[96],stage1_34[116],stage1_33[147],stage1_32[207]}
   );
   gpc606_5 gpc1293 (
      {stage0_32[432], stage0_32[433], stage0_32[434], stage0_32[435], stage0_32[436], stage0_32[437]},
      {stage0_34[258], stage0_34[259], stage0_34[260], stage0_34[261], stage0_34[262], stage0_34[263]},
      {stage1_36[43],stage1_35[97],stage1_34[117],stage1_33[148],stage1_32[208]}
   );
   gpc606_5 gpc1294 (
      {stage0_32[438], stage0_32[439], stage0_32[440], stage0_32[441], stage0_32[442], stage0_32[443]},
      {stage0_34[264], stage0_34[265], stage0_34[266], stage0_34[267], stage0_34[268], stage0_34[269]},
      {stage1_36[44],stage1_35[98],stage1_34[118],stage1_33[149],stage1_32[209]}
   );
   gpc606_5 gpc1295 (
      {stage0_32[444], stage0_32[445], stage0_32[446], stage0_32[447], stage0_32[448], stage0_32[449]},
      {stage0_34[270], stage0_34[271], stage0_34[272], stage0_34[273], stage0_34[274], stage0_34[275]},
      {stage1_36[45],stage1_35[99],stage1_34[119],stage1_33[150],stage1_32[210]}
   );
   gpc606_5 gpc1296 (
      {stage0_32[450], stage0_32[451], stage0_32[452], stage0_32[453], stage0_32[454], stage0_32[455]},
      {stage0_34[276], stage0_34[277], stage0_34[278], stage0_34[279], stage0_34[280], stage0_34[281]},
      {stage1_36[46],stage1_35[100],stage1_34[120],stage1_33[151],stage1_32[211]}
   );
   gpc606_5 gpc1297 (
      {stage0_32[456], stage0_32[457], stage0_32[458], stage0_32[459], stage0_32[460], stage0_32[461]},
      {stage0_34[282], stage0_34[283], stage0_34[284], stage0_34[285], stage0_34[286], stage0_34[287]},
      {stage1_36[47],stage1_35[101],stage1_34[121],stage1_33[152],stage1_32[212]}
   );
   gpc606_5 gpc1298 (
      {stage0_32[462], stage0_32[463], stage0_32[464], stage0_32[465], stage0_32[466], stage0_32[467]},
      {stage0_34[288], stage0_34[289], stage0_34[290], stage0_34[291], stage0_34[292], stage0_34[293]},
      {stage1_36[48],stage1_35[102],stage1_34[122],stage1_33[153],stage1_32[213]}
   );
   gpc606_5 gpc1299 (
      {stage0_32[468], stage0_32[469], stage0_32[470], stage0_32[471], stage0_32[472], stage0_32[473]},
      {stage0_34[294], stage0_34[295], stage0_34[296], stage0_34[297], stage0_34[298], stage0_34[299]},
      {stage1_36[49],stage1_35[103],stage1_34[123],stage1_33[154],stage1_32[214]}
   );
   gpc606_5 gpc1300 (
      {stage0_32[474], stage0_32[475], stage0_32[476], stage0_32[477], stage0_32[478], stage0_32[479]},
      {stage0_34[300], stage0_34[301], stage0_34[302], stage0_34[303], stage0_34[304], stage0_34[305]},
      {stage1_36[50],stage1_35[104],stage1_34[124],stage1_33[155],stage1_32[215]}
   );
   gpc606_5 gpc1301 (
      {stage0_32[480], stage0_32[481], stage0_32[482], stage0_32[483], stage0_32[484], stage0_32[485]},
      {stage0_34[306], stage0_34[307], stage0_34[308], stage0_34[309], stage0_34[310], stage0_34[311]},
      {stage1_36[51],stage1_35[105],stage1_34[125],stage1_33[156],stage1_32[216]}
   );
   gpc606_5 gpc1302 (
      {stage0_33[324], stage0_33[325], stage0_33[326], stage0_33[327], stage0_33[328], stage0_33[329]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[52],stage1_35[106],stage1_34[126],stage1_33[157]}
   );
   gpc606_5 gpc1303 (
      {stage0_33[330], stage0_33[331], stage0_33[332], stage0_33[333], stage0_33[334], stage0_33[335]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[53],stage1_35[107],stage1_34[127],stage1_33[158]}
   );
   gpc606_5 gpc1304 (
      {stage0_33[336], stage0_33[337], stage0_33[338], stage0_33[339], stage0_33[340], stage0_33[341]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[54],stage1_35[108],stage1_34[128],stage1_33[159]}
   );
   gpc606_5 gpc1305 (
      {stage0_33[342], stage0_33[343], stage0_33[344], stage0_33[345], stage0_33[346], stage0_33[347]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[55],stage1_35[109],stage1_34[129],stage1_33[160]}
   );
   gpc606_5 gpc1306 (
      {stage0_33[348], stage0_33[349], stage0_33[350], stage0_33[351], stage0_33[352], stage0_33[353]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[56],stage1_35[110],stage1_34[130],stage1_33[161]}
   );
   gpc606_5 gpc1307 (
      {stage0_33[354], stage0_33[355], stage0_33[356], stage0_33[357], stage0_33[358], stage0_33[359]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[57],stage1_35[111],stage1_34[131],stage1_33[162]}
   );
   gpc606_5 gpc1308 (
      {stage0_33[360], stage0_33[361], stage0_33[362], stage0_33[363], stage0_33[364], stage0_33[365]},
      {stage0_35[36], stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage1_37[6],stage1_36[58],stage1_35[112],stage1_34[132],stage1_33[163]}
   );
   gpc606_5 gpc1309 (
      {stage0_33[366], stage0_33[367], stage0_33[368], stage0_33[369], stage0_33[370], stage0_33[371]},
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46], stage0_35[47]},
      {stage1_37[7],stage1_36[59],stage1_35[113],stage1_34[133],stage1_33[164]}
   );
   gpc606_5 gpc1310 (
      {stage0_33[372], stage0_33[373], stage0_33[374], stage0_33[375], stage0_33[376], stage0_33[377]},
      {stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51], stage0_35[52], stage0_35[53]},
      {stage1_37[8],stage1_36[60],stage1_35[114],stage1_34[134],stage1_33[165]}
   );
   gpc606_5 gpc1311 (
      {stage0_33[378], stage0_33[379], stage0_33[380], stage0_33[381], stage0_33[382], stage0_33[383]},
      {stage0_35[54], stage0_35[55], stage0_35[56], stage0_35[57], stage0_35[58], stage0_35[59]},
      {stage1_37[9],stage1_36[61],stage1_35[115],stage1_34[135],stage1_33[166]}
   );
   gpc606_5 gpc1312 (
      {stage0_33[384], stage0_33[385], stage0_33[386], stage0_33[387], stage0_33[388], stage0_33[389]},
      {stage0_35[60], stage0_35[61], stage0_35[62], stage0_35[63], stage0_35[64], stage0_35[65]},
      {stage1_37[10],stage1_36[62],stage1_35[116],stage1_34[136],stage1_33[167]}
   );
   gpc606_5 gpc1313 (
      {stage0_33[390], stage0_33[391], stage0_33[392], stage0_33[393], stage0_33[394], stage0_33[395]},
      {stage0_35[66], stage0_35[67], stage0_35[68], stage0_35[69], stage0_35[70], stage0_35[71]},
      {stage1_37[11],stage1_36[63],stage1_35[117],stage1_34[137],stage1_33[168]}
   );
   gpc1163_5 gpc1314 (
      {stage0_34[312], stage0_34[313], stage0_34[314]},
      {stage0_35[72], stage0_35[73], stage0_35[74], stage0_35[75], stage0_35[76], stage0_35[77]},
      {stage0_36[0]},
      {stage0_37[0]},
      {stage1_38[0],stage1_37[12],stage1_36[64],stage1_35[118],stage1_34[138]}
   );
   gpc1163_5 gpc1315 (
      {stage0_34[315], stage0_34[316], stage0_34[317]},
      {stage0_35[78], stage0_35[79], stage0_35[80], stage0_35[81], stage0_35[82], stage0_35[83]},
      {stage0_36[1]},
      {stage0_37[1]},
      {stage1_38[1],stage1_37[13],stage1_36[65],stage1_35[119],stage1_34[139]}
   );
   gpc1163_5 gpc1316 (
      {stage0_34[318], stage0_34[319], stage0_34[320]},
      {stage0_35[84], stage0_35[85], stage0_35[86], stage0_35[87], stage0_35[88], stage0_35[89]},
      {stage0_36[2]},
      {stage0_37[2]},
      {stage1_38[2],stage1_37[14],stage1_36[66],stage1_35[120],stage1_34[140]}
   );
   gpc1163_5 gpc1317 (
      {stage0_34[321], stage0_34[322], stage0_34[323]},
      {stage0_35[90], stage0_35[91], stage0_35[92], stage0_35[93], stage0_35[94], stage0_35[95]},
      {stage0_36[3]},
      {stage0_37[3]},
      {stage1_38[3],stage1_37[15],stage1_36[67],stage1_35[121],stage1_34[141]}
   );
   gpc1163_5 gpc1318 (
      {stage0_34[324], stage0_34[325], stage0_34[326]},
      {stage0_35[96], stage0_35[97], stage0_35[98], stage0_35[99], stage0_35[100], stage0_35[101]},
      {stage0_36[4]},
      {stage0_37[4]},
      {stage1_38[4],stage1_37[16],stage1_36[68],stage1_35[122],stage1_34[142]}
   );
   gpc1163_5 gpc1319 (
      {stage0_34[327], stage0_34[328], stage0_34[329]},
      {stage0_35[102], stage0_35[103], stage0_35[104], stage0_35[105], stage0_35[106], stage0_35[107]},
      {stage0_36[5]},
      {stage0_37[5]},
      {stage1_38[5],stage1_37[17],stage1_36[69],stage1_35[123],stage1_34[143]}
   );
   gpc1163_5 gpc1320 (
      {stage0_34[330], stage0_34[331], stage0_34[332]},
      {stage0_35[108], stage0_35[109], stage0_35[110], stage0_35[111], stage0_35[112], stage0_35[113]},
      {stage0_36[6]},
      {stage0_37[6]},
      {stage1_38[6],stage1_37[18],stage1_36[70],stage1_35[124],stage1_34[144]}
   );
   gpc1163_5 gpc1321 (
      {stage0_34[333], stage0_34[334], stage0_34[335]},
      {stage0_35[114], stage0_35[115], stage0_35[116], stage0_35[117], stage0_35[118], stage0_35[119]},
      {stage0_36[7]},
      {stage0_37[7]},
      {stage1_38[7],stage1_37[19],stage1_36[71],stage1_35[125],stage1_34[145]}
   );
   gpc1163_5 gpc1322 (
      {stage0_34[336], stage0_34[337], stage0_34[338]},
      {stage0_35[120], stage0_35[121], stage0_35[122], stage0_35[123], stage0_35[124], stage0_35[125]},
      {stage0_36[8]},
      {stage0_37[8]},
      {stage1_38[8],stage1_37[20],stage1_36[72],stage1_35[126],stage1_34[146]}
   );
   gpc1163_5 gpc1323 (
      {stage0_34[339], stage0_34[340], stage0_34[341]},
      {stage0_35[126], stage0_35[127], stage0_35[128], stage0_35[129], stage0_35[130], stage0_35[131]},
      {stage0_36[9]},
      {stage0_37[9]},
      {stage1_38[9],stage1_37[21],stage1_36[73],stage1_35[127],stage1_34[147]}
   );
   gpc1163_5 gpc1324 (
      {stage0_34[342], stage0_34[343], stage0_34[344]},
      {stage0_35[132], stage0_35[133], stage0_35[134], stage0_35[135], stage0_35[136], stage0_35[137]},
      {stage0_36[10]},
      {stage0_37[10]},
      {stage1_38[10],stage1_37[22],stage1_36[74],stage1_35[128],stage1_34[148]}
   );
   gpc1163_5 gpc1325 (
      {stage0_34[345], stage0_34[346], stage0_34[347]},
      {stage0_35[138], stage0_35[139], stage0_35[140], stage0_35[141], stage0_35[142], stage0_35[143]},
      {stage0_36[11]},
      {stage0_37[11]},
      {stage1_38[11],stage1_37[23],stage1_36[75],stage1_35[129],stage1_34[149]}
   );
   gpc1163_5 gpc1326 (
      {stage0_34[348], stage0_34[349], stage0_34[350]},
      {stage0_35[144], stage0_35[145], stage0_35[146], stage0_35[147], stage0_35[148], stage0_35[149]},
      {stage0_36[12]},
      {stage0_37[12]},
      {stage1_38[12],stage1_37[24],stage1_36[76],stage1_35[130],stage1_34[150]}
   );
   gpc1163_5 gpc1327 (
      {stage0_34[351], stage0_34[352], stage0_34[353]},
      {stage0_35[150], stage0_35[151], stage0_35[152], stage0_35[153], stage0_35[154], stage0_35[155]},
      {stage0_36[13]},
      {stage0_37[13]},
      {stage1_38[13],stage1_37[25],stage1_36[77],stage1_35[131],stage1_34[151]}
   );
   gpc1163_5 gpc1328 (
      {stage0_34[354], stage0_34[355], stage0_34[356]},
      {stage0_35[156], stage0_35[157], stage0_35[158], stage0_35[159], stage0_35[160], stage0_35[161]},
      {stage0_36[14]},
      {stage0_37[14]},
      {stage1_38[14],stage1_37[26],stage1_36[78],stage1_35[132],stage1_34[152]}
   );
   gpc1163_5 gpc1329 (
      {stage0_34[357], stage0_34[358], stage0_34[359]},
      {stage0_35[162], stage0_35[163], stage0_35[164], stage0_35[165], stage0_35[166], stage0_35[167]},
      {stage0_36[15]},
      {stage0_37[15]},
      {stage1_38[15],stage1_37[27],stage1_36[79],stage1_35[133],stage1_34[153]}
   );
   gpc1163_5 gpc1330 (
      {stage0_34[360], stage0_34[361], stage0_34[362]},
      {stage0_35[168], stage0_35[169], stage0_35[170], stage0_35[171], stage0_35[172], stage0_35[173]},
      {stage0_36[16]},
      {stage0_37[16]},
      {stage1_38[16],stage1_37[28],stage1_36[80],stage1_35[134],stage1_34[154]}
   );
   gpc1163_5 gpc1331 (
      {stage0_34[363], stage0_34[364], stage0_34[365]},
      {stage0_35[174], stage0_35[175], stage0_35[176], stage0_35[177], stage0_35[178], stage0_35[179]},
      {stage0_36[17]},
      {stage0_37[17]},
      {stage1_38[17],stage1_37[29],stage1_36[81],stage1_35[135],stage1_34[155]}
   );
   gpc1163_5 gpc1332 (
      {stage0_34[366], stage0_34[367], stage0_34[368]},
      {stage0_35[180], stage0_35[181], stage0_35[182], stage0_35[183], stage0_35[184], stage0_35[185]},
      {stage0_36[18]},
      {stage0_37[18]},
      {stage1_38[18],stage1_37[30],stage1_36[82],stage1_35[136],stage1_34[156]}
   );
   gpc1163_5 gpc1333 (
      {stage0_34[369], stage0_34[370], stage0_34[371]},
      {stage0_35[186], stage0_35[187], stage0_35[188], stage0_35[189], stage0_35[190], stage0_35[191]},
      {stage0_36[19]},
      {stage0_37[19]},
      {stage1_38[19],stage1_37[31],stage1_36[83],stage1_35[137],stage1_34[157]}
   );
   gpc1163_5 gpc1334 (
      {stage0_34[372], stage0_34[373], stage0_34[374]},
      {stage0_35[192], stage0_35[193], stage0_35[194], stage0_35[195], stage0_35[196], stage0_35[197]},
      {stage0_36[20]},
      {stage0_37[20]},
      {stage1_38[20],stage1_37[32],stage1_36[84],stage1_35[138],stage1_34[158]}
   );
   gpc1163_5 gpc1335 (
      {stage0_34[375], stage0_34[376], stage0_34[377]},
      {stage0_35[198], stage0_35[199], stage0_35[200], stage0_35[201], stage0_35[202], stage0_35[203]},
      {stage0_36[21]},
      {stage0_37[21]},
      {stage1_38[21],stage1_37[33],stage1_36[85],stage1_35[139],stage1_34[159]}
   );
   gpc1163_5 gpc1336 (
      {stage0_34[378], stage0_34[379], stage0_34[380]},
      {stage0_35[204], stage0_35[205], stage0_35[206], stage0_35[207], stage0_35[208], stage0_35[209]},
      {stage0_36[22]},
      {stage0_37[22]},
      {stage1_38[22],stage1_37[34],stage1_36[86],stage1_35[140],stage1_34[160]}
   );
   gpc1163_5 gpc1337 (
      {stage0_34[381], stage0_34[382], stage0_34[383]},
      {stage0_35[210], stage0_35[211], stage0_35[212], stage0_35[213], stage0_35[214], stage0_35[215]},
      {stage0_36[23]},
      {stage0_37[23]},
      {stage1_38[23],stage1_37[35],stage1_36[87],stage1_35[141],stage1_34[161]}
   );
   gpc1163_5 gpc1338 (
      {stage0_34[384], stage0_34[385], stage0_34[386]},
      {stage0_35[216], stage0_35[217], stage0_35[218], stage0_35[219], stage0_35[220], stage0_35[221]},
      {stage0_36[24]},
      {stage0_37[24]},
      {stage1_38[24],stage1_37[36],stage1_36[88],stage1_35[142],stage1_34[162]}
   );
   gpc1163_5 gpc1339 (
      {stage0_34[387], stage0_34[388], stage0_34[389]},
      {stage0_35[222], stage0_35[223], stage0_35[224], stage0_35[225], stage0_35[226], stage0_35[227]},
      {stage0_36[25]},
      {stage0_37[25]},
      {stage1_38[25],stage1_37[37],stage1_36[89],stage1_35[143],stage1_34[163]}
   );
   gpc1163_5 gpc1340 (
      {stage0_34[390], stage0_34[391], stage0_34[392]},
      {stage0_35[228], stage0_35[229], stage0_35[230], stage0_35[231], stage0_35[232], stage0_35[233]},
      {stage0_36[26]},
      {stage0_37[26]},
      {stage1_38[26],stage1_37[38],stage1_36[90],stage1_35[144],stage1_34[164]}
   );
   gpc1163_5 gpc1341 (
      {stage0_34[393], stage0_34[394], stage0_34[395]},
      {stage0_35[234], stage0_35[235], stage0_35[236], stage0_35[237], stage0_35[238], stage0_35[239]},
      {stage0_36[27]},
      {stage0_37[27]},
      {stage1_38[27],stage1_37[39],stage1_36[91],stage1_35[145],stage1_34[165]}
   );
   gpc1163_5 gpc1342 (
      {stage0_34[396], stage0_34[397], stage0_34[398]},
      {stage0_35[240], stage0_35[241], stage0_35[242], stage0_35[243], stage0_35[244], stage0_35[245]},
      {stage0_36[28]},
      {stage0_37[28]},
      {stage1_38[28],stage1_37[40],stage1_36[92],stage1_35[146],stage1_34[166]}
   );
   gpc1163_5 gpc1343 (
      {stage0_34[399], stage0_34[400], stage0_34[401]},
      {stage0_35[246], stage0_35[247], stage0_35[248], stage0_35[249], stage0_35[250], stage0_35[251]},
      {stage0_36[29]},
      {stage0_37[29]},
      {stage1_38[29],stage1_37[41],stage1_36[93],stage1_35[147],stage1_34[167]}
   );
   gpc1163_5 gpc1344 (
      {stage0_34[402], stage0_34[403], stage0_34[404]},
      {stage0_35[252], stage0_35[253], stage0_35[254], stage0_35[255], stage0_35[256], stage0_35[257]},
      {stage0_36[30]},
      {stage0_37[30]},
      {stage1_38[30],stage1_37[42],stage1_36[94],stage1_35[148],stage1_34[168]}
   );
   gpc1163_5 gpc1345 (
      {stage0_34[405], stage0_34[406], stage0_34[407]},
      {stage0_35[258], stage0_35[259], stage0_35[260], stage0_35[261], stage0_35[262], stage0_35[263]},
      {stage0_36[31]},
      {stage0_37[31]},
      {stage1_38[31],stage1_37[43],stage1_36[95],stage1_35[149],stage1_34[169]}
   );
   gpc1163_5 gpc1346 (
      {stage0_34[408], stage0_34[409], stage0_34[410]},
      {stage0_35[264], stage0_35[265], stage0_35[266], stage0_35[267], stage0_35[268], stage0_35[269]},
      {stage0_36[32]},
      {stage0_37[32]},
      {stage1_38[32],stage1_37[44],stage1_36[96],stage1_35[150],stage1_34[170]}
   );
   gpc1163_5 gpc1347 (
      {stage0_34[411], stage0_34[412], stage0_34[413]},
      {stage0_35[270], stage0_35[271], stage0_35[272], stage0_35[273], stage0_35[274], stage0_35[275]},
      {stage0_36[33]},
      {stage0_37[33]},
      {stage1_38[33],stage1_37[45],stage1_36[97],stage1_35[151],stage1_34[171]}
   );
   gpc1163_5 gpc1348 (
      {stage0_34[414], stage0_34[415], stage0_34[416]},
      {stage0_35[276], stage0_35[277], stage0_35[278], stage0_35[279], stage0_35[280], stage0_35[281]},
      {stage0_36[34]},
      {stage0_37[34]},
      {stage1_38[34],stage1_37[46],stage1_36[98],stage1_35[152],stage1_34[172]}
   );
   gpc1163_5 gpc1349 (
      {stage0_34[417], stage0_34[418], stage0_34[419]},
      {stage0_35[282], stage0_35[283], stage0_35[284], stage0_35[285], stage0_35[286], stage0_35[287]},
      {stage0_36[35]},
      {stage0_37[35]},
      {stage1_38[35],stage1_37[47],stage1_36[99],stage1_35[153],stage1_34[173]}
   );
   gpc1163_5 gpc1350 (
      {stage0_34[420], stage0_34[421], stage0_34[422]},
      {stage0_35[288], stage0_35[289], stage0_35[290], stage0_35[291], stage0_35[292], stage0_35[293]},
      {stage0_36[36]},
      {stage0_37[36]},
      {stage1_38[36],stage1_37[48],stage1_36[100],stage1_35[154],stage1_34[174]}
   );
   gpc1163_5 gpc1351 (
      {stage0_34[423], stage0_34[424], stage0_34[425]},
      {stage0_35[294], stage0_35[295], stage0_35[296], stage0_35[297], stage0_35[298], stage0_35[299]},
      {stage0_36[37]},
      {stage0_37[37]},
      {stage1_38[37],stage1_37[49],stage1_36[101],stage1_35[155],stage1_34[175]}
   );
   gpc1163_5 gpc1352 (
      {stage0_34[426], stage0_34[427], stage0_34[428]},
      {stage0_35[300], stage0_35[301], stage0_35[302], stage0_35[303], stage0_35[304], stage0_35[305]},
      {stage0_36[38]},
      {stage0_37[38]},
      {stage1_38[38],stage1_37[50],stage1_36[102],stage1_35[156],stage1_34[176]}
   );
   gpc1163_5 gpc1353 (
      {stage0_34[429], stage0_34[430], stage0_34[431]},
      {stage0_35[306], stage0_35[307], stage0_35[308], stage0_35[309], stage0_35[310], stage0_35[311]},
      {stage0_36[39]},
      {stage0_37[39]},
      {stage1_38[39],stage1_37[51],stage1_36[103],stage1_35[157],stage1_34[177]}
   );
   gpc1163_5 gpc1354 (
      {stage0_34[432], stage0_34[433], stage0_34[434]},
      {stage0_35[312], stage0_35[313], stage0_35[314], stage0_35[315], stage0_35[316], stage0_35[317]},
      {stage0_36[40]},
      {stage0_37[40]},
      {stage1_38[40],stage1_37[52],stage1_36[104],stage1_35[158],stage1_34[178]}
   );
   gpc1163_5 gpc1355 (
      {stage0_34[435], stage0_34[436], stage0_34[437]},
      {stage0_35[318], stage0_35[319], stage0_35[320], stage0_35[321], stage0_35[322], stage0_35[323]},
      {stage0_36[41]},
      {stage0_37[41]},
      {stage1_38[41],stage1_37[53],stage1_36[105],stage1_35[159],stage1_34[179]}
   );
   gpc1163_5 gpc1356 (
      {stage0_34[438], stage0_34[439], stage0_34[440]},
      {stage0_35[324], stage0_35[325], stage0_35[326], stage0_35[327], stage0_35[328], stage0_35[329]},
      {stage0_36[42]},
      {stage0_37[42]},
      {stage1_38[42],stage1_37[54],stage1_36[106],stage1_35[160],stage1_34[180]}
   );
   gpc615_5 gpc1357 (
      {stage0_34[441], stage0_34[442], stage0_34[443], stage0_34[444], stage0_34[445]},
      {stage0_35[330]},
      {stage0_36[43], stage0_36[44], stage0_36[45], stage0_36[46], stage0_36[47], stage0_36[48]},
      {stage1_38[43],stage1_37[55],stage1_36[107],stage1_35[161],stage1_34[181]}
   );
   gpc615_5 gpc1358 (
      {stage0_34[446], stage0_34[447], stage0_34[448], stage0_34[449], stage0_34[450]},
      {stage0_35[331]},
      {stage0_36[49], stage0_36[50], stage0_36[51], stage0_36[52], stage0_36[53], stage0_36[54]},
      {stage1_38[44],stage1_37[56],stage1_36[108],stage1_35[162],stage1_34[182]}
   );
   gpc615_5 gpc1359 (
      {stage0_34[451], stage0_34[452], stage0_34[453], stage0_34[454], stage0_34[455]},
      {stage0_35[332]},
      {stage0_36[55], stage0_36[56], stage0_36[57], stage0_36[58], stage0_36[59], stage0_36[60]},
      {stage1_38[45],stage1_37[57],stage1_36[109],stage1_35[163],stage1_34[183]}
   );
   gpc615_5 gpc1360 (
      {stage0_34[456], stage0_34[457], stage0_34[458], stage0_34[459], stage0_34[460]},
      {stage0_35[333]},
      {stage0_36[61], stage0_36[62], stage0_36[63], stage0_36[64], stage0_36[65], stage0_36[66]},
      {stage1_38[46],stage1_37[58],stage1_36[110],stage1_35[164],stage1_34[184]}
   );
   gpc615_5 gpc1361 (
      {stage0_34[461], stage0_34[462], stage0_34[463], stage0_34[464], stage0_34[465]},
      {stage0_35[334]},
      {stage0_36[67], stage0_36[68], stage0_36[69], stage0_36[70], stage0_36[71], stage0_36[72]},
      {stage1_38[47],stage1_37[59],stage1_36[111],stage1_35[165],stage1_34[185]}
   );
   gpc615_5 gpc1362 (
      {stage0_34[466], stage0_34[467], stage0_34[468], stage0_34[469], stage0_34[470]},
      {stage0_35[335]},
      {stage0_36[73], stage0_36[74], stage0_36[75], stage0_36[76], stage0_36[77], stage0_36[78]},
      {stage1_38[48],stage1_37[60],stage1_36[112],stage1_35[166],stage1_34[186]}
   );
   gpc615_5 gpc1363 (
      {stage0_34[471], stage0_34[472], stage0_34[473], stage0_34[474], stage0_34[475]},
      {stage0_35[336]},
      {stage0_36[79], stage0_36[80], stage0_36[81], stage0_36[82], stage0_36[83], stage0_36[84]},
      {stage1_38[49],stage1_37[61],stage1_36[113],stage1_35[167],stage1_34[187]}
   );
   gpc615_5 gpc1364 (
      {stage0_34[476], stage0_34[477], stage0_34[478], stage0_34[479], stage0_34[480]},
      {stage0_35[337]},
      {stage0_36[85], stage0_36[86], stage0_36[87], stage0_36[88], stage0_36[89], stage0_36[90]},
      {stage1_38[50],stage1_37[62],stage1_36[114],stage1_35[168],stage1_34[188]}
   );
   gpc615_5 gpc1365 (
      {stage0_34[481], stage0_34[482], stage0_34[483], stage0_34[484], stage0_34[485]},
      {stage0_35[338]},
      {stage0_36[91], stage0_36[92], stage0_36[93], stage0_36[94], stage0_36[95], stage0_36[96]},
      {stage1_38[51],stage1_37[63],stage1_36[115],stage1_35[169],stage1_34[189]}
   );
   gpc615_5 gpc1366 (
      {stage0_35[339], stage0_35[340], stage0_35[341], stage0_35[342], stage0_35[343]},
      {stage0_36[97]},
      {stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47], stage0_37[48]},
      {stage1_39[0],stage1_38[52],stage1_37[64],stage1_36[116],stage1_35[170]}
   );
   gpc615_5 gpc1367 (
      {stage0_35[344], stage0_35[345], stage0_35[346], stage0_35[347], stage0_35[348]},
      {stage0_36[98]},
      {stage0_37[49], stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53], stage0_37[54]},
      {stage1_39[1],stage1_38[53],stage1_37[65],stage1_36[117],stage1_35[171]}
   );
   gpc615_5 gpc1368 (
      {stage0_35[349], stage0_35[350], stage0_35[351], stage0_35[352], stage0_35[353]},
      {stage0_36[99]},
      {stage0_37[55], stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59], stage0_37[60]},
      {stage1_39[2],stage1_38[54],stage1_37[66],stage1_36[118],stage1_35[172]}
   );
   gpc615_5 gpc1369 (
      {stage0_35[354], stage0_35[355], stage0_35[356], stage0_35[357], stage0_35[358]},
      {stage0_36[100]},
      {stage0_37[61], stage0_37[62], stage0_37[63], stage0_37[64], stage0_37[65], stage0_37[66]},
      {stage1_39[3],stage1_38[55],stage1_37[67],stage1_36[119],stage1_35[173]}
   );
   gpc615_5 gpc1370 (
      {stage0_35[359], stage0_35[360], stage0_35[361], stage0_35[362], stage0_35[363]},
      {stage0_36[101]},
      {stage0_37[67], stage0_37[68], stage0_37[69], stage0_37[70], stage0_37[71], stage0_37[72]},
      {stage1_39[4],stage1_38[56],stage1_37[68],stage1_36[120],stage1_35[174]}
   );
   gpc615_5 gpc1371 (
      {stage0_35[364], stage0_35[365], stage0_35[366], stage0_35[367], stage0_35[368]},
      {stage0_36[102]},
      {stage0_37[73], stage0_37[74], stage0_37[75], stage0_37[76], stage0_37[77], stage0_37[78]},
      {stage1_39[5],stage1_38[57],stage1_37[69],stage1_36[121],stage1_35[175]}
   );
   gpc615_5 gpc1372 (
      {stage0_35[369], stage0_35[370], stage0_35[371], stage0_35[372], stage0_35[373]},
      {stage0_36[103]},
      {stage0_37[79], stage0_37[80], stage0_37[81], stage0_37[82], stage0_37[83], stage0_37[84]},
      {stage1_39[6],stage1_38[58],stage1_37[70],stage1_36[122],stage1_35[176]}
   );
   gpc615_5 gpc1373 (
      {stage0_35[374], stage0_35[375], stage0_35[376], stage0_35[377], stage0_35[378]},
      {stage0_36[104]},
      {stage0_37[85], stage0_37[86], stage0_37[87], stage0_37[88], stage0_37[89], stage0_37[90]},
      {stage1_39[7],stage1_38[59],stage1_37[71],stage1_36[123],stage1_35[177]}
   );
   gpc615_5 gpc1374 (
      {stage0_35[379], stage0_35[380], stage0_35[381], stage0_35[382], stage0_35[383]},
      {stage0_36[105]},
      {stage0_37[91], stage0_37[92], stage0_37[93], stage0_37[94], stage0_37[95], stage0_37[96]},
      {stage1_39[8],stage1_38[60],stage1_37[72],stage1_36[124],stage1_35[178]}
   );
   gpc615_5 gpc1375 (
      {stage0_35[384], stage0_35[385], stage0_35[386], stage0_35[387], stage0_35[388]},
      {stage0_36[106]},
      {stage0_37[97], stage0_37[98], stage0_37[99], stage0_37[100], stage0_37[101], stage0_37[102]},
      {stage1_39[9],stage1_38[61],stage1_37[73],stage1_36[125],stage1_35[179]}
   );
   gpc615_5 gpc1376 (
      {stage0_35[389], stage0_35[390], stage0_35[391], stage0_35[392], stage0_35[393]},
      {stage0_36[107]},
      {stage0_37[103], stage0_37[104], stage0_37[105], stage0_37[106], stage0_37[107], stage0_37[108]},
      {stage1_39[10],stage1_38[62],stage1_37[74],stage1_36[126],stage1_35[180]}
   );
   gpc615_5 gpc1377 (
      {stage0_35[394], stage0_35[395], stage0_35[396], stage0_35[397], stage0_35[398]},
      {stage0_36[108]},
      {stage0_37[109], stage0_37[110], stage0_37[111], stage0_37[112], stage0_37[113], stage0_37[114]},
      {stage1_39[11],stage1_38[63],stage1_37[75],stage1_36[127],stage1_35[181]}
   );
   gpc615_5 gpc1378 (
      {stage0_35[399], stage0_35[400], stage0_35[401], stage0_35[402], stage0_35[403]},
      {stage0_36[109]},
      {stage0_37[115], stage0_37[116], stage0_37[117], stage0_37[118], stage0_37[119], stage0_37[120]},
      {stage1_39[12],stage1_38[64],stage1_37[76],stage1_36[128],stage1_35[182]}
   );
   gpc615_5 gpc1379 (
      {stage0_35[404], stage0_35[405], stage0_35[406], stage0_35[407], stage0_35[408]},
      {stage0_36[110]},
      {stage0_37[121], stage0_37[122], stage0_37[123], stage0_37[124], stage0_37[125], stage0_37[126]},
      {stage1_39[13],stage1_38[65],stage1_37[77],stage1_36[129],stage1_35[183]}
   );
   gpc615_5 gpc1380 (
      {stage0_35[409], stage0_35[410], stage0_35[411], stage0_35[412], stage0_35[413]},
      {stage0_36[111]},
      {stage0_37[127], stage0_37[128], stage0_37[129], stage0_37[130], stage0_37[131], stage0_37[132]},
      {stage1_39[14],stage1_38[66],stage1_37[78],stage1_36[130],stage1_35[184]}
   );
   gpc615_5 gpc1381 (
      {stage0_35[414], stage0_35[415], stage0_35[416], stage0_35[417], stage0_35[418]},
      {stage0_36[112]},
      {stage0_37[133], stage0_37[134], stage0_37[135], stage0_37[136], stage0_37[137], stage0_37[138]},
      {stage1_39[15],stage1_38[67],stage1_37[79],stage1_36[131],stage1_35[185]}
   );
   gpc615_5 gpc1382 (
      {stage0_35[419], stage0_35[420], stage0_35[421], stage0_35[422], stage0_35[423]},
      {stage0_36[113]},
      {stage0_37[139], stage0_37[140], stage0_37[141], stage0_37[142], stage0_37[143], stage0_37[144]},
      {stage1_39[16],stage1_38[68],stage1_37[80],stage1_36[132],stage1_35[186]}
   );
   gpc615_5 gpc1383 (
      {stage0_35[424], stage0_35[425], stage0_35[426], stage0_35[427], stage0_35[428]},
      {stage0_36[114]},
      {stage0_37[145], stage0_37[146], stage0_37[147], stage0_37[148], stage0_37[149], stage0_37[150]},
      {stage1_39[17],stage1_38[69],stage1_37[81],stage1_36[133],stage1_35[187]}
   );
   gpc615_5 gpc1384 (
      {stage0_35[429], stage0_35[430], stage0_35[431], stage0_35[432], stage0_35[433]},
      {stage0_36[115]},
      {stage0_37[151], stage0_37[152], stage0_37[153], stage0_37[154], stage0_37[155], stage0_37[156]},
      {stage1_39[18],stage1_38[70],stage1_37[82],stage1_36[134],stage1_35[188]}
   );
   gpc615_5 gpc1385 (
      {stage0_35[434], stage0_35[435], stage0_35[436], stage0_35[437], stage0_35[438]},
      {stage0_36[116]},
      {stage0_37[157], stage0_37[158], stage0_37[159], stage0_37[160], stage0_37[161], stage0_37[162]},
      {stage1_39[19],stage1_38[71],stage1_37[83],stage1_36[135],stage1_35[189]}
   );
   gpc615_5 gpc1386 (
      {stage0_35[439], stage0_35[440], stage0_35[441], stage0_35[442], stage0_35[443]},
      {stage0_36[117]},
      {stage0_37[163], stage0_37[164], stage0_37[165], stage0_37[166], stage0_37[167], stage0_37[168]},
      {stage1_39[20],stage1_38[72],stage1_37[84],stage1_36[136],stage1_35[190]}
   );
   gpc615_5 gpc1387 (
      {stage0_35[444], stage0_35[445], stage0_35[446], stage0_35[447], stage0_35[448]},
      {stage0_36[118]},
      {stage0_37[169], stage0_37[170], stage0_37[171], stage0_37[172], stage0_37[173], stage0_37[174]},
      {stage1_39[21],stage1_38[73],stage1_37[85],stage1_36[137],stage1_35[191]}
   );
   gpc615_5 gpc1388 (
      {stage0_35[449], stage0_35[450], stage0_35[451], stage0_35[452], stage0_35[453]},
      {stage0_36[119]},
      {stage0_37[175], stage0_37[176], stage0_37[177], stage0_37[178], stage0_37[179], stage0_37[180]},
      {stage1_39[22],stage1_38[74],stage1_37[86],stage1_36[138],stage1_35[192]}
   );
   gpc615_5 gpc1389 (
      {stage0_35[454], stage0_35[455], stage0_35[456], stage0_35[457], stage0_35[458]},
      {stage0_36[120]},
      {stage0_37[181], stage0_37[182], stage0_37[183], stage0_37[184], stage0_37[185], stage0_37[186]},
      {stage1_39[23],stage1_38[75],stage1_37[87],stage1_36[139],stage1_35[193]}
   );
   gpc615_5 gpc1390 (
      {stage0_35[459], stage0_35[460], stage0_35[461], stage0_35[462], stage0_35[463]},
      {stage0_36[121]},
      {stage0_37[187], stage0_37[188], stage0_37[189], stage0_37[190], stage0_37[191], stage0_37[192]},
      {stage1_39[24],stage1_38[76],stage1_37[88],stage1_36[140],stage1_35[194]}
   );
   gpc606_5 gpc1391 (
      {stage0_36[122], stage0_36[123], stage0_36[124], stage0_36[125], stage0_36[126], stage0_36[127]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[25],stage1_38[77],stage1_37[89],stage1_36[141]}
   );
   gpc606_5 gpc1392 (
      {stage0_36[128], stage0_36[129], stage0_36[130], stage0_36[131], stage0_36[132], stage0_36[133]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[26],stage1_38[78],stage1_37[90],stage1_36[142]}
   );
   gpc606_5 gpc1393 (
      {stage0_36[134], stage0_36[135], stage0_36[136], stage0_36[137], stage0_36[138], stage0_36[139]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[27],stage1_38[79],stage1_37[91],stage1_36[143]}
   );
   gpc606_5 gpc1394 (
      {stage0_36[140], stage0_36[141], stage0_36[142], stage0_36[143], stage0_36[144], stage0_36[145]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[28],stage1_38[80],stage1_37[92],stage1_36[144]}
   );
   gpc606_5 gpc1395 (
      {stage0_36[146], stage0_36[147], stage0_36[148], stage0_36[149], stage0_36[150], stage0_36[151]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[29],stage1_38[81],stage1_37[93],stage1_36[145]}
   );
   gpc606_5 gpc1396 (
      {stage0_36[152], stage0_36[153], stage0_36[154], stage0_36[155], stage0_36[156], stage0_36[157]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[30],stage1_38[82],stage1_37[94],stage1_36[146]}
   );
   gpc606_5 gpc1397 (
      {stage0_36[158], stage0_36[159], stage0_36[160], stage0_36[161], stage0_36[162], stage0_36[163]},
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40], stage0_38[41]},
      {stage1_40[6],stage1_39[31],stage1_38[83],stage1_37[95],stage1_36[147]}
   );
   gpc606_5 gpc1398 (
      {stage0_36[164], stage0_36[165], stage0_36[166], stage0_36[167], stage0_36[168], stage0_36[169]},
      {stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45], stage0_38[46], stage0_38[47]},
      {stage1_40[7],stage1_39[32],stage1_38[84],stage1_37[96],stage1_36[148]}
   );
   gpc606_5 gpc1399 (
      {stage0_36[170], stage0_36[171], stage0_36[172], stage0_36[173], stage0_36[174], stage0_36[175]},
      {stage0_38[48], stage0_38[49], stage0_38[50], stage0_38[51], stage0_38[52], stage0_38[53]},
      {stage1_40[8],stage1_39[33],stage1_38[85],stage1_37[97],stage1_36[149]}
   );
   gpc606_5 gpc1400 (
      {stage0_36[176], stage0_36[177], stage0_36[178], stage0_36[179], stage0_36[180], stage0_36[181]},
      {stage0_38[54], stage0_38[55], stage0_38[56], stage0_38[57], stage0_38[58], stage0_38[59]},
      {stage1_40[9],stage1_39[34],stage1_38[86],stage1_37[98],stage1_36[150]}
   );
   gpc606_5 gpc1401 (
      {stage0_36[182], stage0_36[183], stage0_36[184], stage0_36[185], stage0_36[186], stage0_36[187]},
      {stage0_38[60], stage0_38[61], stage0_38[62], stage0_38[63], stage0_38[64], stage0_38[65]},
      {stage1_40[10],stage1_39[35],stage1_38[87],stage1_37[99],stage1_36[151]}
   );
   gpc606_5 gpc1402 (
      {stage0_36[188], stage0_36[189], stage0_36[190], stage0_36[191], stage0_36[192], stage0_36[193]},
      {stage0_38[66], stage0_38[67], stage0_38[68], stage0_38[69], stage0_38[70], stage0_38[71]},
      {stage1_40[11],stage1_39[36],stage1_38[88],stage1_37[100],stage1_36[152]}
   );
   gpc606_5 gpc1403 (
      {stage0_36[194], stage0_36[195], stage0_36[196], stage0_36[197], stage0_36[198], stage0_36[199]},
      {stage0_38[72], stage0_38[73], stage0_38[74], stage0_38[75], stage0_38[76], stage0_38[77]},
      {stage1_40[12],stage1_39[37],stage1_38[89],stage1_37[101],stage1_36[153]}
   );
   gpc606_5 gpc1404 (
      {stage0_36[200], stage0_36[201], stage0_36[202], stage0_36[203], stage0_36[204], stage0_36[205]},
      {stage0_38[78], stage0_38[79], stage0_38[80], stage0_38[81], stage0_38[82], stage0_38[83]},
      {stage1_40[13],stage1_39[38],stage1_38[90],stage1_37[102],stage1_36[154]}
   );
   gpc606_5 gpc1405 (
      {stage0_36[206], stage0_36[207], stage0_36[208], stage0_36[209], stage0_36[210], stage0_36[211]},
      {stage0_38[84], stage0_38[85], stage0_38[86], stage0_38[87], stage0_38[88], stage0_38[89]},
      {stage1_40[14],stage1_39[39],stage1_38[91],stage1_37[103],stage1_36[155]}
   );
   gpc606_5 gpc1406 (
      {stage0_36[212], stage0_36[213], stage0_36[214], stage0_36[215], stage0_36[216], stage0_36[217]},
      {stage0_38[90], stage0_38[91], stage0_38[92], stage0_38[93], stage0_38[94], stage0_38[95]},
      {stage1_40[15],stage1_39[40],stage1_38[92],stage1_37[104],stage1_36[156]}
   );
   gpc606_5 gpc1407 (
      {stage0_36[218], stage0_36[219], stage0_36[220], stage0_36[221], stage0_36[222], stage0_36[223]},
      {stage0_38[96], stage0_38[97], stage0_38[98], stage0_38[99], stage0_38[100], stage0_38[101]},
      {stage1_40[16],stage1_39[41],stage1_38[93],stage1_37[105],stage1_36[157]}
   );
   gpc606_5 gpc1408 (
      {stage0_36[224], stage0_36[225], stage0_36[226], stage0_36[227], stage0_36[228], stage0_36[229]},
      {stage0_38[102], stage0_38[103], stage0_38[104], stage0_38[105], stage0_38[106], stage0_38[107]},
      {stage1_40[17],stage1_39[42],stage1_38[94],stage1_37[106],stage1_36[158]}
   );
   gpc606_5 gpc1409 (
      {stage0_36[230], stage0_36[231], stage0_36[232], stage0_36[233], stage0_36[234], stage0_36[235]},
      {stage0_38[108], stage0_38[109], stage0_38[110], stage0_38[111], stage0_38[112], stage0_38[113]},
      {stage1_40[18],stage1_39[43],stage1_38[95],stage1_37[107],stage1_36[159]}
   );
   gpc606_5 gpc1410 (
      {stage0_36[236], stage0_36[237], stage0_36[238], stage0_36[239], stage0_36[240], stage0_36[241]},
      {stage0_38[114], stage0_38[115], stage0_38[116], stage0_38[117], stage0_38[118], stage0_38[119]},
      {stage1_40[19],stage1_39[44],stage1_38[96],stage1_37[108],stage1_36[160]}
   );
   gpc606_5 gpc1411 (
      {stage0_36[242], stage0_36[243], stage0_36[244], stage0_36[245], stage0_36[246], stage0_36[247]},
      {stage0_38[120], stage0_38[121], stage0_38[122], stage0_38[123], stage0_38[124], stage0_38[125]},
      {stage1_40[20],stage1_39[45],stage1_38[97],stage1_37[109],stage1_36[161]}
   );
   gpc606_5 gpc1412 (
      {stage0_36[248], stage0_36[249], stage0_36[250], stage0_36[251], stage0_36[252], stage0_36[253]},
      {stage0_38[126], stage0_38[127], stage0_38[128], stage0_38[129], stage0_38[130], stage0_38[131]},
      {stage1_40[21],stage1_39[46],stage1_38[98],stage1_37[110],stage1_36[162]}
   );
   gpc606_5 gpc1413 (
      {stage0_36[254], stage0_36[255], stage0_36[256], stage0_36[257], stage0_36[258], stage0_36[259]},
      {stage0_38[132], stage0_38[133], stage0_38[134], stage0_38[135], stage0_38[136], stage0_38[137]},
      {stage1_40[22],stage1_39[47],stage1_38[99],stage1_37[111],stage1_36[163]}
   );
   gpc606_5 gpc1414 (
      {stage0_36[260], stage0_36[261], stage0_36[262], stage0_36[263], stage0_36[264], stage0_36[265]},
      {stage0_38[138], stage0_38[139], stage0_38[140], stage0_38[141], stage0_38[142], stage0_38[143]},
      {stage1_40[23],stage1_39[48],stage1_38[100],stage1_37[112],stage1_36[164]}
   );
   gpc606_5 gpc1415 (
      {stage0_36[266], stage0_36[267], stage0_36[268], stage0_36[269], stage0_36[270], stage0_36[271]},
      {stage0_38[144], stage0_38[145], stage0_38[146], stage0_38[147], stage0_38[148], stage0_38[149]},
      {stage1_40[24],stage1_39[49],stage1_38[101],stage1_37[113],stage1_36[165]}
   );
   gpc606_5 gpc1416 (
      {stage0_36[272], stage0_36[273], stage0_36[274], stage0_36[275], stage0_36[276], stage0_36[277]},
      {stage0_38[150], stage0_38[151], stage0_38[152], stage0_38[153], stage0_38[154], stage0_38[155]},
      {stage1_40[25],stage1_39[50],stage1_38[102],stage1_37[114],stage1_36[166]}
   );
   gpc606_5 gpc1417 (
      {stage0_36[278], stage0_36[279], stage0_36[280], stage0_36[281], stage0_36[282], stage0_36[283]},
      {stage0_38[156], stage0_38[157], stage0_38[158], stage0_38[159], stage0_38[160], stage0_38[161]},
      {stage1_40[26],stage1_39[51],stage1_38[103],stage1_37[115],stage1_36[167]}
   );
   gpc606_5 gpc1418 (
      {stage0_36[284], stage0_36[285], stage0_36[286], stage0_36[287], stage0_36[288], stage0_36[289]},
      {stage0_38[162], stage0_38[163], stage0_38[164], stage0_38[165], stage0_38[166], stage0_38[167]},
      {stage1_40[27],stage1_39[52],stage1_38[104],stage1_37[116],stage1_36[168]}
   );
   gpc606_5 gpc1419 (
      {stage0_36[290], stage0_36[291], stage0_36[292], stage0_36[293], stage0_36[294], stage0_36[295]},
      {stage0_38[168], stage0_38[169], stage0_38[170], stage0_38[171], stage0_38[172], stage0_38[173]},
      {stage1_40[28],stage1_39[53],stage1_38[105],stage1_37[117],stage1_36[169]}
   );
   gpc606_5 gpc1420 (
      {stage0_36[296], stage0_36[297], stage0_36[298], stage0_36[299], stage0_36[300], stage0_36[301]},
      {stage0_38[174], stage0_38[175], stage0_38[176], stage0_38[177], stage0_38[178], stage0_38[179]},
      {stage1_40[29],stage1_39[54],stage1_38[106],stage1_37[118],stage1_36[170]}
   );
   gpc606_5 gpc1421 (
      {stage0_36[302], stage0_36[303], stage0_36[304], stage0_36[305], stage0_36[306], stage0_36[307]},
      {stage0_38[180], stage0_38[181], stage0_38[182], stage0_38[183], stage0_38[184], stage0_38[185]},
      {stage1_40[30],stage1_39[55],stage1_38[107],stage1_37[119],stage1_36[171]}
   );
   gpc606_5 gpc1422 (
      {stage0_36[308], stage0_36[309], stage0_36[310], stage0_36[311], stage0_36[312], stage0_36[313]},
      {stage0_38[186], stage0_38[187], stage0_38[188], stage0_38[189], stage0_38[190], stage0_38[191]},
      {stage1_40[31],stage1_39[56],stage1_38[108],stage1_37[120],stage1_36[172]}
   );
   gpc606_5 gpc1423 (
      {stage0_36[314], stage0_36[315], stage0_36[316], stage0_36[317], stage0_36[318], stage0_36[319]},
      {stage0_38[192], stage0_38[193], stage0_38[194], stage0_38[195], stage0_38[196], stage0_38[197]},
      {stage1_40[32],stage1_39[57],stage1_38[109],stage1_37[121],stage1_36[173]}
   );
   gpc606_5 gpc1424 (
      {stage0_36[320], stage0_36[321], stage0_36[322], stage0_36[323], stage0_36[324], stage0_36[325]},
      {stage0_38[198], stage0_38[199], stage0_38[200], stage0_38[201], stage0_38[202], stage0_38[203]},
      {stage1_40[33],stage1_39[58],stage1_38[110],stage1_37[122],stage1_36[174]}
   );
   gpc606_5 gpc1425 (
      {stage0_36[326], stage0_36[327], stage0_36[328], stage0_36[329], stage0_36[330], stage0_36[331]},
      {stage0_38[204], stage0_38[205], stage0_38[206], stage0_38[207], stage0_38[208], stage0_38[209]},
      {stage1_40[34],stage1_39[59],stage1_38[111],stage1_37[123],stage1_36[175]}
   );
   gpc606_5 gpc1426 (
      {stage0_36[332], stage0_36[333], stage0_36[334], stage0_36[335], stage0_36[336], stage0_36[337]},
      {stage0_38[210], stage0_38[211], stage0_38[212], stage0_38[213], stage0_38[214], stage0_38[215]},
      {stage1_40[35],stage1_39[60],stage1_38[112],stage1_37[124],stage1_36[176]}
   );
   gpc606_5 gpc1427 (
      {stage0_36[338], stage0_36[339], stage0_36[340], stage0_36[341], stage0_36[342], stage0_36[343]},
      {stage0_38[216], stage0_38[217], stage0_38[218], stage0_38[219], stage0_38[220], stage0_38[221]},
      {stage1_40[36],stage1_39[61],stage1_38[113],stage1_37[125],stage1_36[177]}
   );
   gpc606_5 gpc1428 (
      {stage0_36[344], stage0_36[345], stage0_36[346], stage0_36[347], stage0_36[348], stage0_36[349]},
      {stage0_38[222], stage0_38[223], stage0_38[224], stage0_38[225], stage0_38[226], stage0_38[227]},
      {stage1_40[37],stage1_39[62],stage1_38[114],stage1_37[126],stage1_36[178]}
   );
   gpc606_5 gpc1429 (
      {stage0_36[350], stage0_36[351], stage0_36[352], stage0_36[353], stage0_36[354], stage0_36[355]},
      {stage0_38[228], stage0_38[229], stage0_38[230], stage0_38[231], stage0_38[232], stage0_38[233]},
      {stage1_40[38],stage1_39[63],stage1_38[115],stage1_37[127],stage1_36[179]}
   );
   gpc606_5 gpc1430 (
      {stage0_36[356], stage0_36[357], stage0_36[358], stage0_36[359], stage0_36[360], stage0_36[361]},
      {stage0_38[234], stage0_38[235], stage0_38[236], stage0_38[237], stage0_38[238], stage0_38[239]},
      {stage1_40[39],stage1_39[64],stage1_38[116],stage1_37[128],stage1_36[180]}
   );
   gpc606_5 gpc1431 (
      {stage0_36[362], stage0_36[363], stage0_36[364], stage0_36[365], stage0_36[366], stage0_36[367]},
      {stage0_38[240], stage0_38[241], stage0_38[242], stage0_38[243], stage0_38[244], stage0_38[245]},
      {stage1_40[40],stage1_39[65],stage1_38[117],stage1_37[129],stage1_36[181]}
   );
   gpc606_5 gpc1432 (
      {stage0_36[368], stage0_36[369], stage0_36[370], stage0_36[371], stage0_36[372], stage0_36[373]},
      {stage0_38[246], stage0_38[247], stage0_38[248], stage0_38[249], stage0_38[250], stage0_38[251]},
      {stage1_40[41],stage1_39[66],stage1_38[118],stage1_37[130],stage1_36[182]}
   );
   gpc606_5 gpc1433 (
      {stage0_36[374], stage0_36[375], stage0_36[376], stage0_36[377], stage0_36[378], stage0_36[379]},
      {stage0_38[252], stage0_38[253], stage0_38[254], stage0_38[255], stage0_38[256], stage0_38[257]},
      {stage1_40[42],stage1_39[67],stage1_38[119],stage1_37[131],stage1_36[183]}
   );
   gpc606_5 gpc1434 (
      {stage0_36[380], stage0_36[381], stage0_36[382], stage0_36[383], stage0_36[384], stage0_36[385]},
      {stage0_38[258], stage0_38[259], stage0_38[260], stage0_38[261], stage0_38[262], stage0_38[263]},
      {stage1_40[43],stage1_39[68],stage1_38[120],stage1_37[132],stage1_36[184]}
   );
   gpc606_5 gpc1435 (
      {stage0_36[386], stage0_36[387], stage0_36[388], stage0_36[389], stage0_36[390], stage0_36[391]},
      {stage0_38[264], stage0_38[265], stage0_38[266], stage0_38[267], stage0_38[268], stage0_38[269]},
      {stage1_40[44],stage1_39[69],stage1_38[121],stage1_37[133],stage1_36[185]}
   );
   gpc606_5 gpc1436 (
      {stage0_36[392], stage0_36[393], stage0_36[394], stage0_36[395], stage0_36[396], stage0_36[397]},
      {stage0_38[270], stage0_38[271], stage0_38[272], stage0_38[273], stage0_38[274], stage0_38[275]},
      {stage1_40[45],stage1_39[70],stage1_38[122],stage1_37[134],stage1_36[186]}
   );
   gpc606_5 gpc1437 (
      {stage0_36[398], stage0_36[399], stage0_36[400], stage0_36[401], stage0_36[402], stage0_36[403]},
      {stage0_38[276], stage0_38[277], stage0_38[278], stage0_38[279], stage0_38[280], stage0_38[281]},
      {stage1_40[46],stage1_39[71],stage1_38[123],stage1_37[135],stage1_36[187]}
   );
   gpc606_5 gpc1438 (
      {stage0_36[404], stage0_36[405], stage0_36[406], stage0_36[407], stage0_36[408], stage0_36[409]},
      {stage0_38[282], stage0_38[283], stage0_38[284], stage0_38[285], stage0_38[286], stage0_38[287]},
      {stage1_40[47],stage1_39[72],stage1_38[124],stage1_37[136],stage1_36[188]}
   );
   gpc606_5 gpc1439 (
      {stage0_36[410], stage0_36[411], stage0_36[412], stage0_36[413], stage0_36[414], stage0_36[415]},
      {stage0_38[288], stage0_38[289], stage0_38[290], stage0_38[291], stage0_38[292], stage0_38[293]},
      {stage1_40[48],stage1_39[73],stage1_38[125],stage1_37[137],stage1_36[189]}
   );
   gpc606_5 gpc1440 (
      {stage0_36[416], stage0_36[417], stage0_36[418], stage0_36[419], stage0_36[420], stage0_36[421]},
      {stage0_38[294], stage0_38[295], stage0_38[296], stage0_38[297], stage0_38[298], stage0_38[299]},
      {stage1_40[49],stage1_39[74],stage1_38[126],stage1_37[138],stage1_36[190]}
   );
   gpc606_5 gpc1441 (
      {stage0_36[422], stage0_36[423], stage0_36[424], stage0_36[425], stage0_36[426], stage0_36[427]},
      {stage0_38[300], stage0_38[301], stage0_38[302], stage0_38[303], stage0_38[304], stage0_38[305]},
      {stage1_40[50],stage1_39[75],stage1_38[127],stage1_37[139],stage1_36[191]}
   );
   gpc606_5 gpc1442 (
      {stage0_36[428], stage0_36[429], stage0_36[430], stage0_36[431], stage0_36[432], stage0_36[433]},
      {stage0_38[306], stage0_38[307], stage0_38[308], stage0_38[309], stage0_38[310], stage0_38[311]},
      {stage1_40[51],stage1_39[76],stage1_38[128],stage1_37[140],stage1_36[192]}
   );
   gpc606_5 gpc1443 (
      {stage0_36[434], stage0_36[435], stage0_36[436], stage0_36[437], stage0_36[438], stage0_36[439]},
      {stage0_38[312], stage0_38[313], stage0_38[314], stage0_38[315], stage0_38[316], stage0_38[317]},
      {stage1_40[52],stage1_39[77],stage1_38[129],stage1_37[141],stage1_36[193]}
   );
   gpc606_5 gpc1444 (
      {stage0_36[440], stage0_36[441], stage0_36[442], stage0_36[443], stage0_36[444], stage0_36[445]},
      {stage0_38[318], stage0_38[319], stage0_38[320], stage0_38[321], stage0_38[322], stage0_38[323]},
      {stage1_40[53],stage1_39[78],stage1_38[130],stage1_37[142],stage1_36[194]}
   );
   gpc606_5 gpc1445 (
      {stage0_36[446], stage0_36[447], stage0_36[448], stage0_36[449], stage0_36[450], stage0_36[451]},
      {stage0_38[324], stage0_38[325], stage0_38[326], stage0_38[327], stage0_38[328], stage0_38[329]},
      {stage1_40[54],stage1_39[79],stage1_38[131],stage1_37[143],stage1_36[195]}
   );
   gpc606_5 gpc1446 (
      {stage0_36[452], stage0_36[453], stage0_36[454], stage0_36[455], stage0_36[456], stage0_36[457]},
      {stage0_38[330], stage0_38[331], stage0_38[332], stage0_38[333], stage0_38[334], stage0_38[335]},
      {stage1_40[55],stage1_39[80],stage1_38[132],stage1_37[144],stage1_36[196]}
   );
   gpc606_5 gpc1447 (
      {stage0_36[458], stage0_36[459], stage0_36[460], stage0_36[461], stage0_36[462], stage0_36[463]},
      {stage0_38[336], stage0_38[337], stage0_38[338], stage0_38[339], stage0_38[340], stage0_38[341]},
      {stage1_40[56],stage1_39[81],stage1_38[133],stage1_37[145],stage1_36[197]}
   );
   gpc606_5 gpc1448 (
      {stage0_36[464], stage0_36[465], stage0_36[466], stage0_36[467], stage0_36[468], stage0_36[469]},
      {stage0_38[342], stage0_38[343], stage0_38[344], stage0_38[345], stage0_38[346], stage0_38[347]},
      {stage1_40[57],stage1_39[82],stage1_38[134],stage1_37[146],stage1_36[198]}
   );
   gpc606_5 gpc1449 (
      {stage0_36[470], stage0_36[471], stage0_36[472], stage0_36[473], stage0_36[474], stage0_36[475]},
      {stage0_38[348], stage0_38[349], stage0_38[350], stage0_38[351], stage0_38[352], stage0_38[353]},
      {stage1_40[58],stage1_39[83],stage1_38[135],stage1_37[147],stage1_36[199]}
   );
   gpc606_5 gpc1450 (
      {stage0_36[476], stage0_36[477], stage0_36[478], stage0_36[479], stage0_36[480], stage0_36[481]},
      {stage0_38[354], stage0_38[355], stage0_38[356], stage0_38[357], stage0_38[358], stage0_38[359]},
      {stage1_40[59],stage1_39[84],stage1_38[136],stage1_37[148],stage1_36[200]}
   );
   gpc606_5 gpc1451 (
      {stage0_36[482], stage0_36[483], stage0_36[484], stage0_36[485], 1'b0, 1'b0},
      {stage0_38[360], stage0_38[361], stage0_38[362], stage0_38[363], stage0_38[364], stage0_38[365]},
      {stage1_40[60],stage1_39[85],stage1_38[137],stage1_37[149],stage1_36[201]}
   );
   gpc606_5 gpc1452 (
      {stage0_37[193], stage0_37[194], stage0_37[195], stage0_37[196], stage0_37[197], stage0_37[198]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[61],stage1_39[86],stage1_38[138],stage1_37[150]}
   );
   gpc606_5 gpc1453 (
      {stage0_37[199], stage0_37[200], stage0_37[201], stage0_37[202], stage0_37[203], stage0_37[204]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[62],stage1_39[87],stage1_38[139],stage1_37[151]}
   );
   gpc606_5 gpc1454 (
      {stage0_37[205], stage0_37[206], stage0_37[207], stage0_37[208], stage0_37[209], stage0_37[210]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[63],stage1_39[88],stage1_38[140],stage1_37[152]}
   );
   gpc606_5 gpc1455 (
      {stage0_37[211], stage0_37[212], stage0_37[213], stage0_37[214], stage0_37[215], stage0_37[216]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[64],stage1_39[89],stage1_38[141],stage1_37[153]}
   );
   gpc606_5 gpc1456 (
      {stage0_37[217], stage0_37[218], stage0_37[219], stage0_37[220], stage0_37[221], stage0_37[222]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[65],stage1_39[90],stage1_38[142],stage1_37[154]}
   );
   gpc606_5 gpc1457 (
      {stage0_37[223], stage0_37[224], stage0_37[225], stage0_37[226], stage0_37[227], stage0_37[228]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[66],stage1_39[91],stage1_38[143],stage1_37[155]}
   );
   gpc606_5 gpc1458 (
      {stage0_37[229], stage0_37[230], stage0_37[231], stage0_37[232], stage0_37[233], stage0_37[234]},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[67],stage1_39[92],stage1_38[144],stage1_37[156]}
   );
   gpc606_5 gpc1459 (
      {stage0_37[235], stage0_37[236], stage0_37[237], stage0_37[238], stage0_37[239], stage0_37[240]},
      {stage0_39[42], stage0_39[43], stage0_39[44], stage0_39[45], stage0_39[46], stage0_39[47]},
      {stage1_41[7],stage1_40[68],stage1_39[93],stage1_38[145],stage1_37[157]}
   );
   gpc606_5 gpc1460 (
      {stage0_37[241], stage0_37[242], stage0_37[243], stage0_37[244], stage0_37[245], stage0_37[246]},
      {stage0_39[48], stage0_39[49], stage0_39[50], stage0_39[51], stage0_39[52], stage0_39[53]},
      {stage1_41[8],stage1_40[69],stage1_39[94],stage1_38[146],stage1_37[158]}
   );
   gpc606_5 gpc1461 (
      {stage0_37[247], stage0_37[248], stage0_37[249], stage0_37[250], stage0_37[251], stage0_37[252]},
      {stage0_39[54], stage0_39[55], stage0_39[56], stage0_39[57], stage0_39[58], stage0_39[59]},
      {stage1_41[9],stage1_40[70],stage1_39[95],stage1_38[147],stage1_37[159]}
   );
   gpc606_5 gpc1462 (
      {stage0_37[253], stage0_37[254], stage0_37[255], stage0_37[256], stage0_37[257], stage0_37[258]},
      {stage0_39[60], stage0_39[61], stage0_39[62], stage0_39[63], stage0_39[64], stage0_39[65]},
      {stage1_41[10],stage1_40[71],stage1_39[96],stage1_38[148],stage1_37[160]}
   );
   gpc606_5 gpc1463 (
      {stage0_37[259], stage0_37[260], stage0_37[261], stage0_37[262], stage0_37[263], stage0_37[264]},
      {stage0_39[66], stage0_39[67], stage0_39[68], stage0_39[69], stage0_39[70], stage0_39[71]},
      {stage1_41[11],stage1_40[72],stage1_39[97],stage1_38[149],stage1_37[161]}
   );
   gpc606_5 gpc1464 (
      {stage0_37[265], stage0_37[266], stage0_37[267], stage0_37[268], stage0_37[269], stage0_37[270]},
      {stage0_39[72], stage0_39[73], stage0_39[74], stage0_39[75], stage0_39[76], stage0_39[77]},
      {stage1_41[12],stage1_40[73],stage1_39[98],stage1_38[150],stage1_37[162]}
   );
   gpc606_5 gpc1465 (
      {stage0_37[271], stage0_37[272], stage0_37[273], stage0_37[274], stage0_37[275], stage0_37[276]},
      {stage0_39[78], stage0_39[79], stage0_39[80], stage0_39[81], stage0_39[82], stage0_39[83]},
      {stage1_41[13],stage1_40[74],stage1_39[99],stage1_38[151],stage1_37[163]}
   );
   gpc606_5 gpc1466 (
      {stage0_37[277], stage0_37[278], stage0_37[279], stage0_37[280], stage0_37[281], stage0_37[282]},
      {stage0_39[84], stage0_39[85], stage0_39[86], stage0_39[87], stage0_39[88], stage0_39[89]},
      {stage1_41[14],stage1_40[75],stage1_39[100],stage1_38[152],stage1_37[164]}
   );
   gpc606_5 gpc1467 (
      {stage0_37[283], stage0_37[284], stage0_37[285], stage0_37[286], stage0_37[287], stage0_37[288]},
      {stage0_39[90], stage0_39[91], stage0_39[92], stage0_39[93], stage0_39[94], stage0_39[95]},
      {stage1_41[15],stage1_40[76],stage1_39[101],stage1_38[153],stage1_37[165]}
   );
   gpc606_5 gpc1468 (
      {stage0_37[289], stage0_37[290], stage0_37[291], stage0_37[292], stage0_37[293], stage0_37[294]},
      {stage0_39[96], stage0_39[97], stage0_39[98], stage0_39[99], stage0_39[100], stage0_39[101]},
      {stage1_41[16],stage1_40[77],stage1_39[102],stage1_38[154],stage1_37[166]}
   );
   gpc606_5 gpc1469 (
      {stage0_37[295], stage0_37[296], stage0_37[297], stage0_37[298], stage0_37[299], stage0_37[300]},
      {stage0_39[102], stage0_39[103], stage0_39[104], stage0_39[105], stage0_39[106], stage0_39[107]},
      {stage1_41[17],stage1_40[78],stage1_39[103],stage1_38[155],stage1_37[167]}
   );
   gpc606_5 gpc1470 (
      {stage0_37[301], stage0_37[302], stage0_37[303], stage0_37[304], stage0_37[305], stage0_37[306]},
      {stage0_39[108], stage0_39[109], stage0_39[110], stage0_39[111], stage0_39[112], stage0_39[113]},
      {stage1_41[18],stage1_40[79],stage1_39[104],stage1_38[156],stage1_37[168]}
   );
   gpc606_5 gpc1471 (
      {stage0_37[307], stage0_37[308], stage0_37[309], stage0_37[310], stage0_37[311], stage0_37[312]},
      {stage0_39[114], stage0_39[115], stage0_39[116], stage0_39[117], stage0_39[118], stage0_39[119]},
      {stage1_41[19],stage1_40[80],stage1_39[105],stage1_38[157],stage1_37[169]}
   );
   gpc606_5 gpc1472 (
      {stage0_37[313], stage0_37[314], stage0_37[315], stage0_37[316], stage0_37[317], stage0_37[318]},
      {stage0_39[120], stage0_39[121], stage0_39[122], stage0_39[123], stage0_39[124], stage0_39[125]},
      {stage1_41[20],stage1_40[81],stage1_39[106],stage1_38[158],stage1_37[170]}
   );
   gpc606_5 gpc1473 (
      {stage0_37[319], stage0_37[320], stage0_37[321], stage0_37[322], stage0_37[323], stage0_37[324]},
      {stage0_39[126], stage0_39[127], stage0_39[128], stage0_39[129], stage0_39[130], stage0_39[131]},
      {stage1_41[21],stage1_40[82],stage1_39[107],stage1_38[159],stage1_37[171]}
   );
   gpc606_5 gpc1474 (
      {stage0_37[325], stage0_37[326], stage0_37[327], stage0_37[328], stage0_37[329], stage0_37[330]},
      {stage0_39[132], stage0_39[133], stage0_39[134], stage0_39[135], stage0_39[136], stage0_39[137]},
      {stage1_41[22],stage1_40[83],stage1_39[108],stage1_38[160],stage1_37[172]}
   );
   gpc606_5 gpc1475 (
      {stage0_37[331], stage0_37[332], stage0_37[333], stage0_37[334], stage0_37[335], stage0_37[336]},
      {stage0_39[138], stage0_39[139], stage0_39[140], stage0_39[141], stage0_39[142], stage0_39[143]},
      {stage1_41[23],stage1_40[84],stage1_39[109],stage1_38[161],stage1_37[173]}
   );
   gpc606_5 gpc1476 (
      {stage0_37[337], stage0_37[338], stage0_37[339], stage0_37[340], stage0_37[341], stage0_37[342]},
      {stage0_39[144], stage0_39[145], stage0_39[146], stage0_39[147], stage0_39[148], stage0_39[149]},
      {stage1_41[24],stage1_40[85],stage1_39[110],stage1_38[162],stage1_37[174]}
   );
   gpc606_5 gpc1477 (
      {stage0_37[343], stage0_37[344], stage0_37[345], stage0_37[346], stage0_37[347], stage0_37[348]},
      {stage0_39[150], stage0_39[151], stage0_39[152], stage0_39[153], stage0_39[154], stage0_39[155]},
      {stage1_41[25],stage1_40[86],stage1_39[111],stage1_38[163],stage1_37[175]}
   );
   gpc606_5 gpc1478 (
      {stage0_37[349], stage0_37[350], stage0_37[351], stage0_37[352], stage0_37[353], stage0_37[354]},
      {stage0_39[156], stage0_39[157], stage0_39[158], stage0_39[159], stage0_39[160], stage0_39[161]},
      {stage1_41[26],stage1_40[87],stage1_39[112],stage1_38[164],stage1_37[176]}
   );
   gpc615_5 gpc1479 (
      {stage0_38[366], stage0_38[367], stage0_38[368], stage0_38[369], stage0_38[370]},
      {stage0_39[162]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[27],stage1_40[88],stage1_39[113],stage1_38[165]}
   );
   gpc615_5 gpc1480 (
      {stage0_38[371], stage0_38[372], stage0_38[373], stage0_38[374], stage0_38[375]},
      {stage0_39[163]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[28],stage1_40[89],stage1_39[114],stage1_38[166]}
   );
   gpc615_5 gpc1481 (
      {stage0_38[376], stage0_38[377], stage0_38[378], stage0_38[379], stage0_38[380]},
      {stage0_39[164]},
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage1_42[2],stage1_41[29],stage1_40[90],stage1_39[115],stage1_38[167]}
   );
   gpc615_5 gpc1482 (
      {stage0_38[381], stage0_38[382], stage0_38[383], stage0_38[384], stage0_38[385]},
      {stage0_39[165]},
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage1_42[3],stage1_41[30],stage1_40[91],stage1_39[116],stage1_38[168]}
   );
   gpc615_5 gpc1483 (
      {stage0_38[386], stage0_38[387], stage0_38[388], stage0_38[389], stage0_38[390]},
      {stage0_39[166]},
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage1_42[4],stage1_41[31],stage1_40[92],stage1_39[117],stage1_38[169]}
   );
   gpc615_5 gpc1484 (
      {stage0_39[167], stage0_39[168], stage0_39[169], stage0_39[170], stage0_39[171]},
      {stage0_40[30]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[5],stage1_41[32],stage1_40[93],stage1_39[118]}
   );
   gpc615_5 gpc1485 (
      {stage0_39[172], stage0_39[173], stage0_39[174], stage0_39[175], stage0_39[176]},
      {stage0_40[31]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[6],stage1_41[33],stage1_40[94],stage1_39[119]}
   );
   gpc615_5 gpc1486 (
      {stage0_39[177], stage0_39[178], stage0_39[179], stage0_39[180], stage0_39[181]},
      {stage0_40[32]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[7],stage1_41[34],stage1_40[95],stage1_39[120]}
   );
   gpc615_5 gpc1487 (
      {stage0_39[182], stage0_39[183], stage0_39[184], stage0_39[185], stage0_39[186]},
      {stage0_40[33]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[8],stage1_41[35],stage1_40[96],stage1_39[121]}
   );
   gpc615_5 gpc1488 (
      {stage0_39[187], stage0_39[188], stage0_39[189], stage0_39[190], stage0_39[191]},
      {stage0_40[34]},
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage1_43[4],stage1_42[9],stage1_41[36],stage1_40[97],stage1_39[122]}
   );
   gpc615_5 gpc1489 (
      {stage0_39[192], stage0_39[193], stage0_39[194], stage0_39[195], stage0_39[196]},
      {stage0_40[35]},
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage1_43[5],stage1_42[10],stage1_41[37],stage1_40[98],stage1_39[123]}
   );
   gpc615_5 gpc1490 (
      {stage0_39[197], stage0_39[198], stage0_39[199], stage0_39[200], stage0_39[201]},
      {stage0_40[36]},
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage1_43[6],stage1_42[11],stage1_41[38],stage1_40[99],stage1_39[124]}
   );
   gpc615_5 gpc1491 (
      {stage0_39[202], stage0_39[203], stage0_39[204], stage0_39[205], stage0_39[206]},
      {stage0_40[37]},
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage1_43[7],stage1_42[12],stage1_41[39],stage1_40[100],stage1_39[125]}
   );
   gpc615_5 gpc1492 (
      {stage0_39[207], stage0_39[208], stage0_39[209], stage0_39[210], stage0_39[211]},
      {stage0_40[38]},
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage1_43[8],stage1_42[13],stage1_41[40],stage1_40[101],stage1_39[126]}
   );
   gpc615_5 gpc1493 (
      {stage0_39[212], stage0_39[213], stage0_39[214], stage0_39[215], stage0_39[216]},
      {stage0_40[39]},
      {stage0_41[54], stage0_41[55], stage0_41[56], stage0_41[57], stage0_41[58], stage0_41[59]},
      {stage1_43[9],stage1_42[14],stage1_41[41],stage1_40[102],stage1_39[127]}
   );
   gpc615_5 gpc1494 (
      {stage0_39[217], stage0_39[218], stage0_39[219], stage0_39[220], stage0_39[221]},
      {stage0_40[40]},
      {stage0_41[60], stage0_41[61], stage0_41[62], stage0_41[63], stage0_41[64], stage0_41[65]},
      {stage1_43[10],stage1_42[15],stage1_41[42],stage1_40[103],stage1_39[128]}
   );
   gpc615_5 gpc1495 (
      {stage0_39[222], stage0_39[223], stage0_39[224], stage0_39[225], stage0_39[226]},
      {stage0_40[41]},
      {stage0_41[66], stage0_41[67], stage0_41[68], stage0_41[69], stage0_41[70], stage0_41[71]},
      {stage1_43[11],stage1_42[16],stage1_41[43],stage1_40[104],stage1_39[129]}
   );
   gpc615_5 gpc1496 (
      {stage0_39[227], stage0_39[228], stage0_39[229], stage0_39[230], stage0_39[231]},
      {stage0_40[42]},
      {stage0_41[72], stage0_41[73], stage0_41[74], stage0_41[75], stage0_41[76], stage0_41[77]},
      {stage1_43[12],stage1_42[17],stage1_41[44],stage1_40[105],stage1_39[130]}
   );
   gpc615_5 gpc1497 (
      {stage0_39[232], stage0_39[233], stage0_39[234], stage0_39[235], stage0_39[236]},
      {stage0_40[43]},
      {stage0_41[78], stage0_41[79], stage0_41[80], stage0_41[81], stage0_41[82], stage0_41[83]},
      {stage1_43[13],stage1_42[18],stage1_41[45],stage1_40[106],stage1_39[131]}
   );
   gpc615_5 gpc1498 (
      {stage0_39[237], stage0_39[238], stage0_39[239], stage0_39[240], stage0_39[241]},
      {stage0_40[44]},
      {stage0_41[84], stage0_41[85], stage0_41[86], stage0_41[87], stage0_41[88], stage0_41[89]},
      {stage1_43[14],stage1_42[19],stage1_41[46],stage1_40[107],stage1_39[132]}
   );
   gpc615_5 gpc1499 (
      {stage0_39[242], stage0_39[243], stage0_39[244], stage0_39[245], stage0_39[246]},
      {stage0_40[45]},
      {stage0_41[90], stage0_41[91], stage0_41[92], stage0_41[93], stage0_41[94], stage0_41[95]},
      {stage1_43[15],stage1_42[20],stage1_41[47],stage1_40[108],stage1_39[133]}
   );
   gpc615_5 gpc1500 (
      {stage0_39[247], stage0_39[248], stage0_39[249], stage0_39[250], stage0_39[251]},
      {stage0_40[46]},
      {stage0_41[96], stage0_41[97], stage0_41[98], stage0_41[99], stage0_41[100], stage0_41[101]},
      {stage1_43[16],stage1_42[21],stage1_41[48],stage1_40[109],stage1_39[134]}
   );
   gpc615_5 gpc1501 (
      {stage0_39[252], stage0_39[253], stage0_39[254], stage0_39[255], stage0_39[256]},
      {stage0_40[47]},
      {stage0_41[102], stage0_41[103], stage0_41[104], stage0_41[105], stage0_41[106], stage0_41[107]},
      {stage1_43[17],stage1_42[22],stage1_41[49],stage1_40[110],stage1_39[135]}
   );
   gpc615_5 gpc1502 (
      {stage0_39[257], stage0_39[258], stage0_39[259], stage0_39[260], stage0_39[261]},
      {stage0_40[48]},
      {stage0_41[108], stage0_41[109], stage0_41[110], stage0_41[111], stage0_41[112], stage0_41[113]},
      {stage1_43[18],stage1_42[23],stage1_41[50],stage1_40[111],stage1_39[136]}
   );
   gpc615_5 gpc1503 (
      {stage0_39[262], stage0_39[263], stage0_39[264], stage0_39[265], stage0_39[266]},
      {stage0_40[49]},
      {stage0_41[114], stage0_41[115], stage0_41[116], stage0_41[117], stage0_41[118], stage0_41[119]},
      {stage1_43[19],stage1_42[24],stage1_41[51],stage1_40[112],stage1_39[137]}
   );
   gpc615_5 gpc1504 (
      {stage0_39[267], stage0_39[268], stage0_39[269], stage0_39[270], stage0_39[271]},
      {stage0_40[50]},
      {stage0_41[120], stage0_41[121], stage0_41[122], stage0_41[123], stage0_41[124], stage0_41[125]},
      {stage1_43[20],stage1_42[25],stage1_41[52],stage1_40[113],stage1_39[138]}
   );
   gpc615_5 gpc1505 (
      {stage0_39[272], stage0_39[273], stage0_39[274], stage0_39[275], stage0_39[276]},
      {stage0_40[51]},
      {stage0_41[126], stage0_41[127], stage0_41[128], stage0_41[129], stage0_41[130], stage0_41[131]},
      {stage1_43[21],stage1_42[26],stage1_41[53],stage1_40[114],stage1_39[139]}
   );
   gpc615_5 gpc1506 (
      {stage0_39[277], stage0_39[278], stage0_39[279], stage0_39[280], stage0_39[281]},
      {stage0_40[52]},
      {stage0_41[132], stage0_41[133], stage0_41[134], stage0_41[135], stage0_41[136], stage0_41[137]},
      {stage1_43[22],stage1_42[27],stage1_41[54],stage1_40[115],stage1_39[140]}
   );
   gpc615_5 gpc1507 (
      {stage0_39[282], stage0_39[283], stage0_39[284], stage0_39[285], stage0_39[286]},
      {stage0_40[53]},
      {stage0_41[138], stage0_41[139], stage0_41[140], stage0_41[141], stage0_41[142], stage0_41[143]},
      {stage1_43[23],stage1_42[28],stage1_41[55],stage1_40[116],stage1_39[141]}
   );
   gpc615_5 gpc1508 (
      {stage0_39[287], stage0_39[288], stage0_39[289], stage0_39[290], stage0_39[291]},
      {stage0_40[54]},
      {stage0_41[144], stage0_41[145], stage0_41[146], stage0_41[147], stage0_41[148], stage0_41[149]},
      {stage1_43[24],stage1_42[29],stage1_41[56],stage1_40[117],stage1_39[142]}
   );
   gpc615_5 gpc1509 (
      {stage0_39[292], stage0_39[293], stage0_39[294], stage0_39[295], stage0_39[296]},
      {stage0_40[55]},
      {stage0_41[150], stage0_41[151], stage0_41[152], stage0_41[153], stage0_41[154], stage0_41[155]},
      {stage1_43[25],stage1_42[30],stage1_41[57],stage1_40[118],stage1_39[143]}
   );
   gpc615_5 gpc1510 (
      {stage0_39[297], stage0_39[298], stage0_39[299], stage0_39[300], stage0_39[301]},
      {stage0_40[56]},
      {stage0_41[156], stage0_41[157], stage0_41[158], stage0_41[159], stage0_41[160], stage0_41[161]},
      {stage1_43[26],stage1_42[31],stage1_41[58],stage1_40[119],stage1_39[144]}
   );
   gpc615_5 gpc1511 (
      {stage0_39[302], stage0_39[303], stage0_39[304], stage0_39[305], stage0_39[306]},
      {stage0_40[57]},
      {stage0_41[162], stage0_41[163], stage0_41[164], stage0_41[165], stage0_41[166], stage0_41[167]},
      {stage1_43[27],stage1_42[32],stage1_41[59],stage1_40[120],stage1_39[145]}
   );
   gpc615_5 gpc1512 (
      {stage0_39[307], stage0_39[308], stage0_39[309], stage0_39[310], stage0_39[311]},
      {stage0_40[58]},
      {stage0_41[168], stage0_41[169], stage0_41[170], stage0_41[171], stage0_41[172], stage0_41[173]},
      {stage1_43[28],stage1_42[33],stage1_41[60],stage1_40[121],stage1_39[146]}
   );
   gpc615_5 gpc1513 (
      {stage0_39[312], stage0_39[313], stage0_39[314], stage0_39[315], stage0_39[316]},
      {stage0_40[59]},
      {stage0_41[174], stage0_41[175], stage0_41[176], stage0_41[177], stage0_41[178], stage0_41[179]},
      {stage1_43[29],stage1_42[34],stage1_41[61],stage1_40[122],stage1_39[147]}
   );
   gpc615_5 gpc1514 (
      {stage0_39[317], stage0_39[318], stage0_39[319], stage0_39[320], stage0_39[321]},
      {stage0_40[60]},
      {stage0_41[180], stage0_41[181], stage0_41[182], stage0_41[183], stage0_41[184], stage0_41[185]},
      {stage1_43[30],stage1_42[35],stage1_41[62],stage1_40[123],stage1_39[148]}
   );
   gpc615_5 gpc1515 (
      {stage0_39[322], stage0_39[323], stage0_39[324], stage0_39[325], stage0_39[326]},
      {stage0_40[61]},
      {stage0_41[186], stage0_41[187], stage0_41[188], stage0_41[189], stage0_41[190], stage0_41[191]},
      {stage1_43[31],stage1_42[36],stage1_41[63],stage1_40[124],stage1_39[149]}
   );
   gpc615_5 gpc1516 (
      {stage0_39[327], stage0_39[328], stage0_39[329], stage0_39[330], stage0_39[331]},
      {stage0_40[62]},
      {stage0_41[192], stage0_41[193], stage0_41[194], stage0_41[195], stage0_41[196], stage0_41[197]},
      {stage1_43[32],stage1_42[37],stage1_41[64],stage1_40[125],stage1_39[150]}
   );
   gpc615_5 gpc1517 (
      {stage0_39[332], stage0_39[333], stage0_39[334], stage0_39[335], stage0_39[336]},
      {stage0_40[63]},
      {stage0_41[198], stage0_41[199], stage0_41[200], stage0_41[201], stage0_41[202], stage0_41[203]},
      {stage1_43[33],stage1_42[38],stage1_41[65],stage1_40[126],stage1_39[151]}
   );
   gpc615_5 gpc1518 (
      {stage0_39[337], stage0_39[338], stage0_39[339], stage0_39[340], stage0_39[341]},
      {stage0_40[64]},
      {stage0_41[204], stage0_41[205], stage0_41[206], stage0_41[207], stage0_41[208], stage0_41[209]},
      {stage1_43[34],stage1_42[39],stage1_41[66],stage1_40[127],stage1_39[152]}
   );
   gpc615_5 gpc1519 (
      {stage0_39[342], stage0_39[343], stage0_39[344], stage0_39[345], stage0_39[346]},
      {stage0_40[65]},
      {stage0_41[210], stage0_41[211], stage0_41[212], stage0_41[213], stage0_41[214], stage0_41[215]},
      {stage1_43[35],stage1_42[40],stage1_41[67],stage1_40[128],stage1_39[153]}
   );
   gpc615_5 gpc1520 (
      {stage0_39[347], stage0_39[348], stage0_39[349], stage0_39[350], stage0_39[351]},
      {stage0_40[66]},
      {stage0_41[216], stage0_41[217], stage0_41[218], stage0_41[219], stage0_41[220], stage0_41[221]},
      {stage1_43[36],stage1_42[41],stage1_41[68],stage1_40[129],stage1_39[154]}
   );
   gpc615_5 gpc1521 (
      {stage0_39[352], stage0_39[353], stage0_39[354], stage0_39[355], stage0_39[356]},
      {stage0_40[67]},
      {stage0_41[222], stage0_41[223], stage0_41[224], stage0_41[225], stage0_41[226], stage0_41[227]},
      {stage1_43[37],stage1_42[42],stage1_41[69],stage1_40[130],stage1_39[155]}
   );
   gpc615_5 gpc1522 (
      {stage0_39[357], stage0_39[358], stage0_39[359], stage0_39[360], stage0_39[361]},
      {stage0_40[68]},
      {stage0_41[228], stage0_41[229], stage0_41[230], stage0_41[231], stage0_41[232], stage0_41[233]},
      {stage1_43[38],stage1_42[43],stage1_41[70],stage1_40[131],stage1_39[156]}
   );
   gpc615_5 gpc1523 (
      {stage0_39[362], stage0_39[363], stage0_39[364], stage0_39[365], stage0_39[366]},
      {stage0_40[69]},
      {stage0_41[234], stage0_41[235], stage0_41[236], stage0_41[237], stage0_41[238], stage0_41[239]},
      {stage1_43[39],stage1_42[44],stage1_41[71],stage1_40[132],stage1_39[157]}
   );
   gpc615_5 gpc1524 (
      {stage0_39[367], stage0_39[368], stage0_39[369], stage0_39[370], stage0_39[371]},
      {stage0_40[70]},
      {stage0_41[240], stage0_41[241], stage0_41[242], stage0_41[243], stage0_41[244], stage0_41[245]},
      {stage1_43[40],stage1_42[45],stage1_41[72],stage1_40[133],stage1_39[158]}
   );
   gpc615_5 gpc1525 (
      {stage0_39[372], stage0_39[373], stage0_39[374], stage0_39[375], stage0_39[376]},
      {stage0_40[71]},
      {stage0_41[246], stage0_41[247], stage0_41[248], stage0_41[249], stage0_41[250], stage0_41[251]},
      {stage1_43[41],stage1_42[46],stage1_41[73],stage1_40[134],stage1_39[159]}
   );
   gpc615_5 gpc1526 (
      {stage0_39[377], stage0_39[378], stage0_39[379], stage0_39[380], stage0_39[381]},
      {stage0_40[72]},
      {stage0_41[252], stage0_41[253], stage0_41[254], stage0_41[255], stage0_41[256], stage0_41[257]},
      {stage1_43[42],stage1_42[47],stage1_41[74],stage1_40[135],stage1_39[160]}
   );
   gpc615_5 gpc1527 (
      {stage0_39[382], stage0_39[383], stage0_39[384], stage0_39[385], stage0_39[386]},
      {stage0_40[73]},
      {stage0_41[258], stage0_41[259], stage0_41[260], stage0_41[261], stage0_41[262], stage0_41[263]},
      {stage1_43[43],stage1_42[48],stage1_41[75],stage1_40[136],stage1_39[161]}
   );
   gpc615_5 gpc1528 (
      {stage0_39[387], stage0_39[388], stage0_39[389], stage0_39[390], stage0_39[391]},
      {stage0_40[74]},
      {stage0_41[264], stage0_41[265], stage0_41[266], stage0_41[267], stage0_41[268], stage0_41[269]},
      {stage1_43[44],stage1_42[49],stage1_41[76],stage1_40[137],stage1_39[162]}
   );
   gpc615_5 gpc1529 (
      {stage0_39[392], stage0_39[393], stage0_39[394], stage0_39[395], stage0_39[396]},
      {stage0_40[75]},
      {stage0_41[270], stage0_41[271], stage0_41[272], stage0_41[273], stage0_41[274], stage0_41[275]},
      {stage1_43[45],stage1_42[50],stage1_41[77],stage1_40[138],stage1_39[163]}
   );
   gpc615_5 gpc1530 (
      {stage0_39[397], stage0_39[398], stage0_39[399], stage0_39[400], stage0_39[401]},
      {stage0_40[76]},
      {stage0_41[276], stage0_41[277], stage0_41[278], stage0_41[279], stage0_41[280], stage0_41[281]},
      {stage1_43[46],stage1_42[51],stage1_41[78],stage1_40[139],stage1_39[164]}
   );
   gpc615_5 gpc1531 (
      {stage0_39[402], stage0_39[403], stage0_39[404], stage0_39[405], stage0_39[406]},
      {stage0_40[77]},
      {stage0_41[282], stage0_41[283], stage0_41[284], stage0_41[285], stage0_41[286], stage0_41[287]},
      {stage1_43[47],stage1_42[52],stage1_41[79],stage1_40[140],stage1_39[165]}
   );
   gpc615_5 gpc1532 (
      {stage0_39[407], stage0_39[408], stage0_39[409], stage0_39[410], stage0_39[411]},
      {stage0_40[78]},
      {stage0_41[288], stage0_41[289], stage0_41[290], stage0_41[291], stage0_41[292], stage0_41[293]},
      {stage1_43[48],stage1_42[53],stage1_41[80],stage1_40[141],stage1_39[166]}
   );
   gpc615_5 gpc1533 (
      {stage0_39[412], stage0_39[413], stage0_39[414], stage0_39[415], stage0_39[416]},
      {stage0_40[79]},
      {stage0_41[294], stage0_41[295], stage0_41[296], stage0_41[297], stage0_41[298], stage0_41[299]},
      {stage1_43[49],stage1_42[54],stage1_41[81],stage1_40[142],stage1_39[167]}
   );
   gpc615_5 gpc1534 (
      {stage0_39[417], stage0_39[418], stage0_39[419], stage0_39[420], stage0_39[421]},
      {stage0_40[80]},
      {stage0_41[300], stage0_41[301], stage0_41[302], stage0_41[303], stage0_41[304], stage0_41[305]},
      {stage1_43[50],stage1_42[55],stage1_41[82],stage1_40[143],stage1_39[168]}
   );
   gpc615_5 gpc1535 (
      {stage0_39[422], stage0_39[423], stage0_39[424], stage0_39[425], stage0_39[426]},
      {stage0_40[81]},
      {stage0_41[306], stage0_41[307], stage0_41[308], stage0_41[309], stage0_41[310], stage0_41[311]},
      {stage1_43[51],stage1_42[56],stage1_41[83],stage1_40[144],stage1_39[169]}
   );
   gpc615_5 gpc1536 (
      {stage0_39[427], stage0_39[428], stage0_39[429], stage0_39[430], stage0_39[431]},
      {stage0_40[82]},
      {stage0_41[312], stage0_41[313], stage0_41[314], stage0_41[315], stage0_41[316], stage0_41[317]},
      {stage1_43[52],stage1_42[57],stage1_41[84],stage1_40[145],stage1_39[170]}
   );
   gpc615_5 gpc1537 (
      {stage0_39[432], stage0_39[433], stage0_39[434], stage0_39[435], stage0_39[436]},
      {stage0_40[83]},
      {stage0_41[318], stage0_41[319], stage0_41[320], stage0_41[321], stage0_41[322], stage0_41[323]},
      {stage1_43[53],stage1_42[58],stage1_41[85],stage1_40[146],stage1_39[171]}
   );
   gpc615_5 gpc1538 (
      {stage0_39[437], stage0_39[438], stage0_39[439], stage0_39[440], stage0_39[441]},
      {stage0_40[84]},
      {stage0_41[324], stage0_41[325], stage0_41[326], stage0_41[327], stage0_41[328], stage0_41[329]},
      {stage1_43[54],stage1_42[59],stage1_41[86],stage1_40[147],stage1_39[172]}
   );
   gpc615_5 gpc1539 (
      {stage0_39[442], stage0_39[443], stage0_39[444], stage0_39[445], stage0_39[446]},
      {stage0_40[85]},
      {stage0_41[330], stage0_41[331], stage0_41[332], stage0_41[333], stage0_41[334], stage0_41[335]},
      {stage1_43[55],stage1_42[60],stage1_41[87],stage1_40[148],stage1_39[173]}
   );
   gpc606_5 gpc1540 (
      {stage0_40[86], stage0_40[87], stage0_40[88], stage0_40[89], stage0_40[90], stage0_40[91]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[56],stage1_42[61],stage1_41[88],stage1_40[149]}
   );
   gpc606_5 gpc1541 (
      {stage0_40[92], stage0_40[93], stage0_40[94], stage0_40[95], stage0_40[96], stage0_40[97]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[57],stage1_42[62],stage1_41[89],stage1_40[150]}
   );
   gpc606_5 gpc1542 (
      {stage0_40[98], stage0_40[99], stage0_40[100], stage0_40[101], stage0_40[102], stage0_40[103]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[58],stage1_42[63],stage1_41[90],stage1_40[151]}
   );
   gpc606_5 gpc1543 (
      {stage0_40[104], stage0_40[105], stage0_40[106], stage0_40[107], stage0_40[108], stage0_40[109]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[59],stage1_42[64],stage1_41[91],stage1_40[152]}
   );
   gpc606_5 gpc1544 (
      {stage0_40[110], stage0_40[111], stage0_40[112], stage0_40[113], stage0_40[114], stage0_40[115]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[60],stage1_42[65],stage1_41[92],stage1_40[153]}
   );
   gpc606_5 gpc1545 (
      {stage0_40[116], stage0_40[117], stage0_40[118], stage0_40[119], stage0_40[120], stage0_40[121]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[61],stage1_42[66],stage1_41[93],stage1_40[154]}
   );
   gpc606_5 gpc1546 (
      {stage0_40[122], stage0_40[123], stage0_40[124], stage0_40[125], stage0_40[126], stage0_40[127]},
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage1_44[6],stage1_43[62],stage1_42[67],stage1_41[94],stage1_40[155]}
   );
   gpc606_5 gpc1547 (
      {stage0_40[128], stage0_40[129], stage0_40[130], stage0_40[131], stage0_40[132], stage0_40[133]},
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage1_44[7],stage1_43[63],stage1_42[68],stage1_41[95],stage1_40[156]}
   );
   gpc606_5 gpc1548 (
      {stage0_40[134], stage0_40[135], stage0_40[136], stage0_40[137], stage0_40[138], stage0_40[139]},
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage1_44[8],stage1_43[64],stage1_42[69],stage1_41[96],stage1_40[157]}
   );
   gpc606_5 gpc1549 (
      {stage0_40[140], stage0_40[141], stage0_40[142], stage0_40[143], stage0_40[144], stage0_40[145]},
      {stage0_42[54], stage0_42[55], stage0_42[56], stage0_42[57], stage0_42[58], stage0_42[59]},
      {stage1_44[9],stage1_43[65],stage1_42[70],stage1_41[97],stage1_40[158]}
   );
   gpc606_5 gpc1550 (
      {stage0_40[146], stage0_40[147], stage0_40[148], stage0_40[149], stage0_40[150], stage0_40[151]},
      {stage0_42[60], stage0_42[61], stage0_42[62], stage0_42[63], stage0_42[64], stage0_42[65]},
      {stage1_44[10],stage1_43[66],stage1_42[71],stage1_41[98],stage1_40[159]}
   );
   gpc606_5 gpc1551 (
      {stage0_40[152], stage0_40[153], stage0_40[154], stage0_40[155], stage0_40[156], stage0_40[157]},
      {stage0_42[66], stage0_42[67], stage0_42[68], stage0_42[69], stage0_42[70], stage0_42[71]},
      {stage1_44[11],stage1_43[67],stage1_42[72],stage1_41[99],stage1_40[160]}
   );
   gpc606_5 gpc1552 (
      {stage0_40[158], stage0_40[159], stage0_40[160], stage0_40[161], stage0_40[162], stage0_40[163]},
      {stage0_42[72], stage0_42[73], stage0_42[74], stage0_42[75], stage0_42[76], stage0_42[77]},
      {stage1_44[12],stage1_43[68],stage1_42[73],stage1_41[100],stage1_40[161]}
   );
   gpc606_5 gpc1553 (
      {stage0_40[164], stage0_40[165], stage0_40[166], stage0_40[167], stage0_40[168], stage0_40[169]},
      {stage0_42[78], stage0_42[79], stage0_42[80], stage0_42[81], stage0_42[82], stage0_42[83]},
      {stage1_44[13],stage1_43[69],stage1_42[74],stage1_41[101],stage1_40[162]}
   );
   gpc606_5 gpc1554 (
      {stage0_40[170], stage0_40[171], stage0_40[172], stage0_40[173], stage0_40[174], stage0_40[175]},
      {stage0_42[84], stage0_42[85], stage0_42[86], stage0_42[87], stage0_42[88], stage0_42[89]},
      {stage1_44[14],stage1_43[70],stage1_42[75],stage1_41[102],stage1_40[163]}
   );
   gpc606_5 gpc1555 (
      {stage0_40[176], stage0_40[177], stage0_40[178], stage0_40[179], stage0_40[180], stage0_40[181]},
      {stage0_42[90], stage0_42[91], stage0_42[92], stage0_42[93], stage0_42[94], stage0_42[95]},
      {stage1_44[15],stage1_43[71],stage1_42[76],stage1_41[103],stage1_40[164]}
   );
   gpc606_5 gpc1556 (
      {stage0_40[182], stage0_40[183], stage0_40[184], stage0_40[185], stage0_40[186], stage0_40[187]},
      {stage0_42[96], stage0_42[97], stage0_42[98], stage0_42[99], stage0_42[100], stage0_42[101]},
      {stage1_44[16],stage1_43[72],stage1_42[77],stage1_41[104],stage1_40[165]}
   );
   gpc606_5 gpc1557 (
      {stage0_40[188], stage0_40[189], stage0_40[190], stage0_40[191], stage0_40[192], stage0_40[193]},
      {stage0_42[102], stage0_42[103], stage0_42[104], stage0_42[105], stage0_42[106], stage0_42[107]},
      {stage1_44[17],stage1_43[73],stage1_42[78],stage1_41[105],stage1_40[166]}
   );
   gpc606_5 gpc1558 (
      {stage0_40[194], stage0_40[195], stage0_40[196], stage0_40[197], stage0_40[198], stage0_40[199]},
      {stage0_42[108], stage0_42[109], stage0_42[110], stage0_42[111], stage0_42[112], stage0_42[113]},
      {stage1_44[18],stage1_43[74],stage1_42[79],stage1_41[106],stage1_40[167]}
   );
   gpc606_5 gpc1559 (
      {stage0_40[200], stage0_40[201], stage0_40[202], stage0_40[203], stage0_40[204], stage0_40[205]},
      {stage0_42[114], stage0_42[115], stage0_42[116], stage0_42[117], stage0_42[118], stage0_42[119]},
      {stage1_44[19],stage1_43[75],stage1_42[80],stage1_41[107],stage1_40[168]}
   );
   gpc606_5 gpc1560 (
      {stage0_40[206], stage0_40[207], stage0_40[208], stage0_40[209], stage0_40[210], stage0_40[211]},
      {stage0_42[120], stage0_42[121], stage0_42[122], stage0_42[123], stage0_42[124], stage0_42[125]},
      {stage1_44[20],stage1_43[76],stage1_42[81],stage1_41[108],stage1_40[169]}
   );
   gpc606_5 gpc1561 (
      {stage0_40[212], stage0_40[213], stage0_40[214], stage0_40[215], stage0_40[216], stage0_40[217]},
      {stage0_42[126], stage0_42[127], stage0_42[128], stage0_42[129], stage0_42[130], stage0_42[131]},
      {stage1_44[21],stage1_43[77],stage1_42[82],stage1_41[109],stage1_40[170]}
   );
   gpc606_5 gpc1562 (
      {stage0_40[218], stage0_40[219], stage0_40[220], stage0_40[221], stage0_40[222], stage0_40[223]},
      {stage0_42[132], stage0_42[133], stage0_42[134], stage0_42[135], stage0_42[136], stage0_42[137]},
      {stage1_44[22],stage1_43[78],stage1_42[83],stage1_41[110],stage1_40[171]}
   );
   gpc606_5 gpc1563 (
      {stage0_40[224], stage0_40[225], stage0_40[226], stage0_40[227], stage0_40[228], stage0_40[229]},
      {stage0_42[138], stage0_42[139], stage0_42[140], stage0_42[141], stage0_42[142], stage0_42[143]},
      {stage1_44[23],stage1_43[79],stage1_42[84],stage1_41[111],stage1_40[172]}
   );
   gpc606_5 gpc1564 (
      {stage0_40[230], stage0_40[231], stage0_40[232], stage0_40[233], stage0_40[234], stage0_40[235]},
      {stage0_42[144], stage0_42[145], stage0_42[146], stage0_42[147], stage0_42[148], stage0_42[149]},
      {stage1_44[24],stage1_43[80],stage1_42[85],stage1_41[112],stage1_40[173]}
   );
   gpc606_5 gpc1565 (
      {stage0_40[236], stage0_40[237], stage0_40[238], stage0_40[239], stage0_40[240], stage0_40[241]},
      {stage0_42[150], stage0_42[151], stage0_42[152], stage0_42[153], stage0_42[154], stage0_42[155]},
      {stage1_44[25],stage1_43[81],stage1_42[86],stage1_41[113],stage1_40[174]}
   );
   gpc606_5 gpc1566 (
      {stage0_40[242], stage0_40[243], stage0_40[244], stage0_40[245], stage0_40[246], stage0_40[247]},
      {stage0_42[156], stage0_42[157], stage0_42[158], stage0_42[159], stage0_42[160], stage0_42[161]},
      {stage1_44[26],stage1_43[82],stage1_42[87],stage1_41[114],stage1_40[175]}
   );
   gpc606_5 gpc1567 (
      {stage0_40[248], stage0_40[249], stage0_40[250], stage0_40[251], stage0_40[252], stage0_40[253]},
      {stage0_42[162], stage0_42[163], stage0_42[164], stage0_42[165], stage0_42[166], stage0_42[167]},
      {stage1_44[27],stage1_43[83],stage1_42[88],stage1_41[115],stage1_40[176]}
   );
   gpc606_5 gpc1568 (
      {stage0_40[254], stage0_40[255], stage0_40[256], stage0_40[257], stage0_40[258], stage0_40[259]},
      {stage0_42[168], stage0_42[169], stage0_42[170], stage0_42[171], stage0_42[172], stage0_42[173]},
      {stage1_44[28],stage1_43[84],stage1_42[89],stage1_41[116],stage1_40[177]}
   );
   gpc606_5 gpc1569 (
      {stage0_40[260], stage0_40[261], stage0_40[262], stage0_40[263], stage0_40[264], stage0_40[265]},
      {stage0_42[174], stage0_42[175], stage0_42[176], stage0_42[177], stage0_42[178], stage0_42[179]},
      {stage1_44[29],stage1_43[85],stage1_42[90],stage1_41[117],stage1_40[178]}
   );
   gpc606_5 gpc1570 (
      {stage0_40[266], stage0_40[267], stage0_40[268], stage0_40[269], stage0_40[270], stage0_40[271]},
      {stage0_42[180], stage0_42[181], stage0_42[182], stage0_42[183], stage0_42[184], stage0_42[185]},
      {stage1_44[30],stage1_43[86],stage1_42[91],stage1_41[118],stage1_40[179]}
   );
   gpc606_5 gpc1571 (
      {stage0_40[272], stage0_40[273], stage0_40[274], stage0_40[275], stage0_40[276], stage0_40[277]},
      {stage0_42[186], stage0_42[187], stage0_42[188], stage0_42[189], stage0_42[190], stage0_42[191]},
      {stage1_44[31],stage1_43[87],stage1_42[92],stage1_41[119],stage1_40[180]}
   );
   gpc606_5 gpc1572 (
      {stage0_40[278], stage0_40[279], stage0_40[280], stage0_40[281], stage0_40[282], stage0_40[283]},
      {stage0_42[192], stage0_42[193], stage0_42[194], stage0_42[195], stage0_42[196], stage0_42[197]},
      {stage1_44[32],stage1_43[88],stage1_42[93],stage1_41[120],stage1_40[181]}
   );
   gpc606_5 gpc1573 (
      {stage0_40[284], stage0_40[285], stage0_40[286], stage0_40[287], stage0_40[288], stage0_40[289]},
      {stage0_42[198], stage0_42[199], stage0_42[200], stage0_42[201], stage0_42[202], stage0_42[203]},
      {stage1_44[33],stage1_43[89],stage1_42[94],stage1_41[121],stage1_40[182]}
   );
   gpc606_5 gpc1574 (
      {stage0_40[290], stage0_40[291], stage0_40[292], stage0_40[293], stage0_40[294], stage0_40[295]},
      {stage0_42[204], stage0_42[205], stage0_42[206], stage0_42[207], stage0_42[208], stage0_42[209]},
      {stage1_44[34],stage1_43[90],stage1_42[95],stage1_41[122],stage1_40[183]}
   );
   gpc606_5 gpc1575 (
      {stage0_40[296], stage0_40[297], stage0_40[298], stage0_40[299], stage0_40[300], stage0_40[301]},
      {stage0_42[210], stage0_42[211], stage0_42[212], stage0_42[213], stage0_42[214], stage0_42[215]},
      {stage1_44[35],stage1_43[91],stage1_42[96],stage1_41[123],stage1_40[184]}
   );
   gpc606_5 gpc1576 (
      {stage0_40[302], stage0_40[303], stage0_40[304], stage0_40[305], stage0_40[306], stage0_40[307]},
      {stage0_42[216], stage0_42[217], stage0_42[218], stage0_42[219], stage0_42[220], stage0_42[221]},
      {stage1_44[36],stage1_43[92],stage1_42[97],stage1_41[124],stage1_40[185]}
   );
   gpc606_5 gpc1577 (
      {stage0_40[308], stage0_40[309], stage0_40[310], stage0_40[311], stage0_40[312], stage0_40[313]},
      {stage0_42[222], stage0_42[223], stage0_42[224], stage0_42[225], stage0_42[226], stage0_42[227]},
      {stage1_44[37],stage1_43[93],stage1_42[98],stage1_41[125],stage1_40[186]}
   );
   gpc606_5 gpc1578 (
      {stage0_40[314], stage0_40[315], stage0_40[316], stage0_40[317], stage0_40[318], stage0_40[319]},
      {stage0_42[228], stage0_42[229], stage0_42[230], stage0_42[231], stage0_42[232], stage0_42[233]},
      {stage1_44[38],stage1_43[94],stage1_42[99],stage1_41[126],stage1_40[187]}
   );
   gpc606_5 gpc1579 (
      {stage0_40[320], stage0_40[321], stage0_40[322], stage0_40[323], stage0_40[324], stage0_40[325]},
      {stage0_42[234], stage0_42[235], stage0_42[236], stage0_42[237], stage0_42[238], stage0_42[239]},
      {stage1_44[39],stage1_43[95],stage1_42[100],stage1_41[127],stage1_40[188]}
   );
   gpc606_5 gpc1580 (
      {stage0_40[326], stage0_40[327], stage0_40[328], stage0_40[329], stage0_40[330], stage0_40[331]},
      {stage0_42[240], stage0_42[241], stage0_42[242], stage0_42[243], stage0_42[244], stage0_42[245]},
      {stage1_44[40],stage1_43[96],stage1_42[101],stage1_41[128],stage1_40[189]}
   );
   gpc606_5 gpc1581 (
      {stage0_40[332], stage0_40[333], stage0_40[334], stage0_40[335], stage0_40[336], stage0_40[337]},
      {stage0_42[246], stage0_42[247], stage0_42[248], stage0_42[249], stage0_42[250], stage0_42[251]},
      {stage1_44[41],stage1_43[97],stage1_42[102],stage1_41[129],stage1_40[190]}
   );
   gpc606_5 gpc1582 (
      {stage0_40[338], stage0_40[339], stage0_40[340], stage0_40[341], stage0_40[342], stage0_40[343]},
      {stage0_42[252], stage0_42[253], stage0_42[254], stage0_42[255], stage0_42[256], stage0_42[257]},
      {stage1_44[42],stage1_43[98],stage1_42[103],stage1_41[130],stage1_40[191]}
   );
   gpc606_5 gpc1583 (
      {stage0_40[344], stage0_40[345], stage0_40[346], stage0_40[347], stage0_40[348], stage0_40[349]},
      {stage0_42[258], stage0_42[259], stage0_42[260], stage0_42[261], stage0_42[262], stage0_42[263]},
      {stage1_44[43],stage1_43[99],stage1_42[104],stage1_41[131],stage1_40[192]}
   );
   gpc606_5 gpc1584 (
      {stage0_40[350], stage0_40[351], stage0_40[352], stage0_40[353], stage0_40[354], stage0_40[355]},
      {stage0_42[264], stage0_42[265], stage0_42[266], stage0_42[267], stage0_42[268], stage0_42[269]},
      {stage1_44[44],stage1_43[100],stage1_42[105],stage1_41[132],stage1_40[193]}
   );
   gpc606_5 gpc1585 (
      {stage0_40[356], stage0_40[357], stage0_40[358], stage0_40[359], stage0_40[360], stage0_40[361]},
      {stage0_42[270], stage0_42[271], stage0_42[272], stage0_42[273], stage0_42[274], stage0_42[275]},
      {stage1_44[45],stage1_43[101],stage1_42[106],stage1_41[133],stage1_40[194]}
   );
   gpc606_5 gpc1586 (
      {stage0_40[362], stage0_40[363], stage0_40[364], stage0_40[365], stage0_40[366], stage0_40[367]},
      {stage0_42[276], stage0_42[277], stage0_42[278], stage0_42[279], stage0_42[280], stage0_42[281]},
      {stage1_44[46],stage1_43[102],stage1_42[107],stage1_41[134],stage1_40[195]}
   );
   gpc606_5 gpc1587 (
      {stage0_40[368], stage0_40[369], stage0_40[370], stage0_40[371], stage0_40[372], stage0_40[373]},
      {stage0_42[282], stage0_42[283], stage0_42[284], stage0_42[285], stage0_42[286], stage0_42[287]},
      {stage1_44[47],stage1_43[103],stage1_42[108],stage1_41[135],stage1_40[196]}
   );
   gpc606_5 gpc1588 (
      {stage0_40[374], stage0_40[375], stage0_40[376], stage0_40[377], stage0_40[378], stage0_40[379]},
      {stage0_42[288], stage0_42[289], stage0_42[290], stage0_42[291], stage0_42[292], stage0_42[293]},
      {stage1_44[48],stage1_43[104],stage1_42[109],stage1_41[136],stage1_40[197]}
   );
   gpc606_5 gpc1589 (
      {stage0_41[336], stage0_41[337], stage0_41[338], stage0_41[339], stage0_41[340], stage0_41[341]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[49],stage1_43[105],stage1_42[110],stage1_41[137]}
   );
   gpc606_5 gpc1590 (
      {stage0_41[342], stage0_41[343], stage0_41[344], stage0_41[345], stage0_41[346], stage0_41[347]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[50],stage1_43[106],stage1_42[111],stage1_41[138]}
   );
   gpc606_5 gpc1591 (
      {stage0_41[348], stage0_41[349], stage0_41[350], stage0_41[351], stage0_41[352], stage0_41[353]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[51],stage1_43[107],stage1_42[112],stage1_41[139]}
   );
   gpc606_5 gpc1592 (
      {stage0_41[354], stage0_41[355], stage0_41[356], stage0_41[357], stage0_41[358], stage0_41[359]},
      {stage0_43[18], stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23]},
      {stage1_45[3],stage1_44[52],stage1_43[108],stage1_42[113],stage1_41[140]}
   );
   gpc606_5 gpc1593 (
      {stage0_41[360], stage0_41[361], stage0_41[362], stage0_41[363], stage0_41[364], stage0_41[365]},
      {stage0_43[24], stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage1_45[4],stage1_44[53],stage1_43[109],stage1_42[114],stage1_41[141]}
   );
   gpc606_5 gpc1594 (
      {stage0_41[366], stage0_41[367], stage0_41[368], stage0_41[369], stage0_41[370], stage0_41[371]},
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34], stage0_43[35]},
      {stage1_45[5],stage1_44[54],stage1_43[110],stage1_42[115],stage1_41[142]}
   );
   gpc606_5 gpc1595 (
      {stage0_41[372], stage0_41[373], stage0_41[374], stage0_41[375], stage0_41[376], stage0_41[377]},
      {stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39], stage0_43[40], stage0_43[41]},
      {stage1_45[6],stage1_44[55],stage1_43[111],stage1_42[116],stage1_41[143]}
   );
   gpc606_5 gpc1596 (
      {stage0_41[378], stage0_41[379], stage0_41[380], stage0_41[381], stage0_41[382], stage0_41[383]},
      {stage0_43[42], stage0_43[43], stage0_43[44], stage0_43[45], stage0_43[46], stage0_43[47]},
      {stage1_45[7],stage1_44[56],stage1_43[112],stage1_42[117],stage1_41[144]}
   );
   gpc606_5 gpc1597 (
      {stage0_41[384], stage0_41[385], stage0_41[386], stage0_41[387], stage0_41[388], stage0_41[389]},
      {stage0_43[48], stage0_43[49], stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53]},
      {stage1_45[8],stage1_44[57],stage1_43[113],stage1_42[118],stage1_41[145]}
   );
   gpc606_5 gpc1598 (
      {stage0_41[390], stage0_41[391], stage0_41[392], stage0_41[393], stage0_41[394], stage0_41[395]},
      {stage0_43[54], stage0_43[55], stage0_43[56], stage0_43[57], stage0_43[58], stage0_43[59]},
      {stage1_45[9],stage1_44[58],stage1_43[114],stage1_42[119],stage1_41[146]}
   );
   gpc606_5 gpc1599 (
      {stage0_41[396], stage0_41[397], stage0_41[398], stage0_41[399], stage0_41[400], stage0_41[401]},
      {stage0_43[60], stage0_43[61], stage0_43[62], stage0_43[63], stage0_43[64], stage0_43[65]},
      {stage1_45[10],stage1_44[59],stage1_43[115],stage1_42[120],stage1_41[147]}
   );
   gpc606_5 gpc1600 (
      {stage0_41[402], stage0_41[403], stage0_41[404], stage0_41[405], stage0_41[406], stage0_41[407]},
      {stage0_43[66], stage0_43[67], stage0_43[68], stage0_43[69], stage0_43[70], stage0_43[71]},
      {stage1_45[11],stage1_44[60],stage1_43[116],stage1_42[121],stage1_41[148]}
   );
   gpc606_5 gpc1601 (
      {stage0_41[408], stage0_41[409], stage0_41[410], stage0_41[411], stage0_41[412], stage0_41[413]},
      {stage0_43[72], stage0_43[73], stage0_43[74], stage0_43[75], stage0_43[76], stage0_43[77]},
      {stage1_45[12],stage1_44[61],stage1_43[117],stage1_42[122],stage1_41[149]}
   );
   gpc606_5 gpc1602 (
      {stage0_41[414], stage0_41[415], stage0_41[416], stage0_41[417], stage0_41[418], stage0_41[419]},
      {stage0_43[78], stage0_43[79], stage0_43[80], stage0_43[81], stage0_43[82], stage0_43[83]},
      {stage1_45[13],stage1_44[62],stage1_43[118],stage1_42[123],stage1_41[150]}
   );
   gpc606_5 gpc1603 (
      {stage0_41[420], stage0_41[421], stage0_41[422], stage0_41[423], stage0_41[424], stage0_41[425]},
      {stage0_43[84], stage0_43[85], stage0_43[86], stage0_43[87], stage0_43[88], stage0_43[89]},
      {stage1_45[14],stage1_44[63],stage1_43[119],stage1_42[124],stage1_41[151]}
   );
   gpc606_5 gpc1604 (
      {stage0_41[426], stage0_41[427], stage0_41[428], stage0_41[429], stage0_41[430], stage0_41[431]},
      {stage0_43[90], stage0_43[91], stage0_43[92], stage0_43[93], stage0_43[94], stage0_43[95]},
      {stage1_45[15],stage1_44[64],stage1_43[120],stage1_42[125],stage1_41[152]}
   );
   gpc615_5 gpc1605 (
      {stage0_41[432], stage0_41[433], stage0_41[434], stage0_41[435], stage0_41[436]},
      {stage0_42[294]},
      {stage0_43[96], stage0_43[97], stage0_43[98], stage0_43[99], stage0_43[100], stage0_43[101]},
      {stage1_45[16],stage1_44[65],stage1_43[121],stage1_42[126],stage1_41[153]}
   );
   gpc615_5 gpc1606 (
      {stage0_41[437], stage0_41[438], stage0_41[439], stage0_41[440], stage0_41[441]},
      {stage0_42[295]},
      {stage0_43[102], stage0_43[103], stage0_43[104], stage0_43[105], stage0_43[106], stage0_43[107]},
      {stage1_45[17],stage1_44[66],stage1_43[122],stage1_42[127],stage1_41[154]}
   );
   gpc615_5 gpc1607 (
      {stage0_41[442], stage0_41[443], stage0_41[444], stage0_41[445], stage0_41[446]},
      {stage0_42[296]},
      {stage0_43[108], stage0_43[109], stage0_43[110], stage0_43[111], stage0_43[112], stage0_43[113]},
      {stage1_45[18],stage1_44[67],stage1_43[123],stage1_42[128],stage1_41[155]}
   );
   gpc615_5 gpc1608 (
      {stage0_41[447], stage0_41[448], stage0_41[449], stage0_41[450], stage0_41[451]},
      {stage0_42[297]},
      {stage0_43[114], stage0_43[115], stage0_43[116], stage0_43[117], stage0_43[118], stage0_43[119]},
      {stage1_45[19],stage1_44[68],stage1_43[124],stage1_42[129],stage1_41[156]}
   );
   gpc615_5 gpc1609 (
      {stage0_41[452], stage0_41[453], stage0_41[454], stage0_41[455], stage0_41[456]},
      {stage0_42[298]},
      {stage0_43[120], stage0_43[121], stage0_43[122], stage0_43[123], stage0_43[124], stage0_43[125]},
      {stage1_45[20],stage1_44[69],stage1_43[125],stage1_42[130],stage1_41[157]}
   );
   gpc615_5 gpc1610 (
      {stage0_41[457], stage0_41[458], stage0_41[459], stage0_41[460], stage0_41[461]},
      {stage0_42[299]},
      {stage0_43[126], stage0_43[127], stage0_43[128], stage0_43[129], stage0_43[130], stage0_43[131]},
      {stage1_45[21],stage1_44[70],stage1_43[126],stage1_42[131],stage1_41[158]}
   );
   gpc615_5 gpc1611 (
      {stage0_41[462], stage0_41[463], stage0_41[464], stage0_41[465], stage0_41[466]},
      {stage0_42[300]},
      {stage0_43[132], stage0_43[133], stage0_43[134], stage0_43[135], stage0_43[136], stage0_43[137]},
      {stage1_45[22],stage1_44[71],stage1_43[127],stage1_42[132],stage1_41[159]}
   );
   gpc615_5 gpc1612 (
      {stage0_41[467], stage0_41[468], stage0_41[469], stage0_41[470], stage0_41[471]},
      {stage0_42[301]},
      {stage0_43[138], stage0_43[139], stage0_43[140], stage0_43[141], stage0_43[142], stage0_43[143]},
      {stage1_45[23],stage1_44[72],stage1_43[128],stage1_42[133],stage1_41[160]}
   );
   gpc615_5 gpc1613 (
      {stage0_41[472], stage0_41[473], stage0_41[474], stage0_41[475], stage0_41[476]},
      {stage0_42[302]},
      {stage0_43[144], stage0_43[145], stage0_43[146], stage0_43[147], stage0_43[148], stage0_43[149]},
      {stage1_45[24],stage1_44[73],stage1_43[129],stage1_42[134],stage1_41[161]}
   );
   gpc615_5 gpc1614 (
      {stage0_42[303], stage0_42[304], stage0_42[305], stage0_42[306], stage0_42[307]},
      {stage0_43[150]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[25],stage1_44[74],stage1_43[130],stage1_42[135]}
   );
   gpc615_5 gpc1615 (
      {stage0_42[308], stage0_42[309], stage0_42[310], stage0_42[311], stage0_42[312]},
      {stage0_43[151]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[26],stage1_44[75],stage1_43[131],stage1_42[136]}
   );
   gpc615_5 gpc1616 (
      {stage0_42[313], stage0_42[314], stage0_42[315], stage0_42[316], stage0_42[317]},
      {stage0_43[152]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[27],stage1_44[76],stage1_43[132],stage1_42[137]}
   );
   gpc615_5 gpc1617 (
      {stage0_42[318], stage0_42[319], stage0_42[320], stage0_42[321], stage0_42[322]},
      {stage0_43[153]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[28],stage1_44[77],stage1_43[133],stage1_42[138]}
   );
   gpc615_5 gpc1618 (
      {stage0_42[323], stage0_42[324], stage0_42[325], stage0_42[326], stage0_42[327]},
      {stage0_43[154]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[29],stage1_44[78],stage1_43[134],stage1_42[139]}
   );
   gpc615_5 gpc1619 (
      {stage0_42[328], stage0_42[329], stage0_42[330], stage0_42[331], stage0_42[332]},
      {stage0_43[155]},
      {stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33], stage0_44[34], stage0_44[35]},
      {stage1_46[5],stage1_45[30],stage1_44[79],stage1_43[135],stage1_42[140]}
   );
   gpc615_5 gpc1620 (
      {stage0_42[333], stage0_42[334], stage0_42[335], stage0_42[336], stage0_42[337]},
      {stage0_43[156]},
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage1_46[6],stage1_45[31],stage1_44[80],stage1_43[136],stage1_42[141]}
   );
   gpc615_5 gpc1621 (
      {stage0_42[338], stage0_42[339], stage0_42[340], stage0_42[341], stage0_42[342]},
      {stage0_43[157]},
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage1_46[7],stage1_45[32],stage1_44[81],stage1_43[137],stage1_42[142]}
   );
   gpc615_5 gpc1622 (
      {stage0_42[343], stage0_42[344], stage0_42[345], stage0_42[346], stage0_42[347]},
      {stage0_43[158]},
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage1_46[8],stage1_45[33],stage1_44[82],stage1_43[138],stage1_42[143]}
   );
   gpc615_5 gpc1623 (
      {stage0_42[348], stage0_42[349], stage0_42[350], stage0_42[351], stage0_42[352]},
      {stage0_43[159]},
      {stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57], stage0_44[58], stage0_44[59]},
      {stage1_46[9],stage1_45[34],stage1_44[83],stage1_43[139],stage1_42[144]}
   );
   gpc615_5 gpc1624 (
      {stage0_42[353], stage0_42[354], stage0_42[355], stage0_42[356], stage0_42[357]},
      {stage0_43[160]},
      {stage0_44[60], stage0_44[61], stage0_44[62], stage0_44[63], stage0_44[64], stage0_44[65]},
      {stage1_46[10],stage1_45[35],stage1_44[84],stage1_43[140],stage1_42[145]}
   );
   gpc615_5 gpc1625 (
      {stage0_42[358], stage0_42[359], stage0_42[360], stage0_42[361], stage0_42[362]},
      {stage0_43[161]},
      {stage0_44[66], stage0_44[67], stage0_44[68], stage0_44[69], stage0_44[70], stage0_44[71]},
      {stage1_46[11],stage1_45[36],stage1_44[85],stage1_43[141],stage1_42[146]}
   );
   gpc615_5 gpc1626 (
      {stage0_42[363], stage0_42[364], stage0_42[365], stage0_42[366], stage0_42[367]},
      {stage0_43[162]},
      {stage0_44[72], stage0_44[73], stage0_44[74], stage0_44[75], stage0_44[76], stage0_44[77]},
      {stage1_46[12],stage1_45[37],stage1_44[86],stage1_43[142],stage1_42[147]}
   );
   gpc615_5 gpc1627 (
      {stage0_42[368], stage0_42[369], stage0_42[370], stage0_42[371], stage0_42[372]},
      {stage0_43[163]},
      {stage0_44[78], stage0_44[79], stage0_44[80], stage0_44[81], stage0_44[82], stage0_44[83]},
      {stage1_46[13],stage1_45[38],stage1_44[87],stage1_43[143],stage1_42[148]}
   );
   gpc615_5 gpc1628 (
      {stage0_42[373], stage0_42[374], stage0_42[375], stage0_42[376], stage0_42[377]},
      {stage0_43[164]},
      {stage0_44[84], stage0_44[85], stage0_44[86], stage0_44[87], stage0_44[88], stage0_44[89]},
      {stage1_46[14],stage1_45[39],stage1_44[88],stage1_43[144],stage1_42[149]}
   );
   gpc615_5 gpc1629 (
      {stage0_42[378], stage0_42[379], stage0_42[380], stage0_42[381], stage0_42[382]},
      {stage0_43[165]},
      {stage0_44[90], stage0_44[91], stage0_44[92], stage0_44[93], stage0_44[94], stage0_44[95]},
      {stage1_46[15],stage1_45[40],stage1_44[89],stage1_43[145],stage1_42[150]}
   );
   gpc615_5 gpc1630 (
      {stage0_42[383], stage0_42[384], stage0_42[385], stage0_42[386], stage0_42[387]},
      {stage0_43[166]},
      {stage0_44[96], stage0_44[97], stage0_44[98], stage0_44[99], stage0_44[100], stage0_44[101]},
      {stage1_46[16],stage1_45[41],stage1_44[90],stage1_43[146],stage1_42[151]}
   );
   gpc615_5 gpc1631 (
      {stage0_42[388], stage0_42[389], stage0_42[390], stage0_42[391], stage0_42[392]},
      {stage0_43[167]},
      {stage0_44[102], stage0_44[103], stage0_44[104], stage0_44[105], stage0_44[106], stage0_44[107]},
      {stage1_46[17],stage1_45[42],stage1_44[91],stage1_43[147],stage1_42[152]}
   );
   gpc615_5 gpc1632 (
      {stage0_42[393], stage0_42[394], stage0_42[395], stage0_42[396], stage0_42[397]},
      {stage0_43[168]},
      {stage0_44[108], stage0_44[109], stage0_44[110], stage0_44[111], stage0_44[112], stage0_44[113]},
      {stage1_46[18],stage1_45[43],stage1_44[92],stage1_43[148],stage1_42[153]}
   );
   gpc615_5 gpc1633 (
      {stage0_42[398], stage0_42[399], stage0_42[400], stage0_42[401], stage0_42[402]},
      {stage0_43[169]},
      {stage0_44[114], stage0_44[115], stage0_44[116], stage0_44[117], stage0_44[118], stage0_44[119]},
      {stage1_46[19],stage1_45[44],stage1_44[93],stage1_43[149],stage1_42[154]}
   );
   gpc615_5 gpc1634 (
      {stage0_42[403], stage0_42[404], stage0_42[405], stage0_42[406], stage0_42[407]},
      {stage0_43[170]},
      {stage0_44[120], stage0_44[121], stage0_44[122], stage0_44[123], stage0_44[124], stage0_44[125]},
      {stage1_46[20],stage1_45[45],stage1_44[94],stage1_43[150],stage1_42[155]}
   );
   gpc615_5 gpc1635 (
      {stage0_42[408], stage0_42[409], stage0_42[410], stage0_42[411], stage0_42[412]},
      {stage0_43[171]},
      {stage0_44[126], stage0_44[127], stage0_44[128], stage0_44[129], stage0_44[130], stage0_44[131]},
      {stage1_46[21],stage1_45[46],stage1_44[95],stage1_43[151],stage1_42[156]}
   );
   gpc615_5 gpc1636 (
      {stage0_42[413], stage0_42[414], stage0_42[415], stage0_42[416], stage0_42[417]},
      {stage0_43[172]},
      {stage0_44[132], stage0_44[133], stage0_44[134], stage0_44[135], stage0_44[136], stage0_44[137]},
      {stage1_46[22],stage1_45[47],stage1_44[96],stage1_43[152],stage1_42[157]}
   );
   gpc615_5 gpc1637 (
      {stage0_42[418], stage0_42[419], stage0_42[420], stage0_42[421], stage0_42[422]},
      {stage0_43[173]},
      {stage0_44[138], stage0_44[139], stage0_44[140], stage0_44[141], stage0_44[142], stage0_44[143]},
      {stage1_46[23],stage1_45[48],stage1_44[97],stage1_43[153],stage1_42[158]}
   );
   gpc615_5 gpc1638 (
      {stage0_42[423], stage0_42[424], stage0_42[425], stage0_42[426], stage0_42[427]},
      {stage0_43[174]},
      {stage0_44[144], stage0_44[145], stage0_44[146], stage0_44[147], stage0_44[148], stage0_44[149]},
      {stage1_46[24],stage1_45[49],stage1_44[98],stage1_43[154],stage1_42[159]}
   );
   gpc615_5 gpc1639 (
      {stage0_42[428], stage0_42[429], stage0_42[430], stage0_42[431], stage0_42[432]},
      {stage0_43[175]},
      {stage0_44[150], stage0_44[151], stage0_44[152], stage0_44[153], stage0_44[154], stage0_44[155]},
      {stage1_46[25],stage1_45[50],stage1_44[99],stage1_43[155],stage1_42[160]}
   );
   gpc615_5 gpc1640 (
      {stage0_42[433], stage0_42[434], stage0_42[435], stage0_42[436], stage0_42[437]},
      {stage0_43[176]},
      {stage0_44[156], stage0_44[157], stage0_44[158], stage0_44[159], stage0_44[160], stage0_44[161]},
      {stage1_46[26],stage1_45[51],stage1_44[100],stage1_43[156],stage1_42[161]}
   );
   gpc615_5 gpc1641 (
      {stage0_42[438], stage0_42[439], stage0_42[440], stage0_42[441], stage0_42[442]},
      {stage0_43[177]},
      {stage0_44[162], stage0_44[163], stage0_44[164], stage0_44[165], stage0_44[166], stage0_44[167]},
      {stage1_46[27],stage1_45[52],stage1_44[101],stage1_43[157],stage1_42[162]}
   );
   gpc615_5 gpc1642 (
      {stage0_42[443], stage0_42[444], stage0_42[445], stage0_42[446], stage0_42[447]},
      {stage0_43[178]},
      {stage0_44[168], stage0_44[169], stage0_44[170], stage0_44[171], stage0_44[172], stage0_44[173]},
      {stage1_46[28],stage1_45[53],stage1_44[102],stage1_43[158],stage1_42[163]}
   );
   gpc615_5 gpc1643 (
      {stage0_42[448], stage0_42[449], stage0_42[450], stage0_42[451], stage0_42[452]},
      {stage0_43[179]},
      {stage0_44[174], stage0_44[175], stage0_44[176], stage0_44[177], stage0_44[178], stage0_44[179]},
      {stage1_46[29],stage1_45[54],stage1_44[103],stage1_43[159],stage1_42[164]}
   );
   gpc615_5 gpc1644 (
      {stage0_42[453], stage0_42[454], stage0_42[455], stage0_42[456], stage0_42[457]},
      {stage0_43[180]},
      {stage0_44[180], stage0_44[181], stage0_44[182], stage0_44[183], stage0_44[184], stage0_44[185]},
      {stage1_46[30],stage1_45[55],stage1_44[104],stage1_43[160],stage1_42[165]}
   );
   gpc615_5 gpc1645 (
      {stage0_42[458], stage0_42[459], stage0_42[460], stage0_42[461], stage0_42[462]},
      {stage0_43[181]},
      {stage0_44[186], stage0_44[187], stage0_44[188], stage0_44[189], stage0_44[190], stage0_44[191]},
      {stage1_46[31],stage1_45[56],stage1_44[105],stage1_43[161],stage1_42[166]}
   );
   gpc615_5 gpc1646 (
      {stage0_42[463], stage0_42[464], stage0_42[465], stage0_42[466], stage0_42[467]},
      {stage0_43[182]},
      {stage0_44[192], stage0_44[193], stage0_44[194], stage0_44[195], stage0_44[196], stage0_44[197]},
      {stage1_46[32],stage1_45[57],stage1_44[106],stage1_43[162],stage1_42[167]}
   );
   gpc615_5 gpc1647 (
      {stage0_42[468], stage0_42[469], stage0_42[470], stage0_42[471], stage0_42[472]},
      {stage0_43[183]},
      {stage0_44[198], stage0_44[199], stage0_44[200], stage0_44[201], stage0_44[202], stage0_44[203]},
      {stage1_46[33],stage1_45[58],stage1_44[107],stage1_43[163],stage1_42[168]}
   );
   gpc615_5 gpc1648 (
      {stage0_42[473], stage0_42[474], stage0_42[475], stage0_42[476], stage0_42[477]},
      {stage0_43[184]},
      {stage0_44[204], stage0_44[205], stage0_44[206], stage0_44[207], stage0_44[208], stage0_44[209]},
      {stage1_46[34],stage1_45[59],stage1_44[108],stage1_43[164],stage1_42[169]}
   );
   gpc615_5 gpc1649 (
      {stage0_42[478], stage0_42[479], stage0_42[480], stage0_42[481], stage0_42[482]},
      {stage0_43[185]},
      {stage0_44[210], stage0_44[211], stage0_44[212], stage0_44[213], stage0_44[214], stage0_44[215]},
      {stage1_46[35],stage1_45[60],stage1_44[109],stage1_43[165],stage1_42[170]}
   );
   gpc615_5 gpc1650 (
      {stage0_43[186], stage0_43[187], stage0_43[188], stage0_43[189], stage0_43[190]},
      {stage0_44[216]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[36],stage1_45[61],stage1_44[110],stage1_43[166]}
   );
   gpc615_5 gpc1651 (
      {stage0_43[191], stage0_43[192], stage0_43[193], stage0_43[194], stage0_43[195]},
      {stage0_44[217]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[37],stage1_45[62],stage1_44[111],stage1_43[167]}
   );
   gpc615_5 gpc1652 (
      {stage0_43[196], stage0_43[197], stage0_43[198], stage0_43[199], stage0_43[200]},
      {stage0_44[218]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[38],stage1_45[63],stage1_44[112],stage1_43[168]}
   );
   gpc615_5 gpc1653 (
      {stage0_43[201], stage0_43[202], stage0_43[203], stage0_43[204], stage0_43[205]},
      {stage0_44[219]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[39],stage1_45[64],stage1_44[113],stage1_43[169]}
   );
   gpc615_5 gpc1654 (
      {stage0_43[206], stage0_43[207], stage0_43[208], stage0_43[209], stage0_43[210]},
      {stage0_44[220]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[40],stage1_45[65],stage1_44[114],stage1_43[170]}
   );
   gpc615_5 gpc1655 (
      {stage0_43[211], stage0_43[212], stage0_43[213], stage0_43[214], stage0_43[215]},
      {stage0_44[221]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[41],stage1_45[66],stage1_44[115],stage1_43[171]}
   );
   gpc615_5 gpc1656 (
      {stage0_43[216], stage0_43[217], stage0_43[218], stage0_43[219], stage0_43[220]},
      {stage0_44[222]},
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40], stage0_45[41]},
      {stage1_47[6],stage1_46[42],stage1_45[67],stage1_44[116],stage1_43[172]}
   );
   gpc615_5 gpc1657 (
      {stage0_43[221], stage0_43[222], stage0_43[223], stage0_43[224], stage0_43[225]},
      {stage0_44[223]},
      {stage0_45[42], stage0_45[43], stage0_45[44], stage0_45[45], stage0_45[46], stage0_45[47]},
      {stage1_47[7],stage1_46[43],stage1_45[68],stage1_44[117],stage1_43[173]}
   );
   gpc615_5 gpc1658 (
      {stage0_43[226], stage0_43[227], stage0_43[228], stage0_43[229], stage0_43[230]},
      {stage0_44[224]},
      {stage0_45[48], stage0_45[49], stage0_45[50], stage0_45[51], stage0_45[52], stage0_45[53]},
      {stage1_47[8],stage1_46[44],stage1_45[69],stage1_44[118],stage1_43[174]}
   );
   gpc615_5 gpc1659 (
      {stage0_43[231], stage0_43[232], stage0_43[233], stage0_43[234], stage0_43[235]},
      {stage0_44[225]},
      {stage0_45[54], stage0_45[55], stage0_45[56], stage0_45[57], stage0_45[58], stage0_45[59]},
      {stage1_47[9],stage1_46[45],stage1_45[70],stage1_44[119],stage1_43[175]}
   );
   gpc615_5 gpc1660 (
      {stage0_43[236], stage0_43[237], stage0_43[238], stage0_43[239], stage0_43[240]},
      {stage0_44[226]},
      {stage0_45[60], stage0_45[61], stage0_45[62], stage0_45[63], stage0_45[64], stage0_45[65]},
      {stage1_47[10],stage1_46[46],stage1_45[71],stage1_44[120],stage1_43[176]}
   );
   gpc615_5 gpc1661 (
      {stage0_43[241], stage0_43[242], stage0_43[243], stage0_43[244], stage0_43[245]},
      {stage0_44[227]},
      {stage0_45[66], stage0_45[67], stage0_45[68], stage0_45[69], stage0_45[70], stage0_45[71]},
      {stage1_47[11],stage1_46[47],stage1_45[72],stage1_44[121],stage1_43[177]}
   );
   gpc615_5 gpc1662 (
      {stage0_43[246], stage0_43[247], stage0_43[248], stage0_43[249], stage0_43[250]},
      {stage0_44[228]},
      {stage0_45[72], stage0_45[73], stage0_45[74], stage0_45[75], stage0_45[76], stage0_45[77]},
      {stage1_47[12],stage1_46[48],stage1_45[73],stage1_44[122],stage1_43[178]}
   );
   gpc615_5 gpc1663 (
      {stage0_43[251], stage0_43[252], stage0_43[253], stage0_43[254], stage0_43[255]},
      {stage0_44[229]},
      {stage0_45[78], stage0_45[79], stage0_45[80], stage0_45[81], stage0_45[82], stage0_45[83]},
      {stage1_47[13],stage1_46[49],stage1_45[74],stage1_44[123],stage1_43[179]}
   );
   gpc615_5 gpc1664 (
      {stage0_43[256], stage0_43[257], stage0_43[258], stage0_43[259], stage0_43[260]},
      {stage0_44[230]},
      {stage0_45[84], stage0_45[85], stage0_45[86], stage0_45[87], stage0_45[88], stage0_45[89]},
      {stage1_47[14],stage1_46[50],stage1_45[75],stage1_44[124],stage1_43[180]}
   );
   gpc615_5 gpc1665 (
      {stage0_43[261], stage0_43[262], stage0_43[263], stage0_43[264], stage0_43[265]},
      {stage0_44[231]},
      {stage0_45[90], stage0_45[91], stage0_45[92], stage0_45[93], stage0_45[94], stage0_45[95]},
      {stage1_47[15],stage1_46[51],stage1_45[76],stage1_44[125],stage1_43[181]}
   );
   gpc615_5 gpc1666 (
      {stage0_43[266], stage0_43[267], stage0_43[268], stage0_43[269], stage0_43[270]},
      {stage0_44[232]},
      {stage0_45[96], stage0_45[97], stage0_45[98], stage0_45[99], stage0_45[100], stage0_45[101]},
      {stage1_47[16],stage1_46[52],stage1_45[77],stage1_44[126],stage1_43[182]}
   );
   gpc615_5 gpc1667 (
      {stage0_43[271], stage0_43[272], stage0_43[273], stage0_43[274], stage0_43[275]},
      {stage0_44[233]},
      {stage0_45[102], stage0_45[103], stage0_45[104], stage0_45[105], stage0_45[106], stage0_45[107]},
      {stage1_47[17],stage1_46[53],stage1_45[78],stage1_44[127],stage1_43[183]}
   );
   gpc615_5 gpc1668 (
      {stage0_43[276], stage0_43[277], stage0_43[278], stage0_43[279], stage0_43[280]},
      {stage0_44[234]},
      {stage0_45[108], stage0_45[109], stage0_45[110], stage0_45[111], stage0_45[112], stage0_45[113]},
      {stage1_47[18],stage1_46[54],stage1_45[79],stage1_44[128],stage1_43[184]}
   );
   gpc615_5 gpc1669 (
      {stage0_43[281], stage0_43[282], stage0_43[283], stage0_43[284], stage0_43[285]},
      {stage0_44[235]},
      {stage0_45[114], stage0_45[115], stage0_45[116], stage0_45[117], stage0_45[118], stage0_45[119]},
      {stage1_47[19],stage1_46[55],stage1_45[80],stage1_44[129],stage1_43[185]}
   );
   gpc615_5 gpc1670 (
      {stage0_43[286], stage0_43[287], stage0_43[288], stage0_43[289], stage0_43[290]},
      {stage0_44[236]},
      {stage0_45[120], stage0_45[121], stage0_45[122], stage0_45[123], stage0_45[124], stage0_45[125]},
      {stage1_47[20],stage1_46[56],stage1_45[81],stage1_44[130],stage1_43[186]}
   );
   gpc615_5 gpc1671 (
      {stage0_43[291], stage0_43[292], stage0_43[293], stage0_43[294], stage0_43[295]},
      {stage0_44[237]},
      {stage0_45[126], stage0_45[127], stage0_45[128], stage0_45[129], stage0_45[130], stage0_45[131]},
      {stage1_47[21],stage1_46[57],stage1_45[82],stage1_44[131],stage1_43[187]}
   );
   gpc615_5 gpc1672 (
      {stage0_43[296], stage0_43[297], stage0_43[298], stage0_43[299], stage0_43[300]},
      {stage0_44[238]},
      {stage0_45[132], stage0_45[133], stage0_45[134], stage0_45[135], stage0_45[136], stage0_45[137]},
      {stage1_47[22],stage1_46[58],stage1_45[83],stage1_44[132],stage1_43[188]}
   );
   gpc615_5 gpc1673 (
      {stage0_43[301], stage0_43[302], stage0_43[303], stage0_43[304], stage0_43[305]},
      {stage0_44[239]},
      {stage0_45[138], stage0_45[139], stage0_45[140], stage0_45[141], stage0_45[142], stage0_45[143]},
      {stage1_47[23],stage1_46[59],stage1_45[84],stage1_44[133],stage1_43[189]}
   );
   gpc615_5 gpc1674 (
      {stage0_43[306], stage0_43[307], stage0_43[308], stage0_43[309], stage0_43[310]},
      {stage0_44[240]},
      {stage0_45[144], stage0_45[145], stage0_45[146], stage0_45[147], stage0_45[148], stage0_45[149]},
      {stage1_47[24],stage1_46[60],stage1_45[85],stage1_44[134],stage1_43[190]}
   );
   gpc615_5 gpc1675 (
      {stage0_43[311], stage0_43[312], stage0_43[313], stage0_43[314], stage0_43[315]},
      {stage0_44[241]},
      {stage0_45[150], stage0_45[151], stage0_45[152], stage0_45[153], stage0_45[154], stage0_45[155]},
      {stage1_47[25],stage1_46[61],stage1_45[86],stage1_44[135],stage1_43[191]}
   );
   gpc615_5 gpc1676 (
      {stage0_43[316], stage0_43[317], stage0_43[318], stage0_43[319], stage0_43[320]},
      {stage0_44[242]},
      {stage0_45[156], stage0_45[157], stage0_45[158], stage0_45[159], stage0_45[160], stage0_45[161]},
      {stage1_47[26],stage1_46[62],stage1_45[87],stage1_44[136],stage1_43[192]}
   );
   gpc615_5 gpc1677 (
      {stage0_43[321], stage0_43[322], stage0_43[323], stage0_43[324], stage0_43[325]},
      {stage0_44[243]},
      {stage0_45[162], stage0_45[163], stage0_45[164], stage0_45[165], stage0_45[166], stage0_45[167]},
      {stage1_47[27],stage1_46[63],stage1_45[88],stage1_44[137],stage1_43[193]}
   );
   gpc615_5 gpc1678 (
      {stage0_43[326], stage0_43[327], stage0_43[328], stage0_43[329], stage0_43[330]},
      {stage0_44[244]},
      {stage0_45[168], stage0_45[169], stage0_45[170], stage0_45[171], stage0_45[172], stage0_45[173]},
      {stage1_47[28],stage1_46[64],stage1_45[89],stage1_44[138],stage1_43[194]}
   );
   gpc615_5 gpc1679 (
      {stage0_43[331], stage0_43[332], stage0_43[333], stage0_43[334], stage0_43[335]},
      {stage0_44[245]},
      {stage0_45[174], stage0_45[175], stage0_45[176], stage0_45[177], stage0_45[178], stage0_45[179]},
      {stage1_47[29],stage1_46[65],stage1_45[90],stage1_44[139],stage1_43[195]}
   );
   gpc615_5 gpc1680 (
      {stage0_43[336], stage0_43[337], stage0_43[338], stage0_43[339], stage0_43[340]},
      {stage0_44[246]},
      {stage0_45[180], stage0_45[181], stage0_45[182], stage0_45[183], stage0_45[184], stage0_45[185]},
      {stage1_47[30],stage1_46[66],stage1_45[91],stage1_44[140],stage1_43[196]}
   );
   gpc615_5 gpc1681 (
      {stage0_43[341], stage0_43[342], stage0_43[343], stage0_43[344], stage0_43[345]},
      {stage0_44[247]},
      {stage0_45[186], stage0_45[187], stage0_45[188], stage0_45[189], stage0_45[190], stage0_45[191]},
      {stage1_47[31],stage1_46[67],stage1_45[92],stage1_44[141],stage1_43[197]}
   );
   gpc615_5 gpc1682 (
      {stage0_43[346], stage0_43[347], stage0_43[348], stage0_43[349], stage0_43[350]},
      {stage0_44[248]},
      {stage0_45[192], stage0_45[193], stage0_45[194], stage0_45[195], stage0_45[196], stage0_45[197]},
      {stage1_47[32],stage1_46[68],stage1_45[93],stage1_44[142],stage1_43[198]}
   );
   gpc615_5 gpc1683 (
      {stage0_43[351], stage0_43[352], stage0_43[353], stage0_43[354], stage0_43[355]},
      {stage0_44[249]},
      {stage0_45[198], stage0_45[199], stage0_45[200], stage0_45[201], stage0_45[202], stage0_45[203]},
      {stage1_47[33],stage1_46[69],stage1_45[94],stage1_44[143],stage1_43[199]}
   );
   gpc615_5 gpc1684 (
      {stage0_43[356], stage0_43[357], stage0_43[358], stage0_43[359], stage0_43[360]},
      {stage0_44[250]},
      {stage0_45[204], stage0_45[205], stage0_45[206], stage0_45[207], stage0_45[208], stage0_45[209]},
      {stage1_47[34],stage1_46[70],stage1_45[95],stage1_44[144],stage1_43[200]}
   );
   gpc615_5 gpc1685 (
      {stage0_43[361], stage0_43[362], stage0_43[363], stage0_43[364], stage0_43[365]},
      {stage0_44[251]},
      {stage0_45[210], stage0_45[211], stage0_45[212], stage0_45[213], stage0_45[214], stage0_45[215]},
      {stage1_47[35],stage1_46[71],stage1_45[96],stage1_44[145],stage1_43[201]}
   );
   gpc615_5 gpc1686 (
      {stage0_43[366], stage0_43[367], stage0_43[368], stage0_43[369], stage0_43[370]},
      {stage0_44[252]},
      {stage0_45[216], stage0_45[217], stage0_45[218], stage0_45[219], stage0_45[220], stage0_45[221]},
      {stage1_47[36],stage1_46[72],stage1_45[97],stage1_44[146],stage1_43[202]}
   );
   gpc615_5 gpc1687 (
      {stage0_43[371], stage0_43[372], stage0_43[373], stage0_43[374], stage0_43[375]},
      {stage0_44[253]},
      {stage0_45[222], stage0_45[223], stage0_45[224], stage0_45[225], stage0_45[226], stage0_45[227]},
      {stage1_47[37],stage1_46[73],stage1_45[98],stage1_44[147],stage1_43[203]}
   );
   gpc615_5 gpc1688 (
      {stage0_43[376], stage0_43[377], stage0_43[378], stage0_43[379], stage0_43[380]},
      {stage0_44[254]},
      {stage0_45[228], stage0_45[229], stage0_45[230], stage0_45[231], stage0_45[232], stage0_45[233]},
      {stage1_47[38],stage1_46[74],stage1_45[99],stage1_44[148],stage1_43[204]}
   );
   gpc615_5 gpc1689 (
      {stage0_43[381], stage0_43[382], stage0_43[383], stage0_43[384], stage0_43[385]},
      {stage0_44[255]},
      {stage0_45[234], stage0_45[235], stage0_45[236], stage0_45[237], stage0_45[238], stage0_45[239]},
      {stage1_47[39],stage1_46[75],stage1_45[100],stage1_44[149],stage1_43[205]}
   );
   gpc615_5 gpc1690 (
      {stage0_43[386], stage0_43[387], stage0_43[388], stage0_43[389], stage0_43[390]},
      {stage0_44[256]},
      {stage0_45[240], stage0_45[241], stage0_45[242], stage0_45[243], stage0_45[244], stage0_45[245]},
      {stage1_47[40],stage1_46[76],stage1_45[101],stage1_44[150],stage1_43[206]}
   );
   gpc615_5 gpc1691 (
      {stage0_43[391], stage0_43[392], stage0_43[393], stage0_43[394], stage0_43[395]},
      {stage0_44[257]},
      {stage0_45[246], stage0_45[247], stage0_45[248], stage0_45[249], stage0_45[250], stage0_45[251]},
      {stage1_47[41],stage1_46[77],stage1_45[102],stage1_44[151],stage1_43[207]}
   );
   gpc615_5 gpc1692 (
      {stage0_43[396], stage0_43[397], stage0_43[398], stage0_43[399], stage0_43[400]},
      {stage0_44[258]},
      {stage0_45[252], stage0_45[253], stage0_45[254], stage0_45[255], stage0_45[256], stage0_45[257]},
      {stage1_47[42],stage1_46[78],stage1_45[103],stage1_44[152],stage1_43[208]}
   );
   gpc615_5 gpc1693 (
      {stage0_43[401], stage0_43[402], stage0_43[403], stage0_43[404], stage0_43[405]},
      {stage0_44[259]},
      {stage0_45[258], stage0_45[259], stage0_45[260], stage0_45[261], stage0_45[262], stage0_45[263]},
      {stage1_47[43],stage1_46[79],stage1_45[104],stage1_44[153],stage1_43[209]}
   );
   gpc615_5 gpc1694 (
      {stage0_43[406], stage0_43[407], stage0_43[408], stage0_43[409], stage0_43[410]},
      {stage0_44[260]},
      {stage0_45[264], stage0_45[265], stage0_45[266], stage0_45[267], stage0_45[268], stage0_45[269]},
      {stage1_47[44],stage1_46[80],stage1_45[105],stage1_44[154],stage1_43[210]}
   );
   gpc615_5 gpc1695 (
      {stage0_43[411], stage0_43[412], stage0_43[413], stage0_43[414], stage0_43[415]},
      {stage0_44[261]},
      {stage0_45[270], stage0_45[271], stage0_45[272], stage0_45[273], stage0_45[274], stage0_45[275]},
      {stage1_47[45],stage1_46[81],stage1_45[106],stage1_44[155],stage1_43[211]}
   );
   gpc615_5 gpc1696 (
      {stage0_43[416], stage0_43[417], stage0_43[418], stage0_43[419], stage0_43[420]},
      {stage0_44[262]},
      {stage0_45[276], stage0_45[277], stage0_45[278], stage0_45[279], stage0_45[280], stage0_45[281]},
      {stage1_47[46],stage1_46[82],stage1_45[107],stage1_44[156],stage1_43[212]}
   );
   gpc615_5 gpc1697 (
      {stage0_43[421], stage0_43[422], stage0_43[423], stage0_43[424], stage0_43[425]},
      {stage0_44[263]},
      {stage0_45[282], stage0_45[283], stage0_45[284], stage0_45[285], stage0_45[286], stage0_45[287]},
      {stage1_47[47],stage1_46[83],stage1_45[108],stage1_44[157],stage1_43[213]}
   );
   gpc615_5 gpc1698 (
      {stage0_43[426], stage0_43[427], stage0_43[428], stage0_43[429], stage0_43[430]},
      {stage0_44[264]},
      {stage0_45[288], stage0_45[289], stage0_45[290], stage0_45[291], stage0_45[292], stage0_45[293]},
      {stage1_47[48],stage1_46[84],stage1_45[109],stage1_44[158],stage1_43[214]}
   );
   gpc615_5 gpc1699 (
      {stage0_43[431], stage0_43[432], stage0_43[433], stage0_43[434], stage0_43[435]},
      {stage0_44[265]},
      {stage0_45[294], stage0_45[295], stage0_45[296], stage0_45[297], stage0_45[298], stage0_45[299]},
      {stage1_47[49],stage1_46[85],stage1_45[110],stage1_44[159],stage1_43[215]}
   );
   gpc615_5 gpc1700 (
      {stage0_43[436], stage0_43[437], stage0_43[438], stage0_43[439], stage0_43[440]},
      {stage0_44[266]},
      {stage0_45[300], stage0_45[301], stage0_45[302], stage0_45[303], stage0_45[304], stage0_45[305]},
      {stage1_47[50],stage1_46[86],stage1_45[111],stage1_44[160],stage1_43[216]}
   );
   gpc615_5 gpc1701 (
      {stage0_43[441], stage0_43[442], stage0_43[443], stage0_43[444], stage0_43[445]},
      {stage0_44[267]},
      {stage0_45[306], stage0_45[307], stage0_45[308], stage0_45[309], stage0_45[310], stage0_45[311]},
      {stage1_47[51],stage1_46[87],stage1_45[112],stage1_44[161],stage1_43[217]}
   );
   gpc615_5 gpc1702 (
      {stage0_43[446], stage0_43[447], stage0_43[448], stage0_43[449], stage0_43[450]},
      {stage0_44[268]},
      {stage0_45[312], stage0_45[313], stage0_45[314], stage0_45[315], stage0_45[316], stage0_45[317]},
      {stage1_47[52],stage1_46[88],stage1_45[113],stage1_44[162],stage1_43[218]}
   );
   gpc615_5 gpc1703 (
      {stage0_44[269], stage0_44[270], stage0_44[271], stage0_44[272], stage0_44[273]},
      {stage0_45[318]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[53],stage1_46[89],stage1_45[114],stage1_44[163]}
   );
   gpc615_5 gpc1704 (
      {stage0_44[274], stage0_44[275], stage0_44[276], stage0_44[277], stage0_44[278]},
      {stage0_45[319]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[54],stage1_46[90],stage1_45[115],stage1_44[164]}
   );
   gpc615_5 gpc1705 (
      {stage0_44[279], stage0_44[280], stage0_44[281], stage0_44[282], stage0_44[283]},
      {stage0_45[320]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[55],stage1_46[91],stage1_45[116],stage1_44[165]}
   );
   gpc615_5 gpc1706 (
      {stage0_44[284], stage0_44[285], stage0_44[286], stage0_44[287], stage0_44[288]},
      {stage0_45[321]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[56],stage1_46[92],stage1_45[117],stage1_44[166]}
   );
   gpc615_5 gpc1707 (
      {stage0_44[289], stage0_44[290], stage0_44[291], stage0_44[292], stage0_44[293]},
      {stage0_45[322]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[57],stage1_46[93],stage1_45[118],stage1_44[167]}
   );
   gpc615_5 gpc1708 (
      {stage0_44[294], stage0_44[295], stage0_44[296], stage0_44[297], stage0_44[298]},
      {stage0_45[323]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[58],stage1_46[94],stage1_45[119],stage1_44[168]}
   );
   gpc615_5 gpc1709 (
      {stage0_44[299], stage0_44[300], stage0_44[301], stage0_44[302], stage0_44[303]},
      {stage0_45[324]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[59],stage1_46[95],stage1_45[120],stage1_44[169]}
   );
   gpc615_5 gpc1710 (
      {stage0_44[304], stage0_44[305], stage0_44[306], stage0_44[307], stage0_44[308]},
      {stage0_45[325]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[60],stage1_46[96],stage1_45[121],stage1_44[170]}
   );
   gpc615_5 gpc1711 (
      {stage0_44[309], stage0_44[310], stage0_44[311], stage0_44[312], stage0_44[313]},
      {stage0_45[326]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[61],stage1_46[97],stage1_45[122],stage1_44[171]}
   );
   gpc615_5 gpc1712 (
      {stage0_44[314], stage0_44[315], stage0_44[316], stage0_44[317], stage0_44[318]},
      {stage0_45[327]},
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58], stage0_46[59]},
      {stage1_48[9],stage1_47[62],stage1_46[98],stage1_45[123],stage1_44[172]}
   );
   gpc615_5 gpc1713 (
      {stage0_44[319], stage0_44[320], stage0_44[321], stage0_44[322], stage0_44[323]},
      {stage0_45[328]},
      {stage0_46[60], stage0_46[61], stage0_46[62], stage0_46[63], stage0_46[64], stage0_46[65]},
      {stage1_48[10],stage1_47[63],stage1_46[99],stage1_45[124],stage1_44[173]}
   );
   gpc615_5 gpc1714 (
      {stage0_44[324], stage0_44[325], stage0_44[326], stage0_44[327], stage0_44[328]},
      {stage0_45[329]},
      {stage0_46[66], stage0_46[67], stage0_46[68], stage0_46[69], stage0_46[70], stage0_46[71]},
      {stage1_48[11],stage1_47[64],stage1_46[100],stage1_45[125],stage1_44[174]}
   );
   gpc615_5 gpc1715 (
      {stage0_44[329], stage0_44[330], stage0_44[331], stage0_44[332], stage0_44[333]},
      {stage0_45[330]},
      {stage0_46[72], stage0_46[73], stage0_46[74], stage0_46[75], stage0_46[76], stage0_46[77]},
      {stage1_48[12],stage1_47[65],stage1_46[101],stage1_45[126],stage1_44[175]}
   );
   gpc615_5 gpc1716 (
      {stage0_44[334], stage0_44[335], stage0_44[336], stage0_44[337], stage0_44[338]},
      {stage0_45[331]},
      {stage0_46[78], stage0_46[79], stage0_46[80], stage0_46[81], stage0_46[82], stage0_46[83]},
      {stage1_48[13],stage1_47[66],stage1_46[102],stage1_45[127],stage1_44[176]}
   );
   gpc615_5 gpc1717 (
      {stage0_44[339], stage0_44[340], stage0_44[341], stage0_44[342], stage0_44[343]},
      {stage0_45[332]},
      {stage0_46[84], stage0_46[85], stage0_46[86], stage0_46[87], stage0_46[88], stage0_46[89]},
      {stage1_48[14],stage1_47[67],stage1_46[103],stage1_45[128],stage1_44[177]}
   );
   gpc615_5 gpc1718 (
      {stage0_44[344], stage0_44[345], stage0_44[346], stage0_44[347], stage0_44[348]},
      {stage0_45[333]},
      {stage0_46[90], stage0_46[91], stage0_46[92], stage0_46[93], stage0_46[94], stage0_46[95]},
      {stage1_48[15],stage1_47[68],stage1_46[104],stage1_45[129],stage1_44[178]}
   );
   gpc615_5 gpc1719 (
      {stage0_44[349], stage0_44[350], stage0_44[351], stage0_44[352], stage0_44[353]},
      {stage0_45[334]},
      {stage0_46[96], stage0_46[97], stage0_46[98], stage0_46[99], stage0_46[100], stage0_46[101]},
      {stage1_48[16],stage1_47[69],stage1_46[105],stage1_45[130],stage1_44[179]}
   );
   gpc615_5 gpc1720 (
      {stage0_44[354], stage0_44[355], stage0_44[356], stage0_44[357], stage0_44[358]},
      {stage0_45[335]},
      {stage0_46[102], stage0_46[103], stage0_46[104], stage0_46[105], stage0_46[106], stage0_46[107]},
      {stage1_48[17],stage1_47[70],stage1_46[106],stage1_45[131],stage1_44[180]}
   );
   gpc615_5 gpc1721 (
      {stage0_44[359], stage0_44[360], stage0_44[361], stage0_44[362], stage0_44[363]},
      {stage0_45[336]},
      {stage0_46[108], stage0_46[109], stage0_46[110], stage0_46[111], stage0_46[112], stage0_46[113]},
      {stage1_48[18],stage1_47[71],stage1_46[107],stage1_45[132],stage1_44[181]}
   );
   gpc615_5 gpc1722 (
      {stage0_44[364], stage0_44[365], stage0_44[366], stage0_44[367], stage0_44[368]},
      {stage0_45[337]},
      {stage0_46[114], stage0_46[115], stage0_46[116], stage0_46[117], stage0_46[118], stage0_46[119]},
      {stage1_48[19],stage1_47[72],stage1_46[108],stage1_45[133],stage1_44[182]}
   );
   gpc615_5 gpc1723 (
      {stage0_44[369], stage0_44[370], stage0_44[371], stage0_44[372], stage0_44[373]},
      {stage0_45[338]},
      {stage0_46[120], stage0_46[121], stage0_46[122], stage0_46[123], stage0_46[124], stage0_46[125]},
      {stage1_48[20],stage1_47[73],stage1_46[109],stage1_45[134],stage1_44[183]}
   );
   gpc615_5 gpc1724 (
      {stage0_44[374], stage0_44[375], stage0_44[376], stage0_44[377], stage0_44[378]},
      {stage0_45[339]},
      {stage0_46[126], stage0_46[127], stage0_46[128], stage0_46[129], stage0_46[130], stage0_46[131]},
      {stage1_48[21],stage1_47[74],stage1_46[110],stage1_45[135],stage1_44[184]}
   );
   gpc615_5 gpc1725 (
      {stage0_44[379], stage0_44[380], stage0_44[381], stage0_44[382], stage0_44[383]},
      {stage0_45[340]},
      {stage0_46[132], stage0_46[133], stage0_46[134], stage0_46[135], stage0_46[136], stage0_46[137]},
      {stage1_48[22],stage1_47[75],stage1_46[111],stage1_45[136],stage1_44[185]}
   );
   gpc615_5 gpc1726 (
      {stage0_44[384], stage0_44[385], stage0_44[386], stage0_44[387], stage0_44[388]},
      {stage0_45[341]},
      {stage0_46[138], stage0_46[139], stage0_46[140], stage0_46[141], stage0_46[142], stage0_46[143]},
      {stage1_48[23],stage1_47[76],stage1_46[112],stage1_45[137],stage1_44[186]}
   );
   gpc615_5 gpc1727 (
      {stage0_44[389], stage0_44[390], stage0_44[391], stage0_44[392], stage0_44[393]},
      {stage0_45[342]},
      {stage0_46[144], stage0_46[145], stage0_46[146], stage0_46[147], stage0_46[148], stage0_46[149]},
      {stage1_48[24],stage1_47[77],stage1_46[113],stage1_45[138],stage1_44[187]}
   );
   gpc615_5 gpc1728 (
      {stage0_44[394], stage0_44[395], stage0_44[396], stage0_44[397], stage0_44[398]},
      {stage0_45[343]},
      {stage0_46[150], stage0_46[151], stage0_46[152], stage0_46[153], stage0_46[154], stage0_46[155]},
      {stage1_48[25],stage1_47[78],stage1_46[114],stage1_45[139],stage1_44[188]}
   );
   gpc615_5 gpc1729 (
      {stage0_44[399], stage0_44[400], stage0_44[401], stage0_44[402], stage0_44[403]},
      {stage0_45[344]},
      {stage0_46[156], stage0_46[157], stage0_46[158], stage0_46[159], stage0_46[160], stage0_46[161]},
      {stage1_48[26],stage1_47[79],stage1_46[115],stage1_45[140],stage1_44[189]}
   );
   gpc615_5 gpc1730 (
      {stage0_44[404], stage0_44[405], stage0_44[406], stage0_44[407], stage0_44[408]},
      {stage0_45[345]},
      {stage0_46[162], stage0_46[163], stage0_46[164], stage0_46[165], stage0_46[166], stage0_46[167]},
      {stage1_48[27],stage1_47[80],stage1_46[116],stage1_45[141],stage1_44[190]}
   );
   gpc615_5 gpc1731 (
      {stage0_44[409], stage0_44[410], stage0_44[411], stage0_44[412], stage0_44[413]},
      {stage0_45[346]},
      {stage0_46[168], stage0_46[169], stage0_46[170], stage0_46[171], stage0_46[172], stage0_46[173]},
      {stage1_48[28],stage1_47[81],stage1_46[117],stage1_45[142],stage1_44[191]}
   );
   gpc615_5 gpc1732 (
      {stage0_44[414], stage0_44[415], stage0_44[416], stage0_44[417], stage0_44[418]},
      {stage0_45[347]},
      {stage0_46[174], stage0_46[175], stage0_46[176], stage0_46[177], stage0_46[178], stage0_46[179]},
      {stage1_48[29],stage1_47[82],stage1_46[118],stage1_45[143],stage1_44[192]}
   );
   gpc615_5 gpc1733 (
      {stage0_44[419], stage0_44[420], stage0_44[421], stage0_44[422], stage0_44[423]},
      {stage0_45[348]},
      {stage0_46[180], stage0_46[181], stage0_46[182], stage0_46[183], stage0_46[184], stage0_46[185]},
      {stage1_48[30],stage1_47[83],stage1_46[119],stage1_45[144],stage1_44[193]}
   );
   gpc606_5 gpc1734 (
      {stage0_45[349], stage0_45[350], stage0_45[351], stage0_45[352], stage0_45[353], stage0_45[354]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[31],stage1_47[84],stage1_46[120],stage1_45[145]}
   );
   gpc606_5 gpc1735 (
      {stage0_45[355], stage0_45[356], stage0_45[357], stage0_45[358], stage0_45[359], stage0_45[360]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[32],stage1_47[85],stage1_46[121],stage1_45[146]}
   );
   gpc606_5 gpc1736 (
      {stage0_45[361], stage0_45[362], stage0_45[363], stage0_45[364], stage0_45[365], stage0_45[366]},
      {stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17]},
      {stage1_49[2],stage1_48[33],stage1_47[86],stage1_46[122],stage1_45[147]}
   );
   gpc606_5 gpc1737 (
      {stage0_45[367], stage0_45[368], stage0_45[369], stage0_45[370], stage0_45[371], stage0_45[372]},
      {stage0_47[18], stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23]},
      {stage1_49[3],stage1_48[34],stage1_47[87],stage1_46[123],stage1_45[148]}
   );
   gpc606_5 gpc1738 (
      {stage0_45[373], stage0_45[374], stage0_45[375], stage0_45[376], stage0_45[377], stage0_45[378]},
      {stage0_47[24], stage0_47[25], stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29]},
      {stage1_49[4],stage1_48[35],stage1_47[88],stage1_46[124],stage1_45[149]}
   );
   gpc606_5 gpc1739 (
      {stage0_45[379], stage0_45[380], stage0_45[381], stage0_45[382], stage0_45[383], stage0_45[384]},
      {stage0_47[30], stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage1_49[5],stage1_48[36],stage1_47[89],stage1_46[125],stage1_45[150]}
   );
   gpc606_5 gpc1740 (
      {stage0_45[385], stage0_45[386], stage0_45[387], stage0_45[388], stage0_45[389], stage0_45[390]},
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40], stage0_47[41]},
      {stage1_49[6],stage1_48[37],stage1_47[90],stage1_46[126],stage1_45[151]}
   );
   gpc606_5 gpc1741 (
      {stage0_45[391], stage0_45[392], stage0_45[393], stage0_45[394], stage0_45[395], stage0_45[396]},
      {stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45], stage0_47[46], stage0_47[47]},
      {stage1_49[7],stage1_48[38],stage1_47[91],stage1_46[127],stage1_45[152]}
   );
   gpc606_5 gpc1742 (
      {stage0_45[397], stage0_45[398], stage0_45[399], stage0_45[400], stage0_45[401], stage0_45[402]},
      {stage0_47[48], stage0_47[49], stage0_47[50], stage0_47[51], stage0_47[52], stage0_47[53]},
      {stage1_49[8],stage1_48[39],stage1_47[92],stage1_46[128],stage1_45[153]}
   );
   gpc606_5 gpc1743 (
      {stage0_45[403], stage0_45[404], stage0_45[405], stage0_45[406], stage0_45[407], stage0_45[408]},
      {stage0_47[54], stage0_47[55], stage0_47[56], stage0_47[57], stage0_47[58], stage0_47[59]},
      {stage1_49[9],stage1_48[40],stage1_47[93],stage1_46[129],stage1_45[154]}
   );
   gpc606_5 gpc1744 (
      {stage0_45[409], stage0_45[410], stage0_45[411], stage0_45[412], stage0_45[413], stage0_45[414]},
      {stage0_47[60], stage0_47[61], stage0_47[62], stage0_47[63], stage0_47[64], stage0_47[65]},
      {stage1_49[10],stage1_48[41],stage1_47[94],stage1_46[130],stage1_45[155]}
   );
   gpc606_5 gpc1745 (
      {stage0_45[415], stage0_45[416], stage0_45[417], stage0_45[418], stage0_45[419], stage0_45[420]},
      {stage0_47[66], stage0_47[67], stage0_47[68], stage0_47[69], stage0_47[70], stage0_47[71]},
      {stage1_49[11],stage1_48[42],stage1_47[95],stage1_46[131],stage1_45[156]}
   );
   gpc606_5 gpc1746 (
      {stage0_45[421], stage0_45[422], stage0_45[423], stage0_45[424], stage0_45[425], stage0_45[426]},
      {stage0_47[72], stage0_47[73], stage0_47[74], stage0_47[75], stage0_47[76], stage0_47[77]},
      {stage1_49[12],stage1_48[43],stage1_47[96],stage1_46[132],stage1_45[157]}
   );
   gpc606_5 gpc1747 (
      {stage0_45[427], stage0_45[428], stage0_45[429], stage0_45[430], stage0_45[431], stage0_45[432]},
      {stage0_47[78], stage0_47[79], stage0_47[80], stage0_47[81], stage0_47[82], stage0_47[83]},
      {stage1_49[13],stage1_48[44],stage1_47[97],stage1_46[133],stage1_45[158]}
   );
   gpc135_4 gpc1748 (
      {stage0_46[186], stage0_46[187], stage0_46[188], stage0_46[189], stage0_46[190]},
      {stage0_47[84], stage0_47[85], stage0_47[86]},
      {stage0_48[0]},
      {stage1_49[14],stage1_48[45],stage1_47[98],stage1_46[134]}
   );
   gpc135_4 gpc1749 (
      {stage0_46[191], stage0_46[192], stage0_46[193], stage0_46[194], stage0_46[195]},
      {stage0_47[87], stage0_47[88], stage0_47[89]},
      {stage0_48[1]},
      {stage1_49[15],stage1_48[46],stage1_47[99],stage1_46[135]}
   );
   gpc135_4 gpc1750 (
      {stage0_46[196], stage0_46[197], stage0_46[198], stage0_46[199], stage0_46[200]},
      {stage0_47[90], stage0_47[91], stage0_47[92]},
      {stage0_48[2]},
      {stage1_49[16],stage1_48[47],stage1_47[100],stage1_46[136]}
   );
   gpc135_4 gpc1751 (
      {stage0_46[201], stage0_46[202], stage0_46[203], stage0_46[204], stage0_46[205]},
      {stage0_47[93], stage0_47[94], stage0_47[95]},
      {stage0_48[3]},
      {stage1_49[17],stage1_48[48],stage1_47[101],stage1_46[137]}
   );
   gpc135_4 gpc1752 (
      {stage0_46[206], stage0_46[207], stage0_46[208], stage0_46[209], stage0_46[210]},
      {stage0_47[96], stage0_47[97], stage0_47[98]},
      {stage0_48[4]},
      {stage1_49[18],stage1_48[49],stage1_47[102],stage1_46[138]}
   );
   gpc135_4 gpc1753 (
      {stage0_46[211], stage0_46[212], stage0_46[213], stage0_46[214], stage0_46[215]},
      {stage0_47[99], stage0_47[100], stage0_47[101]},
      {stage0_48[5]},
      {stage1_49[19],stage1_48[50],stage1_47[103],stage1_46[139]}
   );
   gpc135_4 gpc1754 (
      {stage0_46[216], stage0_46[217], stage0_46[218], stage0_46[219], stage0_46[220]},
      {stage0_47[102], stage0_47[103], stage0_47[104]},
      {stage0_48[6]},
      {stage1_49[20],stage1_48[51],stage1_47[104],stage1_46[140]}
   );
   gpc135_4 gpc1755 (
      {stage0_46[221], stage0_46[222], stage0_46[223], stage0_46[224], stage0_46[225]},
      {stage0_47[105], stage0_47[106], stage0_47[107]},
      {stage0_48[7]},
      {stage1_49[21],stage1_48[52],stage1_47[105],stage1_46[141]}
   );
   gpc135_4 gpc1756 (
      {stage0_46[226], stage0_46[227], stage0_46[228], stage0_46[229], stage0_46[230]},
      {stage0_47[108], stage0_47[109], stage0_47[110]},
      {stage0_48[8]},
      {stage1_49[22],stage1_48[53],stage1_47[106],stage1_46[142]}
   );
   gpc135_4 gpc1757 (
      {stage0_46[231], stage0_46[232], stage0_46[233], stage0_46[234], stage0_46[235]},
      {stage0_47[111], stage0_47[112], stage0_47[113]},
      {stage0_48[9]},
      {stage1_49[23],stage1_48[54],stage1_47[107],stage1_46[143]}
   );
   gpc615_5 gpc1758 (
      {stage0_46[236], stage0_46[237], stage0_46[238], stage0_46[239], stage0_46[240]},
      {stage0_47[114]},
      {stage0_48[10], stage0_48[11], stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15]},
      {stage1_50[0],stage1_49[24],stage1_48[55],stage1_47[108],stage1_46[144]}
   );
   gpc615_5 gpc1759 (
      {stage0_46[241], stage0_46[242], stage0_46[243], stage0_46[244], stage0_46[245]},
      {stage0_47[115]},
      {stage0_48[16], stage0_48[17], stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21]},
      {stage1_50[1],stage1_49[25],stage1_48[56],stage1_47[109],stage1_46[145]}
   );
   gpc615_5 gpc1760 (
      {stage0_46[246], stage0_46[247], stage0_46[248], stage0_46[249], stage0_46[250]},
      {stage0_47[116]},
      {stage0_48[22], stage0_48[23], stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27]},
      {stage1_50[2],stage1_49[26],stage1_48[57],stage1_47[110],stage1_46[146]}
   );
   gpc615_5 gpc1761 (
      {stage0_46[251], stage0_46[252], stage0_46[253], stage0_46[254], stage0_46[255]},
      {stage0_47[117]},
      {stage0_48[28], stage0_48[29], stage0_48[30], stage0_48[31], stage0_48[32], stage0_48[33]},
      {stage1_50[3],stage1_49[27],stage1_48[58],stage1_47[111],stage1_46[147]}
   );
   gpc615_5 gpc1762 (
      {stage0_46[256], stage0_46[257], stage0_46[258], stage0_46[259], stage0_46[260]},
      {stage0_47[118]},
      {stage0_48[34], stage0_48[35], stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39]},
      {stage1_50[4],stage1_49[28],stage1_48[59],stage1_47[112],stage1_46[148]}
   );
   gpc615_5 gpc1763 (
      {stage0_46[261], stage0_46[262], stage0_46[263], stage0_46[264], stage0_46[265]},
      {stage0_47[119]},
      {stage0_48[40], stage0_48[41], stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45]},
      {stage1_50[5],stage1_49[29],stage1_48[60],stage1_47[113],stage1_46[149]}
   );
   gpc615_5 gpc1764 (
      {stage0_46[266], stage0_46[267], stage0_46[268], stage0_46[269], stage0_46[270]},
      {stage0_47[120]},
      {stage0_48[46], stage0_48[47], stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51]},
      {stage1_50[6],stage1_49[30],stage1_48[61],stage1_47[114],stage1_46[150]}
   );
   gpc615_5 gpc1765 (
      {stage0_46[271], stage0_46[272], stage0_46[273], stage0_46[274], stage0_46[275]},
      {stage0_47[121]},
      {stage0_48[52], stage0_48[53], stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57]},
      {stage1_50[7],stage1_49[31],stage1_48[62],stage1_47[115],stage1_46[151]}
   );
   gpc615_5 gpc1766 (
      {stage0_46[276], stage0_46[277], stage0_46[278], stage0_46[279], stage0_46[280]},
      {stage0_47[122]},
      {stage0_48[58], stage0_48[59], stage0_48[60], stage0_48[61], stage0_48[62], stage0_48[63]},
      {stage1_50[8],stage1_49[32],stage1_48[63],stage1_47[116],stage1_46[152]}
   );
   gpc615_5 gpc1767 (
      {stage0_46[281], stage0_46[282], stage0_46[283], stage0_46[284], stage0_46[285]},
      {stage0_47[123]},
      {stage0_48[64], stage0_48[65], stage0_48[66], stage0_48[67], stage0_48[68], stage0_48[69]},
      {stage1_50[9],stage1_49[33],stage1_48[64],stage1_47[117],stage1_46[153]}
   );
   gpc615_5 gpc1768 (
      {stage0_46[286], stage0_46[287], stage0_46[288], stage0_46[289], stage0_46[290]},
      {stage0_47[124]},
      {stage0_48[70], stage0_48[71], stage0_48[72], stage0_48[73], stage0_48[74], stage0_48[75]},
      {stage1_50[10],stage1_49[34],stage1_48[65],stage1_47[118],stage1_46[154]}
   );
   gpc615_5 gpc1769 (
      {stage0_46[291], stage0_46[292], stage0_46[293], stage0_46[294], stage0_46[295]},
      {stage0_47[125]},
      {stage0_48[76], stage0_48[77], stage0_48[78], stage0_48[79], stage0_48[80], stage0_48[81]},
      {stage1_50[11],stage1_49[35],stage1_48[66],stage1_47[119],stage1_46[155]}
   );
   gpc615_5 gpc1770 (
      {stage0_46[296], stage0_46[297], stage0_46[298], stage0_46[299], stage0_46[300]},
      {stage0_47[126]},
      {stage0_48[82], stage0_48[83], stage0_48[84], stage0_48[85], stage0_48[86], stage0_48[87]},
      {stage1_50[12],stage1_49[36],stage1_48[67],stage1_47[120],stage1_46[156]}
   );
   gpc615_5 gpc1771 (
      {stage0_46[301], stage0_46[302], stage0_46[303], stage0_46[304], stage0_46[305]},
      {stage0_47[127]},
      {stage0_48[88], stage0_48[89], stage0_48[90], stage0_48[91], stage0_48[92], stage0_48[93]},
      {stage1_50[13],stage1_49[37],stage1_48[68],stage1_47[121],stage1_46[157]}
   );
   gpc615_5 gpc1772 (
      {stage0_46[306], stage0_46[307], stage0_46[308], stage0_46[309], stage0_46[310]},
      {stage0_47[128]},
      {stage0_48[94], stage0_48[95], stage0_48[96], stage0_48[97], stage0_48[98], stage0_48[99]},
      {stage1_50[14],stage1_49[38],stage1_48[69],stage1_47[122],stage1_46[158]}
   );
   gpc615_5 gpc1773 (
      {stage0_46[311], stage0_46[312], stage0_46[313], stage0_46[314], stage0_46[315]},
      {stage0_47[129]},
      {stage0_48[100], stage0_48[101], stage0_48[102], stage0_48[103], stage0_48[104], stage0_48[105]},
      {stage1_50[15],stage1_49[39],stage1_48[70],stage1_47[123],stage1_46[159]}
   );
   gpc615_5 gpc1774 (
      {stage0_46[316], stage0_46[317], stage0_46[318], stage0_46[319], stage0_46[320]},
      {stage0_47[130]},
      {stage0_48[106], stage0_48[107], stage0_48[108], stage0_48[109], stage0_48[110], stage0_48[111]},
      {stage1_50[16],stage1_49[40],stage1_48[71],stage1_47[124],stage1_46[160]}
   );
   gpc615_5 gpc1775 (
      {stage0_46[321], stage0_46[322], stage0_46[323], stage0_46[324], stage0_46[325]},
      {stage0_47[131]},
      {stage0_48[112], stage0_48[113], stage0_48[114], stage0_48[115], stage0_48[116], stage0_48[117]},
      {stage1_50[17],stage1_49[41],stage1_48[72],stage1_47[125],stage1_46[161]}
   );
   gpc615_5 gpc1776 (
      {stage0_46[326], stage0_46[327], stage0_46[328], stage0_46[329], stage0_46[330]},
      {stage0_47[132]},
      {stage0_48[118], stage0_48[119], stage0_48[120], stage0_48[121], stage0_48[122], stage0_48[123]},
      {stage1_50[18],stage1_49[42],stage1_48[73],stage1_47[126],stage1_46[162]}
   );
   gpc615_5 gpc1777 (
      {stage0_46[331], stage0_46[332], stage0_46[333], stage0_46[334], stage0_46[335]},
      {stage0_47[133]},
      {stage0_48[124], stage0_48[125], stage0_48[126], stage0_48[127], stage0_48[128], stage0_48[129]},
      {stage1_50[19],stage1_49[43],stage1_48[74],stage1_47[127],stage1_46[163]}
   );
   gpc615_5 gpc1778 (
      {stage0_46[336], stage0_46[337], stage0_46[338], stage0_46[339], stage0_46[340]},
      {stage0_47[134]},
      {stage0_48[130], stage0_48[131], stage0_48[132], stage0_48[133], stage0_48[134], stage0_48[135]},
      {stage1_50[20],stage1_49[44],stage1_48[75],stage1_47[128],stage1_46[164]}
   );
   gpc615_5 gpc1779 (
      {stage0_46[341], stage0_46[342], stage0_46[343], stage0_46[344], stage0_46[345]},
      {stage0_47[135]},
      {stage0_48[136], stage0_48[137], stage0_48[138], stage0_48[139], stage0_48[140], stage0_48[141]},
      {stage1_50[21],stage1_49[45],stage1_48[76],stage1_47[129],stage1_46[165]}
   );
   gpc615_5 gpc1780 (
      {stage0_46[346], stage0_46[347], stage0_46[348], stage0_46[349], stage0_46[350]},
      {stage0_47[136]},
      {stage0_48[142], stage0_48[143], stage0_48[144], stage0_48[145], stage0_48[146], stage0_48[147]},
      {stage1_50[22],stage1_49[46],stage1_48[77],stage1_47[130],stage1_46[166]}
   );
   gpc615_5 gpc1781 (
      {stage0_46[351], stage0_46[352], stage0_46[353], stage0_46[354], stage0_46[355]},
      {stage0_47[137]},
      {stage0_48[148], stage0_48[149], stage0_48[150], stage0_48[151], stage0_48[152], stage0_48[153]},
      {stage1_50[23],stage1_49[47],stage1_48[78],stage1_47[131],stage1_46[167]}
   );
   gpc615_5 gpc1782 (
      {stage0_47[138], stage0_47[139], stage0_47[140], stage0_47[141], stage0_47[142]},
      {stage0_48[154]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[24],stage1_49[48],stage1_48[79],stage1_47[132]}
   );
   gpc615_5 gpc1783 (
      {stage0_47[143], stage0_47[144], stage0_47[145], stage0_47[146], stage0_47[147]},
      {stage0_48[155]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[25],stage1_49[49],stage1_48[80],stage1_47[133]}
   );
   gpc615_5 gpc1784 (
      {stage0_47[148], stage0_47[149], stage0_47[150], stage0_47[151], stage0_47[152]},
      {stage0_48[156]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[26],stage1_49[50],stage1_48[81],stage1_47[134]}
   );
   gpc615_5 gpc1785 (
      {stage0_47[153], stage0_47[154], stage0_47[155], stage0_47[156], stage0_47[157]},
      {stage0_48[157]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[27],stage1_49[51],stage1_48[82],stage1_47[135]}
   );
   gpc615_5 gpc1786 (
      {stage0_47[158], stage0_47[159], stage0_47[160], stage0_47[161], stage0_47[162]},
      {stage0_48[158]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[28],stage1_49[52],stage1_48[83],stage1_47[136]}
   );
   gpc615_5 gpc1787 (
      {stage0_47[163], stage0_47[164], stage0_47[165], stage0_47[166], stage0_47[167]},
      {stage0_48[159]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[29],stage1_49[53],stage1_48[84],stage1_47[137]}
   );
   gpc615_5 gpc1788 (
      {stage0_47[168], stage0_47[169], stage0_47[170], stage0_47[171], stage0_47[172]},
      {stage0_48[160]},
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage1_51[6],stage1_50[30],stage1_49[54],stage1_48[85],stage1_47[138]}
   );
   gpc615_5 gpc1789 (
      {stage0_47[173], stage0_47[174], stage0_47[175], stage0_47[176], stage0_47[177]},
      {stage0_48[161]},
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46], stage0_49[47]},
      {stage1_51[7],stage1_50[31],stage1_49[55],stage1_48[86],stage1_47[139]}
   );
   gpc615_5 gpc1790 (
      {stage0_47[178], stage0_47[179], stage0_47[180], stage0_47[181], stage0_47[182]},
      {stage0_48[162]},
      {stage0_49[48], stage0_49[49], stage0_49[50], stage0_49[51], stage0_49[52], stage0_49[53]},
      {stage1_51[8],stage1_50[32],stage1_49[56],stage1_48[87],stage1_47[140]}
   );
   gpc615_5 gpc1791 (
      {stage0_47[183], stage0_47[184], stage0_47[185], stage0_47[186], stage0_47[187]},
      {stage0_48[163]},
      {stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58], stage0_49[59]},
      {stage1_51[9],stage1_50[33],stage1_49[57],stage1_48[88],stage1_47[141]}
   );
   gpc615_5 gpc1792 (
      {stage0_47[188], stage0_47[189], stage0_47[190], stage0_47[191], stage0_47[192]},
      {stage0_48[164]},
      {stage0_49[60], stage0_49[61], stage0_49[62], stage0_49[63], stage0_49[64], stage0_49[65]},
      {stage1_51[10],stage1_50[34],stage1_49[58],stage1_48[89],stage1_47[142]}
   );
   gpc615_5 gpc1793 (
      {stage0_47[193], stage0_47[194], stage0_47[195], stage0_47[196], stage0_47[197]},
      {stage0_48[165]},
      {stage0_49[66], stage0_49[67], stage0_49[68], stage0_49[69], stage0_49[70], stage0_49[71]},
      {stage1_51[11],stage1_50[35],stage1_49[59],stage1_48[90],stage1_47[143]}
   );
   gpc615_5 gpc1794 (
      {stage0_47[198], stage0_47[199], stage0_47[200], stage0_47[201], stage0_47[202]},
      {stage0_48[166]},
      {stage0_49[72], stage0_49[73], stage0_49[74], stage0_49[75], stage0_49[76], stage0_49[77]},
      {stage1_51[12],stage1_50[36],stage1_49[60],stage1_48[91],stage1_47[144]}
   );
   gpc615_5 gpc1795 (
      {stage0_47[203], stage0_47[204], stage0_47[205], stage0_47[206], stage0_47[207]},
      {stage0_48[167]},
      {stage0_49[78], stage0_49[79], stage0_49[80], stage0_49[81], stage0_49[82], stage0_49[83]},
      {stage1_51[13],stage1_50[37],stage1_49[61],stage1_48[92],stage1_47[145]}
   );
   gpc615_5 gpc1796 (
      {stage0_47[208], stage0_47[209], stage0_47[210], stage0_47[211], stage0_47[212]},
      {stage0_48[168]},
      {stage0_49[84], stage0_49[85], stage0_49[86], stage0_49[87], stage0_49[88], stage0_49[89]},
      {stage1_51[14],stage1_50[38],stage1_49[62],stage1_48[93],stage1_47[146]}
   );
   gpc615_5 gpc1797 (
      {stage0_47[213], stage0_47[214], stage0_47[215], stage0_47[216], stage0_47[217]},
      {stage0_48[169]},
      {stage0_49[90], stage0_49[91], stage0_49[92], stage0_49[93], stage0_49[94], stage0_49[95]},
      {stage1_51[15],stage1_50[39],stage1_49[63],stage1_48[94],stage1_47[147]}
   );
   gpc615_5 gpc1798 (
      {stage0_47[218], stage0_47[219], stage0_47[220], stage0_47[221], stage0_47[222]},
      {stage0_48[170]},
      {stage0_49[96], stage0_49[97], stage0_49[98], stage0_49[99], stage0_49[100], stage0_49[101]},
      {stage1_51[16],stage1_50[40],stage1_49[64],stage1_48[95],stage1_47[148]}
   );
   gpc615_5 gpc1799 (
      {stage0_47[223], stage0_47[224], stage0_47[225], stage0_47[226], stage0_47[227]},
      {stage0_48[171]},
      {stage0_49[102], stage0_49[103], stage0_49[104], stage0_49[105], stage0_49[106], stage0_49[107]},
      {stage1_51[17],stage1_50[41],stage1_49[65],stage1_48[96],stage1_47[149]}
   );
   gpc615_5 gpc1800 (
      {stage0_47[228], stage0_47[229], stage0_47[230], stage0_47[231], stage0_47[232]},
      {stage0_48[172]},
      {stage0_49[108], stage0_49[109], stage0_49[110], stage0_49[111], stage0_49[112], stage0_49[113]},
      {stage1_51[18],stage1_50[42],stage1_49[66],stage1_48[97],stage1_47[150]}
   );
   gpc615_5 gpc1801 (
      {stage0_47[233], stage0_47[234], stage0_47[235], stage0_47[236], stage0_47[237]},
      {stage0_48[173]},
      {stage0_49[114], stage0_49[115], stage0_49[116], stage0_49[117], stage0_49[118], stage0_49[119]},
      {stage1_51[19],stage1_50[43],stage1_49[67],stage1_48[98],stage1_47[151]}
   );
   gpc615_5 gpc1802 (
      {stage0_47[238], stage0_47[239], stage0_47[240], stage0_47[241], stage0_47[242]},
      {stage0_48[174]},
      {stage0_49[120], stage0_49[121], stage0_49[122], stage0_49[123], stage0_49[124], stage0_49[125]},
      {stage1_51[20],stage1_50[44],stage1_49[68],stage1_48[99],stage1_47[152]}
   );
   gpc615_5 gpc1803 (
      {stage0_47[243], stage0_47[244], stage0_47[245], stage0_47[246], stage0_47[247]},
      {stage0_48[175]},
      {stage0_49[126], stage0_49[127], stage0_49[128], stage0_49[129], stage0_49[130], stage0_49[131]},
      {stage1_51[21],stage1_50[45],stage1_49[69],stage1_48[100],stage1_47[153]}
   );
   gpc615_5 gpc1804 (
      {stage0_47[248], stage0_47[249], stage0_47[250], stage0_47[251], stage0_47[252]},
      {stage0_48[176]},
      {stage0_49[132], stage0_49[133], stage0_49[134], stage0_49[135], stage0_49[136], stage0_49[137]},
      {stage1_51[22],stage1_50[46],stage1_49[70],stage1_48[101],stage1_47[154]}
   );
   gpc615_5 gpc1805 (
      {stage0_47[253], stage0_47[254], stage0_47[255], stage0_47[256], stage0_47[257]},
      {stage0_48[177]},
      {stage0_49[138], stage0_49[139], stage0_49[140], stage0_49[141], stage0_49[142], stage0_49[143]},
      {stage1_51[23],stage1_50[47],stage1_49[71],stage1_48[102],stage1_47[155]}
   );
   gpc615_5 gpc1806 (
      {stage0_47[258], stage0_47[259], stage0_47[260], stage0_47[261], stage0_47[262]},
      {stage0_48[178]},
      {stage0_49[144], stage0_49[145], stage0_49[146], stage0_49[147], stage0_49[148], stage0_49[149]},
      {stage1_51[24],stage1_50[48],stage1_49[72],stage1_48[103],stage1_47[156]}
   );
   gpc615_5 gpc1807 (
      {stage0_47[263], stage0_47[264], stage0_47[265], stage0_47[266], stage0_47[267]},
      {stage0_48[179]},
      {stage0_49[150], stage0_49[151], stage0_49[152], stage0_49[153], stage0_49[154], stage0_49[155]},
      {stage1_51[25],stage1_50[49],stage1_49[73],stage1_48[104],stage1_47[157]}
   );
   gpc615_5 gpc1808 (
      {stage0_47[268], stage0_47[269], stage0_47[270], stage0_47[271], stage0_47[272]},
      {stage0_48[180]},
      {stage0_49[156], stage0_49[157], stage0_49[158], stage0_49[159], stage0_49[160], stage0_49[161]},
      {stage1_51[26],stage1_50[50],stage1_49[74],stage1_48[105],stage1_47[158]}
   );
   gpc615_5 gpc1809 (
      {stage0_47[273], stage0_47[274], stage0_47[275], stage0_47[276], stage0_47[277]},
      {stage0_48[181]},
      {stage0_49[162], stage0_49[163], stage0_49[164], stage0_49[165], stage0_49[166], stage0_49[167]},
      {stage1_51[27],stage1_50[51],stage1_49[75],stage1_48[106],stage1_47[159]}
   );
   gpc615_5 gpc1810 (
      {stage0_47[278], stage0_47[279], stage0_47[280], stage0_47[281], stage0_47[282]},
      {stage0_48[182]},
      {stage0_49[168], stage0_49[169], stage0_49[170], stage0_49[171], stage0_49[172], stage0_49[173]},
      {stage1_51[28],stage1_50[52],stage1_49[76],stage1_48[107],stage1_47[160]}
   );
   gpc615_5 gpc1811 (
      {stage0_47[283], stage0_47[284], stage0_47[285], stage0_47[286], stage0_47[287]},
      {stage0_48[183]},
      {stage0_49[174], stage0_49[175], stage0_49[176], stage0_49[177], stage0_49[178], stage0_49[179]},
      {stage1_51[29],stage1_50[53],stage1_49[77],stage1_48[108],stage1_47[161]}
   );
   gpc615_5 gpc1812 (
      {stage0_47[288], stage0_47[289], stage0_47[290], stage0_47[291], stage0_47[292]},
      {stage0_48[184]},
      {stage0_49[180], stage0_49[181], stage0_49[182], stage0_49[183], stage0_49[184], stage0_49[185]},
      {stage1_51[30],stage1_50[54],stage1_49[78],stage1_48[109],stage1_47[162]}
   );
   gpc615_5 gpc1813 (
      {stage0_47[293], stage0_47[294], stage0_47[295], stage0_47[296], stage0_47[297]},
      {stage0_48[185]},
      {stage0_49[186], stage0_49[187], stage0_49[188], stage0_49[189], stage0_49[190], stage0_49[191]},
      {stage1_51[31],stage1_50[55],stage1_49[79],stage1_48[110],stage1_47[163]}
   );
   gpc615_5 gpc1814 (
      {stage0_47[298], stage0_47[299], stage0_47[300], stage0_47[301], stage0_47[302]},
      {stage0_48[186]},
      {stage0_49[192], stage0_49[193], stage0_49[194], stage0_49[195], stage0_49[196], stage0_49[197]},
      {stage1_51[32],stage1_50[56],stage1_49[80],stage1_48[111],stage1_47[164]}
   );
   gpc615_5 gpc1815 (
      {stage0_47[303], stage0_47[304], stage0_47[305], stage0_47[306], stage0_47[307]},
      {stage0_48[187]},
      {stage0_49[198], stage0_49[199], stage0_49[200], stage0_49[201], stage0_49[202], stage0_49[203]},
      {stage1_51[33],stage1_50[57],stage1_49[81],stage1_48[112],stage1_47[165]}
   );
   gpc615_5 gpc1816 (
      {stage0_47[308], stage0_47[309], stage0_47[310], stage0_47[311], stage0_47[312]},
      {stage0_48[188]},
      {stage0_49[204], stage0_49[205], stage0_49[206], stage0_49[207], stage0_49[208], stage0_49[209]},
      {stage1_51[34],stage1_50[58],stage1_49[82],stage1_48[113],stage1_47[166]}
   );
   gpc615_5 gpc1817 (
      {stage0_47[313], stage0_47[314], stage0_47[315], stage0_47[316], stage0_47[317]},
      {stage0_48[189]},
      {stage0_49[210], stage0_49[211], stage0_49[212], stage0_49[213], stage0_49[214], stage0_49[215]},
      {stage1_51[35],stage1_50[59],stage1_49[83],stage1_48[114],stage1_47[167]}
   );
   gpc615_5 gpc1818 (
      {stage0_47[318], stage0_47[319], stage0_47[320], stage0_47[321], stage0_47[322]},
      {stage0_48[190]},
      {stage0_49[216], stage0_49[217], stage0_49[218], stage0_49[219], stage0_49[220], stage0_49[221]},
      {stage1_51[36],stage1_50[60],stage1_49[84],stage1_48[115],stage1_47[168]}
   );
   gpc615_5 gpc1819 (
      {stage0_47[323], stage0_47[324], stage0_47[325], stage0_47[326], stage0_47[327]},
      {stage0_48[191]},
      {stage0_49[222], stage0_49[223], stage0_49[224], stage0_49[225], stage0_49[226], stage0_49[227]},
      {stage1_51[37],stage1_50[61],stage1_49[85],stage1_48[116],stage1_47[169]}
   );
   gpc615_5 gpc1820 (
      {stage0_47[328], stage0_47[329], stage0_47[330], stage0_47[331], stage0_47[332]},
      {stage0_48[192]},
      {stage0_49[228], stage0_49[229], stage0_49[230], stage0_49[231], stage0_49[232], stage0_49[233]},
      {stage1_51[38],stage1_50[62],stage1_49[86],stage1_48[117],stage1_47[170]}
   );
   gpc615_5 gpc1821 (
      {stage0_47[333], stage0_47[334], stage0_47[335], stage0_47[336], stage0_47[337]},
      {stage0_48[193]},
      {stage0_49[234], stage0_49[235], stage0_49[236], stage0_49[237], stage0_49[238], stage0_49[239]},
      {stage1_51[39],stage1_50[63],stage1_49[87],stage1_48[118],stage1_47[171]}
   );
   gpc615_5 gpc1822 (
      {stage0_47[338], stage0_47[339], stage0_47[340], stage0_47[341], stage0_47[342]},
      {stage0_48[194]},
      {stage0_49[240], stage0_49[241], stage0_49[242], stage0_49[243], stage0_49[244], stage0_49[245]},
      {stage1_51[40],stage1_50[64],stage1_49[88],stage1_48[119],stage1_47[172]}
   );
   gpc615_5 gpc1823 (
      {stage0_47[343], stage0_47[344], stage0_47[345], stage0_47[346], stage0_47[347]},
      {stage0_48[195]},
      {stage0_49[246], stage0_49[247], stage0_49[248], stage0_49[249], stage0_49[250], stage0_49[251]},
      {stage1_51[41],stage1_50[65],stage1_49[89],stage1_48[120],stage1_47[173]}
   );
   gpc615_5 gpc1824 (
      {stage0_47[348], stage0_47[349], stage0_47[350], stage0_47[351], stage0_47[352]},
      {stage0_48[196]},
      {stage0_49[252], stage0_49[253], stage0_49[254], stage0_49[255], stage0_49[256], stage0_49[257]},
      {stage1_51[42],stage1_50[66],stage1_49[90],stage1_48[121],stage1_47[174]}
   );
   gpc615_5 gpc1825 (
      {stage0_47[353], stage0_47[354], stage0_47[355], stage0_47[356], stage0_47[357]},
      {stage0_48[197]},
      {stage0_49[258], stage0_49[259], stage0_49[260], stage0_49[261], stage0_49[262], stage0_49[263]},
      {stage1_51[43],stage1_50[67],stage1_49[91],stage1_48[122],stage1_47[175]}
   );
   gpc615_5 gpc1826 (
      {stage0_47[358], stage0_47[359], stage0_47[360], stage0_47[361], stage0_47[362]},
      {stage0_48[198]},
      {stage0_49[264], stage0_49[265], stage0_49[266], stage0_49[267], stage0_49[268], stage0_49[269]},
      {stage1_51[44],stage1_50[68],stage1_49[92],stage1_48[123],stage1_47[176]}
   );
   gpc615_5 gpc1827 (
      {stage0_47[363], stage0_47[364], stage0_47[365], stage0_47[366], stage0_47[367]},
      {stage0_48[199]},
      {stage0_49[270], stage0_49[271], stage0_49[272], stage0_49[273], stage0_49[274], stage0_49[275]},
      {stage1_51[45],stage1_50[69],stage1_49[93],stage1_48[124],stage1_47[177]}
   );
   gpc615_5 gpc1828 (
      {stage0_47[368], stage0_47[369], stage0_47[370], stage0_47[371], stage0_47[372]},
      {stage0_48[200]},
      {stage0_49[276], stage0_49[277], stage0_49[278], stage0_49[279], stage0_49[280], stage0_49[281]},
      {stage1_51[46],stage1_50[70],stage1_49[94],stage1_48[125],stage1_47[178]}
   );
   gpc615_5 gpc1829 (
      {stage0_47[373], stage0_47[374], stage0_47[375], stage0_47[376], stage0_47[377]},
      {stage0_48[201]},
      {stage0_49[282], stage0_49[283], stage0_49[284], stage0_49[285], stage0_49[286], stage0_49[287]},
      {stage1_51[47],stage1_50[71],stage1_49[95],stage1_48[126],stage1_47[179]}
   );
   gpc615_5 gpc1830 (
      {stage0_47[378], stage0_47[379], stage0_47[380], stage0_47[381], stage0_47[382]},
      {stage0_48[202]},
      {stage0_49[288], stage0_49[289], stage0_49[290], stage0_49[291], stage0_49[292], stage0_49[293]},
      {stage1_51[48],stage1_50[72],stage1_49[96],stage1_48[127],stage1_47[180]}
   );
   gpc615_5 gpc1831 (
      {stage0_47[383], stage0_47[384], stage0_47[385], stage0_47[386], stage0_47[387]},
      {stage0_48[203]},
      {stage0_49[294], stage0_49[295], stage0_49[296], stage0_49[297], stage0_49[298], stage0_49[299]},
      {stage1_51[49],stage1_50[73],stage1_49[97],stage1_48[128],stage1_47[181]}
   );
   gpc615_5 gpc1832 (
      {stage0_47[388], stage0_47[389], stage0_47[390], stage0_47[391], stage0_47[392]},
      {stage0_48[204]},
      {stage0_49[300], stage0_49[301], stage0_49[302], stage0_49[303], stage0_49[304], stage0_49[305]},
      {stage1_51[50],stage1_50[74],stage1_49[98],stage1_48[129],stage1_47[182]}
   );
   gpc615_5 gpc1833 (
      {stage0_47[393], stage0_47[394], stage0_47[395], stage0_47[396], stage0_47[397]},
      {stage0_48[205]},
      {stage0_49[306], stage0_49[307], stage0_49[308], stage0_49[309], stage0_49[310], stage0_49[311]},
      {stage1_51[51],stage1_50[75],stage1_49[99],stage1_48[130],stage1_47[183]}
   );
   gpc615_5 gpc1834 (
      {stage0_47[398], stage0_47[399], stage0_47[400], stage0_47[401], stage0_47[402]},
      {stage0_48[206]},
      {stage0_49[312], stage0_49[313], stage0_49[314], stage0_49[315], stage0_49[316], stage0_49[317]},
      {stage1_51[52],stage1_50[76],stage1_49[100],stage1_48[131],stage1_47[184]}
   );
   gpc615_5 gpc1835 (
      {stage0_47[403], stage0_47[404], stage0_47[405], stage0_47[406], stage0_47[407]},
      {stage0_48[207]},
      {stage0_49[318], stage0_49[319], stage0_49[320], stage0_49[321], stage0_49[322], stage0_49[323]},
      {stage1_51[53],stage1_50[77],stage1_49[101],stage1_48[132],stage1_47[185]}
   );
   gpc615_5 gpc1836 (
      {stage0_47[408], stage0_47[409], stage0_47[410], stage0_47[411], stage0_47[412]},
      {stage0_48[208]},
      {stage0_49[324], stage0_49[325], stage0_49[326], stage0_49[327], stage0_49[328], stage0_49[329]},
      {stage1_51[54],stage1_50[78],stage1_49[102],stage1_48[133],stage1_47[186]}
   );
   gpc615_5 gpc1837 (
      {stage0_47[413], stage0_47[414], stage0_47[415], stage0_47[416], stage0_47[417]},
      {stage0_48[209]},
      {stage0_49[330], stage0_49[331], stage0_49[332], stage0_49[333], stage0_49[334], stage0_49[335]},
      {stage1_51[55],stage1_50[79],stage1_49[103],stage1_48[134],stage1_47[187]}
   );
   gpc615_5 gpc1838 (
      {stage0_47[418], stage0_47[419], stage0_47[420], stage0_47[421], stage0_47[422]},
      {stage0_48[210]},
      {stage0_49[336], stage0_49[337], stage0_49[338], stage0_49[339], stage0_49[340], stage0_49[341]},
      {stage1_51[56],stage1_50[80],stage1_49[104],stage1_48[135],stage1_47[188]}
   );
   gpc615_5 gpc1839 (
      {stage0_47[423], stage0_47[424], stage0_47[425], stage0_47[426], stage0_47[427]},
      {stage0_48[211]},
      {stage0_49[342], stage0_49[343], stage0_49[344], stage0_49[345], stage0_49[346], stage0_49[347]},
      {stage1_51[57],stage1_50[81],stage1_49[105],stage1_48[136],stage1_47[189]}
   );
   gpc615_5 gpc1840 (
      {stage0_47[428], stage0_47[429], stage0_47[430], stage0_47[431], stage0_47[432]},
      {stage0_48[212]},
      {stage0_49[348], stage0_49[349], stage0_49[350], stage0_49[351], stage0_49[352], stage0_49[353]},
      {stage1_51[58],stage1_50[82],stage1_49[106],stage1_48[137],stage1_47[190]}
   );
   gpc615_5 gpc1841 (
      {stage0_47[433], stage0_47[434], stage0_47[435], stage0_47[436], stage0_47[437]},
      {stage0_48[213]},
      {stage0_49[354], stage0_49[355], stage0_49[356], stage0_49[357], stage0_49[358], stage0_49[359]},
      {stage1_51[59],stage1_50[83],stage1_49[107],stage1_48[138],stage1_47[191]}
   );
   gpc615_5 gpc1842 (
      {stage0_47[438], stage0_47[439], stage0_47[440], stage0_47[441], stage0_47[442]},
      {stage0_48[214]},
      {stage0_49[360], stage0_49[361], stage0_49[362], stage0_49[363], stage0_49[364], stage0_49[365]},
      {stage1_51[60],stage1_50[84],stage1_49[108],stage1_48[139],stage1_47[192]}
   );
   gpc606_5 gpc1843 (
      {stage0_48[215], stage0_48[216], stage0_48[217], stage0_48[218], stage0_48[219], stage0_48[220]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[61],stage1_50[85],stage1_49[109],stage1_48[140]}
   );
   gpc606_5 gpc1844 (
      {stage0_48[221], stage0_48[222], stage0_48[223], stage0_48[224], stage0_48[225], stage0_48[226]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[62],stage1_50[86],stage1_49[110],stage1_48[141]}
   );
   gpc606_5 gpc1845 (
      {stage0_48[227], stage0_48[228], stage0_48[229], stage0_48[230], stage0_48[231], stage0_48[232]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[63],stage1_50[87],stage1_49[111],stage1_48[142]}
   );
   gpc606_5 gpc1846 (
      {stage0_48[233], stage0_48[234], stage0_48[235], stage0_48[236], stage0_48[237], stage0_48[238]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[64],stage1_50[88],stage1_49[112],stage1_48[143]}
   );
   gpc606_5 gpc1847 (
      {stage0_48[239], stage0_48[240], stage0_48[241], stage0_48[242], stage0_48[243], stage0_48[244]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[65],stage1_50[89],stage1_49[113],stage1_48[144]}
   );
   gpc606_5 gpc1848 (
      {stage0_48[245], stage0_48[246], stage0_48[247], stage0_48[248], stage0_48[249], stage0_48[250]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[66],stage1_50[90],stage1_49[114],stage1_48[145]}
   );
   gpc606_5 gpc1849 (
      {stage0_48[251], stage0_48[252], stage0_48[253], stage0_48[254], stage0_48[255], stage0_48[256]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[67],stage1_50[91],stage1_49[115],stage1_48[146]}
   );
   gpc606_5 gpc1850 (
      {stage0_48[257], stage0_48[258], stage0_48[259], stage0_48[260], stage0_48[261], stage0_48[262]},
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46], stage0_50[47]},
      {stage1_52[7],stage1_51[68],stage1_50[92],stage1_49[116],stage1_48[147]}
   );
   gpc606_5 gpc1851 (
      {stage0_48[263], stage0_48[264], stage0_48[265], stage0_48[266], stage0_48[267], stage0_48[268]},
      {stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51], stage0_50[52], stage0_50[53]},
      {stage1_52[8],stage1_51[69],stage1_50[93],stage1_49[117],stage1_48[148]}
   );
   gpc606_5 gpc1852 (
      {stage0_48[269], stage0_48[270], stage0_48[271], stage0_48[272], stage0_48[273], stage0_48[274]},
      {stage0_50[54], stage0_50[55], stage0_50[56], stage0_50[57], stage0_50[58], stage0_50[59]},
      {stage1_52[9],stage1_51[70],stage1_50[94],stage1_49[118],stage1_48[149]}
   );
   gpc606_5 gpc1853 (
      {stage0_48[275], stage0_48[276], stage0_48[277], stage0_48[278], stage0_48[279], stage0_48[280]},
      {stage0_50[60], stage0_50[61], stage0_50[62], stage0_50[63], stage0_50[64], stage0_50[65]},
      {stage1_52[10],stage1_51[71],stage1_50[95],stage1_49[119],stage1_48[150]}
   );
   gpc606_5 gpc1854 (
      {stage0_48[281], stage0_48[282], stage0_48[283], stage0_48[284], stage0_48[285], stage0_48[286]},
      {stage0_50[66], stage0_50[67], stage0_50[68], stage0_50[69], stage0_50[70], stage0_50[71]},
      {stage1_52[11],stage1_51[72],stage1_50[96],stage1_49[120],stage1_48[151]}
   );
   gpc606_5 gpc1855 (
      {stage0_48[287], stage0_48[288], stage0_48[289], stage0_48[290], stage0_48[291], stage0_48[292]},
      {stage0_50[72], stage0_50[73], stage0_50[74], stage0_50[75], stage0_50[76], stage0_50[77]},
      {stage1_52[12],stage1_51[73],stage1_50[97],stage1_49[121],stage1_48[152]}
   );
   gpc615_5 gpc1856 (
      {stage0_48[293], stage0_48[294], stage0_48[295], stage0_48[296], stage0_48[297]},
      {stage0_49[366]},
      {stage0_50[78], stage0_50[79], stage0_50[80], stage0_50[81], stage0_50[82], stage0_50[83]},
      {stage1_52[13],stage1_51[74],stage1_50[98],stage1_49[122],stage1_48[153]}
   );
   gpc615_5 gpc1857 (
      {stage0_48[298], stage0_48[299], stage0_48[300], stage0_48[301], stage0_48[302]},
      {stage0_49[367]},
      {stage0_50[84], stage0_50[85], stage0_50[86], stage0_50[87], stage0_50[88], stage0_50[89]},
      {stage1_52[14],stage1_51[75],stage1_50[99],stage1_49[123],stage1_48[154]}
   );
   gpc615_5 gpc1858 (
      {stage0_48[303], stage0_48[304], stage0_48[305], stage0_48[306], stage0_48[307]},
      {stage0_49[368]},
      {stage0_50[90], stage0_50[91], stage0_50[92], stage0_50[93], stage0_50[94], stage0_50[95]},
      {stage1_52[15],stage1_51[76],stage1_50[100],stage1_49[124],stage1_48[155]}
   );
   gpc615_5 gpc1859 (
      {stage0_48[308], stage0_48[309], stage0_48[310], stage0_48[311], stage0_48[312]},
      {stage0_49[369]},
      {stage0_50[96], stage0_50[97], stage0_50[98], stage0_50[99], stage0_50[100], stage0_50[101]},
      {stage1_52[16],stage1_51[77],stage1_50[101],stage1_49[125],stage1_48[156]}
   );
   gpc615_5 gpc1860 (
      {stage0_48[313], stage0_48[314], stage0_48[315], stage0_48[316], stage0_48[317]},
      {stage0_49[370]},
      {stage0_50[102], stage0_50[103], stage0_50[104], stage0_50[105], stage0_50[106], stage0_50[107]},
      {stage1_52[17],stage1_51[78],stage1_50[102],stage1_49[126],stage1_48[157]}
   );
   gpc615_5 gpc1861 (
      {stage0_48[318], stage0_48[319], stage0_48[320], stage0_48[321], stage0_48[322]},
      {stage0_49[371]},
      {stage0_50[108], stage0_50[109], stage0_50[110], stage0_50[111], stage0_50[112], stage0_50[113]},
      {stage1_52[18],stage1_51[79],stage1_50[103],stage1_49[127],stage1_48[158]}
   );
   gpc615_5 gpc1862 (
      {stage0_48[323], stage0_48[324], stage0_48[325], stage0_48[326], stage0_48[327]},
      {stage0_49[372]},
      {stage0_50[114], stage0_50[115], stage0_50[116], stage0_50[117], stage0_50[118], stage0_50[119]},
      {stage1_52[19],stage1_51[80],stage1_50[104],stage1_49[128],stage1_48[159]}
   );
   gpc615_5 gpc1863 (
      {stage0_48[328], stage0_48[329], stage0_48[330], stage0_48[331], stage0_48[332]},
      {stage0_49[373]},
      {stage0_50[120], stage0_50[121], stage0_50[122], stage0_50[123], stage0_50[124], stage0_50[125]},
      {stage1_52[20],stage1_51[81],stage1_50[105],stage1_49[129],stage1_48[160]}
   );
   gpc615_5 gpc1864 (
      {stage0_48[333], stage0_48[334], stage0_48[335], stage0_48[336], stage0_48[337]},
      {stage0_49[374]},
      {stage0_50[126], stage0_50[127], stage0_50[128], stage0_50[129], stage0_50[130], stage0_50[131]},
      {stage1_52[21],stage1_51[82],stage1_50[106],stage1_49[130],stage1_48[161]}
   );
   gpc615_5 gpc1865 (
      {stage0_48[338], stage0_48[339], stage0_48[340], stage0_48[341], stage0_48[342]},
      {stage0_49[375]},
      {stage0_50[132], stage0_50[133], stage0_50[134], stage0_50[135], stage0_50[136], stage0_50[137]},
      {stage1_52[22],stage1_51[83],stage1_50[107],stage1_49[131],stage1_48[162]}
   );
   gpc615_5 gpc1866 (
      {stage0_48[343], stage0_48[344], stage0_48[345], stage0_48[346], stage0_48[347]},
      {stage0_49[376]},
      {stage0_50[138], stage0_50[139], stage0_50[140], stage0_50[141], stage0_50[142], stage0_50[143]},
      {stage1_52[23],stage1_51[84],stage1_50[108],stage1_49[132],stage1_48[163]}
   );
   gpc615_5 gpc1867 (
      {stage0_48[348], stage0_48[349], stage0_48[350], stage0_48[351], stage0_48[352]},
      {stage0_49[377]},
      {stage0_50[144], stage0_50[145], stage0_50[146], stage0_50[147], stage0_50[148], stage0_50[149]},
      {stage1_52[24],stage1_51[85],stage1_50[109],stage1_49[133],stage1_48[164]}
   );
   gpc615_5 gpc1868 (
      {stage0_48[353], stage0_48[354], stage0_48[355], stage0_48[356], stage0_48[357]},
      {stage0_49[378]},
      {stage0_50[150], stage0_50[151], stage0_50[152], stage0_50[153], stage0_50[154], stage0_50[155]},
      {stage1_52[25],stage1_51[86],stage1_50[110],stage1_49[134],stage1_48[165]}
   );
   gpc615_5 gpc1869 (
      {stage0_48[358], stage0_48[359], stage0_48[360], stage0_48[361], stage0_48[362]},
      {stage0_49[379]},
      {stage0_50[156], stage0_50[157], stage0_50[158], stage0_50[159], stage0_50[160], stage0_50[161]},
      {stage1_52[26],stage1_51[87],stage1_50[111],stage1_49[135],stage1_48[166]}
   );
   gpc615_5 gpc1870 (
      {stage0_48[363], stage0_48[364], stage0_48[365], stage0_48[366], stage0_48[367]},
      {stage0_49[380]},
      {stage0_50[162], stage0_50[163], stage0_50[164], stage0_50[165], stage0_50[166], stage0_50[167]},
      {stage1_52[27],stage1_51[88],stage1_50[112],stage1_49[136],stage1_48[167]}
   );
   gpc615_5 gpc1871 (
      {stage0_48[368], stage0_48[369], stage0_48[370], stage0_48[371], stage0_48[372]},
      {stage0_49[381]},
      {stage0_50[168], stage0_50[169], stage0_50[170], stage0_50[171], stage0_50[172], stage0_50[173]},
      {stage1_52[28],stage1_51[89],stage1_50[113],stage1_49[137],stage1_48[168]}
   );
   gpc615_5 gpc1872 (
      {stage0_48[373], stage0_48[374], stage0_48[375], stage0_48[376], stage0_48[377]},
      {stage0_49[382]},
      {stage0_50[174], stage0_50[175], stage0_50[176], stage0_50[177], stage0_50[178], stage0_50[179]},
      {stage1_52[29],stage1_51[90],stage1_50[114],stage1_49[138],stage1_48[169]}
   );
   gpc615_5 gpc1873 (
      {stage0_48[378], stage0_48[379], stage0_48[380], stage0_48[381], stage0_48[382]},
      {stage0_49[383]},
      {stage0_50[180], stage0_50[181], stage0_50[182], stage0_50[183], stage0_50[184], stage0_50[185]},
      {stage1_52[30],stage1_51[91],stage1_50[115],stage1_49[139],stage1_48[170]}
   );
   gpc615_5 gpc1874 (
      {stage0_48[383], stage0_48[384], stage0_48[385], stage0_48[386], stage0_48[387]},
      {stage0_49[384]},
      {stage0_50[186], stage0_50[187], stage0_50[188], stage0_50[189], stage0_50[190], stage0_50[191]},
      {stage1_52[31],stage1_51[92],stage1_50[116],stage1_49[140],stage1_48[171]}
   );
   gpc615_5 gpc1875 (
      {stage0_48[388], stage0_48[389], stage0_48[390], stage0_48[391], stage0_48[392]},
      {stage0_49[385]},
      {stage0_50[192], stage0_50[193], stage0_50[194], stage0_50[195], stage0_50[196], stage0_50[197]},
      {stage1_52[32],stage1_51[93],stage1_50[117],stage1_49[141],stage1_48[172]}
   );
   gpc615_5 gpc1876 (
      {stage0_48[393], stage0_48[394], stage0_48[395], stage0_48[396], stage0_48[397]},
      {stage0_49[386]},
      {stage0_50[198], stage0_50[199], stage0_50[200], stage0_50[201], stage0_50[202], stage0_50[203]},
      {stage1_52[33],stage1_51[94],stage1_50[118],stage1_49[142],stage1_48[173]}
   );
   gpc615_5 gpc1877 (
      {stage0_48[398], stage0_48[399], stage0_48[400], stage0_48[401], stage0_48[402]},
      {stage0_49[387]},
      {stage0_50[204], stage0_50[205], stage0_50[206], stage0_50[207], stage0_50[208], stage0_50[209]},
      {stage1_52[34],stage1_51[95],stage1_50[119],stage1_49[143],stage1_48[174]}
   );
   gpc615_5 gpc1878 (
      {stage0_48[403], stage0_48[404], stage0_48[405], stage0_48[406], stage0_48[407]},
      {stage0_49[388]},
      {stage0_50[210], stage0_50[211], stage0_50[212], stage0_50[213], stage0_50[214], stage0_50[215]},
      {stage1_52[35],stage1_51[96],stage1_50[120],stage1_49[144],stage1_48[175]}
   );
   gpc615_5 gpc1879 (
      {stage0_48[408], stage0_48[409], stage0_48[410], stage0_48[411], stage0_48[412]},
      {stage0_49[389]},
      {stage0_50[216], stage0_50[217], stage0_50[218], stage0_50[219], stage0_50[220], stage0_50[221]},
      {stage1_52[36],stage1_51[97],stage1_50[121],stage1_49[145],stage1_48[176]}
   );
   gpc615_5 gpc1880 (
      {stage0_48[413], stage0_48[414], stage0_48[415], stage0_48[416], stage0_48[417]},
      {stage0_49[390]},
      {stage0_50[222], stage0_50[223], stage0_50[224], stage0_50[225], stage0_50[226], stage0_50[227]},
      {stage1_52[37],stage1_51[98],stage1_50[122],stage1_49[146],stage1_48[177]}
   );
   gpc615_5 gpc1881 (
      {stage0_48[418], stage0_48[419], stage0_48[420], stage0_48[421], stage0_48[422]},
      {stage0_49[391]},
      {stage0_50[228], stage0_50[229], stage0_50[230], stage0_50[231], stage0_50[232], stage0_50[233]},
      {stage1_52[38],stage1_51[99],stage1_50[123],stage1_49[147],stage1_48[178]}
   );
   gpc615_5 gpc1882 (
      {stage0_48[423], stage0_48[424], stage0_48[425], stage0_48[426], stage0_48[427]},
      {stage0_49[392]},
      {stage0_50[234], stage0_50[235], stage0_50[236], stage0_50[237], stage0_50[238], stage0_50[239]},
      {stage1_52[39],stage1_51[100],stage1_50[124],stage1_49[148],stage1_48[179]}
   );
   gpc615_5 gpc1883 (
      {stage0_48[428], stage0_48[429], stage0_48[430], stage0_48[431], stage0_48[432]},
      {stage0_49[393]},
      {stage0_50[240], stage0_50[241], stage0_50[242], stage0_50[243], stage0_50[244], stage0_50[245]},
      {stage1_52[40],stage1_51[101],stage1_50[125],stage1_49[149],stage1_48[180]}
   );
   gpc615_5 gpc1884 (
      {stage0_48[433], stage0_48[434], stage0_48[435], stage0_48[436], stage0_48[437]},
      {stage0_49[394]},
      {stage0_50[246], stage0_50[247], stage0_50[248], stage0_50[249], stage0_50[250], stage0_50[251]},
      {stage1_52[41],stage1_51[102],stage1_50[126],stage1_49[150],stage1_48[181]}
   );
   gpc615_5 gpc1885 (
      {stage0_48[438], stage0_48[439], stage0_48[440], stage0_48[441], stage0_48[442]},
      {stage0_49[395]},
      {stage0_50[252], stage0_50[253], stage0_50[254], stage0_50[255], stage0_50[256], stage0_50[257]},
      {stage1_52[42],stage1_51[103],stage1_50[127],stage1_49[151],stage1_48[182]}
   );
   gpc615_5 gpc1886 (
      {stage0_48[443], stage0_48[444], stage0_48[445], stage0_48[446], stage0_48[447]},
      {stage0_49[396]},
      {stage0_50[258], stage0_50[259], stage0_50[260], stage0_50[261], stage0_50[262], stage0_50[263]},
      {stage1_52[43],stage1_51[104],stage1_50[128],stage1_49[152],stage1_48[183]}
   );
   gpc615_5 gpc1887 (
      {stage0_48[448], stage0_48[449], stage0_48[450], stage0_48[451], stage0_48[452]},
      {stage0_49[397]},
      {stage0_50[264], stage0_50[265], stage0_50[266], stage0_50[267], stage0_50[268], stage0_50[269]},
      {stage1_52[44],stage1_51[105],stage1_50[129],stage1_49[153],stage1_48[184]}
   );
   gpc615_5 gpc1888 (
      {stage0_48[453], stage0_48[454], stage0_48[455], stage0_48[456], stage0_48[457]},
      {stage0_49[398]},
      {stage0_50[270], stage0_50[271], stage0_50[272], stage0_50[273], stage0_50[274], stage0_50[275]},
      {stage1_52[45],stage1_51[106],stage1_50[130],stage1_49[154],stage1_48[185]}
   );
   gpc615_5 gpc1889 (
      {stage0_48[458], stage0_48[459], stage0_48[460], stage0_48[461], stage0_48[462]},
      {stage0_49[399]},
      {stage0_50[276], stage0_50[277], stage0_50[278], stage0_50[279], stage0_50[280], stage0_50[281]},
      {stage1_52[46],stage1_51[107],stage1_50[131],stage1_49[155],stage1_48[186]}
   );
   gpc615_5 gpc1890 (
      {stage0_48[463], stage0_48[464], stage0_48[465], stage0_48[466], stage0_48[467]},
      {stage0_49[400]},
      {stage0_50[282], stage0_50[283], stage0_50[284], stage0_50[285], stage0_50[286], stage0_50[287]},
      {stage1_52[47],stage1_51[108],stage1_50[132],stage1_49[156],stage1_48[187]}
   );
   gpc615_5 gpc1891 (
      {stage0_48[468], stage0_48[469], stage0_48[470], stage0_48[471], stage0_48[472]},
      {stage0_49[401]},
      {stage0_50[288], stage0_50[289], stage0_50[290], stage0_50[291], stage0_50[292], stage0_50[293]},
      {stage1_52[48],stage1_51[109],stage1_50[133],stage1_49[157],stage1_48[188]}
   );
   gpc615_5 gpc1892 (
      {stage0_48[473], stage0_48[474], stage0_48[475], stage0_48[476], stage0_48[477]},
      {stage0_49[402]},
      {stage0_50[294], stage0_50[295], stage0_50[296], stage0_50[297], stage0_50[298], stage0_50[299]},
      {stage1_52[49],stage1_51[110],stage1_50[134],stage1_49[158],stage1_48[189]}
   );
   gpc606_5 gpc1893 (
      {stage0_49[403], stage0_49[404], stage0_49[405], stage0_49[406], stage0_49[407], stage0_49[408]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[50],stage1_51[111],stage1_50[135],stage1_49[159]}
   );
   gpc606_5 gpc1894 (
      {stage0_49[409], stage0_49[410], stage0_49[411], stage0_49[412], stage0_49[413], stage0_49[414]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[51],stage1_51[112],stage1_50[136],stage1_49[160]}
   );
   gpc606_5 gpc1895 (
      {stage0_49[415], stage0_49[416], stage0_49[417], stage0_49[418], stage0_49[419], stage0_49[420]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[52],stage1_51[113],stage1_50[137],stage1_49[161]}
   );
   gpc606_5 gpc1896 (
      {stage0_49[421], stage0_49[422], stage0_49[423], stage0_49[424], stage0_49[425], stage0_49[426]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[53],stage1_51[114],stage1_50[138],stage1_49[162]}
   );
   gpc606_5 gpc1897 (
      {stage0_49[427], stage0_49[428], stage0_49[429], stage0_49[430], stage0_49[431], stage0_49[432]},
      {stage0_51[24], stage0_51[25], stage0_51[26], stage0_51[27], stage0_51[28], stage0_51[29]},
      {stage1_53[4],stage1_52[54],stage1_51[115],stage1_50[139],stage1_49[163]}
   );
   gpc606_5 gpc1898 (
      {stage0_49[433], stage0_49[434], stage0_49[435], stage0_49[436], stage0_49[437], stage0_49[438]},
      {stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33], stage0_51[34], stage0_51[35]},
      {stage1_53[5],stage1_52[55],stage1_51[116],stage1_50[140],stage1_49[164]}
   );
   gpc606_5 gpc1899 (
      {stage0_49[439], stage0_49[440], stage0_49[441], stage0_49[442], stage0_49[443], stage0_49[444]},
      {stage0_51[36], stage0_51[37], stage0_51[38], stage0_51[39], stage0_51[40], stage0_51[41]},
      {stage1_53[6],stage1_52[56],stage1_51[117],stage1_50[141],stage1_49[165]}
   );
   gpc606_5 gpc1900 (
      {stage0_49[445], stage0_49[446], stage0_49[447], stage0_49[448], stage0_49[449], stage0_49[450]},
      {stage0_51[42], stage0_51[43], stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47]},
      {stage1_53[7],stage1_52[57],stage1_51[118],stage1_50[142],stage1_49[166]}
   );
   gpc606_5 gpc1901 (
      {stage0_49[451], stage0_49[452], stage0_49[453], stage0_49[454], stage0_49[455], stage0_49[456]},
      {stage0_51[48], stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage1_53[8],stage1_52[58],stage1_51[119],stage1_50[143],stage1_49[167]}
   );
   gpc606_5 gpc1902 (
      {stage0_49[457], stage0_49[458], stage0_49[459], stage0_49[460], stage0_49[461], stage0_49[462]},
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58], stage0_51[59]},
      {stage1_53[9],stage1_52[59],stage1_51[120],stage1_50[144],stage1_49[168]}
   );
   gpc606_5 gpc1903 (
      {stage0_49[463], stage0_49[464], stage0_49[465], stage0_49[466], stage0_49[467], stage0_49[468]},
      {stage0_51[60], stage0_51[61], stage0_51[62], stage0_51[63], stage0_51[64], stage0_51[65]},
      {stage1_53[10],stage1_52[60],stage1_51[121],stage1_50[145],stage1_49[169]}
   );
   gpc606_5 gpc1904 (
      {stage0_49[469], stage0_49[470], stage0_49[471], stage0_49[472], stage0_49[473], stage0_49[474]},
      {stage0_51[66], stage0_51[67], stage0_51[68], stage0_51[69], stage0_51[70], stage0_51[71]},
      {stage1_53[11],stage1_52[61],stage1_51[122],stage1_50[146],stage1_49[170]}
   );
   gpc606_5 gpc1905 (
      {stage0_49[475], stage0_49[476], stage0_49[477], stage0_49[478], stage0_49[479], stage0_49[480]},
      {stage0_51[72], stage0_51[73], stage0_51[74], stage0_51[75], stage0_51[76], stage0_51[77]},
      {stage1_53[12],stage1_52[62],stage1_51[123],stage1_50[147],stage1_49[171]}
   );
   gpc615_5 gpc1906 (
      {stage0_49[481], stage0_49[482], stage0_49[483], stage0_49[484], stage0_49[485]},
      {stage0_50[300]},
      {stage0_51[78], stage0_51[79], stage0_51[80], stage0_51[81], stage0_51[82], stage0_51[83]},
      {stage1_53[13],stage1_52[63],stage1_51[124],stage1_50[148],stage1_49[172]}
   );
   gpc615_5 gpc1907 (
      {stage0_50[301], stage0_50[302], stage0_50[303], stage0_50[304], stage0_50[305]},
      {stage0_51[84]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[14],stage1_52[64],stage1_51[125],stage1_50[149]}
   );
   gpc615_5 gpc1908 (
      {stage0_50[306], stage0_50[307], stage0_50[308], stage0_50[309], stage0_50[310]},
      {stage0_51[85]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[15],stage1_52[65],stage1_51[126],stage1_50[150]}
   );
   gpc615_5 gpc1909 (
      {stage0_50[311], stage0_50[312], stage0_50[313], stage0_50[314], stage0_50[315]},
      {stage0_51[86]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[16],stage1_52[66],stage1_51[127],stage1_50[151]}
   );
   gpc615_5 gpc1910 (
      {stage0_50[316], stage0_50[317], stage0_50[318], stage0_50[319], stage0_50[320]},
      {stage0_51[87]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[17],stage1_52[67],stage1_51[128],stage1_50[152]}
   );
   gpc615_5 gpc1911 (
      {stage0_50[321], stage0_50[322], stage0_50[323], stage0_50[324], stage0_50[325]},
      {stage0_51[88]},
      {stage0_52[24], stage0_52[25], stage0_52[26], stage0_52[27], stage0_52[28], stage0_52[29]},
      {stage1_54[4],stage1_53[18],stage1_52[68],stage1_51[129],stage1_50[153]}
   );
   gpc615_5 gpc1912 (
      {stage0_50[326], stage0_50[327], stage0_50[328], stage0_50[329], stage0_50[330]},
      {stage0_51[89]},
      {stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35]},
      {stage1_54[5],stage1_53[19],stage1_52[69],stage1_51[130],stage1_50[154]}
   );
   gpc615_5 gpc1913 (
      {stage0_50[331], stage0_50[332], stage0_50[333], stage0_50[334], stage0_50[335]},
      {stage0_51[90]},
      {stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage1_54[6],stage1_53[20],stage1_52[70],stage1_51[131],stage1_50[155]}
   );
   gpc615_5 gpc1914 (
      {stage0_50[336], stage0_50[337], stage0_50[338], stage0_50[339], stage0_50[340]},
      {stage0_51[91]},
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46], stage0_52[47]},
      {stage1_54[7],stage1_53[21],stage1_52[71],stage1_51[132],stage1_50[156]}
   );
   gpc615_5 gpc1915 (
      {stage0_50[341], stage0_50[342], stage0_50[343], stage0_50[344], stage0_50[345]},
      {stage0_51[92]},
      {stage0_52[48], stage0_52[49], stage0_52[50], stage0_52[51], stage0_52[52], stage0_52[53]},
      {stage1_54[8],stage1_53[22],stage1_52[72],stage1_51[133],stage1_50[157]}
   );
   gpc615_5 gpc1916 (
      {stage0_50[346], stage0_50[347], stage0_50[348], stage0_50[349], stage0_50[350]},
      {stage0_51[93]},
      {stage0_52[54], stage0_52[55], stage0_52[56], stage0_52[57], stage0_52[58], stage0_52[59]},
      {stage1_54[9],stage1_53[23],stage1_52[73],stage1_51[134],stage1_50[158]}
   );
   gpc615_5 gpc1917 (
      {stage0_50[351], stage0_50[352], stage0_50[353], stage0_50[354], stage0_50[355]},
      {stage0_51[94]},
      {stage0_52[60], stage0_52[61], stage0_52[62], stage0_52[63], stage0_52[64], stage0_52[65]},
      {stage1_54[10],stage1_53[24],stage1_52[74],stage1_51[135],stage1_50[159]}
   );
   gpc615_5 gpc1918 (
      {stage0_50[356], stage0_50[357], stage0_50[358], stage0_50[359], stage0_50[360]},
      {stage0_51[95]},
      {stage0_52[66], stage0_52[67], stage0_52[68], stage0_52[69], stage0_52[70], stage0_52[71]},
      {stage1_54[11],stage1_53[25],stage1_52[75],stage1_51[136],stage1_50[160]}
   );
   gpc615_5 gpc1919 (
      {stage0_50[361], stage0_50[362], stage0_50[363], stage0_50[364], stage0_50[365]},
      {stage0_51[96]},
      {stage0_52[72], stage0_52[73], stage0_52[74], stage0_52[75], stage0_52[76], stage0_52[77]},
      {stage1_54[12],stage1_53[26],stage1_52[76],stage1_51[137],stage1_50[161]}
   );
   gpc615_5 gpc1920 (
      {stage0_50[366], stage0_50[367], stage0_50[368], stage0_50[369], stage0_50[370]},
      {stage0_51[97]},
      {stage0_52[78], stage0_52[79], stage0_52[80], stage0_52[81], stage0_52[82], stage0_52[83]},
      {stage1_54[13],stage1_53[27],stage1_52[77],stage1_51[138],stage1_50[162]}
   );
   gpc615_5 gpc1921 (
      {stage0_50[371], stage0_50[372], stage0_50[373], stage0_50[374], stage0_50[375]},
      {stage0_51[98]},
      {stage0_52[84], stage0_52[85], stage0_52[86], stage0_52[87], stage0_52[88], stage0_52[89]},
      {stage1_54[14],stage1_53[28],stage1_52[78],stage1_51[139],stage1_50[163]}
   );
   gpc615_5 gpc1922 (
      {stage0_50[376], stage0_50[377], stage0_50[378], stage0_50[379], stage0_50[380]},
      {stage0_51[99]},
      {stage0_52[90], stage0_52[91], stage0_52[92], stage0_52[93], stage0_52[94], stage0_52[95]},
      {stage1_54[15],stage1_53[29],stage1_52[79],stage1_51[140],stage1_50[164]}
   );
   gpc615_5 gpc1923 (
      {stage0_50[381], stage0_50[382], stage0_50[383], stage0_50[384], stage0_50[385]},
      {stage0_51[100]},
      {stage0_52[96], stage0_52[97], stage0_52[98], stage0_52[99], stage0_52[100], stage0_52[101]},
      {stage1_54[16],stage1_53[30],stage1_52[80],stage1_51[141],stage1_50[165]}
   );
   gpc615_5 gpc1924 (
      {stage0_50[386], stage0_50[387], stage0_50[388], stage0_50[389], stage0_50[390]},
      {stage0_51[101]},
      {stage0_52[102], stage0_52[103], stage0_52[104], stage0_52[105], stage0_52[106], stage0_52[107]},
      {stage1_54[17],stage1_53[31],stage1_52[81],stage1_51[142],stage1_50[166]}
   );
   gpc615_5 gpc1925 (
      {stage0_50[391], stage0_50[392], stage0_50[393], stage0_50[394], stage0_50[395]},
      {stage0_51[102]},
      {stage0_52[108], stage0_52[109], stage0_52[110], stage0_52[111], stage0_52[112], stage0_52[113]},
      {stage1_54[18],stage1_53[32],stage1_52[82],stage1_51[143],stage1_50[167]}
   );
   gpc615_5 gpc1926 (
      {stage0_50[396], stage0_50[397], stage0_50[398], stage0_50[399], stage0_50[400]},
      {stage0_51[103]},
      {stage0_52[114], stage0_52[115], stage0_52[116], stage0_52[117], stage0_52[118], stage0_52[119]},
      {stage1_54[19],stage1_53[33],stage1_52[83],stage1_51[144],stage1_50[168]}
   );
   gpc615_5 gpc1927 (
      {stage0_50[401], stage0_50[402], stage0_50[403], stage0_50[404], stage0_50[405]},
      {stage0_51[104]},
      {stage0_52[120], stage0_52[121], stage0_52[122], stage0_52[123], stage0_52[124], stage0_52[125]},
      {stage1_54[20],stage1_53[34],stage1_52[84],stage1_51[145],stage1_50[169]}
   );
   gpc615_5 gpc1928 (
      {stage0_50[406], stage0_50[407], stage0_50[408], stage0_50[409], stage0_50[410]},
      {stage0_51[105]},
      {stage0_52[126], stage0_52[127], stage0_52[128], stage0_52[129], stage0_52[130], stage0_52[131]},
      {stage1_54[21],stage1_53[35],stage1_52[85],stage1_51[146],stage1_50[170]}
   );
   gpc615_5 gpc1929 (
      {stage0_50[411], stage0_50[412], stage0_50[413], stage0_50[414], stage0_50[415]},
      {stage0_51[106]},
      {stage0_52[132], stage0_52[133], stage0_52[134], stage0_52[135], stage0_52[136], stage0_52[137]},
      {stage1_54[22],stage1_53[36],stage1_52[86],stage1_51[147],stage1_50[171]}
   );
   gpc615_5 gpc1930 (
      {stage0_50[416], stage0_50[417], stage0_50[418], stage0_50[419], stage0_50[420]},
      {stage0_51[107]},
      {stage0_52[138], stage0_52[139], stage0_52[140], stage0_52[141], stage0_52[142], stage0_52[143]},
      {stage1_54[23],stage1_53[37],stage1_52[87],stage1_51[148],stage1_50[172]}
   );
   gpc615_5 gpc1931 (
      {stage0_50[421], stage0_50[422], stage0_50[423], stage0_50[424], stage0_50[425]},
      {stage0_51[108]},
      {stage0_52[144], stage0_52[145], stage0_52[146], stage0_52[147], stage0_52[148], stage0_52[149]},
      {stage1_54[24],stage1_53[38],stage1_52[88],stage1_51[149],stage1_50[173]}
   );
   gpc615_5 gpc1932 (
      {stage0_50[426], stage0_50[427], stage0_50[428], stage0_50[429], stage0_50[430]},
      {stage0_51[109]},
      {stage0_52[150], stage0_52[151], stage0_52[152], stage0_52[153], stage0_52[154], stage0_52[155]},
      {stage1_54[25],stage1_53[39],stage1_52[89],stage1_51[150],stage1_50[174]}
   );
   gpc615_5 gpc1933 (
      {stage0_50[431], stage0_50[432], stage0_50[433], stage0_50[434], stage0_50[435]},
      {stage0_51[110]},
      {stage0_52[156], stage0_52[157], stage0_52[158], stage0_52[159], stage0_52[160], stage0_52[161]},
      {stage1_54[26],stage1_53[40],stage1_52[90],stage1_51[151],stage1_50[175]}
   );
   gpc615_5 gpc1934 (
      {stage0_50[436], stage0_50[437], stage0_50[438], stage0_50[439], stage0_50[440]},
      {stage0_51[111]},
      {stage0_52[162], stage0_52[163], stage0_52[164], stage0_52[165], stage0_52[166], stage0_52[167]},
      {stage1_54[27],stage1_53[41],stage1_52[91],stage1_51[152],stage1_50[176]}
   );
   gpc615_5 gpc1935 (
      {stage0_50[441], stage0_50[442], stage0_50[443], stage0_50[444], stage0_50[445]},
      {stage0_51[112]},
      {stage0_52[168], stage0_52[169], stage0_52[170], stage0_52[171], stage0_52[172], stage0_52[173]},
      {stage1_54[28],stage1_53[42],stage1_52[92],stage1_51[153],stage1_50[177]}
   );
   gpc615_5 gpc1936 (
      {stage0_50[446], stage0_50[447], stage0_50[448], stage0_50[449], stage0_50[450]},
      {stage0_51[113]},
      {stage0_52[174], stage0_52[175], stage0_52[176], stage0_52[177], stage0_52[178], stage0_52[179]},
      {stage1_54[29],stage1_53[43],stage1_52[93],stage1_51[154],stage1_50[178]}
   );
   gpc615_5 gpc1937 (
      {stage0_50[451], stage0_50[452], stage0_50[453], stage0_50[454], stage0_50[455]},
      {stage0_51[114]},
      {stage0_52[180], stage0_52[181], stage0_52[182], stage0_52[183], stage0_52[184], stage0_52[185]},
      {stage1_54[30],stage1_53[44],stage1_52[94],stage1_51[155],stage1_50[179]}
   );
   gpc615_5 gpc1938 (
      {stage0_50[456], stage0_50[457], stage0_50[458], stage0_50[459], stage0_50[460]},
      {stage0_51[115]},
      {stage0_52[186], stage0_52[187], stage0_52[188], stage0_52[189], stage0_52[190], stage0_52[191]},
      {stage1_54[31],stage1_53[45],stage1_52[95],stage1_51[156],stage1_50[180]}
   );
   gpc615_5 gpc1939 (
      {stage0_50[461], stage0_50[462], stage0_50[463], stage0_50[464], stage0_50[465]},
      {stage0_51[116]},
      {stage0_52[192], stage0_52[193], stage0_52[194], stage0_52[195], stage0_52[196], stage0_52[197]},
      {stage1_54[32],stage1_53[46],stage1_52[96],stage1_51[157],stage1_50[181]}
   );
   gpc615_5 gpc1940 (
      {stage0_50[466], stage0_50[467], stage0_50[468], stage0_50[469], stage0_50[470]},
      {stage0_51[117]},
      {stage0_52[198], stage0_52[199], stage0_52[200], stage0_52[201], stage0_52[202], stage0_52[203]},
      {stage1_54[33],stage1_53[47],stage1_52[97],stage1_51[158],stage1_50[182]}
   );
   gpc615_5 gpc1941 (
      {stage0_50[471], stage0_50[472], stage0_50[473], stage0_50[474], stage0_50[475]},
      {stage0_51[118]},
      {stage0_52[204], stage0_52[205], stage0_52[206], stage0_52[207], stage0_52[208], stage0_52[209]},
      {stage1_54[34],stage1_53[48],stage1_52[98],stage1_51[159],stage1_50[183]}
   );
   gpc615_5 gpc1942 (
      {stage0_50[476], stage0_50[477], stage0_50[478], stage0_50[479], stage0_50[480]},
      {stage0_51[119]},
      {stage0_52[210], stage0_52[211], stage0_52[212], stage0_52[213], stage0_52[214], stage0_52[215]},
      {stage1_54[35],stage1_53[49],stage1_52[99],stage1_51[160],stage1_50[184]}
   );
   gpc615_5 gpc1943 (
      {stage0_51[120], stage0_51[121], stage0_51[122], stage0_51[123], stage0_51[124]},
      {stage0_52[216]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[36],stage1_53[50],stage1_52[100],stage1_51[161]}
   );
   gpc615_5 gpc1944 (
      {stage0_51[125], stage0_51[126], stage0_51[127], stage0_51[128], stage0_51[129]},
      {stage0_52[217]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[37],stage1_53[51],stage1_52[101],stage1_51[162]}
   );
   gpc615_5 gpc1945 (
      {stage0_51[130], stage0_51[131], stage0_51[132], stage0_51[133], stage0_51[134]},
      {stage0_52[218]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[38],stage1_53[52],stage1_52[102],stage1_51[163]}
   );
   gpc615_5 gpc1946 (
      {stage0_51[135], stage0_51[136], stage0_51[137], stage0_51[138], stage0_51[139]},
      {stage0_52[219]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[39],stage1_53[53],stage1_52[103],stage1_51[164]}
   );
   gpc615_5 gpc1947 (
      {stage0_51[140], stage0_51[141], stage0_51[142], stage0_51[143], stage0_51[144]},
      {stage0_52[220]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[40],stage1_53[54],stage1_52[104],stage1_51[165]}
   );
   gpc615_5 gpc1948 (
      {stage0_51[145], stage0_51[146], stage0_51[147], stage0_51[148], stage0_51[149]},
      {stage0_52[221]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[41],stage1_53[55],stage1_52[105],stage1_51[166]}
   );
   gpc615_5 gpc1949 (
      {stage0_51[150], stage0_51[151], stage0_51[152], stage0_51[153], stage0_51[154]},
      {stage0_52[222]},
      {stage0_53[36], stage0_53[37], stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41]},
      {stage1_55[6],stage1_54[42],stage1_53[56],stage1_52[106],stage1_51[167]}
   );
   gpc615_5 gpc1950 (
      {stage0_51[155], stage0_51[156], stage0_51[157], stage0_51[158], stage0_51[159]},
      {stage0_52[223]},
      {stage0_53[42], stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage1_55[7],stage1_54[43],stage1_53[57],stage1_52[107],stage1_51[168]}
   );
   gpc615_5 gpc1951 (
      {stage0_51[160], stage0_51[161], stage0_51[162], stage0_51[163], stage0_51[164]},
      {stage0_52[224]},
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52], stage0_53[53]},
      {stage1_55[8],stage1_54[44],stage1_53[58],stage1_52[108],stage1_51[169]}
   );
   gpc615_5 gpc1952 (
      {stage0_51[165], stage0_51[166], stage0_51[167], stage0_51[168], stage0_51[169]},
      {stage0_52[225]},
      {stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57], stage0_53[58], stage0_53[59]},
      {stage1_55[9],stage1_54[45],stage1_53[59],stage1_52[109],stage1_51[170]}
   );
   gpc615_5 gpc1953 (
      {stage0_51[170], stage0_51[171], stage0_51[172], stage0_51[173], stage0_51[174]},
      {stage0_52[226]},
      {stage0_53[60], stage0_53[61], stage0_53[62], stage0_53[63], stage0_53[64], stage0_53[65]},
      {stage1_55[10],stage1_54[46],stage1_53[60],stage1_52[110],stage1_51[171]}
   );
   gpc615_5 gpc1954 (
      {stage0_51[175], stage0_51[176], stage0_51[177], stage0_51[178], stage0_51[179]},
      {stage0_52[227]},
      {stage0_53[66], stage0_53[67], stage0_53[68], stage0_53[69], stage0_53[70], stage0_53[71]},
      {stage1_55[11],stage1_54[47],stage1_53[61],stage1_52[111],stage1_51[172]}
   );
   gpc615_5 gpc1955 (
      {stage0_51[180], stage0_51[181], stage0_51[182], stage0_51[183], stage0_51[184]},
      {stage0_52[228]},
      {stage0_53[72], stage0_53[73], stage0_53[74], stage0_53[75], stage0_53[76], stage0_53[77]},
      {stage1_55[12],stage1_54[48],stage1_53[62],stage1_52[112],stage1_51[173]}
   );
   gpc615_5 gpc1956 (
      {stage0_51[185], stage0_51[186], stage0_51[187], stage0_51[188], stage0_51[189]},
      {stage0_52[229]},
      {stage0_53[78], stage0_53[79], stage0_53[80], stage0_53[81], stage0_53[82], stage0_53[83]},
      {stage1_55[13],stage1_54[49],stage1_53[63],stage1_52[113],stage1_51[174]}
   );
   gpc615_5 gpc1957 (
      {stage0_51[190], stage0_51[191], stage0_51[192], stage0_51[193], stage0_51[194]},
      {stage0_52[230]},
      {stage0_53[84], stage0_53[85], stage0_53[86], stage0_53[87], stage0_53[88], stage0_53[89]},
      {stage1_55[14],stage1_54[50],stage1_53[64],stage1_52[114],stage1_51[175]}
   );
   gpc615_5 gpc1958 (
      {stage0_51[195], stage0_51[196], stage0_51[197], stage0_51[198], stage0_51[199]},
      {stage0_52[231]},
      {stage0_53[90], stage0_53[91], stage0_53[92], stage0_53[93], stage0_53[94], stage0_53[95]},
      {stage1_55[15],stage1_54[51],stage1_53[65],stage1_52[115],stage1_51[176]}
   );
   gpc615_5 gpc1959 (
      {stage0_51[200], stage0_51[201], stage0_51[202], stage0_51[203], stage0_51[204]},
      {stage0_52[232]},
      {stage0_53[96], stage0_53[97], stage0_53[98], stage0_53[99], stage0_53[100], stage0_53[101]},
      {stage1_55[16],stage1_54[52],stage1_53[66],stage1_52[116],stage1_51[177]}
   );
   gpc615_5 gpc1960 (
      {stage0_51[205], stage0_51[206], stage0_51[207], stage0_51[208], stage0_51[209]},
      {stage0_52[233]},
      {stage0_53[102], stage0_53[103], stage0_53[104], stage0_53[105], stage0_53[106], stage0_53[107]},
      {stage1_55[17],stage1_54[53],stage1_53[67],stage1_52[117],stage1_51[178]}
   );
   gpc615_5 gpc1961 (
      {stage0_51[210], stage0_51[211], stage0_51[212], stage0_51[213], stage0_51[214]},
      {stage0_52[234]},
      {stage0_53[108], stage0_53[109], stage0_53[110], stage0_53[111], stage0_53[112], stage0_53[113]},
      {stage1_55[18],stage1_54[54],stage1_53[68],stage1_52[118],stage1_51[179]}
   );
   gpc615_5 gpc1962 (
      {stage0_51[215], stage0_51[216], stage0_51[217], stage0_51[218], stage0_51[219]},
      {stage0_52[235]},
      {stage0_53[114], stage0_53[115], stage0_53[116], stage0_53[117], stage0_53[118], stage0_53[119]},
      {stage1_55[19],stage1_54[55],stage1_53[69],stage1_52[119],stage1_51[180]}
   );
   gpc615_5 gpc1963 (
      {stage0_51[220], stage0_51[221], stage0_51[222], stage0_51[223], stage0_51[224]},
      {stage0_52[236]},
      {stage0_53[120], stage0_53[121], stage0_53[122], stage0_53[123], stage0_53[124], stage0_53[125]},
      {stage1_55[20],stage1_54[56],stage1_53[70],stage1_52[120],stage1_51[181]}
   );
   gpc615_5 gpc1964 (
      {stage0_51[225], stage0_51[226], stage0_51[227], stage0_51[228], stage0_51[229]},
      {stage0_52[237]},
      {stage0_53[126], stage0_53[127], stage0_53[128], stage0_53[129], stage0_53[130], stage0_53[131]},
      {stage1_55[21],stage1_54[57],stage1_53[71],stage1_52[121],stage1_51[182]}
   );
   gpc615_5 gpc1965 (
      {stage0_51[230], stage0_51[231], stage0_51[232], stage0_51[233], stage0_51[234]},
      {stage0_52[238]},
      {stage0_53[132], stage0_53[133], stage0_53[134], stage0_53[135], stage0_53[136], stage0_53[137]},
      {stage1_55[22],stage1_54[58],stage1_53[72],stage1_52[122],stage1_51[183]}
   );
   gpc615_5 gpc1966 (
      {stage0_51[235], stage0_51[236], stage0_51[237], stage0_51[238], stage0_51[239]},
      {stage0_52[239]},
      {stage0_53[138], stage0_53[139], stage0_53[140], stage0_53[141], stage0_53[142], stage0_53[143]},
      {stage1_55[23],stage1_54[59],stage1_53[73],stage1_52[123],stage1_51[184]}
   );
   gpc615_5 gpc1967 (
      {stage0_51[240], stage0_51[241], stage0_51[242], stage0_51[243], stage0_51[244]},
      {stage0_52[240]},
      {stage0_53[144], stage0_53[145], stage0_53[146], stage0_53[147], stage0_53[148], stage0_53[149]},
      {stage1_55[24],stage1_54[60],stage1_53[74],stage1_52[124],stage1_51[185]}
   );
   gpc615_5 gpc1968 (
      {stage0_51[245], stage0_51[246], stage0_51[247], stage0_51[248], stage0_51[249]},
      {stage0_52[241]},
      {stage0_53[150], stage0_53[151], stage0_53[152], stage0_53[153], stage0_53[154], stage0_53[155]},
      {stage1_55[25],stage1_54[61],stage1_53[75],stage1_52[125],stage1_51[186]}
   );
   gpc615_5 gpc1969 (
      {stage0_51[250], stage0_51[251], stage0_51[252], stage0_51[253], stage0_51[254]},
      {stage0_52[242]},
      {stage0_53[156], stage0_53[157], stage0_53[158], stage0_53[159], stage0_53[160], stage0_53[161]},
      {stage1_55[26],stage1_54[62],stage1_53[76],stage1_52[126],stage1_51[187]}
   );
   gpc615_5 gpc1970 (
      {stage0_51[255], stage0_51[256], stage0_51[257], stage0_51[258], stage0_51[259]},
      {stage0_52[243]},
      {stage0_53[162], stage0_53[163], stage0_53[164], stage0_53[165], stage0_53[166], stage0_53[167]},
      {stage1_55[27],stage1_54[63],stage1_53[77],stage1_52[127],stage1_51[188]}
   );
   gpc615_5 gpc1971 (
      {stage0_51[260], stage0_51[261], stage0_51[262], stage0_51[263], stage0_51[264]},
      {stage0_52[244]},
      {stage0_53[168], stage0_53[169], stage0_53[170], stage0_53[171], stage0_53[172], stage0_53[173]},
      {stage1_55[28],stage1_54[64],stage1_53[78],stage1_52[128],stage1_51[189]}
   );
   gpc615_5 gpc1972 (
      {stage0_51[265], stage0_51[266], stage0_51[267], stage0_51[268], stage0_51[269]},
      {stage0_52[245]},
      {stage0_53[174], stage0_53[175], stage0_53[176], stage0_53[177], stage0_53[178], stage0_53[179]},
      {stage1_55[29],stage1_54[65],stage1_53[79],stage1_52[129],stage1_51[190]}
   );
   gpc615_5 gpc1973 (
      {stage0_51[270], stage0_51[271], stage0_51[272], stage0_51[273], stage0_51[274]},
      {stage0_52[246]},
      {stage0_53[180], stage0_53[181], stage0_53[182], stage0_53[183], stage0_53[184], stage0_53[185]},
      {stage1_55[30],stage1_54[66],stage1_53[80],stage1_52[130],stage1_51[191]}
   );
   gpc615_5 gpc1974 (
      {stage0_51[275], stage0_51[276], stage0_51[277], stage0_51[278], stage0_51[279]},
      {stage0_52[247]},
      {stage0_53[186], stage0_53[187], stage0_53[188], stage0_53[189], stage0_53[190], stage0_53[191]},
      {stage1_55[31],stage1_54[67],stage1_53[81],stage1_52[131],stage1_51[192]}
   );
   gpc615_5 gpc1975 (
      {stage0_51[280], stage0_51[281], stage0_51[282], stage0_51[283], stage0_51[284]},
      {stage0_52[248]},
      {stage0_53[192], stage0_53[193], stage0_53[194], stage0_53[195], stage0_53[196], stage0_53[197]},
      {stage1_55[32],stage1_54[68],stage1_53[82],stage1_52[132],stage1_51[193]}
   );
   gpc615_5 gpc1976 (
      {stage0_51[285], stage0_51[286], stage0_51[287], stage0_51[288], stage0_51[289]},
      {stage0_52[249]},
      {stage0_53[198], stage0_53[199], stage0_53[200], stage0_53[201], stage0_53[202], stage0_53[203]},
      {stage1_55[33],stage1_54[69],stage1_53[83],stage1_52[133],stage1_51[194]}
   );
   gpc615_5 gpc1977 (
      {stage0_51[290], stage0_51[291], stage0_51[292], stage0_51[293], stage0_51[294]},
      {stage0_52[250]},
      {stage0_53[204], stage0_53[205], stage0_53[206], stage0_53[207], stage0_53[208], stage0_53[209]},
      {stage1_55[34],stage1_54[70],stage1_53[84],stage1_52[134],stage1_51[195]}
   );
   gpc615_5 gpc1978 (
      {stage0_51[295], stage0_51[296], stage0_51[297], stage0_51[298], stage0_51[299]},
      {stage0_52[251]},
      {stage0_53[210], stage0_53[211], stage0_53[212], stage0_53[213], stage0_53[214], stage0_53[215]},
      {stage1_55[35],stage1_54[71],stage1_53[85],stage1_52[135],stage1_51[196]}
   );
   gpc615_5 gpc1979 (
      {stage0_51[300], stage0_51[301], stage0_51[302], stage0_51[303], stage0_51[304]},
      {stage0_52[252]},
      {stage0_53[216], stage0_53[217], stage0_53[218], stage0_53[219], stage0_53[220], stage0_53[221]},
      {stage1_55[36],stage1_54[72],stage1_53[86],stage1_52[136],stage1_51[197]}
   );
   gpc615_5 gpc1980 (
      {stage0_51[305], stage0_51[306], stage0_51[307], stage0_51[308], stage0_51[309]},
      {stage0_52[253]},
      {stage0_53[222], stage0_53[223], stage0_53[224], stage0_53[225], stage0_53[226], stage0_53[227]},
      {stage1_55[37],stage1_54[73],stage1_53[87],stage1_52[137],stage1_51[198]}
   );
   gpc615_5 gpc1981 (
      {stage0_51[310], stage0_51[311], stage0_51[312], stage0_51[313], stage0_51[314]},
      {stage0_52[254]},
      {stage0_53[228], stage0_53[229], stage0_53[230], stage0_53[231], stage0_53[232], stage0_53[233]},
      {stage1_55[38],stage1_54[74],stage1_53[88],stage1_52[138],stage1_51[199]}
   );
   gpc615_5 gpc1982 (
      {stage0_51[315], stage0_51[316], stage0_51[317], stage0_51[318], stage0_51[319]},
      {stage0_52[255]},
      {stage0_53[234], stage0_53[235], stage0_53[236], stage0_53[237], stage0_53[238], stage0_53[239]},
      {stage1_55[39],stage1_54[75],stage1_53[89],stage1_52[139],stage1_51[200]}
   );
   gpc615_5 gpc1983 (
      {stage0_51[320], stage0_51[321], stage0_51[322], stage0_51[323], stage0_51[324]},
      {stage0_52[256]},
      {stage0_53[240], stage0_53[241], stage0_53[242], stage0_53[243], stage0_53[244], stage0_53[245]},
      {stage1_55[40],stage1_54[76],stage1_53[90],stage1_52[140],stage1_51[201]}
   );
   gpc615_5 gpc1984 (
      {stage0_51[325], stage0_51[326], stage0_51[327], stage0_51[328], stage0_51[329]},
      {stage0_52[257]},
      {stage0_53[246], stage0_53[247], stage0_53[248], stage0_53[249], stage0_53[250], stage0_53[251]},
      {stage1_55[41],stage1_54[77],stage1_53[91],stage1_52[141],stage1_51[202]}
   );
   gpc615_5 gpc1985 (
      {stage0_51[330], stage0_51[331], stage0_51[332], stage0_51[333], stage0_51[334]},
      {stage0_52[258]},
      {stage0_53[252], stage0_53[253], stage0_53[254], stage0_53[255], stage0_53[256], stage0_53[257]},
      {stage1_55[42],stage1_54[78],stage1_53[92],stage1_52[142],stage1_51[203]}
   );
   gpc615_5 gpc1986 (
      {stage0_51[335], stage0_51[336], stage0_51[337], stage0_51[338], stage0_51[339]},
      {stage0_52[259]},
      {stage0_53[258], stage0_53[259], stage0_53[260], stage0_53[261], stage0_53[262], stage0_53[263]},
      {stage1_55[43],stage1_54[79],stage1_53[93],stage1_52[143],stage1_51[204]}
   );
   gpc615_5 gpc1987 (
      {stage0_51[340], stage0_51[341], stage0_51[342], stage0_51[343], stage0_51[344]},
      {stage0_52[260]},
      {stage0_53[264], stage0_53[265], stage0_53[266], stage0_53[267], stage0_53[268], stage0_53[269]},
      {stage1_55[44],stage1_54[80],stage1_53[94],stage1_52[144],stage1_51[205]}
   );
   gpc615_5 gpc1988 (
      {stage0_51[345], stage0_51[346], stage0_51[347], stage0_51[348], stage0_51[349]},
      {stage0_52[261]},
      {stage0_53[270], stage0_53[271], stage0_53[272], stage0_53[273], stage0_53[274], stage0_53[275]},
      {stage1_55[45],stage1_54[81],stage1_53[95],stage1_52[145],stage1_51[206]}
   );
   gpc615_5 gpc1989 (
      {stage0_51[350], stage0_51[351], stage0_51[352], stage0_51[353], stage0_51[354]},
      {stage0_52[262]},
      {stage0_53[276], stage0_53[277], stage0_53[278], stage0_53[279], stage0_53[280], stage0_53[281]},
      {stage1_55[46],stage1_54[82],stage1_53[96],stage1_52[146],stage1_51[207]}
   );
   gpc615_5 gpc1990 (
      {stage0_51[355], stage0_51[356], stage0_51[357], stage0_51[358], stage0_51[359]},
      {stage0_52[263]},
      {stage0_53[282], stage0_53[283], stage0_53[284], stage0_53[285], stage0_53[286], stage0_53[287]},
      {stage1_55[47],stage1_54[83],stage1_53[97],stage1_52[147],stage1_51[208]}
   );
   gpc615_5 gpc1991 (
      {stage0_51[360], stage0_51[361], stage0_51[362], stage0_51[363], stage0_51[364]},
      {stage0_52[264]},
      {stage0_53[288], stage0_53[289], stage0_53[290], stage0_53[291], stage0_53[292], stage0_53[293]},
      {stage1_55[48],stage1_54[84],stage1_53[98],stage1_52[148],stage1_51[209]}
   );
   gpc615_5 gpc1992 (
      {stage0_51[365], stage0_51[366], stage0_51[367], stage0_51[368], stage0_51[369]},
      {stage0_52[265]},
      {stage0_53[294], stage0_53[295], stage0_53[296], stage0_53[297], stage0_53[298], stage0_53[299]},
      {stage1_55[49],stage1_54[85],stage1_53[99],stage1_52[149],stage1_51[210]}
   );
   gpc615_5 gpc1993 (
      {stage0_51[370], stage0_51[371], stage0_51[372], stage0_51[373], stage0_51[374]},
      {stage0_52[266]},
      {stage0_53[300], stage0_53[301], stage0_53[302], stage0_53[303], stage0_53[304], stage0_53[305]},
      {stage1_55[50],stage1_54[86],stage1_53[100],stage1_52[150],stage1_51[211]}
   );
   gpc615_5 gpc1994 (
      {stage0_51[375], stage0_51[376], stage0_51[377], stage0_51[378], stage0_51[379]},
      {stage0_52[267]},
      {stage0_53[306], stage0_53[307], stage0_53[308], stage0_53[309], stage0_53[310], stage0_53[311]},
      {stage1_55[51],stage1_54[87],stage1_53[101],stage1_52[151],stage1_51[212]}
   );
   gpc615_5 gpc1995 (
      {stage0_51[380], stage0_51[381], stage0_51[382], stage0_51[383], stage0_51[384]},
      {stage0_52[268]},
      {stage0_53[312], stage0_53[313], stage0_53[314], stage0_53[315], stage0_53[316], stage0_53[317]},
      {stage1_55[52],stage1_54[88],stage1_53[102],stage1_52[152],stage1_51[213]}
   );
   gpc615_5 gpc1996 (
      {stage0_51[385], stage0_51[386], stage0_51[387], stage0_51[388], stage0_51[389]},
      {stage0_52[269]},
      {stage0_53[318], stage0_53[319], stage0_53[320], stage0_53[321], stage0_53[322], stage0_53[323]},
      {stage1_55[53],stage1_54[89],stage1_53[103],stage1_52[153],stage1_51[214]}
   );
   gpc615_5 gpc1997 (
      {stage0_51[390], stage0_51[391], stage0_51[392], stage0_51[393], stage0_51[394]},
      {stage0_52[270]},
      {stage0_53[324], stage0_53[325], stage0_53[326], stage0_53[327], stage0_53[328], stage0_53[329]},
      {stage1_55[54],stage1_54[90],stage1_53[104],stage1_52[154],stage1_51[215]}
   );
   gpc615_5 gpc1998 (
      {stage0_51[395], stage0_51[396], stage0_51[397], stage0_51[398], stage0_51[399]},
      {stage0_52[271]},
      {stage0_53[330], stage0_53[331], stage0_53[332], stage0_53[333], stage0_53[334], stage0_53[335]},
      {stage1_55[55],stage1_54[91],stage1_53[105],stage1_52[155],stage1_51[216]}
   );
   gpc615_5 gpc1999 (
      {stage0_51[400], stage0_51[401], stage0_51[402], stage0_51[403], stage0_51[404]},
      {stage0_52[272]},
      {stage0_53[336], stage0_53[337], stage0_53[338], stage0_53[339], stage0_53[340], stage0_53[341]},
      {stage1_55[56],stage1_54[92],stage1_53[106],stage1_52[156],stage1_51[217]}
   );
   gpc615_5 gpc2000 (
      {stage0_51[405], stage0_51[406], stage0_51[407], stage0_51[408], stage0_51[409]},
      {stage0_52[273]},
      {stage0_53[342], stage0_53[343], stage0_53[344], stage0_53[345], stage0_53[346], stage0_53[347]},
      {stage1_55[57],stage1_54[93],stage1_53[107],stage1_52[157],stage1_51[218]}
   );
   gpc615_5 gpc2001 (
      {stage0_51[410], stage0_51[411], stage0_51[412], stage0_51[413], stage0_51[414]},
      {stage0_52[274]},
      {stage0_53[348], stage0_53[349], stage0_53[350], stage0_53[351], stage0_53[352], stage0_53[353]},
      {stage1_55[58],stage1_54[94],stage1_53[108],stage1_52[158],stage1_51[219]}
   );
   gpc615_5 gpc2002 (
      {stage0_51[415], stage0_51[416], stage0_51[417], stage0_51[418], stage0_51[419]},
      {stage0_52[275]},
      {stage0_53[354], stage0_53[355], stage0_53[356], stage0_53[357], stage0_53[358], stage0_53[359]},
      {stage1_55[59],stage1_54[95],stage1_53[109],stage1_52[159],stage1_51[220]}
   );
   gpc615_5 gpc2003 (
      {stage0_51[420], stage0_51[421], stage0_51[422], stage0_51[423], stage0_51[424]},
      {stage0_52[276]},
      {stage0_53[360], stage0_53[361], stage0_53[362], stage0_53[363], stage0_53[364], stage0_53[365]},
      {stage1_55[60],stage1_54[96],stage1_53[110],stage1_52[160],stage1_51[221]}
   );
   gpc615_5 gpc2004 (
      {stage0_51[425], stage0_51[426], stage0_51[427], stage0_51[428], stage0_51[429]},
      {stage0_52[277]},
      {stage0_53[366], stage0_53[367], stage0_53[368], stage0_53[369], stage0_53[370], stage0_53[371]},
      {stage1_55[61],stage1_54[97],stage1_53[111],stage1_52[161],stage1_51[222]}
   );
   gpc615_5 gpc2005 (
      {stage0_51[430], stage0_51[431], stage0_51[432], stage0_51[433], stage0_51[434]},
      {stage0_52[278]},
      {stage0_53[372], stage0_53[373], stage0_53[374], stage0_53[375], stage0_53[376], stage0_53[377]},
      {stage1_55[62],stage1_54[98],stage1_53[112],stage1_52[162],stage1_51[223]}
   );
   gpc606_5 gpc2006 (
      {stage0_52[279], stage0_52[280], stage0_52[281], stage0_52[282], stage0_52[283], stage0_52[284]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[63],stage1_54[99],stage1_53[113],stage1_52[163]}
   );
   gpc606_5 gpc2007 (
      {stage0_52[285], stage0_52[286], stage0_52[287], stage0_52[288], stage0_52[289], stage0_52[290]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[64],stage1_54[100],stage1_53[114],stage1_52[164]}
   );
   gpc606_5 gpc2008 (
      {stage0_52[291], stage0_52[292], stage0_52[293], stage0_52[294], stage0_52[295], stage0_52[296]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[65],stage1_54[101],stage1_53[115],stage1_52[165]}
   );
   gpc606_5 gpc2009 (
      {stage0_52[297], stage0_52[298], stage0_52[299], stage0_52[300], stage0_52[301], stage0_52[302]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[66],stage1_54[102],stage1_53[116],stage1_52[166]}
   );
   gpc606_5 gpc2010 (
      {stage0_52[303], stage0_52[304], stage0_52[305], stage0_52[306], stage0_52[307], stage0_52[308]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[67],stage1_54[103],stage1_53[117],stage1_52[167]}
   );
   gpc606_5 gpc2011 (
      {stage0_52[309], stage0_52[310], stage0_52[311], stage0_52[312], stage0_52[313], stage0_52[314]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[68],stage1_54[104],stage1_53[118],stage1_52[168]}
   );
   gpc606_5 gpc2012 (
      {stage0_52[315], stage0_52[316], stage0_52[317], stage0_52[318], stage0_52[319], stage0_52[320]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[69],stage1_54[105],stage1_53[119],stage1_52[169]}
   );
   gpc606_5 gpc2013 (
      {stage0_52[321], stage0_52[322], stage0_52[323], stage0_52[324], stage0_52[325], stage0_52[326]},
      {stage0_54[42], stage0_54[43], stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47]},
      {stage1_56[7],stage1_55[70],stage1_54[106],stage1_53[120],stage1_52[170]}
   );
   gpc606_5 gpc2014 (
      {stage0_52[327], stage0_52[328], stage0_52[329], stage0_52[330], stage0_52[331], stage0_52[332]},
      {stage0_54[48], stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage1_56[8],stage1_55[71],stage1_54[107],stage1_53[121],stage1_52[171]}
   );
   gpc606_5 gpc2015 (
      {stage0_52[333], stage0_52[334], stage0_52[335], stage0_52[336], stage0_52[337], stage0_52[338]},
      {stage0_54[54], stage0_54[55], stage0_54[56], stage0_54[57], stage0_54[58], stage0_54[59]},
      {stage1_56[9],stage1_55[72],stage1_54[108],stage1_53[122],stage1_52[172]}
   );
   gpc606_5 gpc2016 (
      {stage0_52[339], stage0_52[340], stage0_52[341], stage0_52[342], stage0_52[343], stage0_52[344]},
      {stage0_54[60], stage0_54[61], stage0_54[62], stage0_54[63], stage0_54[64], stage0_54[65]},
      {stage1_56[10],stage1_55[73],stage1_54[109],stage1_53[123],stage1_52[173]}
   );
   gpc606_5 gpc2017 (
      {stage0_52[345], stage0_52[346], stage0_52[347], stage0_52[348], stage0_52[349], stage0_52[350]},
      {stage0_54[66], stage0_54[67], stage0_54[68], stage0_54[69], stage0_54[70], stage0_54[71]},
      {stage1_56[11],stage1_55[74],stage1_54[110],stage1_53[124],stage1_52[174]}
   );
   gpc606_5 gpc2018 (
      {stage0_52[351], stage0_52[352], stage0_52[353], stage0_52[354], stage0_52[355], stage0_52[356]},
      {stage0_54[72], stage0_54[73], stage0_54[74], stage0_54[75], stage0_54[76], stage0_54[77]},
      {stage1_56[12],stage1_55[75],stage1_54[111],stage1_53[125],stage1_52[175]}
   );
   gpc606_5 gpc2019 (
      {stage0_52[357], stage0_52[358], stage0_52[359], stage0_52[360], stage0_52[361], stage0_52[362]},
      {stage0_54[78], stage0_54[79], stage0_54[80], stage0_54[81], stage0_54[82], stage0_54[83]},
      {stage1_56[13],stage1_55[76],stage1_54[112],stage1_53[126],stage1_52[176]}
   );
   gpc606_5 gpc2020 (
      {stage0_52[363], stage0_52[364], stage0_52[365], stage0_52[366], stage0_52[367], stage0_52[368]},
      {stage0_54[84], stage0_54[85], stage0_54[86], stage0_54[87], stage0_54[88], stage0_54[89]},
      {stage1_56[14],stage1_55[77],stage1_54[113],stage1_53[127],stage1_52[177]}
   );
   gpc606_5 gpc2021 (
      {stage0_52[369], stage0_52[370], stage0_52[371], stage0_52[372], stage0_52[373], stage0_52[374]},
      {stage0_54[90], stage0_54[91], stage0_54[92], stage0_54[93], stage0_54[94], stage0_54[95]},
      {stage1_56[15],stage1_55[78],stage1_54[114],stage1_53[128],stage1_52[178]}
   );
   gpc606_5 gpc2022 (
      {stage0_52[375], stage0_52[376], stage0_52[377], stage0_52[378], stage0_52[379], stage0_52[380]},
      {stage0_54[96], stage0_54[97], stage0_54[98], stage0_54[99], stage0_54[100], stage0_54[101]},
      {stage1_56[16],stage1_55[79],stage1_54[115],stage1_53[129],stage1_52[179]}
   );
   gpc606_5 gpc2023 (
      {stage0_52[381], stage0_52[382], stage0_52[383], stage0_52[384], stage0_52[385], stage0_52[386]},
      {stage0_54[102], stage0_54[103], stage0_54[104], stage0_54[105], stage0_54[106], stage0_54[107]},
      {stage1_56[17],stage1_55[80],stage1_54[116],stage1_53[130],stage1_52[180]}
   );
   gpc606_5 gpc2024 (
      {stage0_52[387], stage0_52[388], stage0_52[389], stage0_52[390], stage0_52[391], stage0_52[392]},
      {stage0_54[108], stage0_54[109], stage0_54[110], stage0_54[111], stage0_54[112], stage0_54[113]},
      {stage1_56[18],stage1_55[81],stage1_54[117],stage1_53[131],stage1_52[181]}
   );
   gpc606_5 gpc2025 (
      {stage0_52[393], stage0_52[394], stage0_52[395], stage0_52[396], stage0_52[397], stage0_52[398]},
      {stage0_54[114], stage0_54[115], stage0_54[116], stage0_54[117], stage0_54[118], stage0_54[119]},
      {stage1_56[19],stage1_55[82],stage1_54[118],stage1_53[132],stage1_52[182]}
   );
   gpc606_5 gpc2026 (
      {stage0_52[399], stage0_52[400], stage0_52[401], stage0_52[402], stage0_52[403], stage0_52[404]},
      {stage0_54[120], stage0_54[121], stage0_54[122], stage0_54[123], stage0_54[124], stage0_54[125]},
      {stage1_56[20],stage1_55[83],stage1_54[119],stage1_53[133],stage1_52[183]}
   );
   gpc606_5 gpc2027 (
      {stage0_52[405], stage0_52[406], stage0_52[407], stage0_52[408], stage0_52[409], stage0_52[410]},
      {stage0_54[126], stage0_54[127], stage0_54[128], stage0_54[129], stage0_54[130], stage0_54[131]},
      {stage1_56[21],stage1_55[84],stage1_54[120],stage1_53[134],stage1_52[184]}
   );
   gpc606_5 gpc2028 (
      {stage0_52[411], stage0_52[412], stage0_52[413], stage0_52[414], stage0_52[415], stage0_52[416]},
      {stage0_54[132], stage0_54[133], stage0_54[134], stage0_54[135], stage0_54[136], stage0_54[137]},
      {stage1_56[22],stage1_55[85],stage1_54[121],stage1_53[135],stage1_52[185]}
   );
   gpc606_5 gpc2029 (
      {stage0_52[417], stage0_52[418], stage0_52[419], stage0_52[420], stage0_52[421], stage0_52[422]},
      {stage0_54[138], stage0_54[139], stage0_54[140], stage0_54[141], stage0_54[142], stage0_54[143]},
      {stage1_56[23],stage1_55[86],stage1_54[122],stage1_53[136],stage1_52[186]}
   );
   gpc606_5 gpc2030 (
      {stage0_52[423], stage0_52[424], stage0_52[425], stage0_52[426], stage0_52[427], stage0_52[428]},
      {stage0_54[144], stage0_54[145], stage0_54[146], stage0_54[147], stage0_54[148], stage0_54[149]},
      {stage1_56[24],stage1_55[87],stage1_54[123],stage1_53[137],stage1_52[187]}
   );
   gpc606_5 gpc2031 (
      {stage0_52[429], stage0_52[430], stage0_52[431], stage0_52[432], stage0_52[433], stage0_52[434]},
      {stage0_54[150], stage0_54[151], stage0_54[152], stage0_54[153], stage0_54[154], stage0_54[155]},
      {stage1_56[25],stage1_55[88],stage1_54[124],stage1_53[138],stage1_52[188]}
   );
   gpc606_5 gpc2032 (
      {stage0_52[435], stage0_52[436], stage0_52[437], stage0_52[438], stage0_52[439], stage0_52[440]},
      {stage0_54[156], stage0_54[157], stage0_54[158], stage0_54[159], stage0_54[160], stage0_54[161]},
      {stage1_56[26],stage1_55[89],stage1_54[125],stage1_53[139],stage1_52[189]}
   );
   gpc606_5 gpc2033 (
      {stage0_52[441], stage0_52[442], stage0_52[443], stage0_52[444], stage0_52[445], stage0_52[446]},
      {stage0_54[162], stage0_54[163], stage0_54[164], stage0_54[165], stage0_54[166], stage0_54[167]},
      {stage1_56[27],stage1_55[90],stage1_54[126],stage1_53[140],stage1_52[190]}
   );
   gpc615_5 gpc2034 (
      {stage0_52[447], stage0_52[448], stage0_52[449], stage0_52[450], stage0_52[451]},
      {stage0_53[378]},
      {stage0_54[168], stage0_54[169], stage0_54[170], stage0_54[171], stage0_54[172], stage0_54[173]},
      {stage1_56[28],stage1_55[91],stage1_54[127],stage1_53[141],stage1_52[191]}
   );
   gpc615_5 gpc2035 (
      {stage0_52[452], stage0_52[453], stage0_52[454], stage0_52[455], stage0_52[456]},
      {stage0_53[379]},
      {stage0_54[174], stage0_54[175], stage0_54[176], stage0_54[177], stage0_54[178], stage0_54[179]},
      {stage1_56[29],stage1_55[92],stage1_54[128],stage1_53[142],stage1_52[192]}
   );
   gpc615_5 gpc2036 (
      {stage0_52[457], stage0_52[458], stage0_52[459], stage0_52[460], stage0_52[461]},
      {stage0_53[380]},
      {stage0_54[180], stage0_54[181], stage0_54[182], stage0_54[183], stage0_54[184], stage0_54[185]},
      {stage1_56[30],stage1_55[93],stage1_54[129],stage1_53[143],stage1_52[193]}
   );
   gpc615_5 gpc2037 (
      {stage0_52[462], stage0_52[463], stage0_52[464], stage0_52[465], stage0_52[466]},
      {stage0_53[381]},
      {stage0_54[186], stage0_54[187], stage0_54[188], stage0_54[189], stage0_54[190], stage0_54[191]},
      {stage1_56[31],stage1_55[94],stage1_54[130],stage1_53[144],stage1_52[194]}
   );
   gpc615_5 gpc2038 (
      {stage0_52[467], stage0_52[468], stage0_52[469], stage0_52[470], stage0_52[471]},
      {stage0_53[382]},
      {stage0_54[192], stage0_54[193], stage0_54[194], stage0_54[195], stage0_54[196], stage0_54[197]},
      {stage1_56[32],stage1_55[95],stage1_54[131],stage1_53[145],stage1_52[195]}
   );
   gpc615_5 gpc2039 (
      {stage0_52[472], stage0_52[473], stage0_52[474], stage0_52[475], stage0_52[476]},
      {stage0_53[383]},
      {stage0_54[198], stage0_54[199], stage0_54[200], stage0_54[201], stage0_54[202], stage0_54[203]},
      {stage1_56[33],stage1_55[96],stage1_54[132],stage1_53[146],stage1_52[196]}
   );
   gpc615_5 gpc2040 (
      {stage0_52[477], stage0_52[478], stage0_52[479], stage0_52[480], stage0_52[481]},
      {stage0_53[384]},
      {stage0_54[204], stage0_54[205], stage0_54[206], stage0_54[207], stage0_54[208], stage0_54[209]},
      {stage1_56[34],stage1_55[97],stage1_54[133],stage1_53[147],stage1_52[197]}
   );
   gpc615_5 gpc2041 (
      {stage0_52[482], stage0_52[483], stage0_52[484], stage0_52[485], 1'b0},
      {stage0_53[385]},
      {stage0_54[210], stage0_54[211], stage0_54[212], stage0_54[213], stage0_54[214], stage0_54[215]},
      {stage1_56[35],stage1_55[98],stage1_54[134],stage1_53[148],stage1_52[198]}
   );
   gpc615_5 gpc2042 (
      {stage0_53[386], stage0_53[387], stage0_53[388], stage0_53[389], stage0_53[390]},
      {stage0_54[216]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[36],stage1_55[99],stage1_54[135],stage1_53[149]}
   );
   gpc615_5 gpc2043 (
      {stage0_53[391], stage0_53[392], stage0_53[393], stage0_53[394], stage0_53[395]},
      {stage0_54[217]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[37],stage1_55[100],stage1_54[136],stage1_53[150]}
   );
   gpc615_5 gpc2044 (
      {stage0_53[396], stage0_53[397], stage0_53[398], stage0_53[399], stage0_53[400]},
      {stage0_54[218]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[38],stage1_55[101],stage1_54[137],stage1_53[151]}
   );
   gpc615_5 gpc2045 (
      {stage0_53[401], stage0_53[402], stage0_53[403], stage0_53[404], stage0_53[405]},
      {stage0_54[219]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[39],stage1_55[102],stage1_54[138],stage1_53[152]}
   );
   gpc615_5 gpc2046 (
      {stage0_53[406], stage0_53[407], stage0_53[408], stage0_53[409], stage0_53[410]},
      {stage0_54[220]},
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage1_57[4],stage1_56[40],stage1_55[103],stage1_54[139],stage1_53[153]}
   );
   gpc615_5 gpc2047 (
      {stage0_53[411], stage0_53[412], stage0_53[413], stage0_53[414], stage0_53[415]},
      {stage0_54[221]},
      {stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33], stage0_55[34], stage0_55[35]},
      {stage1_57[5],stage1_56[41],stage1_55[104],stage1_54[140],stage1_53[154]}
   );
   gpc615_5 gpc2048 (
      {stage0_53[416], stage0_53[417], stage0_53[418], stage0_53[419], stage0_53[420]},
      {stage0_54[222]},
      {stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39], stage0_55[40], stage0_55[41]},
      {stage1_57[6],stage1_56[42],stage1_55[105],stage1_54[141],stage1_53[155]}
   );
   gpc615_5 gpc2049 (
      {stage0_53[421], stage0_53[422], stage0_53[423], stage0_53[424], stage0_53[425]},
      {stage0_54[223]},
      {stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45], stage0_55[46], stage0_55[47]},
      {stage1_57[7],stage1_56[43],stage1_55[106],stage1_54[142],stage1_53[156]}
   );
   gpc615_5 gpc2050 (
      {stage0_53[426], stage0_53[427], stage0_53[428], stage0_53[429], stage0_53[430]},
      {stage0_54[224]},
      {stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51], stage0_55[52], stage0_55[53]},
      {stage1_57[8],stage1_56[44],stage1_55[107],stage1_54[143],stage1_53[157]}
   );
   gpc615_5 gpc2051 (
      {stage0_53[431], stage0_53[432], stage0_53[433], stage0_53[434], stage0_53[435]},
      {stage0_54[225]},
      {stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57], stage0_55[58], stage0_55[59]},
      {stage1_57[9],stage1_56[45],stage1_55[108],stage1_54[144],stage1_53[158]}
   );
   gpc615_5 gpc2052 (
      {stage0_53[436], stage0_53[437], stage0_53[438], stage0_53[439], stage0_53[440]},
      {stage0_54[226]},
      {stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63], stage0_55[64], stage0_55[65]},
      {stage1_57[10],stage1_56[46],stage1_55[109],stage1_54[145],stage1_53[159]}
   );
   gpc615_5 gpc2053 (
      {stage0_53[441], stage0_53[442], stage0_53[443], stage0_53[444], stage0_53[445]},
      {stage0_54[227]},
      {stage0_55[66], stage0_55[67], stage0_55[68], stage0_55[69], stage0_55[70], stage0_55[71]},
      {stage1_57[11],stage1_56[47],stage1_55[110],stage1_54[146],stage1_53[160]}
   );
   gpc615_5 gpc2054 (
      {stage0_53[446], stage0_53[447], stage0_53[448], stage0_53[449], stage0_53[450]},
      {stage0_54[228]},
      {stage0_55[72], stage0_55[73], stage0_55[74], stage0_55[75], stage0_55[76], stage0_55[77]},
      {stage1_57[12],stage1_56[48],stage1_55[111],stage1_54[147],stage1_53[161]}
   );
   gpc615_5 gpc2055 (
      {stage0_53[451], stage0_53[452], stage0_53[453], stage0_53[454], stage0_53[455]},
      {stage0_54[229]},
      {stage0_55[78], stage0_55[79], stage0_55[80], stage0_55[81], stage0_55[82], stage0_55[83]},
      {stage1_57[13],stage1_56[49],stage1_55[112],stage1_54[148],stage1_53[162]}
   );
   gpc615_5 gpc2056 (
      {stage0_53[456], stage0_53[457], stage0_53[458], stage0_53[459], stage0_53[460]},
      {stage0_54[230]},
      {stage0_55[84], stage0_55[85], stage0_55[86], stage0_55[87], stage0_55[88], stage0_55[89]},
      {stage1_57[14],stage1_56[50],stage1_55[113],stage1_54[149],stage1_53[163]}
   );
   gpc615_5 gpc2057 (
      {stage0_53[461], stage0_53[462], stage0_53[463], stage0_53[464], stage0_53[465]},
      {stage0_54[231]},
      {stage0_55[90], stage0_55[91], stage0_55[92], stage0_55[93], stage0_55[94], stage0_55[95]},
      {stage1_57[15],stage1_56[51],stage1_55[114],stage1_54[150],stage1_53[164]}
   );
   gpc615_5 gpc2058 (
      {stage0_53[466], stage0_53[467], stage0_53[468], stage0_53[469], stage0_53[470]},
      {stage0_54[232]},
      {stage0_55[96], stage0_55[97], stage0_55[98], stage0_55[99], stage0_55[100], stage0_55[101]},
      {stage1_57[16],stage1_56[52],stage1_55[115],stage1_54[151],stage1_53[165]}
   );
   gpc615_5 gpc2059 (
      {stage0_53[471], stage0_53[472], stage0_53[473], stage0_53[474], stage0_53[475]},
      {stage0_54[233]},
      {stage0_55[102], stage0_55[103], stage0_55[104], stage0_55[105], stage0_55[106], stage0_55[107]},
      {stage1_57[17],stage1_56[53],stage1_55[116],stage1_54[152],stage1_53[166]}
   );
   gpc615_5 gpc2060 (
      {stage0_53[476], stage0_53[477], stage0_53[478], stage0_53[479], stage0_53[480]},
      {stage0_54[234]},
      {stage0_55[108], stage0_55[109], stage0_55[110], stage0_55[111], stage0_55[112], stage0_55[113]},
      {stage1_57[18],stage1_56[54],stage1_55[117],stage1_54[153],stage1_53[167]}
   );
   gpc615_5 gpc2061 (
      {stage0_53[481], stage0_53[482], stage0_53[483], stage0_53[484], stage0_53[485]},
      {stage0_54[235]},
      {stage0_55[114], stage0_55[115], stage0_55[116], stage0_55[117], stage0_55[118], stage0_55[119]},
      {stage1_57[19],stage1_56[55],stage1_55[118],stage1_54[154],stage1_53[168]}
   );
   gpc117_4 gpc2062 (
      {stage0_54[236], stage0_54[237], stage0_54[238], stage0_54[239], stage0_54[240], stage0_54[241], stage0_54[242]},
      {stage0_55[120]},
      {stage0_56[0]},
      {stage1_57[20],stage1_56[56],stage1_55[119],stage1_54[155]}
   );
   gpc615_5 gpc2063 (
      {stage0_54[243], stage0_54[244], stage0_54[245], stage0_54[246], stage0_54[247]},
      {stage0_55[121]},
      {stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5], stage0_56[6]},
      {stage1_58[0],stage1_57[21],stage1_56[57],stage1_55[120],stage1_54[156]}
   );
   gpc615_5 gpc2064 (
      {stage0_54[248], stage0_54[249], stage0_54[250], stage0_54[251], stage0_54[252]},
      {stage0_55[122]},
      {stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11], stage0_56[12]},
      {stage1_58[1],stage1_57[22],stage1_56[58],stage1_55[121],stage1_54[157]}
   );
   gpc615_5 gpc2065 (
      {stage0_54[253], stage0_54[254], stage0_54[255], stage0_54[256], stage0_54[257]},
      {stage0_55[123]},
      {stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17], stage0_56[18]},
      {stage1_58[2],stage1_57[23],stage1_56[59],stage1_55[122],stage1_54[158]}
   );
   gpc615_5 gpc2066 (
      {stage0_54[258], stage0_54[259], stage0_54[260], stage0_54[261], stage0_54[262]},
      {stage0_55[124]},
      {stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23], stage0_56[24]},
      {stage1_58[3],stage1_57[24],stage1_56[60],stage1_55[123],stage1_54[159]}
   );
   gpc615_5 gpc2067 (
      {stage0_54[263], stage0_54[264], stage0_54[265], stage0_54[266], stage0_54[267]},
      {stage0_55[125]},
      {stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29], stage0_56[30]},
      {stage1_58[4],stage1_57[25],stage1_56[61],stage1_55[124],stage1_54[160]}
   );
   gpc615_5 gpc2068 (
      {stage0_54[268], stage0_54[269], stage0_54[270], stage0_54[271], stage0_54[272]},
      {stage0_55[126]},
      {stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35], stage0_56[36]},
      {stage1_58[5],stage1_57[26],stage1_56[62],stage1_55[125],stage1_54[161]}
   );
   gpc615_5 gpc2069 (
      {stage0_54[273], stage0_54[274], stage0_54[275], stage0_54[276], stage0_54[277]},
      {stage0_55[127]},
      {stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41], stage0_56[42]},
      {stage1_58[6],stage1_57[27],stage1_56[63],stage1_55[126],stage1_54[162]}
   );
   gpc615_5 gpc2070 (
      {stage0_54[278], stage0_54[279], stage0_54[280], stage0_54[281], stage0_54[282]},
      {stage0_55[128]},
      {stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46], stage0_56[47], stage0_56[48]},
      {stage1_58[7],stage1_57[28],stage1_56[64],stage1_55[127],stage1_54[163]}
   );
   gpc615_5 gpc2071 (
      {stage0_54[283], stage0_54[284], stage0_54[285], stage0_54[286], stage0_54[287]},
      {stage0_55[129]},
      {stage0_56[49], stage0_56[50], stage0_56[51], stage0_56[52], stage0_56[53], stage0_56[54]},
      {stage1_58[8],stage1_57[29],stage1_56[65],stage1_55[128],stage1_54[164]}
   );
   gpc615_5 gpc2072 (
      {stage0_54[288], stage0_54[289], stage0_54[290], stage0_54[291], stage0_54[292]},
      {stage0_55[130]},
      {stage0_56[55], stage0_56[56], stage0_56[57], stage0_56[58], stage0_56[59], stage0_56[60]},
      {stage1_58[9],stage1_57[30],stage1_56[66],stage1_55[129],stage1_54[165]}
   );
   gpc615_5 gpc2073 (
      {stage0_54[293], stage0_54[294], stage0_54[295], stage0_54[296], stage0_54[297]},
      {stage0_55[131]},
      {stage0_56[61], stage0_56[62], stage0_56[63], stage0_56[64], stage0_56[65], stage0_56[66]},
      {stage1_58[10],stage1_57[31],stage1_56[67],stage1_55[130],stage1_54[166]}
   );
   gpc615_5 gpc2074 (
      {stage0_54[298], stage0_54[299], stage0_54[300], stage0_54[301], stage0_54[302]},
      {stage0_55[132]},
      {stage0_56[67], stage0_56[68], stage0_56[69], stage0_56[70], stage0_56[71], stage0_56[72]},
      {stage1_58[11],stage1_57[32],stage1_56[68],stage1_55[131],stage1_54[167]}
   );
   gpc615_5 gpc2075 (
      {stage0_54[303], stage0_54[304], stage0_54[305], stage0_54[306], stage0_54[307]},
      {stage0_55[133]},
      {stage0_56[73], stage0_56[74], stage0_56[75], stage0_56[76], stage0_56[77], stage0_56[78]},
      {stage1_58[12],stage1_57[33],stage1_56[69],stage1_55[132],stage1_54[168]}
   );
   gpc615_5 gpc2076 (
      {stage0_54[308], stage0_54[309], stage0_54[310], stage0_54[311], stage0_54[312]},
      {stage0_55[134]},
      {stage0_56[79], stage0_56[80], stage0_56[81], stage0_56[82], stage0_56[83], stage0_56[84]},
      {stage1_58[13],stage1_57[34],stage1_56[70],stage1_55[133],stage1_54[169]}
   );
   gpc615_5 gpc2077 (
      {stage0_54[313], stage0_54[314], stage0_54[315], stage0_54[316], stage0_54[317]},
      {stage0_55[135]},
      {stage0_56[85], stage0_56[86], stage0_56[87], stage0_56[88], stage0_56[89], stage0_56[90]},
      {stage1_58[14],stage1_57[35],stage1_56[71],stage1_55[134],stage1_54[170]}
   );
   gpc615_5 gpc2078 (
      {stage0_54[318], stage0_54[319], stage0_54[320], stage0_54[321], stage0_54[322]},
      {stage0_55[136]},
      {stage0_56[91], stage0_56[92], stage0_56[93], stage0_56[94], stage0_56[95], stage0_56[96]},
      {stage1_58[15],stage1_57[36],stage1_56[72],stage1_55[135],stage1_54[171]}
   );
   gpc615_5 gpc2079 (
      {stage0_54[323], stage0_54[324], stage0_54[325], stage0_54[326], stage0_54[327]},
      {stage0_55[137]},
      {stage0_56[97], stage0_56[98], stage0_56[99], stage0_56[100], stage0_56[101], stage0_56[102]},
      {stage1_58[16],stage1_57[37],stage1_56[73],stage1_55[136],stage1_54[172]}
   );
   gpc615_5 gpc2080 (
      {stage0_54[328], stage0_54[329], stage0_54[330], stage0_54[331], stage0_54[332]},
      {stage0_55[138]},
      {stage0_56[103], stage0_56[104], stage0_56[105], stage0_56[106], stage0_56[107], stage0_56[108]},
      {stage1_58[17],stage1_57[38],stage1_56[74],stage1_55[137],stage1_54[173]}
   );
   gpc615_5 gpc2081 (
      {stage0_54[333], stage0_54[334], stage0_54[335], stage0_54[336], stage0_54[337]},
      {stage0_55[139]},
      {stage0_56[109], stage0_56[110], stage0_56[111], stage0_56[112], stage0_56[113], stage0_56[114]},
      {stage1_58[18],stage1_57[39],stage1_56[75],stage1_55[138],stage1_54[174]}
   );
   gpc615_5 gpc2082 (
      {stage0_54[338], stage0_54[339], stage0_54[340], stage0_54[341], stage0_54[342]},
      {stage0_55[140]},
      {stage0_56[115], stage0_56[116], stage0_56[117], stage0_56[118], stage0_56[119], stage0_56[120]},
      {stage1_58[19],stage1_57[40],stage1_56[76],stage1_55[139],stage1_54[175]}
   );
   gpc615_5 gpc2083 (
      {stage0_54[343], stage0_54[344], stage0_54[345], stage0_54[346], stage0_54[347]},
      {stage0_55[141]},
      {stage0_56[121], stage0_56[122], stage0_56[123], stage0_56[124], stage0_56[125], stage0_56[126]},
      {stage1_58[20],stage1_57[41],stage1_56[77],stage1_55[140],stage1_54[176]}
   );
   gpc615_5 gpc2084 (
      {stage0_54[348], stage0_54[349], stage0_54[350], stage0_54[351], stage0_54[352]},
      {stage0_55[142]},
      {stage0_56[127], stage0_56[128], stage0_56[129], stage0_56[130], stage0_56[131], stage0_56[132]},
      {stage1_58[21],stage1_57[42],stage1_56[78],stage1_55[141],stage1_54[177]}
   );
   gpc615_5 gpc2085 (
      {stage0_54[353], stage0_54[354], stage0_54[355], stage0_54[356], stage0_54[357]},
      {stage0_55[143]},
      {stage0_56[133], stage0_56[134], stage0_56[135], stage0_56[136], stage0_56[137], stage0_56[138]},
      {stage1_58[22],stage1_57[43],stage1_56[79],stage1_55[142],stage1_54[178]}
   );
   gpc615_5 gpc2086 (
      {stage0_54[358], stage0_54[359], stage0_54[360], stage0_54[361], stage0_54[362]},
      {stage0_55[144]},
      {stage0_56[139], stage0_56[140], stage0_56[141], stage0_56[142], stage0_56[143], stage0_56[144]},
      {stage1_58[23],stage1_57[44],stage1_56[80],stage1_55[143],stage1_54[179]}
   );
   gpc615_5 gpc2087 (
      {stage0_54[363], stage0_54[364], stage0_54[365], stage0_54[366], stage0_54[367]},
      {stage0_55[145]},
      {stage0_56[145], stage0_56[146], stage0_56[147], stage0_56[148], stage0_56[149], stage0_56[150]},
      {stage1_58[24],stage1_57[45],stage1_56[81],stage1_55[144],stage1_54[180]}
   );
   gpc615_5 gpc2088 (
      {stage0_54[368], stage0_54[369], stage0_54[370], stage0_54[371], stage0_54[372]},
      {stage0_55[146]},
      {stage0_56[151], stage0_56[152], stage0_56[153], stage0_56[154], stage0_56[155], stage0_56[156]},
      {stage1_58[25],stage1_57[46],stage1_56[82],stage1_55[145],stage1_54[181]}
   );
   gpc615_5 gpc2089 (
      {stage0_54[373], stage0_54[374], stage0_54[375], stage0_54[376], stage0_54[377]},
      {stage0_55[147]},
      {stage0_56[157], stage0_56[158], stage0_56[159], stage0_56[160], stage0_56[161], stage0_56[162]},
      {stage1_58[26],stage1_57[47],stage1_56[83],stage1_55[146],stage1_54[182]}
   );
   gpc615_5 gpc2090 (
      {stage0_54[378], stage0_54[379], stage0_54[380], stage0_54[381], stage0_54[382]},
      {stage0_55[148]},
      {stage0_56[163], stage0_56[164], stage0_56[165], stage0_56[166], stage0_56[167], stage0_56[168]},
      {stage1_58[27],stage1_57[48],stage1_56[84],stage1_55[147],stage1_54[183]}
   );
   gpc615_5 gpc2091 (
      {stage0_54[383], stage0_54[384], stage0_54[385], stage0_54[386], stage0_54[387]},
      {stage0_55[149]},
      {stage0_56[169], stage0_56[170], stage0_56[171], stage0_56[172], stage0_56[173], stage0_56[174]},
      {stage1_58[28],stage1_57[49],stage1_56[85],stage1_55[148],stage1_54[184]}
   );
   gpc615_5 gpc2092 (
      {stage0_54[388], stage0_54[389], stage0_54[390], stage0_54[391], stage0_54[392]},
      {stage0_55[150]},
      {stage0_56[175], stage0_56[176], stage0_56[177], stage0_56[178], stage0_56[179], stage0_56[180]},
      {stage1_58[29],stage1_57[50],stage1_56[86],stage1_55[149],stage1_54[185]}
   );
   gpc615_5 gpc2093 (
      {stage0_54[393], stage0_54[394], stage0_54[395], stage0_54[396], stage0_54[397]},
      {stage0_55[151]},
      {stage0_56[181], stage0_56[182], stage0_56[183], stage0_56[184], stage0_56[185], stage0_56[186]},
      {stage1_58[30],stage1_57[51],stage1_56[87],stage1_55[150],stage1_54[186]}
   );
   gpc615_5 gpc2094 (
      {stage0_54[398], stage0_54[399], stage0_54[400], stage0_54[401], stage0_54[402]},
      {stage0_55[152]},
      {stage0_56[187], stage0_56[188], stage0_56[189], stage0_56[190], stage0_56[191], stage0_56[192]},
      {stage1_58[31],stage1_57[52],stage1_56[88],stage1_55[151],stage1_54[187]}
   );
   gpc615_5 gpc2095 (
      {stage0_54[403], stage0_54[404], stage0_54[405], stage0_54[406], stage0_54[407]},
      {stage0_55[153]},
      {stage0_56[193], stage0_56[194], stage0_56[195], stage0_56[196], stage0_56[197], stage0_56[198]},
      {stage1_58[32],stage1_57[53],stage1_56[89],stage1_55[152],stage1_54[188]}
   );
   gpc615_5 gpc2096 (
      {stage0_54[408], stage0_54[409], stage0_54[410], stage0_54[411], stage0_54[412]},
      {stage0_55[154]},
      {stage0_56[199], stage0_56[200], stage0_56[201], stage0_56[202], stage0_56[203], stage0_56[204]},
      {stage1_58[33],stage1_57[54],stage1_56[90],stage1_55[153],stage1_54[189]}
   );
   gpc615_5 gpc2097 (
      {stage0_54[413], stage0_54[414], stage0_54[415], stage0_54[416], stage0_54[417]},
      {stage0_55[155]},
      {stage0_56[205], stage0_56[206], stage0_56[207], stage0_56[208], stage0_56[209], stage0_56[210]},
      {stage1_58[34],stage1_57[55],stage1_56[91],stage1_55[154],stage1_54[190]}
   );
   gpc615_5 gpc2098 (
      {stage0_54[418], stage0_54[419], stage0_54[420], stage0_54[421], stage0_54[422]},
      {stage0_55[156]},
      {stage0_56[211], stage0_56[212], stage0_56[213], stage0_56[214], stage0_56[215], stage0_56[216]},
      {stage1_58[35],stage1_57[56],stage1_56[92],stage1_55[155],stage1_54[191]}
   );
   gpc615_5 gpc2099 (
      {stage0_54[423], stage0_54[424], stage0_54[425], stage0_54[426], stage0_54[427]},
      {stage0_55[157]},
      {stage0_56[217], stage0_56[218], stage0_56[219], stage0_56[220], stage0_56[221], stage0_56[222]},
      {stage1_58[36],stage1_57[57],stage1_56[93],stage1_55[156],stage1_54[192]}
   );
   gpc615_5 gpc2100 (
      {stage0_54[428], stage0_54[429], stage0_54[430], stage0_54[431], stage0_54[432]},
      {stage0_55[158]},
      {stage0_56[223], stage0_56[224], stage0_56[225], stage0_56[226], stage0_56[227], stage0_56[228]},
      {stage1_58[37],stage1_57[58],stage1_56[94],stage1_55[157],stage1_54[193]}
   );
   gpc615_5 gpc2101 (
      {stage0_54[433], stage0_54[434], stage0_54[435], stage0_54[436], stage0_54[437]},
      {stage0_55[159]},
      {stage0_56[229], stage0_56[230], stage0_56[231], stage0_56[232], stage0_56[233], stage0_56[234]},
      {stage1_58[38],stage1_57[59],stage1_56[95],stage1_55[158],stage1_54[194]}
   );
   gpc615_5 gpc2102 (
      {stage0_54[438], stage0_54[439], stage0_54[440], stage0_54[441], stage0_54[442]},
      {stage0_55[160]},
      {stage0_56[235], stage0_56[236], stage0_56[237], stage0_56[238], stage0_56[239], stage0_56[240]},
      {stage1_58[39],stage1_57[60],stage1_56[96],stage1_55[159],stage1_54[195]}
   );
   gpc615_5 gpc2103 (
      {stage0_54[443], stage0_54[444], stage0_54[445], stage0_54[446], stage0_54[447]},
      {stage0_55[161]},
      {stage0_56[241], stage0_56[242], stage0_56[243], stage0_56[244], stage0_56[245], stage0_56[246]},
      {stage1_58[40],stage1_57[61],stage1_56[97],stage1_55[160],stage1_54[196]}
   );
   gpc615_5 gpc2104 (
      {stage0_54[448], stage0_54[449], stage0_54[450], stage0_54[451], stage0_54[452]},
      {stage0_55[162]},
      {stage0_56[247], stage0_56[248], stage0_56[249], stage0_56[250], stage0_56[251], stage0_56[252]},
      {stage1_58[41],stage1_57[62],stage1_56[98],stage1_55[161],stage1_54[197]}
   );
   gpc606_5 gpc2105 (
      {stage0_55[163], stage0_55[164], stage0_55[165], stage0_55[166], stage0_55[167], stage0_55[168]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[42],stage1_57[63],stage1_56[99],stage1_55[162]}
   );
   gpc606_5 gpc2106 (
      {stage0_55[169], stage0_55[170], stage0_55[171], stage0_55[172], stage0_55[173], stage0_55[174]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[43],stage1_57[64],stage1_56[100],stage1_55[163]}
   );
   gpc606_5 gpc2107 (
      {stage0_55[175], stage0_55[176], stage0_55[177], stage0_55[178], stage0_55[179], stage0_55[180]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[44],stage1_57[65],stage1_56[101],stage1_55[164]}
   );
   gpc606_5 gpc2108 (
      {stage0_55[181], stage0_55[182], stage0_55[183], stage0_55[184], stage0_55[185], stage0_55[186]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[45],stage1_57[66],stage1_56[102],stage1_55[165]}
   );
   gpc606_5 gpc2109 (
      {stage0_55[187], stage0_55[188], stage0_55[189], stage0_55[190], stage0_55[191], stage0_55[192]},
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage1_59[4],stage1_58[46],stage1_57[67],stage1_56[103],stage1_55[166]}
   );
   gpc606_5 gpc2110 (
      {stage0_55[193], stage0_55[194], stage0_55[195], stage0_55[196], stage0_55[197], stage0_55[198]},
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage1_59[5],stage1_58[47],stage1_57[68],stage1_56[104],stage1_55[167]}
   );
   gpc606_5 gpc2111 (
      {stage0_55[199], stage0_55[200], stage0_55[201], stage0_55[202], stage0_55[203], stage0_55[204]},
      {stage0_57[36], stage0_57[37], stage0_57[38], stage0_57[39], stage0_57[40], stage0_57[41]},
      {stage1_59[6],stage1_58[48],stage1_57[69],stage1_56[105],stage1_55[168]}
   );
   gpc606_5 gpc2112 (
      {stage0_55[205], stage0_55[206], stage0_55[207], stage0_55[208], stage0_55[209], stage0_55[210]},
      {stage0_57[42], stage0_57[43], stage0_57[44], stage0_57[45], stage0_57[46], stage0_57[47]},
      {stage1_59[7],stage1_58[49],stage1_57[70],stage1_56[106],stage1_55[169]}
   );
   gpc606_5 gpc2113 (
      {stage0_55[211], stage0_55[212], stage0_55[213], stage0_55[214], stage0_55[215], stage0_55[216]},
      {stage0_57[48], stage0_57[49], stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53]},
      {stage1_59[8],stage1_58[50],stage1_57[71],stage1_56[107],stage1_55[170]}
   );
   gpc606_5 gpc2114 (
      {stage0_55[217], stage0_55[218], stage0_55[219], stage0_55[220], stage0_55[221], stage0_55[222]},
      {stage0_57[54], stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage1_59[9],stage1_58[51],stage1_57[72],stage1_56[108],stage1_55[171]}
   );
   gpc606_5 gpc2115 (
      {stage0_55[223], stage0_55[224], stage0_55[225], stage0_55[226], stage0_55[227], stage0_55[228]},
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], stage0_57[64], stage0_57[65]},
      {stage1_59[10],stage1_58[52],stage1_57[73],stage1_56[109],stage1_55[172]}
   );
   gpc606_5 gpc2116 (
      {stage0_55[229], stage0_55[230], stage0_55[231], stage0_55[232], stage0_55[233], stage0_55[234]},
      {stage0_57[66], stage0_57[67], stage0_57[68], stage0_57[69], stage0_57[70], stage0_57[71]},
      {stage1_59[11],stage1_58[53],stage1_57[74],stage1_56[110],stage1_55[173]}
   );
   gpc606_5 gpc2117 (
      {stage0_55[235], stage0_55[236], stage0_55[237], stage0_55[238], stage0_55[239], stage0_55[240]},
      {stage0_57[72], stage0_57[73], stage0_57[74], stage0_57[75], stage0_57[76], stage0_57[77]},
      {stage1_59[12],stage1_58[54],stage1_57[75],stage1_56[111],stage1_55[174]}
   );
   gpc606_5 gpc2118 (
      {stage0_55[241], stage0_55[242], stage0_55[243], stage0_55[244], stage0_55[245], stage0_55[246]},
      {stage0_57[78], stage0_57[79], stage0_57[80], stage0_57[81], stage0_57[82], stage0_57[83]},
      {stage1_59[13],stage1_58[55],stage1_57[76],stage1_56[112],stage1_55[175]}
   );
   gpc606_5 gpc2119 (
      {stage0_55[247], stage0_55[248], stage0_55[249], stage0_55[250], stage0_55[251], stage0_55[252]},
      {stage0_57[84], stage0_57[85], stage0_57[86], stage0_57[87], stage0_57[88], stage0_57[89]},
      {stage1_59[14],stage1_58[56],stage1_57[77],stage1_56[113],stage1_55[176]}
   );
   gpc606_5 gpc2120 (
      {stage0_55[253], stage0_55[254], stage0_55[255], stage0_55[256], stage0_55[257], stage0_55[258]},
      {stage0_57[90], stage0_57[91], stage0_57[92], stage0_57[93], stage0_57[94], stage0_57[95]},
      {stage1_59[15],stage1_58[57],stage1_57[78],stage1_56[114],stage1_55[177]}
   );
   gpc606_5 gpc2121 (
      {stage0_55[259], stage0_55[260], stage0_55[261], stage0_55[262], stage0_55[263], stage0_55[264]},
      {stage0_57[96], stage0_57[97], stage0_57[98], stage0_57[99], stage0_57[100], stage0_57[101]},
      {stage1_59[16],stage1_58[58],stage1_57[79],stage1_56[115],stage1_55[178]}
   );
   gpc606_5 gpc2122 (
      {stage0_55[265], stage0_55[266], stage0_55[267], stage0_55[268], stage0_55[269], stage0_55[270]},
      {stage0_57[102], stage0_57[103], stage0_57[104], stage0_57[105], stage0_57[106], stage0_57[107]},
      {stage1_59[17],stage1_58[59],stage1_57[80],stage1_56[116],stage1_55[179]}
   );
   gpc606_5 gpc2123 (
      {stage0_55[271], stage0_55[272], stage0_55[273], stage0_55[274], stage0_55[275], stage0_55[276]},
      {stage0_57[108], stage0_57[109], stage0_57[110], stage0_57[111], stage0_57[112], stage0_57[113]},
      {stage1_59[18],stage1_58[60],stage1_57[81],stage1_56[117],stage1_55[180]}
   );
   gpc606_5 gpc2124 (
      {stage0_55[277], stage0_55[278], stage0_55[279], stage0_55[280], stage0_55[281], stage0_55[282]},
      {stage0_57[114], stage0_57[115], stage0_57[116], stage0_57[117], stage0_57[118], stage0_57[119]},
      {stage1_59[19],stage1_58[61],stage1_57[82],stage1_56[118],stage1_55[181]}
   );
   gpc606_5 gpc2125 (
      {stage0_55[283], stage0_55[284], stage0_55[285], stage0_55[286], stage0_55[287], stage0_55[288]},
      {stage0_57[120], stage0_57[121], stage0_57[122], stage0_57[123], stage0_57[124], stage0_57[125]},
      {stage1_59[20],stage1_58[62],stage1_57[83],stage1_56[119],stage1_55[182]}
   );
   gpc606_5 gpc2126 (
      {stage0_55[289], stage0_55[290], stage0_55[291], stage0_55[292], stage0_55[293], stage0_55[294]},
      {stage0_57[126], stage0_57[127], stage0_57[128], stage0_57[129], stage0_57[130], stage0_57[131]},
      {stage1_59[21],stage1_58[63],stage1_57[84],stage1_56[120],stage1_55[183]}
   );
   gpc606_5 gpc2127 (
      {stage0_55[295], stage0_55[296], stage0_55[297], stage0_55[298], stage0_55[299], stage0_55[300]},
      {stage0_57[132], stage0_57[133], stage0_57[134], stage0_57[135], stage0_57[136], stage0_57[137]},
      {stage1_59[22],stage1_58[64],stage1_57[85],stage1_56[121],stage1_55[184]}
   );
   gpc606_5 gpc2128 (
      {stage0_55[301], stage0_55[302], stage0_55[303], stage0_55[304], stage0_55[305], stage0_55[306]},
      {stage0_57[138], stage0_57[139], stage0_57[140], stage0_57[141], stage0_57[142], stage0_57[143]},
      {stage1_59[23],stage1_58[65],stage1_57[86],stage1_56[122],stage1_55[185]}
   );
   gpc606_5 gpc2129 (
      {stage0_55[307], stage0_55[308], stage0_55[309], stage0_55[310], stage0_55[311], stage0_55[312]},
      {stage0_57[144], stage0_57[145], stage0_57[146], stage0_57[147], stage0_57[148], stage0_57[149]},
      {stage1_59[24],stage1_58[66],stage1_57[87],stage1_56[123],stage1_55[186]}
   );
   gpc606_5 gpc2130 (
      {stage0_55[313], stage0_55[314], stage0_55[315], stage0_55[316], stage0_55[317], stage0_55[318]},
      {stage0_57[150], stage0_57[151], stage0_57[152], stage0_57[153], stage0_57[154], stage0_57[155]},
      {stage1_59[25],stage1_58[67],stage1_57[88],stage1_56[124],stage1_55[187]}
   );
   gpc606_5 gpc2131 (
      {stage0_55[319], stage0_55[320], stage0_55[321], stage0_55[322], stage0_55[323], stage0_55[324]},
      {stage0_57[156], stage0_57[157], stage0_57[158], stage0_57[159], stage0_57[160], stage0_57[161]},
      {stage1_59[26],stage1_58[68],stage1_57[89],stage1_56[125],stage1_55[188]}
   );
   gpc606_5 gpc2132 (
      {stage0_55[325], stage0_55[326], stage0_55[327], stage0_55[328], stage0_55[329], stage0_55[330]},
      {stage0_57[162], stage0_57[163], stage0_57[164], stage0_57[165], stage0_57[166], stage0_57[167]},
      {stage1_59[27],stage1_58[69],stage1_57[90],stage1_56[126],stage1_55[189]}
   );
   gpc606_5 gpc2133 (
      {stage0_55[331], stage0_55[332], stage0_55[333], stage0_55[334], stage0_55[335], stage0_55[336]},
      {stage0_57[168], stage0_57[169], stage0_57[170], stage0_57[171], stage0_57[172], stage0_57[173]},
      {stage1_59[28],stage1_58[70],stage1_57[91],stage1_56[127],stage1_55[190]}
   );
   gpc606_5 gpc2134 (
      {stage0_55[337], stage0_55[338], stage0_55[339], stage0_55[340], stage0_55[341], stage0_55[342]},
      {stage0_57[174], stage0_57[175], stage0_57[176], stage0_57[177], stage0_57[178], stage0_57[179]},
      {stage1_59[29],stage1_58[71],stage1_57[92],stage1_56[128],stage1_55[191]}
   );
   gpc606_5 gpc2135 (
      {stage0_55[343], stage0_55[344], stage0_55[345], stage0_55[346], stage0_55[347], stage0_55[348]},
      {stage0_57[180], stage0_57[181], stage0_57[182], stage0_57[183], stage0_57[184], stage0_57[185]},
      {stage1_59[30],stage1_58[72],stage1_57[93],stage1_56[129],stage1_55[192]}
   );
   gpc606_5 gpc2136 (
      {stage0_55[349], stage0_55[350], stage0_55[351], stage0_55[352], stage0_55[353], stage0_55[354]},
      {stage0_57[186], stage0_57[187], stage0_57[188], stage0_57[189], stage0_57[190], stage0_57[191]},
      {stage1_59[31],stage1_58[73],stage1_57[94],stage1_56[130],stage1_55[193]}
   );
   gpc606_5 gpc2137 (
      {stage0_55[355], stage0_55[356], stage0_55[357], stage0_55[358], stage0_55[359], stage0_55[360]},
      {stage0_57[192], stage0_57[193], stage0_57[194], stage0_57[195], stage0_57[196], stage0_57[197]},
      {stage1_59[32],stage1_58[74],stage1_57[95],stage1_56[131],stage1_55[194]}
   );
   gpc606_5 gpc2138 (
      {stage0_55[361], stage0_55[362], stage0_55[363], stage0_55[364], stage0_55[365], stage0_55[366]},
      {stage0_57[198], stage0_57[199], stage0_57[200], stage0_57[201], stage0_57[202], stage0_57[203]},
      {stage1_59[33],stage1_58[75],stage1_57[96],stage1_56[132],stage1_55[195]}
   );
   gpc606_5 gpc2139 (
      {stage0_55[367], stage0_55[368], stage0_55[369], stage0_55[370], stage0_55[371], stage0_55[372]},
      {stage0_57[204], stage0_57[205], stage0_57[206], stage0_57[207], stage0_57[208], stage0_57[209]},
      {stage1_59[34],stage1_58[76],stage1_57[97],stage1_56[133],stage1_55[196]}
   );
   gpc606_5 gpc2140 (
      {stage0_55[373], stage0_55[374], stage0_55[375], stage0_55[376], stage0_55[377], stage0_55[378]},
      {stage0_57[210], stage0_57[211], stage0_57[212], stage0_57[213], stage0_57[214], stage0_57[215]},
      {stage1_59[35],stage1_58[77],stage1_57[98],stage1_56[134],stage1_55[197]}
   );
   gpc606_5 gpc2141 (
      {stage0_55[379], stage0_55[380], stage0_55[381], stage0_55[382], stage0_55[383], stage0_55[384]},
      {stage0_57[216], stage0_57[217], stage0_57[218], stage0_57[219], stage0_57[220], stage0_57[221]},
      {stage1_59[36],stage1_58[78],stage1_57[99],stage1_56[135],stage1_55[198]}
   );
   gpc606_5 gpc2142 (
      {stage0_55[385], stage0_55[386], stage0_55[387], stage0_55[388], stage0_55[389], stage0_55[390]},
      {stage0_57[222], stage0_57[223], stage0_57[224], stage0_57[225], stage0_57[226], stage0_57[227]},
      {stage1_59[37],stage1_58[79],stage1_57[100],stage1_56[136],stage1_55[199]}
   );
   gpc606_5 gpc2143 (
      {stage0_55[391], stage0_55[392], stage0_55[393], stage0_55[394], stage0_55[395], stage0_55[396]},
      {stage0_57[228], stage0_57[229], stage0_57[230], stage0_57[231], stage0_57[232], stage0_57[233]},
      {stage1_59[38],stage1_58[80],stage1_57[101],stage1_56[137],stage1_55[200]}
   );
   gpc606_5 gpc2144 (
      {stage0_55[397], stage0_55[398], stage0_55[399], stage0_55[400], stage0_55[401], stage0_55[402]},
      {stage0_57[234], stage0_57[235], stage0_57[236], stage0_57[237], stage0_57[238], stage0_57[239]},
      {stage1_59[39],stage1_58[81],stage1_57[102],stage1_56[138],stage1_55[201]}
   );
   gpc606_5 gpc2145 (
      {stage0_55[403], stage0_55[404], stage0_55[405], stage0_55[406], stage0_55[407], stage0_55[408]},
      {stage0_57[240], stage0_57[241], stage0_57[242], stage0_57[243], stage0_57[244], stage0_57[245]},
      {stage1_59[40],stage1_58[82],stage1_57[103],stage1_56[139],stage1_55[202]}
   );
   gpc606_5 gpc2146 (
      {stage0_55[409], stage0_55[410], stage0_55[411], stage0_55[412], stage0_55[413], stage0_55[414]},
      {stage0_57[246], stage0_57[247], stage0_57[248], stage0_57[249], stage0_57[250], stage0_57[251]},
      {stage1_59[41],stage1_58[83],stage1_57[104],stage1_56[140],stage1_55[203]}
   );
   gpc615_5 gpc2147 (
      {stage0_55[415], stage0_55[416], stage0_55[417], stage0_55[418], stage0_55[419]},
      {stage0_56[253]},
      {stage0_57[252], stage0_57[253], stage0_57[254], stage0_57[255], stage0_57[256], stage0_57[257]},
      {stage1_59[42],stage1_58[84],stage1_57[105],stage1_56[141],stage1_55[204]}
   );
   gpc615_5 gpc2148 (
      {stage0_55[420], stage0_55[421], stage0_55[422], stage0_55[423], stage0_55[424]},
      {stage0_56[254]},
      {stage0_57[258], stage0_57[259], stage0_57[260], stage0_57[261], stage0_57[262], stage0_57[263]},
      {stage1_59[43],stage1_58[85],stage1_57[106],stage1_56[142],stage1_55[205]}
   );
   gpc606_5 gpc2149 (
      {stage0_56[255], stage0_56[256], stage0_56[257], stage0_56[258], stage0_56[259], stage0_56[260]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[44],stage1_58[86],stage1_57[107],stage1_56[143]}
   );
   gpc606_5 gpc2150 (
      {stage0_56[261], stage0_56[262], stage0_56[263], stage0_56[264], stage0_56[265], stage0_56[266]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[45],stage1_58[87],stage1_57[108],stage1_56[144]}
   );
   gpc606_5 gpc2151 (
      {stage0_56[267], stage0_56[268], stage0_56[269], stage0_56[270], stage0_56[271], stage0_56[272]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[46],stage1_58[88],stage1_57[109],stage1_56[145]}
   );
   gpc606_5 gpc2152 (
      {stage0_56[273], stage0_56[274], stage0_56[275], stage0_56[276], stage0_56[277], stage0_56[278]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[47],stage1_58[89],stage1_57[110],stage1_56[146]}
   );
   gpc606_5 gpc2153 (
      {stage0_56[279], stage0_56[280], stage0_56[281], stage0_56[282], stage0_56[283], stage0_56[284]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[48],stage1_58[90],stage1_57[111],stage1_56[147]}
   );
   gpc606_5 gpc2154 (
      {stage0_56[285], stage0_56[286], stage0_56[287], stage0_56[288], stage0_56[289], stage0_56[290]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[49],stage1_58[91],stage1_57[112],stage1_56[148]}
   );
   gpc606_5 gpc2155 (
      {stage0_56[291], stage0_56[292], stage0_56[293], stage0_56[294], stage0_56[295], stage0_56[296]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[50],stage1_58[92],stage1_57[113],stage1_56[149]}
   );
   gpc606_5 gpc2156 (
      {stage0_56[297], stage0_56[298], stage0_56[299], stage0_56[300], stage0_56[301], stage0_56[302]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[51],stage1_58[93],stage1_57[114],stage1_56[150]}
   );
   gpc606_5 gpc2157 (
      {stage0_56[303], stage0_56[304], stage0_56[305], stage0_56[306], stage0_56[307], stage0_56[308]},
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage1_60[8],stage1_59[52],stage1_58[94],stage1_57[115],stage1_56[151]}
   );
   gpc606_5 gpc2158 (
      {stage0_56[309], stage0_56[310], stage0_56[311], stage0_56[312], stage0_56[313], stage0_56[314]},
      {stage0_58[54], stage0_58[55], stage0_58[56], stage0_58[57], stage0_58[58], stage0_58[59]},
      {stage1_60[9],stage1_59[53],stage1_58[95],stage1_57[116],stage1_56[152]}
   );
   gpc606_5 gpc2159 (
      {stage0_56[315], stage0_56[316], stage0_56[317], stage0_56[318], stage0_56[319], stage0_56[320]},
      {stage0_58[60], stage0_58[61], stage0_58[62], stage0_58[63], stage0_58[64], stage0_58[65]},
      {stage1_60[10],stage1_59[54],stage1_58[96],stage1_57[117],stage1_56[153]}
   );
   gpc615_5 gpc2160 (
      {stage0_56[321], stage0_56[322], stage0_56[323], stage0_56[324], stage0_56[325]},
      {stage0_57[264]},
      {stage0_58[66], stage0_58[67], stage0_58[68], stage0_58[69], stage0_58[70], stage0_58[71]},
      {stage1_60[11],stage1_59[55],stage1_58[97],stage1_57[118],stage1_56[154]}
   );
   gpc615_5 gpc2161 (
      {stage0_56[326], stage0_56[327], stage0_56[328], stage0_56[329], stage0_56[330]},
      {stage0_57[265]},
      {stage0_58[72], stage0_58[73], stage0_58[74], stage0_58[75], stage0_58[76], stage0_58[77]},
      {stage1_60[12],stage1_59[56],stage1_58[98],stage1_57[119],stage1_56[155]}
   );
   gpc615_5 gpc2162 (
      {stage0_56[331], stage0_56[332], stage0_56[333], stage0_56[334], stage0_56[335]},
      {stage0_57[266]},
      {stage0_58[78], stage0_58[79], stage0_58[80], stage0_58[81], stage0_58[82], stage0_58[83]},
      {stage1_60[13],stage1_59[57],stage1_58[99],stage1_57[120],stage1_56[156]}
   );
   gpc615_5 gpc2163 (
      {stage0_56[336], stage0_56[337], stage0_56[338], stage0_56[339], stage0_56[340]},
      {stage0_57[267]},
      {stage0_58[84], stage0_58[85], stage0_58[86], stage0_58[87], stage0_58[88], stage0_58[89]},
      {stage1_60[14],stage1_59[58],stage1_58[100],stage1_57[121],stage1_56[157]}
   );
   gpc615_5 gpc2164 (
      {stage0_56[341], stage0_56[342], stage0_56[343], stage0_56[344], stage0_56[345]},
      {stage0_57[268]},
      {stage0_58[90], stage0_58[91], stage0_58[92], stage0_58[93], stage0_58[94], stage0_58[95]},
      {stage1_60[15],stage1_59[59],stage1_58[101],stage1_57[122],stage1_56[158]}
   );
   gpc615_5 gpc2165 (
      {stage0_56[346], stage0_56[347], stage0_56[348], stage0_56[349], stage0_56[350]},
      {stage0_57[269]},
      {stage0_58[96], stage0_58[97], stage0_58[98], stage0_58[99], stage0_58[100], stage0_58[101]},
      {stage1_60[16],stage1_59[60],stage1_58[102],stage1_57[123],stage1_56[159]}
   );
   gpc615_5 gpc2166 (
      {stage0_56[351], stage0_56[352], stage0_56[353], stage0_56[354], stage0_56[355]},
      {stage0_57[270]},
      {stage0_58[102], stage0_58[103], stage0_58[104], stage0_58[105], stage0_58[106], stage0_58[107]},
      {stage1_60[17],stage1_59[61],stage1_58[103],stage1_57[124],stage1_56[160]}
   );
   gpc615_5 gpc2167 (
      {stage0_56[356], stage0_56[357], stage0_56[358], stage0_56[359], stage0_56[360]},
      {stage0_57[271]},
      {stage0_58[108], stage0_58[109], stage0_58[110], stage0_58[111], stage0_58[112], stage0_58[113]},
      {stage1_60[18],stage1_59[62],stage1_58[104],stage1_57[125],stage1_56[161]}
   );
   gpc615_5 gpc2168 (
      {stage0_56[361], stage0_56[362], stage0_56[363], stage0_56[364], stage0_56[365]},
      {stage0_57[272]},
      {stage0_58[114], stage0_58[115], stage0_58[116], stage0_58[117], stage0_58[118], stage0_58[119]},
      {stage1_60[19],stage1_59[63],stage1_58[105],stage1_57[126],stage1_56[162]}
   );
   gpc615_5 gpc2169 (
      {stage0_56[366], stage0_56[367], stage0_56[368], stage0_56[369], stage0_56[370]},
      {stage0_57[273]},
      {stage0_58[120], stage0_58[121], stage0_58[122], stage0_58[123], stage0_58[124], stage0_58[125]},
      {stage1_60[20],stage1_59[64],stage1_58[106],stage1_57[127],stage1_56[163]}
   );
   gpc615_5 gpc2170 (
      {stage0_56[371], stage0_56[372], stage0_56[373], stage0_56[374], stage0_56[375]},
      {stage0_57[274]},
      {stage0_58[126], stage0_58[127], stage0_58[128], stage0_58[129], stage0_58[130], stage0_58[131]},
      {stage1_60[21],stage1_59[65],stage1_58[107],stage1_57[128],stage1_56[164]}
   );
   gpc615_5 gpc2171 (
      {stage0_56[376], stage0_56[377], stage0_56[378], stage0_56[379], stage0_56[380]},
      {stage0_57[275]},
      {stage0_58[132], stage0_58[133], stage0_58[134], stage0_58[135], stage0_58[136], stage0_58[137]},
      {stage1_60[22],stage1_59[66],stage1_58[108],stage1_57[129],stage1_56[165]}
   );
   gpc615_5 gpc2172 (
      {stage0_56[381], stage0_56[382], stage0_56[383], stage0_56[384], stage0_56[385]},
      {stage0_57[276]},
      {stage0_58[138], stage0_58[139], stage0_58[140], stage0_58[141], stage0_58[142], stage0_58[143]},
      {stage1_60[23],stage1_59[67],stage1_58[109],stage1_57[130],stage1_56[166]}
   );
   gpc615_5 gpc2173 (
      {stage0_56[386], stage0_56[387], stage0_56[388], stage0_56[389], stage0_56[390]},
      {stage0_57[277]},
      {stage0_58[144], stage0_58[145], stage0_58[146], stage0_58[147], stage0_58[148], stage0_58[149]},
      {stage1_60[24],stage1_59[68],stage1_58[110],stage1_57[131],stage1_56[167]}
   );
   gpc615_5 gpc2174 (
      {stage0_56[391], stage0_56[392], stage0_56[393], stage0_56[394], stage0_56[395]},
      {stage0_57[278]},
      {stage0_58[150], stage0_58[151], stage0_58[152], stage0_58[153], stage0_58[154], stage0_58[155]},
      {stage1_60[25],stage1_59[69],stage1_58[111],stage1_57[132],stage1_56[168]}
   );
   gpc615_5 gpc2175 (
      {stage0_56[396], stage0_56[397], stage0_56[398], stage0_56[399], stage0_56[400]},
      {stage0_57[279]},
      {stage0_58[156], stage0_58[157], stage0_58[158], stage0_58[159], stage0_58[160], stage0_58[161]},
      {stage1_60[26],stage1_59[70],stage1_58[112],stage1_57[133],stage1_56[169]}
   );
   gpc615_5 gpc2176 (
      {stage0_56[401], stage0_56[402], stage0_56[403], stage0_56[404], stage0_56[405]},
      {stage0_57[280]},
      {stage0_58[162], stage0_58[163], stage0_58[164], stage0_58[165], stage0_58[166], stage0_58[167]},
      {stage1_60[27],stage1_59[71],stage1_58[113],stage1_57[134],stage1_56[170]}
   );
   gpc615_5 gpc2177 (
      {stage0_56[406], stage0_56[407], stage0_56[408], stage0_56[409], stage0_56[410]},
      {stage0_57[281]},
      {stage0_58[168], stage0_58[169], stage0_58[170], stage0_58[171], stage0_58[172], stage0_58[173]},
      {stage1_60[28],stage1_59[72],stage1_58[114],stage1_57[135],stage1_56[171]}
   );
   gpc615_5 gpc2178 (
      {stage0_56[411], stage0_56[412], stage0_56[413], stage0_56[414], stage0_56[415]},
      {stage0_57[282]},
      {stage0_58[174], stage0_58[175], stage0_58[176], stage0_58[177], stage0_58[178], stage0_58[179]},
      {stage1_60[29],stage1_59[73],stage1_58[115],stage1_57[136],stage1_56[172]}
   );
   gpc615_5 gpc2179 (
      {stage0_56[416], stage0_56[417], stage0_56[418], stage0_56[419], stage0_56[420]},
      {stage0_57[283]},
      {stage0_58[180], stage0_58[181], stage0_58[182], stage0_58[183], stage0_58[184], stage0_58[185]},
      {stage1_60[30],stage1_59[74],stage1_58[116],stage1_57[137],stage1_56[173]}
   );
   gpc615_5 gpc2180 (
      {stage0_56[421], stage0_56[422], stage0_56[423], stage0_56[424], stage0_56[425]},
      {stage0_57[284]},
      {stage0_58[186], stage0_58[187], stage0_58[188], stage0_58[189], stage0_58[190], stage0_58[191]},
      {stage1_60[31],stage1_59[75],stage1_58[117],stage1_57[138],stage1_56[174]}
   );
   gpc615_5 gpc2181 (
      {stage0_56[426], stage0_56[427], stage0_56[428], stage0_56[429], stage0_56[430]},
      {stage0_57[285]},
      {stage0_58[192], stage0_58[193], stage0_58[194], stage0_58[195], stage0_58[196], stage0_58[197]},
      {stage1_60[32],stage1_59[76],stage1_58[118],stage1_57[139],stage1_56[175]}
   );
   gpc615_5 gpc2182 (
      {stage0_56[431], stage0_56[432], stage0_56[433], stage0_56[434], stage0_56[435]},
      {stage0_57[286]},
      {stage0_58[198], stage0_58[199], stage0_58[200], stage0_58[201], stage0_58[202], stage0_58[203]},
      {stage1_60[33],stage1_59[77],stage1_58[119],stage1_57[140],stage1_56[176]}
   );
   gpc615_5 gpc2183 (
      {stage0_56[436], stage0_56[437], stage0_56[438], stage0_56[439], stage0_56[440]},
      {stage0_57[287]},
      {stage0_58[204], stage0_58[205], stage0_58[206], stage0_58[207], stage0_58[208], stage0_58[209]},
      {stage1_60[34],stage1_59[78],stage1_58[120],stage1_57[141],stage1_56[177]}
   );
   gpc615_5 gpc2184 (
      {stage0_56[441], stage0_56[442], stage0_56[443], stage0_56[444], stage0_56[445]},
      {stage0_57[288]},
      {stage0_58[210], stage0_58[211], stage0_58[212], stage0_58[213], stage0_58[214], stage0_58[215]},
      {stage1_60[35],stage1_59[79],stage1_58[121],stage1_57[142],stage1_56[178]}
   );
   gpc615_5 gpc2185 (
      {stage0_56[446], stage0_56[447], stage0_56[448], stage0_56[449], stage0_56[450]},
      {stage0_57[289]},
      {stage0_58[216], stage0_58[217], stage0_58[218], stage0_58[219], stage0_58[220], stage0_58[221]},
      {stage1_60[36],stage1_59[80],stage1_58[122],stage1_57[143],stage1_56[179]}
   );
   gpc615_5 gpc2186 (
      {stage0_56[451], stage0_56[452], stage0_56[453], stage0_56[454], stage0_56[455]},
      {stage0_57[290]},
      {stage0_58[222], stage0_58[223], stage0_58[224], stage0_58[225], stage0_58[226], stage0_58[227]},
      {stage1_60[37],stage1_59[81],stage1_58[123],stage1_57[144],stage1_56[180]}
   );
   gpc615_5 gpc2187 (
      {stage0_56[456], stage0_56[457], stage0_56[458], stage0_56[459], stage0_56[460]},
      {stage0_57[291]},
      {stage0_58[228], stage0_58[229], stage0_58[230], stage0_58[231], stage0_58[232], stage0_58[233]},
      {stage1_60[38],stage1_59[82],stage1_58[124],stage1_57[145],stage1_56[181]}
   );
   gpc615_5 gpc2188 (
      {stage0_56[461], stage0_56[462], stage0_56[463], stage0_56[464], stage0_56[465]},
      {stage0_57[292]},
      {stage0_58[234], stage0_58[235], stage0_58[236], stage0_58[237], stage0_58[238], stage0_58[239]},
      {stage1_60[39],stage1_59[83],stage1_58[125],stage1_57[146],stage1_56[182]}
   );
   gpc615_5 gpc2189 (
      {stage0_56[466], stage0_56[467], stage0_56[468], stage0_56[469], stage0_56[470]},
      {stage0_57[293]},
      {stage0_58[240], stage0_58[241], stage0_58[242], stage0_58[243], stage0_58[244], stage0_58[245]},
      {stage1_60[40],stage1_59[84],stage1_58[126],stage1_57[147],stage1_56[183]}
   );
   gpc615_5 gpc2190 (
      {stage0_56[471], stage0_56[472], stage0_56[473], stage0_56[474], stage0_56[475]},
      {stage0_57[294]},
      {stage0_58[246], stage0_58[247], stage0_58[248], stage0_58[249], stage0_58[250], stage0_58[251]},
      {stage1_60[41],stage1_59[85],stage1_58[127],stage1_57[148],stage1_56[184]}
   );
   gpc615_5 gpc2191 (
      {stage0_56[476], stage0_56[477], stage0_56[478], stage0_56[479], stage0_56[480]},
      {stage0_57[295]},
      {stage0_58[252], stage0_58[253], stage0_58[254], stage0_58[255], stage0_58[256], stage0_58[257]},
      {stage1_60[42],stage1_59[86],stage1_58[128],stage1_57[149],stage1_56[185]}
   );
   gpc615_5 gpc2192 (
      {stage0_56[481], stage0_56[482], stage0_56[483], stage0_56[484], stage0_56[485]},
      {stage0_57[296]},
      {stage0_58[258], stage0_58[259], stage0_58[260], stage0_58[261], stage0_58[262], stage0_58[263]},
      {stage1_60[43],stage1_59[87],stage1_58[129],stage1_57[150],stage1_56[186]}
   );
   gpc615_5 gpc2193 (
      {stage0_57[297], stage0_57[298], stage0_57[299], stage0_57[300], stage0_57[301]},
      {stage0_58[264]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[44],stage1_59[88],stage1_58[130],stage1_57[151]}
   );
   gpc615_5 gpc2194 (
      {stage0_57[302], stage0_57[303], stage0_57[304], stage0_57[305], stage0_57[306]},
      {stage0_58[265]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[45],stage1_59[89],stage1_58[131],stage1_57[152]}
   );
   gpc615_5 gpc2195 (
      {stage0_57[307], stage0_57[308], stage0_57[309], stage0_57[310], stage0_57[311]},
      {stage0_58[266]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[46],stage1_59[90],stage1_58[132],stage1_57[153]}
   );
   gpc615_5 gpc2196 (
      {stage0_57[312], stage0_57[313], stage0_57[314], stage0_57[315], stage0_57[316]},
      {stage0_58[267]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[47],stage1_59[91],stage1_58[133],stage1_57[154]}
   );
   gpc615_5 gpc2197 (
      {stage0_57[317], stage0_57[318], stage0_57[319], stage0_57[320], stage0_57[321]},
      {stage0_58[268]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[48],stage1_59[92],stage1_58[134],stage1_57[155]}
   );
   gpc615_5 gpc2198 (
      {stage0_57[322], stage0_57[323], stage0_57[324], stage0_57[325], stage0_57[326]},
      {stage0_58[269]},
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage1_61[5],stage1_60[49],stage1_59[93],stage1_58[135],stage1_57[156]}
   );
   gpc615_5 gpc2199 (
      {stage0_57[327], stage0_57[328], stage0_57[329], stage0_57[330], stage0_57[331]},
      {stage0_58[270]},
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage1_61[6],stage1_60[50],stage1_59[94],stage1_58[136],stage1_57[157]}
   );
   gpc615_5 gpc2200 (
      {stage0_57[332], stage0_57[333], stage0_57[334], stage0_57[335], stage0_57[336]},
      {stage0_58[271]},
      {stage0_59[42], stage0_59[43], stage0_59[44], stage0_59[45], stage0_59[46], stage0_59[47]},
      {stage1_61[7],stage1_60[51],stage1_59[95],stage1_58[137],stage1_57[158]}
   );
   gpc615_5 gpc2201 (
      {stage0_57[337], stage0_57[338], stage0_57[339], stage0_57[340], stage0_57[341]},
      {stage0_58[272]},
      {stage0_59[48], stage0_59[49], stage0_59[50], stage0_59[51], stage0_59[52], stage0_59[53]},
      {stage1_61[8],stage1_60[52],stage1_59[96],stage1_58[138],stage1_57[159]}
   );
   gpc615_5 gpc2202 (
      {stage0_57[342], stage0_57[343], stage0_57[344], stage0_57[345], stage0_57[346]},
      {stage0_58[273]},
      {stage0_59[54], stage0_59[55], stage0_59[56], stage0_59[57], stage0_59[58], stage0_59[59]},
      {stage1_61[9],stage1_60[53],stage1_59[97],stage1_58[139],stage1_57[160]}
   );
   gpc615_5 gpc2203 (
      {stage0_57[347], stage0_57[348], stage0_57[349], stage0_57[350], stage0_57[351]},
      {stage0_58[274]},
      {stage0_59[60], stage0_59[61], stage0_59[62], stage0_59[63], stage0_59[64], stage0_59[65]},
      {stage1_61[10],stage1_60[54],stage1_59[98],stage1_58[140],stage1_57[161]}
   );
   gpc615_5 gpc2204 (
      {stage0_57[352], stage0_57[353], stage0_57[354], stage0_57[355], stage0_57[356]},
      {stage0_58[275]},
      {stage0_59[66], stage0_59[67], stage0_59[68], stage0_59[69], stage0_59[70], stage0_59[71]},
      {stage1_61[11],stage1_60[55],stage1_59[99],stage1_58[141],stage1_57[162]}
   );
   gpc615_5 gpc2205 (
      {stage0_57[357], stage0_57[358], stage0_57[359], stage0_57[360], stage0_57[361]},
      {stage0_58[276]},
      {stage0_59[72], stage0_59[73], stage0_59[74], stage0_59[75], stage0_59[76], stage0_59[77]},
      {stage1_61[12],stage1_60[56],stage1_59[100],stage1_58[142],stage1_57[163]}
   );
   gpc615_5 gpc2206 (
      {stage0_57[362], stage0_57[363], stage0_57[364], stage0_57[365], stage0_57[366]},
      {stage0_58[277]},
      {stage0_59[78], stage0_59[79], stage0_59[80], stage0_59[81], stage0_59[82], stage0_59[83]},
      {stage1_61[13],stage1_60[57],stage1_59[101],stage1_58[143],stage1_57[164]}
   );
   gpc615_5 gpc2207 (
      {stage0_57[367], stage0_57[368], stage0_57[369], stage0_57[370], stage0_57[371]},
      {stage0_58[278]},
      {stage0_59[84], stage0_59[85], stage0_59[86], stage0_59[87], stage0_59[88], stage0_59[89]},
      {stage1_61[14],stage1_60[58],stage1_59[102],stage1_58[144],stage1_57[165]}
   );
   gpc615_5 gpc2208 (
      {stage0_57[372], stage0_57[373], stage0_57[374], stage0_57[375], stage0_57[376]},
      {stage0_58[279]},
      {stage0_59[90], stage0_59[91], stage0_59[92], stage0_59[93], stage0_59[94], stage0_59[95]},
      {stage1_61[15],stage1_60[59],stage1_59[103],stage1_58[145],stage1_57[166]}
   );
   gpc615_5 gpc2209 (
      {stage0_57[377], stage0_57[378], stage0_57[379], stage0_57[380], stage0_57[381]},
      {stage0_58[280]},
      {stage0_59[96], stage0_59[97], stage0_59[98], stage0_59[99], stage0_59[100], stage0_59[101]},
      {stage1_61[16],stage1_60[60],stage1_59[104],stage1_58[146],stage1_57[167]}
   );
   gpc615_5 gpc2210 (
      {stage0_57[382], stage0_57[383], stage0_57[384], stage0_57[385], stage0_57[386]},
      {stage0_58[281]},
      {stage0_59[102], stage0_59[103], stage0_59[104], stage0_59[105], stage0_59[106], stage0_59[107]},
      {stage1_61[17],stage1_60[61],stage1_59[105],stage1_58[147],stage1_57[168]}
   );
   gpc615_5 gpc2211 (
      {stage0_57[387], stage0_57[388], stage0_57[389], stage0_57[390], stage0_57[391]},
      {stage0_58[282]},
      {stage0_59[108], stage0_59[109], stage0_59[110], stage0_59[111], stage0_59[112], stage0_59[113]},
      {stage1_61[18],stage1_60[62],stage1_59[106],stage1_58[148],stage1_57[169]}
   );
   gpc615_5 gpc2212 (
      {stage0_57[392], stage0_57[393], stage0_57[394], stage0_57[395], stage0_57[396]},
      {stage0_58[283]},
      {stage0_59[114], stage0_59[115], stage0_59[116], stage0_59[117], stage0_59[118], stage0_59[119]},
      {stage1_61[19],stage1_60[63],stage1_59[107],stage1_58[149],stage1_57[170]}
   );
   gpc615_5 gpc2213 (
      {stage0_57[397], stage0_57[398], stage0_57[399], stage0_57[400], stage0_57[401]},
      {stage0_58[284]},
      {stage0_59[120], stage0_59[121], stage0_59[122], stage0_59[123], stage0_59[124], stage0_59[125]},
      {stage1_61[20],stage1_60[64],stage1_59[108],stage1_58[150],stage1_57[171]}
   );
   gpc615_5 gpc2214 (
      {stage0_57[402], stage0_57[403], stage0_57[404], stage0_57[405], stage0_57[406]},
      {stage0_58[285]},
      {stage0_59[126], stage0_59[127], stage0_59[128], stage0_59[129], stage0_59[130], stage0_59[131]},
      {stage1_61[21],stage1_60[65],stage1_59[109],stage1_58[151],stage1_57[172]}
   );
   gpc615_5 gpc2215 (
      {stage0_57[407], stage0_57[408], stage0_57[409], stage0_57[410], stage0_57[411]},
      {stage0_58[286]},
      {stage0_59[132], stage0_59[133], stage0_59[134], stage0_59[135], stage0_59[136], stage0_59[137]},
      {stage1_61[22],stage1_60[66],stage1_59[110],stage1_58[152],stage1_57[173]}
   );
   gpc615_5 gpc2216 (
      {stage0_57[412], stage0_57[413], stage0_57[414], stage0_57[415], stage0_57[416]},
      {stage0_58[287]},
      {stage0_59[138], stage0_59[139], stage0_59[140], stage0_59[141], stage0_59[142], stage0_59[143]},
      {stage1_61[23],stage1_60[67],stage1_59[111],stage1_58[153],stage1_57[174]}
   );
   gpc615_5 gpc2217 (
      {stage0_57[417], stage0_57[418], stage0_57[419], stage0_57[420], stage0_57[421]},
      {stage0_58[288]},
      {stage0_59[144], stage0_59[145], stage0_59[146], stage0_59[147], stage0_59[148], stage0_59[149]},
      {stage1_61[24],stage1_60[68],stage1_59[112],stage1_58[154],stage1_57[175]}
   );
   gpc615_5 gpc2218 (
      {stage0_57[422], stage0_57[423], stage0_57[424], stage0_57[425], stage0_57[426]},
      {stage0_58[289]},
      {stage0_59[150], stage0_59[151], stage0_59[152], stage0_59[153], stage0_59[154], stage0_59[155]},
      {stage1_61[25],stage1_60[69],stage1_59[113],stage1_58[155],stage1_57[176]}
   );
   gpc615_5 gpc2219 (
      {stage0_57[427], stage0_57[428], stage0_57[429], stage0_57[430], stage0_57[431]},
      {stage0_58[290]},
      {stage0_59[156], stage0_59[157], stage0_59[158], stage0_59[159], stage0_59[160], stage0_59[161]},
      {stage1_61[26],stage1_60[70],stage1_59[114],stage1_58[156],stage1_57[177]}
   );
   gpc615_5 gpc2220 (
      {stage0_57[432], stage0_57[433], stage0_57[434], stage0_57[435], stage0_57[436]},
      {stage0_58[291]},
      {stage0_59[162], stage0_59[163], stage0_59[164], stage0_59[165], stage0_59[166], stage0_59[167]},
      {stage1_61[27],stage1_60[71],stage1_59[115],stage1_58[157],stage1_57[178]}
   );
   gpc615_5 gpc2221 (
      {stage0_57[437], stage0_57[438], stage0_57[439], stage0_57[440], stage0_57[441]},
      {stage0_58[292]},
      {stage0_59[168], stage0_59[169], stage0_59[170], stage0_59[171], stage0_59[172], stage0_59[173]},
      {stage1_61[28],stage1_60[72],stage1_59[116],stage1_58[158],stage1_57[179]}
   );
   gpc615_5 gpc2222 (
      {stage0_57[442], stage0_57[443], stage0_57[444], stage0_57[445], stage0_57[446]},
      {stage0_58[293]},
      {stage0_59[174], stage0_59[175], stage0_59[176], stage0_59[177], stage0_59[178], stage0_59[179]},
      {stage1_61[29],stage1_60[73],stage1_59[117],stage1_58[159],stage1_57[180]}
   );
   gpc615_5 gpc2223 (
      {stage0_57[447], stage0_57[448], stage0_57[449], stage0_57[450], stage0_57[451]},
      {stage0_58[294]},
      {stage0_59[180], stage0_59[181], stage0_59[182], stage0_59[183], stage0_59[184], stage0_59[185]},
      {stage1_61[30],stage1_60[74],stage1_59[118],stage1_58[160],stage1_57[181]}
   );
   gpc615_5 gpc2224 (
      {stage0_57[452], stage0_57[453], stage0_57[454], stage0_57[455], stage0_57[456]},
      {stage0_58[295]},
      {stage0_59[186], stage0_59[187], stage0_59[188], stage0_59[189], stage0_59[190], stage0_59[191]},
      {stage1_61[31],stage1_60[75],stage1_59[119],stage1_58[161],stage1_57[182]}
   );
   gpc615_5 gpc2225 (
      {stage0_57[457], stage0_57[458], stage0_57[459], stage0_57[460], stage0_57[461]},
      {stage0_58[296]},
      {stage0_59[192], stage0_59[193], stage0_59[194], stage0_59[195], stage0_59[196], stage0_59[197]},
      {stage1_61[32],stage1_60[76],stage1_59[120],stage1_58[162],stage1_57[183]}
   );
   gpc615_5 gpc2226 (
      {stage0_57[462], stage0_57[463], stage0_57[464], stage0_57[465], stage0_57[466]},
      {stage0_58[297]},
      {stage0_59[198], stage0_59[199], stage0_59[200], stage0_59[201], stage0_59[202], stage0_59[203]},
      {stage1_61[33],stage1_60[77],stage1_59[121],stage1_58[163],stage1_57[184]}
   );
   gpc615_5 gpc2227 (
      {stage0_57[467], stage0_57[468], stage0_57[469], stage0_57[470], stage0_57[471]},
      {stage0_58[298]},
      {stage0_59[204], stage0_59[205], stage0_59[206], stage0_59[207], stage0_59[208], stage0_59[209]},
      {stage1_61[34],stage1_60[78],stage1_59[122],stage1_58[164],stage1_57[185]}
   );
   gpc615_5 gpc2228 (
      {stage0_57[472], stage0_57[473], stage0_57[474], stage0_57[475], stage0_57[476]},
      {stage0_58[299]},
      {stage0_59[210], stage0_59[211], stage0_59[212], stage0_59[213], stage0_59[214], stage0_59[215]},
      {stage1_61[35],stage1_60[79],stage1_59[123],stage1_58[165],stage1_57[186]}
   );
   gpc615_5 gpc2229 (
      {stage0_57[477], stage0_57[478], stage0_57[479], stage0_57[480], stage0_57[481]},
      {stage0_58[300]},
      {stage0_59[216], stage0_59[217], stage0_59[218], stage0_59[219], stage0_59[220], stage0_59[221]},
      {stage1_61[36],stage1_60[80],stage1_59[124],stage1_58[166],stage1_57[187]}
   );
   gpc615_5 gpc2230 (
      {stage0_57[482], stage0_57[483], stage0_57[484], stage0_57[485], 1'b0},
      {stage0_58[301]},
      {stage0_59[222], stage0_59[223], stage0_59[224], stage0_59[225], stage0_59[226], stage0_59[227]},
      {stage1_61[37],stage1_60[81],stage1_59[125],stage1_58[167],stage1_57[188]}
   );
   gpc7_3 gpc2231 (
      {stage0_58[302], stage0_58[303], stage0_58[304], stage0_58[305], stage0_58[306], stage0_58[307], stage0_58[308]},
      {stage1_60[82],stage1_59[126],stage1_58[168]}
   );
   gpc7_3 gpc2232 (
      {stage0_58[309], stage0_58[310], stage0_58[311], stage0_58[312], stage0_58[313], stage0_58[314], stage0_58[315]},
      {stage1_60[83],stage1_59[127],stage1_58[169]}
   );
   gpc7_3 gpc2233 (
      {stage0_58[316], stage0_58[317], stage0_58[318], stage0_58[319], stage0_58[320], stage0_58[321], stage0_58[322]},
      {stage1_60[84],stage1_59[128],stage1_58[170]}
   );
   gpc7_3 gpc2234 (
      {stage0_58[323], stage0_58[324], stage0_58[325], stage0_58[326], stage0_58[327], stage0_58[328], stage0_58[329]},
      {stage1_60[85],stage1_59[129],stage1_58[171]}
   );
   gpc7_3 gpc2235 (
      {stage0_58[330], stage0_58[331], stage0_58[332], stage0_58[333], stage0_58[334], stage0_58[335], stage0_58[336]},
      {stage1_60[86],stage1_59[130],stage1_58[172]}
   );
   gpc7_3 gpc2236 (
      {stage0_58[337], stage0_58[338], stage0_58[339], stage0_58[340], stage0_58[341], stage0_58[342], stage0_58[343]},
      {stage1_60[87],stage1_59[131],stage1_58[173]}
   );
   gpc606_5 gpc2237 (
      {stage0_58[344], stage0_58[345], stage0_58[346], stage0_58[347], stage0_58[348], stage0_58[349]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[38],stage1_60[88],stage1_59[132],stage1_58[174]}
   );
   gpc606_5 gpc2238 (
      {stage0_58[350], stage0_58[351], stage0_58[352], stage0_58[353], stage0_58[354], stage0_58[355]},
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage1_62[1],stage1_61[39],stage1_60[89],stage1_59[133],stage1_58[175]}
   );
   gpc606_5 gpc2239 (
      {stage0_58[356], stage0_58[357], stage0_58[358], stage0_58[359], stage0_58[360], stage0_58[361]},
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage1_62[2],stage1_61[40],stage1_60[90],stage1_59[134],stage1_58[176]}
   );
   gpc606_5 gpc2240 (
      {stage0_58[362], stage0_58[363], stage0_58[364], stage0_58[365], stage0_58[366], stage0_58[367]},
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage1_62[3],stage1_61[41],stage1_60[91],stage1_59[135],stage1_58[177]}
   );
   gpc606_5 gpc2241 (
      {stage0_58[368], stage0_58[369], stage0_58[370], stage0_58[371], stage0_58[372], stage0_58[373]},
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage1_62[4],stage1_61[42],stage1_60[92],stage1_59[136],stage1_58[178]}
   );
   gpc606_5 gpc2242 (
      {stage0_58[374], stage0_58[375], stage0_58[376], stage0_58[377], stage0_58[378], stage0_58[379]},
      {stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33], stage0_60[34], stage0_60[35]},
      {stage1_62[5],stage1_61[43],stage1_60[93],stage1_59[137],stage1_58[179]}
   );
   gpc606_5 gpc2243 (
      {stage0_58[380], stage0_58[381], stage0_58[382], stage0_58[383], stage0_58[384], stage0_58[385]},
      {stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41]},
      {stage1_62[6],stage1_61[44],stage1_60[94],stage1_59[138],stage1_58[180]}
   );
   gpc606_5 gpc2244 (
      {stage0_58[386], stage0_58[387], stage0_58[388], stage0_58[389], stage0_58[390], stage0_58[391]},
      {stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47]},
      {stage1_62[7],stage1_61[45],stage1_60[95],stage1_59[139],stage1_58[181]}
   );
   gpc606_5 gpc2245 (
      {stage0_58[392], stage0_58[393], stage0_58[394], stage0_58[395], stage0_58[396], stage0_58[397]},
      {stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53]},
      {stage1_62[8],stage1_61[46],stage1_60[96],stage1_59[140],stage1_58[182]}
   );
   gpc606_5 gpc2246 (
      {stage0_58[398], stage0_58[399], stage0_58[400], stage0_58[401], stage0_58[402], stage0_58[403]},
      {stage0_60[54], stage0_60[55], stage0_60[56], stage0_60[57], stage0_60[58], stage0_60[59]},
      {stage1_62[9],stage1_61[47],stage1_60[97],stage1_59[141],stage1_58[183]}
   );
   gpc606_5 gpc2247 (
      {stage0_58[404], stage0_58[405], stage0_58[406], stage0_58[407], stage0_58[408], stage0_58[409]},
      {stage0_60[60], stage0_60[61], stage0_60[62], stage0_60[63], stage0_60[64], stage0_60[65]},
      {stage1_62[10],stage1_61[48],stage1_60[98],stage1_59[142],stage1_58[184]}
   );
   gpc606_5 gpc2248 (
      {stage0_58[410], stage0_58[411], stage0_58[412], stage0_58[413], stage0_58[414], stage0_58[415]},
      {stage0_60[66], stage0_60[67], stage0_60[68], stage0_60[69], stage0_60[70], stage0_60[71]},
      {stage1_62[11],stage1_61[49],stage1_60[99],stage1_59[143],stage1_58[185]}
   );
   gpc606_5 gpc2249 (
      {stage0_58[416], stage0_58[417], stage0_58[418], stage0_58[419], stage0_58[420], stage0_58[421]},
      {stage0_60[72], stage0_60[73], stage0_60[74], stage0_60[75], stage0_60[76], stage0_60[77]},
      {stage1_62[12],stage1_61[50],stage1_60[100],stage1_59[144],stage1_58[186]}
   );
   gpc606_5 gpc2250 (
      {stage0_58[422], stage0_58[423], stage0_58[424], stage0_58[425], stage0_58[426], stage0_58[427]},
      {stage0_60[78], stage0_60[79], stage0_60[80], stage0_60[81], stage0_60[82], stage0_60[83]},
      {stage1_62[13],stage1_61[51],stage1_60[101],stage1_59[145],stage1_58[187]}
   );
   gpc606_5 gpc2251 (
      {stage0_58[428], stage0_58[429], stage0_58[430], stage0_58[431], stage0_58[432], stage0_58[433]},
      {stage0_60[84], stage0_60[85], stage0_60[86], stage0_60[87], stage0_60[88], stage0_60[89]},
      {stage1_62[14],stage1_61[52],stage1_60[102],stage1_59[146],stage1_58[188]}
   );
   gpc606_5 gpc2252 (
      {stage0_58[434], stage0_58[435], stage0_58[436], stage0_58[437], stage0_58[438], stage0_58[439]},
      {stage0_60[90], stage0_60[91], stage0_60[92], stage0_60[93], stage0_60[94], stage0_60[95]},
      {stage1_62[15],stage1_61[53],stage1_60[103],stage1_59[147],stage1_58[189]}
   );
   gpc615_5 gpc2253 (
      {stage0_58[440], stage0_58[441], stage0_58[442], stage0_58[443], stage0_58[444]},
      {stage0_59[228]},
      {stage0_60[96], stage0_60[97], stage0_60[98], stage0_60[99], stage0_60[100], stage0_60[101]},
      {stage1_62[16],stage1_61[54],stage1_60[104],stage1_59[148],stage1_58[190]}
   );
   gpc615_5 gpc2254 (
      {stage0_58[445], stage0_58[446], stage0_58[447], stage0_58[448], stage0_58[449]},
      {stage0_59[229]},
      {stage0_60[102], stage0_60[103], stage0_60[104], stage0_60[105], stage0_60[106], stage0_60[107]},
      {stage1_62[17],stage1_61[55],stage1_60[105],stage1_59[149],stage1_58[191]}
   );
   gpc615_5 gpc2255 (
      {stage0_58[450], stage0_58[451], stage0_58[452], stage0_58[453], stage0_58[454]},
      {stage0_59[230]},
      {stage0_60[108], stage0_60[109], stage0_60[110], stage0_60[111], stage0_60[112], stage0_60[113]},
      {stage1_62[18],stage1_61[56],stage1_60[106],stage1_59[150],stage1_58[192]}
   );
   gpc615_5 gpc2256 (
      {stage0_58[455], stage0_58[456], stage0_58[457], stage0_58[458], stage0_58[459]},
      {stage0_59[231]},
      {stage0_60[114], stage0_60[115], stage0_60[116], stage0_60[117], stage0_60[118], stage0_60[119]},
      {stage1_62[19],stage1_61[57],stage1_60[107],stage1_59[151],stage1_58[193]}
   );
   gpc117_4 gpc2257 (
      {stage0_59[232], stage0_59[233], stage0_59[234], stage0_59[235], stage0_59[236], stage0_59[237], stage0_59[238]},
      {stage0_60[120]},
      {stage0_61[0]},
      {stage1_62[20],stage1_61[58],stage1_60[108],stage1_59[152]}
   );
   gpc117_4 gpc2258 (
      {stage0_59[239], stage0_59[240], stage0_59[241], stage0_59[242], stage0_59[243], stage0_59[244], stage0_59[245]},
      {stage0_60[121]},
      {stage0_61[1]},
      {stage1_62[21],stage1_61[59],stage1_60[109],stage1_59[153]}
   );
   gpc117_4 gpc2259 (
      {stage0_59[246], stage0_59[247], stage0_59[248], stage0_59[249], stage0_59[250], stage0_59[251], stage0_59[252]},
      {stage0_60[122]},
      {stage0_61[2]},
      {stage1_62[22],stage1_61[60],stage1_60[110],stage1_59[154]}
   );
   gpc117_4 gpc2260 (
      {stage0_59[253], stage0_59[254], stage0_59[255], stage0_59[256], stage0_59[257], stage0_59[258], stage0_59[259]},
      {stage0_60[123]},
      {stage0_61[3]},
      {stage1_62[23],stage1_61[61],stage1_60[111],stage1_59[155]}
   );
   gpc117_4 gpc2261 (
      {stage0_59[260], stage0_59[261], stage0_59[262], stage0_59[263], stage0_59[264], stage0_59[265], stage0_59[266]},
      {stage0_60[124]},
      {stage0_61[4]},
      {stage1_62[24],stage1_61[62],stage1_60[112],stage1_59[156]}
   );
   gpc117_4 gpc2262 (
      {stage0_59[267], stage0_59[268], stage0_59[269], stage0_59[270], stage0_59[271], stage0_59[272], stage0_59[273]},
      {stage0_60[125]},
      {stage0_61[5]},
      {stage1_62[25],stage1_61[63],stage1_60[113],stage1_59[157]}
   );
   gpc117_4 gpc2263 (
      {stage0_59[274], stage0_59[275], stage0_59[276], stage0_59[277], stage0_59[278], stage0_59[279], stage0_59[280]},
      {stage0_60[126]},
      {stage0_61[6]},
      {stage1_62[26],stage1_61[64],stage1_60[114],stage1_59[158]}
   );
   gpc117_4 gpc2264 (
      {stage0_59[281], stage0_59[282], stage0_59[283], stage0_59[284], stage0_59[285], stage0_59[286], stage0_59[287]},
      {stage0_60[127]},
      {stage0_61[7]},
      {stage1_62[27],stage1_61[65],stage1_60[115],stage1_59[159]}
   );
   gpc117_4 gpc2265 (
      {stage0_59[288], stage0_59[289], stage0_59[290], stage0_59[291], stage0_59[292], stage0_59[293], stage0_59[294]},
      {stage0_60[128]},
      {stage0_61[8]},
      {stage1_62[28],stage1_61[66],stage1_60[116],stage1_59[160]}
   );
   gpc117_4 gpc2266 (
      {stage0_59[295], stage0_59[296], stage0_59[297], stage0_59[298], stage0_59[299], stage0_59[300], stage0_59[301]},
      {stage0_60[129]},
      {stage0_61[9]},
      {stage1_62[29],stage1_61[67],stage1_60[117],stage1_59[161]}
   );
   gpc117_4 gpc2267 (
      {stage0_59[302], stage0_59[303], stage0_59[304], stage0_59[305], stage0_59[306], stage0_59[307], stage0_59[308]},
      {stage0_60[130]},
      {stage0_61[10]},
      {stage1_62[30],stage1_61[68],stage1_60[118],stage1_59[162]}
   );
   gpc117_4 gpc2268 (
      {stage0_59[309], stage0_59[310], stage0_59[311], stage0_59[312], stage0_59[313], stage0_59[314], stage0_59[315]},
      {stage0_60[131]},
      {stage0_61[11]},
      {stage1_62[31],stage1_61[69],stage1_60[119],stage1_59[163]}
   );
   gpc117_4 gpc2269 (
      {stage0_59[316], stage0_59[317], stage0_59[318], stage0_59[319], stage0_59[320], stage0_59[321], stage0_59[322]},
      {stage0_60[132]},
      {stage0_61[12]},
      {stage1_62[32],stage1_61[70],stage1_60[120],stage1_59[164]}
   );
   gpc117_4 gpc2270 (
      {stage0_59[323], stage0_59[324], stage0_59[325], stage0_59[326], stage0_59[327], stage0_59[328], stage0_59[329]},
      {stage0_60[133]},
      {stage0_61[13]},
      {stage1_62[33],stage1_61[71],stage1_60[121],stage1_59[165]}
   );
   gpc117_4 gpc2271 (
      {stage0_59[330], stage0_59[331], stage0_59[332], stage0_59[333], stage0_59[334], stage0_59[335], stage0_59[336]},
      {stage0_60[134]},
      {stage0_61[14]},
      {stage1_62[34],stage1_61[72],stage1_60[122],stage1_59[166]}
   );
   gpc606_5 gpc2272 (
      {stage0_59[337], stage0_59[338], stage0_59[339], stage0_59[340], stage0_59[341], stage0_59[342]},
      {stage0_61[15], stage0_61[16], stage0_61[17], stage0_61[18], stage0_61[19], stage0_61[20]},
      {stage1_63[0],stage1_62[35],stage1_61[73],stage1_60[123],stage1_59[167]}
   );
   gpc606_5 gpc2273 (
      {stage0_59[343], stage0_59[344], stage0_59[345], stage0_59[346], stage0_59[347], stage0_59[348]},
      {stage0_61[21], stage0_61[22], stage0_61[23], stage0_61[24], stage0_61[25], stage0_61[26]},
      {stage1_63[1],stage1_62[36],stage1_61[74],stage1_60[124],stage1_59[168]}
   );
   gpc606_5 gpc2274 (
      {stage0_59[349], stage0_59[350], stage0_59[351], stage0_59[352], stage0_59[353], stage0_59[354]},
      {stage0_61[27], stage0_61[28], stage0_61[29], stage0_61[30], stage0_61[31], stage0_61[32]},
      {stage1_63[2],stage1_62[37],stage1_61[75],stage1_60[125],stage1_59[169]}
   );
   gpc606_5 gpc2275 (
      {stage0_59[355], stage0_59[356], stage0_59[357], stage0_59[358], stage0_59[359], stage0_59[360]},
      {stage0_61[33], stage0_61[34], stage0_61[35], stage0_61[36], stage0_61[37], stage0_61[38]},
      {stage1_63[3],stage1_62[38],stage1_61[76],stage1_60[126],stage1_59[170]}
   );
   gpc606_5 gpc2276 (
      {stage0_59[361], stage0_59[362], stage0_59[363], stage0_59[364], stage0_59[365], stage0_59[366]},
      {stage0_61[39], stage0_61[40], stage0_61[41], stage0_61[42], stage0_61[43], stage0_61[44]},
      {stage1_63[4],stage1_62[39],stage1_61[77],stage1_60[127],stage1_59[171]}
   );
   gpc606_5 gpc2277 (
      {stage0_59[367], stage0_59[368], stage0_59[369], stage0_59[370], stage0_59[371], stage0_59[372]},
      {stage0_61[45], stage0_61[46], stage0_61[47], stage0_61[48], stage0_61[49], stage0_61[50]},
      {stage1_63[5],stage1_62[40],stage1_61[78],stage1_60[128],stage1_59[172]}
   );
   gpc606_5 gpc2278 (
      {stage0_59[373], stage0_59[374], stage0_59[375], stage0_59[376], stage0_59[377], stage0_59[378]},
      {stage0_61[51], stage0_61[52], stage0_61[53], stage0_61[54], stage0_61[55], stage0_61[56]},
      {stage1_63[6],stage1_62[41],stage1_61[79],stage1_60[129],stage1_59[173]}
   );
   gpc606_5 gpc2279 (
      {stage0_59[379], stage0_59[380], stage0_59[381], stage0_59[382], stage0_59[383], stage0_59[384]},
      {stage0_61[57], stage0_61[58], stage0_61[59], stage0_61[60], stage0_61[61], stage0_61[62]},
      {stage1_63[7],stage1_62[42],stage1_61[80],stage1_60[130],stage1_59[174]}
   );
   gpc606_5 gpc2280 (
      {stage0_59[385], stage0_59[386], stage0_59[387], stage0_59[388], stage0_59[389], stage0_59[390]},
      {stage0_61[63], stage0_61[64], stage0_61[65], stage0_61[66], stage0_61[67], stage0_61[68]},
      {stage1_63[8],stage1_62[43],stage1_61[81],stage1_60[131],stage1_59[175]}
   );
   gpc606_5 gpc2281 (
      {stage0_59[391], stage0_59[392], stage0_59[393], stage0_59[394], stage0_59[395], stage0_59[396]},
      {stage0_61[69], stage0_61[70], stage0_61[71], stage0_61[72], stage0_61[73], stage0_61[74]},
      {stage1_63[9],stage1_62[44],stage1_61[82],stage1_60[132],stage1_59[176]}
   );
   gpc606_5 gpc2282 (
      {stage0_59[397], stage0_59[398], stage0_59[399], stage0_59[400], stage0_59[401], stage0_59[402]},
      {stage0_61[75], stage0_61[76], stage0_61[77], stage0_61[78], stage0_61[79], stage0_61[80]},
      {stage1_63[10],stage1_62[45],stage1_61[83],stage1_60[133],stage1_59[177]}
   );
   gpc606_5 gpc2283 (
      {stage0_59[403], stage0_59[404], stage0_59[405], stage0_59[406], stage0_59[407], stage0_59[408]},
      {stage0_61[81], stage0_61[82], stage0_61[83], stage0_61[84], stage0_61[85], stage0_61[86]},
      {stage1_63[11],stage1_62[46],stage1_61[84],stage1_60[134],stage1_59[178]}
   );
   gpc606_5 gpc2284 (
      {stage0_59[409], stage0_59[410], stage0_59[411], stage0_59[412], stage0_59[413], stage0_59[414]},
      {stage0_61[87], stage0_61[88], stage0_61[89], stage0_61[90], stage0_61[91], stage0_61[92]},
      {stage1_63[12],stage1_62[47],stage1_61[85],stage1_60[135],stage1_59[179]}
   );
   gpc606_5 gpc2285 (
      {stage0_59[415], stage0_59[416], stage0_59[417], stage0_59[418], stage0_59[419], stage0_59[420]},
      {stage0_61[93], stage0_61[94], stage0_61[95], stage0_61[96], stage0_61[97], stage0_61[98]},
      {stage1_63[13],stage1_62[48],stage1_61[86],stage1_60[136],stage1_59[180]}
   );
   gpc606_5 gpc2286 (
      {stage0_59[421], stage0_59[422], stage0_59[423], stage0_59[424], stage0_59[425], stage0_59[426]},
      {stage0_61[99], stage0_61[100], stage0_61[101], stage0_61[102], stage0_61[103], stage0_61[104]},
      {stage1_63[14],stage1_62[49],stage1_61[87],stage1_60[137],stage1_59[181]}
   );
   gpc606_5 gpc2287 (
      {stage0_59[427], stage0_59[428], stage0_59[429], stage0_59[430], stage0_59[431], stage0_59[432]},
      {stage0_61[105], stage0_61[106], stage0_61[107], stage0_61[108], stage0_61[109], stage0_61[110]},
      {stage1_63[15],stage1_62[50],stage1_61[88],stage1_60[138],stage1_59[182]}
   );
   gpc606_5 gpc2288 (
      {stage0_59[433], stage0_59[434], stage0_59[435], stage0_59[436], stage0_59[437], stage0_59[438]},
      {stage0_61[111], stage0_61[112], stage0_61[113], stage0_61[114], stage0_61[115], stage0_61[116]},
      {stage1_63[16],stage1_62[51],stage1_61[89],stage1_60[139],stage1_59[183]}
   );
   gpc606_5 gpc2289 (
      {stage0_59[439], stage0_59[440], stage0_59[441], stage0_59[442], stage0_59[443], stage0_59[444]},
      {stage0_61[117], stage0_61[118], stage0_61[119], stage0_61[120], stage0_61[121], stage0_61[122]},
      {stage1_63[17],stage1_62[52],stage1_61[90],stage1_60[140],stage1_59[184]}
   );
   gpc606_5 gpc2290 (
      {stage0_59[445], stage0_59[446], stage0_59[447], stage0_59[448], stage0_59[449], stage0_59[450]},
      {stage0_61[123], stage0_61[124], stage0_61[125], stage0_61[126], stage0_61[127], stage0_61[128]},
      {stage1_63[18],stage1_62[53],stage1_61[91],stage1_60[141],stage1_59[185]}
   );
   gpc606_5 gpc2291 (
      {stage0_59[451], stage0_59[452], stage0_59[453], stage0_59[454], stage0_59[455], stage0_59[456]},
      {stage0_61[129], stage0_61[130], stage0_61[131], stage0_61[132], stage0_61[133], stage0_61[134]},
      {stage1_63[19],stage1_62[54],stage1_61[92],stage1_60[142],stage1_59[186]}
   );
   gpc606_5 gpc2292 (
      {stage0_59[457], stage0_59[458], stage0_59[459], stage0_59[460], stage0_59[461], stage0_59[462]},
      {stage0_61[135], stage0_61[136], stage0_61[137], stage0_61[138], stage0_61[139], stage0_61[140]},
      {stage1_63[20],stage1_62[55],stage1_61[93],stage1_60[143],stage1_59[187]}
   );
   gpc606_5 gpc2293 (
      {stage0_59[463], stage0_59[464], stage0_59[465], stage0_59[466], stage0_59[467], stage0_59[468]},
      {stage0_61[141], stage0_61[142], stage0_61[143], stage0_61[144], stage0_61[145], stage0_61[146]},
      {stage1_63[21],stage1_62[56],stage1_61[94],stage1_60[144],stage1_59[188]}
   );
   gpc606_5 gpc2294 (
      {stage0_60[135], stage0_60[136], stage0_60[137], stage0_60[138], stage0_60[139], stage0_60[140]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[22],stage1_62[57],stage1_61[95],stage1_60[145]}
   );
   gpc615_5 gpc2295 (
      {stage0_60[141], stage0_60[142], stage0_60[143], stage0_60[144], stage0_60[145]},
      {stage0_61[147]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[23],stage1_62[58],stage1_61[96],stage1_60[146]}
   );
   gpc615_5 gpc2296 (
      {stage0_60[146], stage0_60[147], stage0_60[148], stage0_60[149], stage0_60[150]},
      {stage0_61[148]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[24],stage1_62[59],stage1_61[97],stage1_60[147]}
   );
   gpc615_5 gpc2297 (
      {stage0_60[151], stage0_60[152], stage0_60[153], stage0_60[154], stage0_60[155]},
      {stage0_61[149]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[25],stage1_62[60],stage1_61[98],stage1_60[148]}
   );
   gpc615_5 gpc2298 (
      {stage0_60[156], stage0_60[157], stage0_60[158], stage0_60[159], stage0_60[160]},
      {stage0_61[150]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[26],stage1_62[61],stage1_61[99],stage1_60[149]}
   );
   gpc615_5 gpc2299 (
      {stage0_60[161], stage0_60[162], stage0_60[163], stage0_60[164], stage0_60[165]},
      {stage0_61[151]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[27],stage1_62[62],stage1_61[100],stage1_60[150]}
   );
   gpc615_5 gpc2300 (
      {stage0_60[166], stage0_60[167], stage0_60[168], stage0_60[169], stage0_60[170]},
      {stage0_61[152]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[28],stage1_62[63],stage1_61[101],stage1_60[151]}
   );
   gpc615_5 gpc2301 (
      {stage0_60[171], stage0_60[172], stage0_60[173], stage0_60[174], stage0_60[175]},
      {stage0_61[153]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[29],stage1_62[64],stage1_61[102],stage1_60[152]}
   );
   gpc615_5 gpc2302 (
      {stage0_60[176], stage0_60[177], stage0_60[178], stage0_60[179], stage0_60[180]},
      {stage0_61[154]},
      {stage0_62[48], stage0_62[49], stage0_62[50], stage0_62[51], stage0_62[52], stage0_62[53]},
      {stage1_64[8],stage1_63[30],stage1_62[65],stage1_61[103],stage1_60[153]}
   );
   gpc615_5 gpc2303 (
      {stage0_60[181], stage0_60[182], stage0_60[183], stage0_60[184], stage0_60[185]},
      {stage0_61[155]},
      {stage0_62[54], stage0_62[55], stage0_62[56], stage0_62[57], stage0_62[58], stage0_62[59]},
      {stage1_64[9],stage1_63[31],stage1_62[66],stage1_61[104],stage1_60[154]}
   );
   gpc615_5 gpc2304 (
      {stage0_60[186], stage0_60[187], stage0_60[188], stage0_60[189], stage0_60[190]},
      {stage0_61[156]},
      {stage0_62[60], stage0_62[61], stage0_62[62], stage0_62[63], stage0_62[64], stage0_62[65]},
      {stage1_64[10],stage1_63[32],stage1_62[67],stage1_61[105],stage1_60[155]}
   );
   gpc615_5 gpc2305 (
      {stage0_60[191], stage0_60[192], stage0_60[193], stage0_60[194], stage0_60[195]},
      {stage0_61[157]},
      {stage0_62[66], stage0_62[67], stage0_62[68], stage0_62[69], stage0_62[70], stage0_62[71]},
      {stage1_64[11],stage1_63[33],stage1_62[68],stage1_61[106],stage1_60[156]}
   );
   gpc615_5 gpc2306 (
      {stage0_60[196], stage0_60[197], stage0_60[198], stage0_60[199], stage0_60[200]},
      {stage0_61[158]},
      {stage0_62[72], stage0_62[73], stage0_62[74], stage0_62[75], stage0_62[76], stage0_62[77]},
      {stage1_64[12],stage1_63[34],stage1_62[69],stage1_61[107],stage1_60[157]}
   );
   gpc615_5 gpc2307 (
      {stage0_60[201], stage0_60[202], stage0_60[203], stage0_60[204], stage0_60[205]},
      {stage0_61[159]},
      {stage0_62[78], stage0_62[79], stage0_62[80], stage0_62[81], stage0_62[82], stage0_62[83]},
      {stage1_64[13],stage1_63[35],stage1_62[70],stage1_61[108],stage1_60[158]}
   );
   gpc615_5 gpc2308 (
      {stage0_60[206], stage0_60[207], stage0_60[208], stage0_60[209], stage0_60[210]},
      {stage0_61[160]},
      {stage0_62[84], stage0_62[85], stage0_62[86], stage0_62[87], stage0_62[88], stage0_62[89]},
      {stage1_64[14],stage1_63[36],stage1_62[71],stage1_61[109],stage1_60[159]}
   );
   gpc615_5 gpc2309 (
      {stage0_60[211], stage0_60[212], stage0_60[213], stage0_60[214], stage0_60[215]},
      {stage0_61[161]},
      {stage0_62[90], stage0_62[91], stage0_62[92], stage0_62[93], stage0_62[94], stage0_62[95]},
      {stage1_64[15],stage1_63[37],stage1_62[72],stage1_61[110],stage1_60[160]}
   );
   gpc615_5 gpc2310 (
      {stage0_60[216], stage0_60[217], stage0_60[218], stage0_60[219], stage0_60[220]},
      {stage0_61[162]},
      {stage0_62[96], stage0_62[97], stage0_62[98], stage0_62[99], stage0_62[100], stage0_62[101]},
      {stage1_64[16],stage1_63[38],stage1_62[73],stage1_61[111],stage1_60[161]}
   );
   gpc615_5 gpc2311 (
      {stage0_60[221], stage0_60[222], stage0_60[223], stage0_60[224], stage0_60[225]},
      {stage0_61[163]},
      {stage0_62[102], stage0_62[103], stage0_62[104], stage0_62[105], stage0_62[106], stage0_62[107]},
      {stage1_64[17],stage1_63[39],stage1_62[74],stage1_61[112],stage1_60[162]}
   );
   gpc615_5 gpc2312 (
      {stage0_60[226], stage0_60[227], stage0_60[228], stage0_60[229], stage0_60[230]},
      {stage0_61[164]},
      {stage0_62[108], stage0_62[109], stage0_62[110], stage0_62[111], stage0_62[112], stage0_62[113]},
      {stage1_64[18],stage1_63[40],stage1_62[75],stage1_61[113],stage1_60[163]}
   );
   gpc615_5 gpc2313 (
      {stage0_60[231], stage0_60[232], stage0_60[233], stage0_60[234], stage0_60[235]},
      {stage0_61[165]},
      {stage0_62[114], stage0_62[115], stage0_62[116], stage0_62[117], stage0_62[118], stage0_62[119]},
      {stage1_64[19],stage1_63[41],stage1_62[76],stage1_61[114],stage1_60[164]}
   );
   gpc615_5 gpc2314 (
      {stage0_60[236], stage0_60[237], stage0_60[238], stage0_60[239], stage0_60[240]},
      {stage0_61[166]},
      {stage0_62[120], stage0_62[121], stage0_62[122], stage0_62[123], stage0_62[124], stage0_62[125]},
      {stage1_64[20],stage1_63[42],stage1_62[77],stage1_61[115],stage1_60[165]}
   );
   gpc615_5 gpc2315 (
      {stage0_60[241], stage0_60[242], stage0_60[243], stage0_60[244], stage0_60[245]},
      {stage0_61[167]},
      {stage0_62[126], stage0_62[127], stage0_62[128], stage0_62[129], stage0_62[130], stage0_62[131]},
      {stage1_64[21],stage1_63[43],stage1_62[78],stage1_61[116],stage1_60[166]}
   );
   gpc615_5 gpc2316 (
      {stage0_60[246], stage0_60[247], stage0_60[248], stage0_60[249], stage0_60[250]},
      {stage0_61[168]},
      {stage0_62[132], stage0_62[133], stage0_62[134], stage0_62[135], stage0_62[136], stage0_62[137]},
      {stage1_64[22],stage1_63[44],stage1_62[79],stage1_61[117],stage1_60[167]}
   );
   gpc615_5 gpc2317 (
      {stage0_60[251], stage0_60[252], stage0_60[253], stage0_60[254], stage0_60[255]},
      {stage0_61[169]},
      {stage0_62[138], stage0_62[139], stage0_62[140], stage0_62[141], stage0_62[142], stage0_62[143]},
      {stage1_64[23],stage1_63[45],stage1_62[80],stage1_61[118],stage1_60[168]}
   );
   gpc615_5 gpc2318 (
      {stage0_60[256], stage0_60[257], stage0_60[258], stage0_60[259], stage0_60[260]},
      {stage0_61[170]},
      {stage0_62[144], stage0_62[145], stage0_62[146], stage0_62[147], stage0_62[148], stage0_62[149]},
      {stage1_64[24],stage1_63[46],stage1_62[81],stage1_61[119],stage1_60[169]}
   );
   gpc615_5 gpc2319 (
      {stage0_60[261], stage0_60[262], stage0_60[263], stage0_60[264], stage0_60[265]},
      {stage0_61[171]},
      {stage0_62[150], stage0_62[151], stage0_62[152], stage0_62[153], stage0_62[154], stage0_62[155]},
      {stage1_64[25],stage1_63[47],stage1_62[82],stage1_61[120],stage1_60[170]}
   );
   gpc615_5 gpc2320 (
      {stage0_60[266], stage0_60[267], stage0_60[268], stage0_60[269], stage0_60[270]},
      {stage0_61[172]},
      {stage0_62[156], stage0_62[157], stage0_62[158], stage0_62[159], stage0_62[160], stage0_62[161]},
      {stage1_64[26],stage1_63[48],stage1_62[83],stage1_61[121],stage1_60[171]}
   );
   gpc615_5 gpc2321 (
      {stage0_60[271], stage0_60[272], stage0_60[273], stage0_60[274], stage0_60[275]},
      {stage0_61[173]},
      {stage0_62[162], stage0_62[163], stage0_62[164], stage0_62[165], stage0_62[166], stage0_62[167]},
      {stage1_64[27],stage1_63[49],stage1_62[84],stage1_61[122],stage1_60[172]}
   );
   gpc615_5 gpc2322 (
      {stage0_60[276], stage0_60[277], stage0_60[278], stage0_60[279], stage0_60[280]},
      {stage0_61[174]},
      {stage0_62[168], stage0_62[169], stage0_62[170], stage0_62[171], stage0_62[172], stage0_62[173]},
      {stage1_64[28],stage1_63[50],stage1_62[85],stage1_61[123],stage1_60[173]}
   );
   gpc615_5 gpc2323 (
      {stage0_60[281], stage0_60[282], stage0_60[283], stage0_60[284], stage0_60[285]},
      {stage0_61[175]},
      {stage0_62[174], stage0_62[175], stage0_62[176], stage0_62[177], stage0_62[178], stage0_62[179]},
      {stage1_64[29],stage1_63[51],stage1_62[86],stage1_61[124],stage1_60[174]}
   );
   gpc615_5 gpc2324 (
      {stage0_60[286], stage0_60[287], stage0_60[288], stage0_60[289], stage0_60[290]},
      {stage0_61[176]},
      {stage0_62[180], stage0_62[181], stage0_62[182], stage0_62[183], stage0_62[184], stage0_62[185]},
      {stage1_64[30],stage1_63[52],stage1_62[87],stage1_61[125],stage1_60[175]}
   );
   gpc615_5 gpc2325 (
      {stage0_60[291], stage0_60[292], stage0_60[293], stage0_60[294], stage0_60[295]},
      {stage0_61[177]},
      {stage0_62[186], stage0_62[187], stage0_62[188], stage0_62[189], stage0_62[190], stage0_62[191]},
      {stage1_64[31],stage1_63[53],stage1_62[88],stage1_61[126],stage1_60[176]}
   );
   gpc615_5 gpc2326 (
      {stage0_60[296], stage0_60[297], stage0_60[298], stage0_60[299], stage0_60[300]},
      {stage0_61[178]},
      {stage0_62[192], stage0_62[193], stage0_62[194], stage0_62[195], stage0_62[196], stage0_62[197]},
      {stage1_64[32],stage1_63[54],stage1_62[89],stage1_61[127],stage1_60[177]}
   );
   gpc615_5 gpc2327 (
      {stage0_60[301], stage0_60[302], stage0_60[303], stage0_60[304], stage0_60[305]},
      {stage0_61[179]},
      {stage0_62[198], stage0_62[199], stage0_62[200], stage0_62[201], stage0_62[202], stage0_62[203]},
      {stage1_64[33],stage1_63[55],stage1_62[90],stage1_61[128],stage1_60[178]}
   );
   gpc615_5 gpc2328 (
      {stage0_60[306], stage0_60[307], stage0_60[308], stage0_60[309], stage0_60[310]},
      {stage0_61[180]},
      {stage0_62[204], stage0_62[205], stage0_62[206], stage0_62[207], stage0_62[208], stage0_62[209]},
      {stage1_64[34],stage1_63[56],stage1_62[91],stage1_61[129],stage1_60[179]}
   );
   gpc615_5 gpc2329 (
      {stage0_60[311], stage0_60[312], stage0_60[313], stage0_60[314], stage0_60[315]},
      {stage0_61[181]},
      {stage0_62[210], stage0_62[211], stage0_62[212], stage0_62[213], stage0_62[214], stage0_62[215]},
      {stage1_64[35],stage1_63[57],stage1_62[92],stage1_61[130],stage1_60[180]}
   );
   gpc615_5 gpc2330 (
      {stage0_60[316], stage0_60[317], stage0_60[318], stage0_60[319], stage0_60[320]},
      {stage0_61[182]},
      {stage0_62[216], stage0_62[217], stage0_62[218], stage0_62[219], stage0_62[220], stage0_62[221]},
      {stage1_64[36],stage1_63[58],stage1_62[93],stage1_61[131],stage1_60[181]}
   );
   gpc615_5 gpc2331 (
      {stage0_60[321], stage0_60[322], stage0_60[323], stage0_60[324], stage0_60[325]},
      {stage0_61[183]},
      {stage0_62[222], stage0_62[223], stage0_62[224], stage0_62[225], stage0_62[226], stage0_62[227]},
      {stage1_64[37],stage1_63[59],stage1_62[94],stage1_61[132],stage1_60[182]}
   );
   gpc615_5 gpc2332 (
      {stage0_60[326], stage0_60[327], stage0_60[328], stage0_60[329], stage0_60[330]},
      {stage0_61[184]},
      {stage0_62[228], stage0_62[229], stage0_62[230], stage0_62[231], stage0_62[232], stage0_62[233]},
      {stage1_64[38],stage1_63[60],stage1_62[95],stage1_61[133],stage1_60[183]}
   );
   gpc615_5 gpc2333 (
      {stage0_60[331], stage0_60[332], stage0_60[333], stage0_60[334], stage0_60[335]},
      {stage0_61[185]},
      {stage0_62[234], stage0_62[235], stage0_62[236], stage0_62[237], stage0_62[238], stage0_62[239]},
      {stage1_64[39],stage1_63[61],stage1_62[96],stage1_61[134],stage1_60[184]}
   );
   gpc615_5 gpc2334 (
      {stage0_60[336], stage0_60[337], stage0_60[338], stage0_60[339], stage0_60[340]},
      {stage0_61[186]},
      {stage0_62[240], stage0_62[241], stage0_62[242], stage0_62[243], stage0_62[244], stage0_62[245]},
      {stage1_64[40],stage1_63[62],stage1_62[97],stage1_61[135],stage1_60[185]}
   );
   gpc615_5 gpc2335 (
      {stage0_60[341], stage0_60[342], stage0_60[343], stage0_60[344], stage0_60[345]},
      {stage0_61[187]},
      {stage0_62[246], stage0_62[247], stage0_62[248], stage0_62[249], stage0_62[250], stage0_62[251]},
      {stage1_64[41],stage1_63[63],stage1_62[98],stage1_61[136],stage1_60[186]}
   );
   gpc615_5 gpc2336 (
      {stage0_60[346], stage0_60[347], stage0_60[348], stage0_60[349], stage0_60[350]},
      {stage0_61[188]},
      {stage0_62[252], stage0_62[253], stage0_62[254], stage0_62[255], stage0_62[256], stage0_62[257]},
      {stage1_64[42],stage1_63[64],stage1_62[99],stage1_61[137],stage1_60[187]}
   );
   gpc615_5 gpc2337 (
      {stage0_60[351], stage0_60[352], stage0_60[353], stage0_60[354], stage0_60[355]},
      {stage0_61[189]},
      {stage0_62[258], stage0_62[259], stage0_62[260], stage0_62[261], stage0_62[262], stage0_62[263]},
      {stage1_64[43],stage1_63[65],stage1_62[100],stage1_61[138],stage1_60[188]}
   );
   gpc615_5 gpc2338 (
      {stage0_60[356], stage0_60[357], stage0_60[358], stage0_60[359], stage0_60[360]},
      {stage0_61[190]},
      {stage0_62[264], stage0_62[265], stage0_62[266], stage0_62[267], stage0_62[268], stage0_62[269]},
      {stage1_64[44],stage1_63[66],stage1_62[101],stage1_61[139],stage1_60[189]}
   );
   gpc615_5 gpc2339 (
      {stage0_60[361], stage0_60[362], stage0_60[363], stage0_60[364], stage0_60[365]},
      {stage0_61[191]},
      {stage0_62[270], stage0_62[271], stage0_62[272], stage0_62[273], stage0_62[274], stage0_62[275]},
      {stage1_64[45],stage1_63[67],stage1_62[102],stage1_61[140],stage1_60[190]}
   );
   gpc615_5 gpc2340 (
      {stage0_60[366], stage0_60[367], stage0_60[368], stage0_60[369], stage0_60[370]},
      {stage0_61[192]},
      {stage0_62[276], stage0_62[277], stage0_62[278], stage0_62[279], stage0_62[280], stage0_62[281]},
      {stage1_64[46],stage1_63[68],stage1_62[103],stage1_61[141],stage1_60[191]}
   );
   gpc615_5 gpc2341 (
      {stage0_60[371], stage0_60[372], stage0_60[373], stage0_60[374], stage0_60[375]},
      {stage0_61[193]},
      {stage0_62[282], stage0_62[283], stage0_62[284], stage0_62[285], stage0_62[286], stage0_62[287]},
      {stage1_64[47],stage1_63[69],stage1_62[104],stage1_61[142],stage1_60[192]}
   );
   gpc615_5 gpc2342 (
      {stage0_60[376], stage0_60[377], stage0_60[378], stage0_60[379], stage0_60[380]},
      {stage0_61[194]},
      {stage0_62[288], stage0_62[289], stage0_62[290], stage0_62[291], stage0_62[292], stage0_62[293]},
      {stage1_64[48],stage1_63[70],stage1_62[105],stage1_61[143],stage1_60[193]}
   );
   gpc615_5 gpc2343 (
      {stage0_60[381], stage0_60[382], stage0_60[383], stage0_60[384], stage0_60[385]},
      {stage0_61[195]},
      {stage0_62[294], stage0_62[295], stage0_62[296], stage0_62[297], stage0_62[298], stage0_62[299]},
      {stage1_64[49],stage1_63[71],stage1_62[106],stage1_61[144],stage1_60[194]}
   );
   gpc615_5 gpc2344 (
      {stage0_60[386], stage0_60[387], stage0_60[388], stage0_60[389], stage0_60[390]},
      {stage0_61[196]},
      {stage0_62[300], stage0_62[301], stage0_62[302], stage0_62[303], stage0_62[304], stage0_62[305]},
      {stage1_64[50],stage1_63[72],stage1_62[107],stage1_61[145],stage1_60[195]}
   );
   gpc615_5 gpc2345 (
      {stage0_60[391], stage0_60[392], stage0_60[393], stage0_60[394], stage0_60[395]},
      {stage0_61[197]},
      {stage0_62[306], stage0_62[307], stage0_62[308], stage0_62[309], stage0_62[310], stage0_62[311]},
      {stage1_64[51],stage1_63[73],stage1_62[108],stage1_61[146],stage1_60[196]}
   );
   gpc615_5 gpc2346 (
      {stage0_60[396], stage0_60[397], stage0_60[398], stage0_60[399], stage0_60[400]},
      {stage0_61[198]},
      {stage0_62[312], stage0_62[313], stage0_62[314], stage0_62[315], stage0_62[316], stage0_62[317]},
      {stage1_64[52],stage1_63[74],stage1_62[109],stage1_61[147],stage1_60[197]}
   );
   gpc615_5 gpc2347 (
      {stage0_60[401], stage0_60[402], stage0_60[403], stage0_60[404], stage0_60[405]},
      {stage0_61[199]},
      {stage0_62[318], stage0_62[319], stage0_62[320], stage0_62[321], stage0_62[322], stage0_62[323]},
      {stage1_64[53],stage1_63[75],stage1_62[110],stage1_61[148],stage1_60[198]}
   );
   gpc615_5 gpc2348 (
      {stage0_60[406], stage0_60[407], stage0_60[408], stage0_60[409], stage0_60[410]},
      {stage0_61[200]},
      {stage0_62[324], stage0_62[325], stage0_62[326], stage0_62[327], stage0_62[328], stage0_62[329]},
      {stage1_64[54],stage1_63[76],stage1_62[111],stage1_61[149],stage1_60[199]}
   );
   gpc615_5 gpc2349 (
      {stage0_60[411], stage0_60[412], stage0_60[413], stage0_60[414], stage0_60[415]},
      {stage0_61[201]},
      {stage0_62[330], stage0_62[331], stage0_62[332], stage0_62[333], stage0_62[334], stage0_62[335]},
      {stage1_64[55],stage1_63[77],stage1_62[112],stage1_61[150],stage1_60[200]}
   );
   gpc615_5 gpc2350 (
      {stage0_60[416], stage0_60[417], stage0_60[418], stage0_60[419], stage0_60[420]},
      {stage0_61[202]},
      {stage0_62[336], stage0_62[337], stage0_62[338], stage0_62[339], stage0_62[340], stage0_62[341]},
      {stage1_64[56],stage1_63[78],stage1_62[113],stage1_61[151],stage1_60[201]}
   );
   gpc615_5 gpc2351 (
      {stage0_60[421], stage0_60[422], stage0_60[423], stage0_60[424], stage0_60[425]},
      {stage0_61[203]},
      {stage0_62[342], stage0_62[343], stage0_62[344], stage0_62[345], stage0_62[346], stage0_62[347]},
      {stage1_64[57],stage1_63[79],stage1_62[114],stage1_61[152],stage1_60[202]}
   );
   gpc615_5 gpc2352 (
      {stage0_60[426], stage0_60[427], stage0_60[428], stage0_60[429], stage0_60[430]},
      {stage0_61[204]},
      {stage0_62[348], stage0_62[349], stage0_62[350], stage0_62[351], stage0_62[352], stage0_62[353]},
      {stage1_64[58],stage1_63[80],stage1_62[115],stage1_61[153],stage1_60[203]}
   );
   gpc615_5 gpc2353 (
      {stage0_60[431], stage0_60[432], stage0_60[433], stage0_60[434], stage0_60[435]},
      {stage0_61[205]},
      {stage0_62[354], stage0_62[355], stage0_62[356], stage0_62[357], stage0_62[358], stage0_62[359]},
      {stage1_64[59],stage1_63[81],stage1_62[116],stage1_61[154],stage1_60[204]}
   );
   gpc615_5 gpc2354 (
      {stage0_60[436], stage0_60[437], stage0_60[438], stage0_60[439], stage0_60[440]},
      {stage0_61[206]},
      {stage0_62[360], stage0_62[361], stage0_62[362], stage0_62[363], stage0_62[364], stage0_62[365]},
      {stage1_64[60],stage1_63[82],stage1_62[117],stage1_61[155],stage1_60[205]}
   );
   gpc615_5 gpc2355 (
      {stage0_60[441], stage0_60[442], stage0_60[443], stage0_60[444], stage0_60[445]},
      {stage0_61[207]},
      {stage0_62[366], stage0_62[367], stage0_62[368], stage0_62[369], stage0_62[370], stage0_62[371]},
      {stage1_64[61],stage1_63[83],stage1_62[118],stage1_61[156],stage1_60[206]}
   );
   gpc615_5 gpc2356 (
      {stage0_60[446], stage0_60[447], stage0_60[448], stage0_60[449], stage0_60[450]},
      {stage0_61[208]},
      {stage0_62[372], stage0_62[373], stage0_62[374], stage0_62[375], stage0_62[376], stage0_62[377]},
      {stage1_64[62],stage1_63[84],stage1_62[119],stage1_61[157],stage1_60[207]}
   );
   gpc615_5 gpc2357 (
      {stage0_60[451], stage0_60[452], stage0_60[453], stage0_60[454], stage0_60[455]},
      {stage0_61[209]},
      {stage0_62[378], stage0_62[379], stage0_62[380], stage0_62[381], stage0_62[382], stage0_62[383]},
      {stage1_64[63],stage1_63[85],stage1_62[120],stage1_61[158],stage1_60[208]}
   );
   gpc615_5 gpc2358 (
      {stage0_60[456], stage0_60[457], stage0_60[458], stage0_60[459], stage0_60[460]},
      {stage0_61[210]},
      {stage0_62[384], stage0_62[385], stage0_62[386], stage0_62[387], stage0_62[388], stage0_62[389]},
      {stage1_64[64],stage1_63[86],stage1_62[121],stage1_61[159],stage1_60[209]}
   );
   gpc615_5 gpc2359 (
      {stage0_60[461], stage0_60[462], stage0_60[463], stage0_60[464], stage0_60[465]},
      {stage0_61[211]},
      {stage0_62[390], stage0_62[391], stage0_62[392], stage0_62[393], stage0_62[394], stage0_62[395]},
      {stage1_64[65],stage1_63[87],stage1_62[122],stage1_61[160],stage1_60[210]}
   );
   gpc615_5 gpc2360 (
      {stage0_60[466], stage0_60[467], stage0_60[468], stage0_60[469], stage0_60[470]},
      {stage0_61[212]},
      {stage0_62[396], stage0_62[397], stage0_62[398], stage0_62[399], stage0_62[400], stage0_62[401]},
      {stage1_64[66],stage1_63[88],stage1_62[123],stage1_61[161],stage1_60[211]}
   );
   gpc615_5 gpc2361 (
      {stage0_60[471], stage0_60[472], stage0_60[473], stage0_60[474], stage0_60[475]},
      {stage0_61[213]},
      {stage0_62[402], stage0_62[403], stage0_62[404], stage0_62[405], stage0_62[406], stage0_62[407]},
      {stage1_64[67],stage1_63[89],stage1_62[124],stage1_61[162],stage1_60[212]}
   );
   gpc615_5 gpc2362 (
      {stage0_60[476], stage0_60[477], stage0_60[478], stage0_60[479], stage0_60[480]},
      {stage0_61[214]},
      {stage0_62[408], stage0_62[409], stage0_62[410], stage0_62[411], stage0_62[412], stage0_62[413]},
      {stage1_64[68],stage1_63[90],stage1_62[125],stage1_61[163],stage1_60[213]}
   );
   gpc615_5 gpc2363 (
      {stage0_60[481], stage0_60[482], stage0_60[483], stage0_60[484], stage0_60[485]},
      {stage0_61[215]},
      {stage0_62[414], stage0_62[415], stage0_62[416], stage0_62[417], stage0_62[418], stage0_62[419]},
      {stage1_64[69],stage1_63[91],stage1_62[126],stage1_61[164],stage1_60[214]}
   );
   gpc615_5 gpc2364 (
      {stage0_61[216], stage0_61[217], stage0_61[218], stage0_61[219], stage0_61[220]},
      {stage0_62[420]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[70],stage1_63[92],stage1_62[127],stage1_61[165]}
   );
   gpc615_5 gpc2365 (
      {stage0_61[221], stage0_61[222], stage0_61[223], stage0_61[224], stage0_61[225]},
      {stage0_62[421]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[71],stage1_63[93],stage1_62[128],stage1_61[166]}
   );
   gpc615_5 gpc2366 (
      {stage0_61[226], stage0_61[227], stage0_61[228], stage0_61[229], stage0_61[230]},
      {stage0_62[422]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[72],stage1_63[94],stage1_62[129],stage1_61[167]}
   );
   gpc615_5 gpc2367 (
      {stage0_61[231], stage0_61[232], stage0_61[233], stage0_61[234], stage0_61[235]},
      {stage0_62[423]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[73],stage1_63[95],stage1_62[130],stage1_61[168]}
   );
   gpc615_5 gpc2368 (
      {stage0_61[236], stage0_61[237], stage0_61[238], stage0_61[239], stage0_61[240]},
      {stage0_62[424]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[74],stage1_63[96],stage1_62[131],stage1_61[169]}
   );
   gpc615_5 gpc2369 (
      {stage0_61[241], stage0_61[242], stage0_61[243], stage0_61[244], stage0_61[245]},
      {stage0_62[425]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[75],stage1_63[97],stage1_62[132],stage1_61[170]}
   );
   gpc615_5 gpc2370 (
      {stage0_61[246], stage0_61[247], stage0_61[248], stage0_61[249], stage0_61[250]},
      {stage0_62[426]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[76],stage1_63[98],stage1_62[133],stage1_61[171]}
   );
   gpc615_5 gpc2371 (
      {stage0_61[251], stage0_61[252], stage0_61[253], stage0_61[254], stage0_61[255]},
      {stage0_62[427]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[77],stage1_63[99],stage1_62[134],stage1_61[172]}
   );
   gpc615_5 gpc2372 (
      {stage0_61[256], stage0_61[257], stage0_61[258], stage0_61[259], stage0_61[260]},
      {stage0_62[428]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[78],stage1_63[100],stage1_62[135],stage1_61[173]}
   );
   gpc615_5 gpc2373 (
      {stage0_61[261], stage0_61[262], stage0_61[263], stage0_61[264], stage0_61[265]},
      {stage0_62[429]},
      {stage0_63[54], stage0_63[55], stage0_63[56], stage0_63[57], stage0_63[58], stage0_63[59]},
      {stage1_65[9],stage1_64[79],stage1_63[101],stage1_62[136],stage1_61[174]}
   );
   gpc615_5 gpc2374 (
      {stage0_61[266], stage0_61[267], stage0_61[268], stage0_61[269], stage0_61[270]},
      {stage0_62[430]},
      {stage0_63[60], stage0_63[61], stage0_63[62], stage0_63[63], stage0_63[64], stage0_63[65]},
      {stage1_65[10],stage1_64[80],stage1_63[102],stage1_62[137],stage1_61[175]}
   );
   gpc615_5 gpc2375 (
      {stage0_61[271], stage0_61[272], stage0_61[273], stage0_61[274], stage0_61[275]},
      {stage0_62[431]},
      {stage0_63[66], stage0_63[67], stage0_63[68], stage0_63[69], stage0_63[70], stage0_63[71]},
      {stage1_65[11],stage1_64[81],stage1_63[103],stage1_62[138],stage1_61[176]}
   );
   gpc615_5 gpc2376 (
      {stage0_61[276], stage0_61[277], stage0_61[278], stage0_61[279], stage0_61[280]},
      {stage0_62[432]},
      {stage0_63[72], stage0_63[73], stage0_63[74], stage0_63[75], stage0_63[76], stage0_63[77]},
      {stage1_65[12],stage1_64[82],stage1_63[104],stage1_62[139],stage1_61[177]}
   );
   gpc615_5 gpc2377 (
      {stage0_61[281], stage0_61[282], stage0_61[283], stage0_61[284], stage0_61[285]},
      {stage0_62[433]},
      {stage0_63[78], stage0_63[79], stage0_63[80], stage0_63[81], stage0_63[82], stage0_63[83]},
      {stage1_65[13],stage1_64[83],stage1_63[105],stage1_62[140],stage1_61[178]}
   );
   gpc615_5 gpc2378 (
      {stage0_61[286], stage0_61[287], stage0_61[288], stage0_61[289], stage0_61[290]},
      {stage0_62[434]},
      {stage0_63[84], stage0_63[85], stage0_63[86], stage0_63[87], stage0_63[88], stage0_63[89]},
      {stage1_65[14],stage1_64[84],stage1_63[106],stage1_62[141],stage1_61[179]}
   );
   gpc615_5 gpc2379 (
      {stage0_61[291], stage0_61[292], stage0_61[293], stage0_61[294], stage0_61[295]},
      {stage0_62[435]},
      {stage0_63[90], stage0_63[91], stage0_63[92], stage0_63[93], stage0_63[94], stage0_63[95]},
      {stage1_65[15],stage1_64[85],stage1_63[107],stage1_62[142],stage1_61[180]}
   );
   gpc615_5 gpc2380 (
      {stage0_61[296], stage0_61[297], stage0_61[298], stage0_61[299], stage0_61[300]},
      {stage0_62[436]},
      {stage0_63[96], stage0_63[97], stage0_63[98], stage0_63[99], stage0_63[100], stage0_63[101]},
      {stage1_65[16],stage1_64[86],stage1_63[108],stage1_62[143],stage1_61[181]}
   );
   gpc615_5 gpc2381 (
      {stage0_61[301], stage0_61[302], stage0_61[303], stage0_61[304], stage0_61[305]},
      {stage0_62[437]},
      {stage0_63[102], stage0_63[103], stage0_63[104], stage0_63[105], stage0_63[106], stage0_63[107]},
      {stage1_65[17],stage1_64[87],stage1_63[109],stage1_62[144],stage1_61[182]}
   );
   gpc615_5 gpc2382 (
      {stage0_61[306], stage0_61[307], stage0_61[308], stage0_61[309], stage0_61[310]},
      {stage0_62[438]},
      {stage0_63[108], stage0_63[109], stage0_63[110], stage0_63[111], stage0_63[112], stage0_63[113]},
      {stage1_65[18],stage1_64[88],stage1_63[110],stage1_62[145],stage1_61[183]}
   );
   gpc615_5 gpc2383 (
      {stage0_61[311], stage0_61[312], stage0_61[313], stage0_61[314], stage0_61[315]},
      {stage0_62[439]},
      {stage0_63[114], stage0_63[115], stage0_63[116], stage0_63[117], stage0_63[118], stage0_63[119]},
      {stage1_65[19],stage1_64[89],stage1_63[111],stage1_62[146],stage1_61[184]}
   );
   gpc615_5 gpc2384 (
      {stage0_61[316], stage0_61[317], stage0_61[318], stage0_61[319], stage0_61[320]},
      {stage0_62[440]},
      {stage0_63[120], stage0_63[121], stage0_63[122], stage0_63[123], stage0_63[124], stage0_63[125]},
      {stage1_65[20],stage1_64[90],stage1_63[112],stage1_62[147],stage1_61[185]}
   );
   gpc615_5 gpc2385 (
      {stage0_61[321], stage0_61[322], stage0_61[323], stage0_61[324], stage0_61[325]},
      {stage0_62[441]},
      {stage0_63[126], stage0_63[127], stage0_63[128], stage0_63[129], stage0_63[130], stage0_63[131]},
      {stage1_65[21],stage1_64[91],stage1_63[113],stage1_62[148],stage1_61[186]}
   );
   gpc615_5 gpc2386 (
      {stage0_61[326], stage0_61[327], stage0_61[328], stage0_61[329], stage0_61[330]},
      {stage0_62[442]},
      {stage0_63[132], stage0_63[133], stage0_63[134], stage0_63[135], stage0_63[136], stage0_63[137]},
      {stage1_65[22],stage1_64[92],stage1_63[114],stage1_62[149],stage1_61[187]}
   );
   gpc615_5 gpc2387 (
      {stage0_61[331], stage0_61[332], stage0_61[333], stage0_61[334], stage0_61[335]},
      {stage0_62[443]},
      {stage0_63[138], stage0_63[139], stage0_63[140], stage0_63[141], stage0_63[142], stage0_63[143]},
      {stage1_65[23],stage1_64[93],stage1_63[115],stage1_62[150],stage1_61[188]}
   );
   gpc615_5 gpc2388 (
      {stage0_61[336], stage0_61[337], stage0_61[338], stage0_61[339], stage0_61[340]},
      {stage0_62[444]},
      {stage0_63[144], stage0_63[145], stage0_63[146], stage0_63[147], stage0_63[148], stage0_63[149]},
      {stage1_65[24],stage1_64[94],stage1_63[116],stage1_62[151],stage1_61[189]}
   );
   gpc615_5 gpc2389 (
      {stage0_61[341], stage0_61[342], stage0_61[343], stage0_61[344], stage0_61[345]},
      {stage0_62[445]},
      {stage0_63[150], stage0_63[151], stage0_63[152], stage0_63[153], stage0_63[154], stage0_63[155]},
      {stage1_65[25],stage1_64[95],stage1_63[117],stage1_62[152],stage1_61[190]}
   );
   gpc615_5 gpc2390 (
      {stage0_61[346], stage0_61[347], stage0_61[348], stage0_61[349], stage0_61[350]},
      {stage0_62[446]},
      {stage0_63[156], stage0_63[157], stage0_63[158], stage0_63[159], stage0_63[160], stage0_63[161]},
      {stage1_65[26],stage1_64[96],stage1_63[118],stage1_62[153],stage1_61[191]}
   );
   gpc615_5 gpc2391 (
      {stage0_61[351], stage0_61[352], stage0_61[353], stage0_61[354], stage0_61[355]},
      {stage0_62[447]},
      {stage0_63[162], stage0_63[163], stage0_63[164], stage0_63[165], stage0_63[166], stage0_63[167]},
      {stage1_65[27],stage1_64[97],stage1_63[119],stage1_62[154],stage1_61[192]}
   );
   gpc615_5 gpc2392 (
      {stage0_61[356], stage0_61[357], stage0_61[358], stage0_61[359], stage0_61[360]},
      {stage0_62[448]},
      {stage0_63[168], stage0_63[169], stage0_63[170], stage0_63[171], stage0_63[172], stage0_63[173]},
      {stage1_65[28],stage1_64[98],stage1_63[120],stage1_62[155],stage1_61[193]}
   );
   gpc615_5 gpc2393 (
      {stage0_61[361], stage0_61[362], stage0_61[363], stage0_61[364], stage0_61[365]},
      {stage0_62[449]},
      {stage0_63[174], stage0_63[175], stage0_63[176], stage0_63[177], stage0_63[178], stage0_63[179]},
      {stage1_65[29],stage1_64[99],stage1_63[121],stage1_62[156],stage1_61[194]}
   );
   gpc615_5 gpc2394 (
      {stage0_61[366], stage0_61[367], stage0_61[368], stage0_61[369], stage0_61[370]},
      {stage0_62[450]},
      {stage0_63[180], stage0_63[181], stage0_63[182], stage0_63[183], stage0_63[184], stage0_63[185]},
      {stage1_65[30],stage1_64[100],stage1_63[122],stage1_62[157],stage1_61[195]}
   );
   gpc615_5 gpc2395 (
      {stage0_61[371], stage0_61[372], stage0_61[373], stage0_61[374], stage0_61[375]},
      {stage0_62[451]},
      {stage0_63[186], stage0_63[187], stage0_63[188], stage0_63[189], stage0_63[190], stage0_63[191]},
      {stage1_65[31],stage1_64[101],stage1_63[123],stage1_62[158],stage1_61[196]}
   );
   gpc615_5 gpc2396 (
      {stage0_61[376], stage0_61[377], stage0_61[378], stage0_61[379], stage0_61[380]},
      {stage0_62[452]},
      {stage0_63[192], stage0_63[193], stage0_63[194], stage0_63[195], stage0_63[196], stage0_63[197]},
      {stage1_65[32],stage1_64[102],stage1_63[124],stage1_62[159],stage1_61[197]}
   );
   gpc615_5 gpc2397 (
      {stage0_61[381], stage0_61[382], stage0_61[383], stage0_61[384], stage0_61[385]},
      {stage0_62[453]},
      {stage0_63[198], stage0_63[199], stage0_63[200], stage0_63[201], stage0_63[202], stage0_63[203]},
      {stage1_65[33],stage1_64[103],stage1_63[125],stage1_62[160],stage1_61[198]}
   );
   gpc615_5 gpc2398 (
      {stage0_61[386], stage0_61[387], stage0_61[388], stage0_61[389], stage0_61[390]},
      {stage0_62[454]},
      {stage0_63[204], stage0_63[205], stage0_63[206], stage0_63[207], stage0_63[208], stage0_63[209]},
      {stage1_65[34],stage1_64[104],stage1_63[126],stage1_62[161],stage1_61[199]}
   );
   gpc615_5 gpc2399 (
      {stage0_61[391], stage0_61[392], stage0_61[393], stage0_61[394], stage0_61[395]},
      {stage0_62[455]},
      {stage0_63[210], stage0_63[211], stage0_63[212], stage0_63[213], stage0_63[214], stage0_63[215]},
      {stage1_65[35],stage1_64[105],stage1_63[127],stage1_62[162],stage1_61[200]}
   );
   gpc615_5 gpc2400 (
      {stage0_61[396], stage0_61[397], stage0_61[398], stage0_61[399], stage0_61[400]},
      {stage0_62[456]},
      {stage0_63[216], stage0_63[217], stage0_63[218], stage0_63[219], stage0_63[220], stage0_63[221]},
      {stage1_65[36],stage1_64[106],stage1_63[128],stage1_62[163],stage1_61[201]}
   );
   gpc615_5 gpc2401 (
      {stage0_61[401], stage0_61[402], stage0_61[403], stage0_61[404], stage0_61[405]},
      {stage0_62[457]},
      {stage0_63[222], stage0_63[223], stage0_63[224], stage0_63[225], stage0_63[226], stage0_63[227]},
      {stage1_65[37],stage1_64[107],stage1_63[129],stage1_62[164],stage1_61[202]}
   );
   gpc615_5 gpc2402 (
      {stage0_61[406], stage0_61[407], stage0_61[408], stage0_61[409], stage0_61[410]},
      {stage0_62[458]},
      {stage0_63[228], stage0_63[229], stage0_63[230], stage0_63[231], stage0_63[232], stage0_63[233]},
      {stage1_65[38],stage1_64[108],stage1_63[130],stage1_62[165],stage1_61[203]}
   );
   gpc615_5 gpc2403 (
      {stage0_61[411], stage0_61[412], stage0_61[413], stage0_61[414], stage0_61[415]},
      {stage0_62[459]},
      {stage0_63[234], stage0_63[235], stage0_63[236], stage0_63[237], stage0_63[238], stage0_63[239]},
      {stage1_65[39],stage1_64[109],stage1_63[131],stage1_62[166],stage1_61[204]}
   );
   gpc615_5 gpc2404 (
      {stage0_61[416], stage0_61[417], stage0_61[418], stage0_61[419], stage0_61[420]},
      {stage0_62[460]},
      {stage0_63[240], stage0_63[241], stage0_63[242], stage0_63[243], stage0_63[244], stage0_63[245]},
      {stage1_65[40],stage1_64[110],stage1_63[132],stage1_62[167],stage1_61[205]}
   );
   gpc615_5 gpc2405 (
      {stage0_61[421], stage0_61[422], stage0_61[423], stage0_61[424], stage0_61[425]},
      {stage0_62[461]},
      {stage0_63[246], stage0_63[247], stage0_63[248], stage0_63[249], stage0_63[250], stage0_63[251]},
      {stage1_65[41],stage1_64[111],stage1_63[133],stage1_62[168],stage1_61[206]}
   );
   gpc615_5 gpc2406 (
      {stage0_61[426], stage0_61[427], stage0_61[428], stage0_61[429], stage0_61[430]},
      {stage0_62[462]},
      {stage0_63[252], stage0_63[253], stage0_63[254], stage0_63[255], stage0_63[256], stage0_63[257]},
      {stage1_65[42],stage1_64[112],stage1_63[134],stage1_62[169],stage1_61[207]}
   );
   gpc615_5 gpc2407 (
      {stage0_61[431], stage0_61[432], stage0_61[433], stage0_61[434], stage0_61[435]},
      {stage0_62[463]},
      {stage0_63[258], stage0_63[259], stage0_63[260], stage0_63[261], stage0_63[262], stage0_63[263]},
      {stage1_65[43],stage1_64[113],stage1_63[135],stage1_62[170],stage1_61[208]}
   );
   gpc615_5 gpc2408 (
      {stage0_61[436], stage0_61[437], stage0_61[438], stage0_61[439], stage0_61[440]},
      {stage0_62[464]},
      {stage0_63[264], stage0_63[265], stage0_63[266], stage0_63[267], stage0_63[268], stage0_63[269]},
      {stage1_65[44],stage1_64[114],stage1_63[136],stage1_62[171],stage1_61[209]}
   );
   gpc615_5 gpc2409 (
      {stage0_61[441], stage0_61[442], stage0_61[443], stage0_61[444], stage0_61[445]},
      {stage0_62[465]},
      {stage0_63[270], stage0_63[271], stage0_63[272], stage0_63[273], stage0_63[274], stage0_63[275]},
      {stage1_65[45],stage1_64[115],stage1_63[137],stage1_62[172],stage1_61[210]}
   );
   gpc615_5 gpc2410 (
      {stage0_61[446], stage0_61[447], stage0_61[448], stage0_61[449], stage0_61[450]},
      {stage0_62[466]},
      {stage0_63[276], stage0_63[277], stage0_63[278], stage0_63[279], stage0_63[280], stage0_63[281]},
      {stage1_65[46],stage1_64[116],stage1_63[138],stage1_62[173],stage1_61[211]}
   );
   gpc615_5 gpc2411 (
      {stage0_61[451], stage0_61[452], stage0_61[453], stage0_61[454], stage0_61[455]},
      {stage0_62[467]},
      {stage0_63[282], stage0_63[283], stage0_63[284], stage0_63[285], stage0_63[286], stage0_63[287]},
      {stage1_65[47],stage1_64[117],stage1_63[139],stage1_62[174],stage1_61[212]}
   );
   gpc615_5 gpc2412 (
      {stage0_61[456], stage0_61[457], stage0_61[458], stage0_61[459], stage0_61[460]},
      {stage0_62[468]},
      {stage0_63[288], stage0_63[289], stage0_63[290], stage0_63[291], stage0_63[292], stage0_63[293]},
      {stage1_65[48],stage1_64[118],stage1_63[140],stage1_62[175],stage1_61[213]}
   );
   gpc615_5 gpc2413 (
      {stage0_61[461], stage0_61[462], stage0_61[463], stage0_61[464], stage0_61[465]},
      {stage0_62[469]},
      {stage0_63[294], stage0_63[295], stage0_63[296], stage0_63[297], stage0_63[298], stage0_63[299]},
      {stage1_65[49],stage1_64[119],stage1_63[141],stage1_62[176],stage1_61[214]}
   );
   gpc615_5 gpc2414 (
      {stage0_61[466], stage0_61[467], stage0_61[468], stage0_61[469], stage0_61[470]},
      {stage0_62[470]},
      {stage0_63[300], stage0_63[301], stage0_63[302], stage0_63[303], stage0_63[304], stage0_63[305]},
      {stage1_65[50],stage1_64[120],stage1_63[142],stage1_62[177],stage1_61[215]}
   );
   gpc615_5 gpc2415 (
      {stage0_61[471], stage0_61[472], stage0_61[473], stage0_61[474], stage0_61[475]},
      {stage0_62[471]},
      {stage0_63[306], stage0_63[307], stage0_63[308], stage0_63[309], stage0_63[310], stage0_63[311]},
      {stage1_65[51],stage1_64[121],stage1_63[143],stage1_62[178],stage1_61[216]}
   );
   gpc615_5 gpc2416 (
      {stage0_61[476], stage0_61[477], stage0_61[478], stage0_61[479], stage0_61[480]},
      {stage0_62[472]},
      {stage0_63[312], stage0_63[313], stage0_63[314], stage0_63[315], stage0_63[316], stage0_63[317]},
      {stage1_65[52],stage1_64[122],stage1_63[144],stage1_62[179],stage1_61[217]}
   );
   gpc615_5 gpc2417 (
      {stage0_61[481], stage0_61[482], stage0_61[483], stage0_61[484], stage0_61[485]},
      {stage0_62[473]},
      {stage0_63[318], stage0_63[319], stage0_63[320], stage0_63[321], stage0_63[322], stage0_63[323]},
      {stage1_65[53],stage1_64[123],stage1_63[145],stage1_62[180],stage1_61[218]}
   );
   gpc1_1 gpc2418 (
      {stage0_0[448]},
      {stage1_0[87]}
   );
   gpc1_1 gpc2419 (
      {stage0_0[449]},
      {stage1_0[88]}
   );
   gpc1_1 gpc2420 (
      {stage0_0[450]},
      {stage1_0[89]}
   );
   gpc1_1 gpc2421 (
      {stage0_0[451]},
      {stage1_0[90]}
   );
   gpc1_1 gpc2422 (
      {stage0_0[452]},
      {stage1_0[91]}
   );
   gpc1_1 gpc2423 (
      {stage0_0[453]},
      {stage1_0[92]}
   );
   gpc1_1 gpc2424 (
      {stage0_0[454]},
      {stage1_0[93]}
   );
   gpc1_1 gpc2425 (
      {stage0_0[455]},
      {stage1_0[94]}
   );
   gpc1_1 gpc2426 (
      {stage0_0[456]},
      {stage1_0[95]}
   );
   gpc1_1 gpc2427 (
      {stage0_0[457]},
      {stage1_0[96]}
   );
   gpc1_1 gpc2428 (
      {stage0_0[458]},
      {stage1_0[97]}
   );
   gpc1_1 gpc2429 (
      {stage0_0[459]},
      {stage1_0[98]}
   );
   gpc1_1 gpc2430 (
      {stage0_0[460]},
      {stage1_0[99]}
   );
   gpc1_1 gpc2431 (
      {stage0_0[461]},
      {stage1_0[100]}
   );
   gpc1_1 gpc2432 (
      {stage0_0[462]},
      {stage1_0[101]}
   );
   gpc1_1 gpc2433 (
      {stage0_0[463]},
      {stage1_0[102]}
   );
   gpc1_1 gpc2434 (
      {stage0_0[464]},
      {stage1_0[103]}
   );
   gpc1_1 gpc2435 (
      {stage0_0[465]},
      {stage1_0[104]}
   );
   gpc1_1 gpc2436 (
      {stage0_0[466]},
      {stage1_0[105]}
   );
   gpc1_1 gpc2437 (
      {stage0_0[467]},
      {stage1_0[106]}
   );
   gpc1_1 gpc2438 (
      {stage0_0[468]},
      {stage1_0[107]}
   );
   gpc1_1 gpc2439 (
      {stage0_0[469]},
      {stage1_0[108]}
   );
   gpc1_1 gpc2440 (
      {stage0_0[470]},
      {stage1_0[109]}
   );
   gpc1_1 gpc2441 (
      {stage0_0[471]},
      {stage1_0[110]}
   );
   gpc1_1 gpc2442 (
      {stage0_0[472]},
      {stage1_0[111]}
   );
   gpc1_1 gpc2443 (
      {stage0_0[473]},
      {stage1_0[112]}
   );
   gpc1_1 gpc2444 (
      {stage0_0[474]},
      {stage1_0[113]}
   );
   gpc1_1 gpc2445 (
      {stage0_0[475]},
      {stage1_0[114]}
   );
   gpc1_1 gpc2446 (
      {stage0_0[476]},
      {stage1_0[115]}
   );
   gpc1_1 gpc2447 (
      {stage0_0[477]},
      {stage1_0[116]}
   );
   gpc1_1 gpc2448 (
      {stage0_0[478]},
      {stage1_0[117]}
   );
   gpc1_1 gpc2449 (
      {stage0_0[479]},
      {stage1_0[118]}
   );
   gpc1_1 gpc2450 (
      {stage0_0[480]},
      {stage1_0[119]}
   );
   gpc1_1 gpc2451 (
      {stage0_0[481]},
      {stage1_0[120]}
   );
   gpc1_1 gpc2452 (
      {stage0_0[482]},
      {stage1_0[121]}
   );
   gpc1_1 gpc2453 (
      {stage0_0[483]},
      {stage1_0[122]}
   );
   gpc1_1 gpc2454 (
      {stage0_0[484]},
      {stage1_0[123]}
   );
   gpc1_1 gpc2455 (
      {stage0_0[485]},
      {stage1_0[124]}
   );
   gpc1_1 gpc2456 (
      {stage0_1[439]},
      {stage1_1[129]}
   );
   gpc1_1 gpc2457 (
      {stage0_1[440]},
      {stage1_1[130]}
   );
   gpc1_1 gpc2458 (
      {stage0_1[441]},
      {stage1_1[131]}
   );
   gpc1_1 gpc2459 (
      {stage0_1[442]},
      {stage1_1[132]}
   );
   gpc1_1 gpc2460 (
      {stage0_1[443]},
      {stage1_1[133]}
   );
   gpc1_1 gpc2461 (
      {stage0_1[444]},
      {stage1_1[134]}
   );
   gpc1_1 gpc2462 (
      {stage0_1[445]},
      {stage1_1[135]}
   );
   gpc1_1 gpc2463 (
      {stage0_1[446]},
      {stage1_1[136]}
   );
   gpc1_1 gpc2464 (
      {stage0_1[447]},
      {stage1_1[137]}
   );
   gpc1_1 gpc2465 (
      {stage0_1[448]},
      {stage1_1[138]}
   );
   gpc1_1 gpc2466 (
      {stage0_1[449]},
      {stage1_1[139]}
   );
   gpc1_1 gpc2467 (
      {stage0_1[450]},
      {stage1_1[140]}
   );
   gpc1_1 gpc2468 (
      {stage0_1[451]},
      {stage1_1[141]}
   );
   gpc1_1 gpc2469 (
      {stage0_1[452]},
      {stage1_1[142]}
   );
   gpc1_1 gpc2470 (
      {stage0_1[453]},
      {stage1_1[143]}
   );
   gpc1_1 gpc2471 (
      {stage0_1[454]},
      {stage1_1[144]}
   );
   gpc1_1 gpc2472 (
      {stage0_1[455]},
      {stage1_1[145]}
   );
   gpc1_1 gpc2473 (
      {stage0_1[456]},
      {stage1_1[146]}
   );
   gpc1_1 gpc2474 (
      {stage0_1[457]},
      {stage1_1[147]}
   );
   gpc1_1 gpc2475 (
      {stage0_1[458]},
      {stage1_1[148]}
   );
   gpc1_1 gpc2476 (
      {stage0_1[459]},
      {stage1_1[149]}
   );
   gpc1_1 gpc2477 (
      {stage0_1[460]},
      {stage1_1[150]}
   );
   gpc1_1 gpc2478 (
      {stage0_1[461]},
      {stage1_1[151]}
   );
   gpc1_1 gpc2479 (
      {stage0_1[462]},
      {stage1_1[152]}
   );
   gpc1_1 gpc2480 (
      {stage0_1[463]},
      {stage1_1[153]}
   );
   gpc1_1 gpc2481 (
      {stage0_1[464]},
      {stage1_1[154]}
   );
   gpc1_1 gpc2482 (
      {stage0_1[465]},
      {stage1_1[155]}
   );
   gpc1_1 gpc2483 (
      {stage0_1[466]},
      {stage1_1[156]}
   );
   gpc1_1 gpc2484 (
      {stage0_1[467]},
      {stage1_1[157]}
   );
   gpc1_1 gpc2485 (
      {stage0_1[468]},
      {stage1_1[158]}
   );
   gpc1_1 gpc2486 (
      {stage0_1[469]},
      {stage1_1[159]}
   );
   gpc1_1 gpc2487 (
      {stage0_1[470]},
      {stage1_1[160]}
   );
   gpc1_1 gpc2488 (
      {stage0_1[471]},
      {stage1_1[161]}
   );
   gpc1_1 gpc2489 (
      {stage0_1[472]},
      {stage1_1[162]}
   );
   gpc1_1 gpc2490 (
      {stage0_1[473]},
      {stage1_1[163]}
   );
   gpc1_1 gpc2491 (
      {stage0_1[474]},
      {stage1_1[164]}
   );
   gpc1_1 gpc2492 (
      {stage0_1[475]},
      {stage1_1[165]}
   );
   gpc1_1 gpc2493 (
      {stage0_1[476]},
      {stage1_1[166]}
   );
   gpc1_1 gpc2494 (
      {stage0_1[477]},
      {stage1_1[167]}
   );
   gpc1_1 gpc2495 (
      {stage0_1[478]},
      {stage1_1[168]}
   );
   gpc1_1 gpc2496 (
      {stage0_1[479]},
      {stage1_1[169]}
   );
   gpc1_1 gpc2497 (
      {stage0_1[480]},
      {stage1_1[170]}
   );
   gpc1_1 gpc2498 (
      {stage0_1[481]},
      {stage1_1[171]}
   );
   gpc1_1 gpc2499 (
      {stage0_1[482]},
      {stage1_1[172]}
   );
   gpc1_1 gpc2500 (
      {stage0_1[483]},
      {stage1_1[173]}
   );
   gpc1_1 gpc2501 (
      {stage0_1[484]},
      {stage1_1[174]}
   );
   gpc1_1 gpc2502 (
      {stage0_1[485]},
      {stage1_1[175]}
   );
   gpc1_1 gpc2503 (
      {stage0_3[466]},
      {stage1_3[195]}
   );
   gpc1_1 gpc2504 (
      {stage0_3[467]},
      {stage1_3[196]}
   );
   gpc1_1 gpc2505 (
      {stage0_3[468]},
      {stage1_3[197]}
   );
   gpc1_1 gpc2506 (
      {stage0_3[469]},
      {stage1_3[198]}
   );
   gpc1_1 gpc2507 (
      {stage0_3[470]},
      {stage1_3[199]}
   );
   gpc1_1 gpc2508 (
      {stage0_3[471]},
      {stage1_3[200]}
   );
   gpc1_1 gpc2509 (
      {stage0_3[472]},
      {stage1_3[201]}
   );
   gpc1_1 gpc2510 (
      {stage0_3[473]},
      {stage1_3[202]}
   );
   gpc1_1 gpc2511 (
      {stage0_3[474]},
      {stage1_3[203]}
   );
   gpc1_1 gpc2512 (
      {stage0_3[475]},
      {stage1_3[204]}
   );
   gpc1_1 gpc2513 (
      {stage0_3[476]},
      {stage1_3[205]}
   );
   gpc1_1 gpc2514 (
      {stage0_3[477]},
      {stage1_3[206]}
   );
   gpc1_1 gpc2515 (
      {stage0_3[478]},
      {stage1_3[207]}
   );
   gpc1_1 gpc2516 (
      {stage0_3[479]},
      {stage1_3[208]}
   );
   gpc1_1 gpc2517 (
      {stage0_3[480]},
      {stage1_3[209]}
   );
   gpc1_1 gpc2518 (
      {stage0_3[481]},
      {stage1_3[210]}
   );
   gpc1_1 gpc2519 (
      {stage0_3[482]},
      {stage1_3[211]}
   );
   gpc1_1 gpc2520 (
      {stage0_3[483]},
      {stage1_3[212]}
   );
   gpc1_1 gpc2521 (
      {stage0_3[484]},
      {stage1_3[213]}
   );
   gpc1_1 gpc2522 (
      {stage0_3[485]},
      {stage1_3[214]}
   );
   gpc1_1 gpc2523 (
      {stage0_6[466]},
      {stage1_6[194]}
   );
   gpc1_1 gpc2524 (
      {stage0_6[467]},
      {stage1_6[195]}
   );
   gpc1_1 gpc2525 (
      {stage0_6[468]},
      {stage1_6[196]}
   );
   gpc1_1 gpc2526 (
      {stage0_6[469]},
      {stage1_6[197]}
   );
   gpc1_1 gpc2527 (
      {stage0_6[470]},
      {stage1_6[198]}
   );
   gpc1_1 gpc2528 (
      {stage0_6[471]},
      {stage1_6[199]}
   );
   gpc1_1 gpc2529 (
      {stage0_6[472]},
      {stage1_6[200]}
   );
   gpc1_1 gpc2530 (
      {stage0_6[473]},
      {stage1_6[201]}
   );
   gpc1_1 gpc2531 (
      {stage0_6[474]},
      {stage1_6[202]}
   );
   gpc1_1 gpc2532 (
      {stage0_6[475]},
      {stage1_6[203]}
   );
   gpc1_1 gpc2533 (
      {stage0_6[476]},
      {stage1_6[204]}
   );
   gpc1_1 gpc2534 (
      {stage0_6[477]},
      {stage1_6[205]}
   );
   gpc1_1 gpc2535 (
      {stage0_6[478]},
      {stage1_6[206]}
   );
   gpc1_1 gpc2536 (
      {stage0_6[479]},
      {stage1_6[207]}
   );
   gpc1_1 gpc2537 (
      {stage0_6[480]},
      {stage1_6[208]}
   );
   gpc1_1 gpc2538 (
      {stage0_6[481]},
      {stage1_6[209]}
   );
   gpc1_1 gpc2539 (
      {stage0_6[482]},
      {stage1_6[210]}
   );
   gpc1_1 gpc2540 (
      {stage0_6[483]},
      {stage1_6[211]}
   );
   gpc1_1 gpc2541 (
      {stage0_6[484]},
      {stage1_6[212]}
   );
   gpc1_1 gpc2542 (
      {stage0_6[485]},
      {stage1_6[213]}
   );
   gpc1_1 gpc2543 (
      {stage0_7[462]},
      {stage1_7[197]}
   );
   gpc1_1 gpc2544 (
      {stage0_7[463]},
      {stage1_7[198]}
   );
   gpc1_1 gpc2545 (
      {stage0_7[464]},
      {stage1_7[199]}
   );
   gpc1_1 gpc2546 (
      {stage0_7[465]},
      {stage1_7[200]}
   );
   gpc1_1 gpc2547 (
      {stage0_7[466]},
      {stage1_7[201]}
   );
   gpc1_1 gpc2548 (
      {stage0_7[467]},
      {stage1_7[202]}
   );
   gpc1_1 gpc2549 (
      {stage0_7[468]},
      {stage1_7[203]}
   );
   gpc1_1 gpc2550 (
      {stage0_7[469]},
      {stage1_7[204]}
   );
   gpc1_1 gpc2551 (
      {stage0_7[470]},
      {stage1_7[205]}
   );
   gpc1_1 gpc2552 (
      {stage0_7[471]},
      {stage1_7[206]}
   );
   gpc1_1 gpc2553 (
      {stage0_7[472]},
      {stage1_7[207]}
   );
   gpc1_1 gpc2554 (
      {stage0_7[473]},
      {stage1_7[208]}
   );
   gpc1_1 gpc2555 (
      {stage0_7[474]},
      {stage1_7[209]}
   );
   gpc1_1 gpc2556 (
      {stage0_7[475]},
      {stage1_7[210]}
   );
   gpc1_1 gpc2557 (
      {stage0_7[476]},
      {stage1_7[211]}
   );
   gpc1_1 gpc2558 (
      {stage0_7[477]},
      {stage1_7[212]}
   );
   gpc1_1 gpc2559 (
      {stage0_7[478]},
      {stage1_7[213]}
   );
   gpc1_1 gpc2560 (
      {stage0_7[479]},
      {stage1_7[214]}
   );
   gpc1_1 gpc2561 (
      {stage0_7[480]},
      {stage1_7[215]}
   );
   gpc1_1 gpc2562 (
      {stage0_7[481]},
      {stage1_7[216]}
   );
   gpc1_1 gpc2563 (
      {stage0_7[482]},
      {stage1_7[217]}
   );
   gpc1_1 gpc2564 (
      {stage0_7[483]},
      {stage1_7[218]}
   );
   gpc1_1 gpc2565 (
      {stage0_7[484]},
      {stage1_7[219]}
   );
   gpc1_1 gpc2566 (
      {stage0_7[485]},
      {stage1_7[220]}
   );
   gpc1_1 gpc2567 (
      {stage0_8[476]},
      {stage1_8[196]}
   );
   gpc1_1 gpc2568 (
      {stage0_8[477]},
      {stage1_8[197]}
   );
   gpc1_1 gpc2569 (
      {stage0_8[478]},
      {stage1_8[198]}
   );
   gpc1_1 gpc2570 (
      {stage0_8[479]},
      {stage1_8[199]}
   );
   gpc1_1 gpc2571 (
      {stage0_8[480]},
      {stage1_8[200]}
   );
   gpc1_1 gpc2572 (
      {stage0_8[481]},
      {stage1_8[201]}
   );
   gpc1_1 gpc2573 (
      {stage0_8[482]},
      {stage1_8[202]}
   );
   gpc1_1 gpc2574 (
      {stage0_8[483]},
      {stage1_8[203]}
   );
   gpc1_1 gpc2575 (
      {stage0_8[484]},
      {stage1_8[204]}
   );
   gpc1_1 gpc2576 (
      {stage0_8[485]},
      {stage1_8[205]}
   );
   gpc1_1 gpc2577 (
      {stage0_9[468]},
      {stage1_9[196]}
   );
   gpc1_1 gpc2578 (
      {stage0_9[469]},
      {stage1_9[197]}
   );
   gpc1_1 gpc2579 (
      {stage0_9[470]},
      {stage1_9[198]}
   );
   gpc1_1 gpc2580 (
      {stage0_9[471]},
      {stage1_9[199]}
   );
   gpc1_1 gpc2581 (
      {stage0_9[472]},
      {stage1_9[200]}
   );
   gpc1_1 gpc2582 (
      {stage0_9[473]},
      {stage1_9[201]}
   );
   gpc1_1 gpc2583 (
      {stage0_9[474]},
      {stage1_9[202]}
   );
   gpc1_1 gpc2584 (
      {stage0_9[475]},
      {stage1_9[203]}
   );
   gpc1_1 gpc2585 (
      {stage0_9[476]},
      {stage1_9[204]}
   );
   gpc1_1 gpc2586 (
      {stage0_9[477]},
      {stage1_9[205]}
   );
   gpc1_1 gpc2587 (
      {stage0_9[478]},
      {stage1_9[206]}
   );
   gpc1_1 gpc2588 (
      {stage0_9[479]},
      {stage1_9[207]}
   );
   gpc1_1 gpc2589 (
      {stage0_9[480]},
      {stage1_9[208]}
   );
   gpc1_1 gpc2590 (
      {stage0_9[481]},
      {stage1_9[209]}
   );
   gpc1_1 gpc2591 (
      {stage0_9[482]},
      {stage1_9[210]}
   );
   gpc1_1 gpc2592 (
      {stage0_9[483]},
      {stage1_9[211]}
   );
   gpc1_1 gpc2593 (
      {stage0_9[484]},
      {stage1_9[212]}
   );
   gpc1_1 gpc2594 (
      {stage0_9[485]},
      {stage1_9[213]}
   );
   gpc1_1 gpc2595 (
      {stage0_10[384]},
      {stage1_10[183]}
   );
   gpc1_1 gpc2596 (
      {stage0_10[385]},
      {stage1_10[184]}
   );
   gpc1_1 gpc2597 (
      {stage0_10[386]},
      {stage1_10[185]}
   );
   gpc1_1 gpc2598 (
      {stage0_10[387]},
      {stage1_10[186]}
   );
   gpc1_1 gpc2599 (
      {stage0_10[388]},
      {stage1_10[187]}
   );
   gpc1_1 gpc2600 (
      {stage0_10[389]},
      {stage1_10[188]}
   );
   gpc1_1 gpc2601 (
      {stage0_10[390]},
      {stage1_10[189]}
   );
   gpc1_1 gpc2602 (
      {stage0_10[391]},
      {stage1_10[190]}
   );
   gpc1_1 gpc2603 (
      {stage0_10[392]},
      {stage1_10[191]}
   );
   gpc1_1 gpc2604 (
      {stage0_10[393]},
      {stage1_10[192]}
   );
   gpc1_1 gpc2605 (
      {stage0_10[394]},
      {stage1_10[193]}
   );
   gpc1_1 gpc2606 (
      {stage0_10[395]},
      {stage1_10[194]}
   );
   gpc1_1 gpc2607 (
      {stage0_10[396]},
      {stage1_10[195]}
   );
   gpc1_1 gpc2608 (
      {stage0_10[397]},
      {stage1_10[196]}
   );
   gpc1_1 gpc2609 (
      {stage0_10[398]},
      {stage1_10[197]}
   );
   gpc1_1 gpc2610 (
      {stage0_10[399]},
      {stage1_10[198]}
   );
   gpc1_1 gpc2611 (
      {stage0_10[400]},
      {stage1_10[199]}
   );
   gpc1_1 gpc2612 (
      {stage0_10[401]},
      {stage1_10[200]}
   );
   gpc1_1 gpc2613 (
      {stage0_10[402]},
      {stage1_10[201]}
   );
   gpc1_1 gpc2614 (
      {stage0_10[403]},
      {stage1_10[202]}
   );
   gpc1_1 gpc2615 (
      {stage0_10[404]},
      {stage1_10[203]}
   );
   gpc1_1 gpc2616 (
      {stage0_10[405]},
      {stage1_10[204]}
   );
   gpc1_1 gpc2617 (
      {stage0_10[406]},
      {stage1_10[205]}
   );
   gpc1_1 gpc2618 (
      {stage0_10[407]},
      {stage1_10[206]}
   );
   gpc1_1 gpc2619 (
      {stage0_10[408]},
      {stage1_10[207]}
   );
   gpc1_1 gpc2620 (
      {stage0_10[409]},
      {stage1_10[208]}
   );
   gpc1_1 gpc2621 (
      {stage0_10[410]},
      {stage1_10[209]}
   );
   gpc1_1 gpc2622 (
      {stage0_10[411]},
      {stage1_10[210]}
   );
   gpc1_1 gpc2623 (
      {stage0_10[412]},
      {stage1_10[211]}
   );
   gpc1_1 gpc2624 (
      {stage0_10[413]},
      {stage1_10[212]}
   );
   gpc1_1 gpc2625 (
      {stage0_10[414]},
      {stage1_10[213]}
   );
   gpc1_1 gpc2626 (
      {stage0_10[415]},
      {stage1_10[214]}
   );
   gpc1_1 gpc2627 (
      {stage0_10[416]},
      {stage1_10[215]}
   );
   gpc1_1 gpc2628 (
      {stage0_10[417]},
      {stage1_10[216]}
   );
   gpc1_1 gpc2629 (
      {stage0_10[418]},
      {stage1_10[217]}
   );
   gpc1_1 gpc2630 (
      {stage0_10[419]},
      {stage1_10[218]}
   );
   gpc1_1 gpc2631 (
      {stage0_10[420]},
      {stage1_10[219]}
   );
   gpc1_1 gpc2632 (
      {stage0_10[421]},
      {stage1_10[220]}
   );
   gpc1_1 gpc2633 (
      {stage0_10[422]},
      {stage1_10[221]}
   );
   gpc1_1 gpc2634 (
      {stage0_10[423]},
      {stage1_10[222]}
   );
   gpc1_1 gpc2635 (
      {stage0_10[424]},
      {stage1_10[223]}
   );
   gpc1_1 gpc2636 (
      {stage0_10[425]},
      {stage1_10[224]}
   );
   gpc1_1 gpc2637 (
      {stage0_10[426]},
      {stage1_10[225]}
   );
   gpc1_1 gpc2638 (
      {stage0_10[427]},
      {stage1_10[226]}
   );
   gpc1_1 gpc2639 (
      {stage0_10[428]},
      {stage1_10[227]}
   );
   gpc1_1 gpc2640 (
      {stage0_10[429]},
      {stage1_10[228]}
   );
   gpc1_1 gpc2641 (
      {stage0_10[430]},
      {stage1_10[229]}
   );
   gpc1_1 gpc2642 (
      {stage0_10[431]},
      {stage1_10[230]}
   );
   gpc1_1 gpc2643 (
      {stage0_10[432]},
      {stage1_10[231]}
   );
   gpc1_1 gpc2644 (
      {stage0_10[433]},
      {stage1_10[232]}
   );
   gpc1_1 gpc2645 (
      {stage0_10[434]},
      {stage1_10[233]}
   );
   gpc1_1 gpc2646 (
      {stage0_10[435]},
      {stage1_10[234]}
   );
   gpc1_1 gpc2647 (
      {stage0_10[436]},
      {stage1_10[235]}
   );
   gpc1_1 gpc2648 (
      {stage0_10[437]},
      {stage1_10[236]}
   );
   gpc1_1 gpc2649 (
      {stage0_10[438]},
      {stage1_10[237]}
   );
   gpc1_1 gpc2650 (
      {stage0_10[439]},
      {stage1_10[238]}
   );
   gpc1_1 gpc2651 (
      {stage0_10[440]},
      {stage1_10[239]}
   );
   gpc1_1 gpc2652 (
      {stage0_10[441]},
      {stage1_10[240]}
   );
   gpc1_1 gpc2653 (
      {stage0_10[442]},
      {stage1_10[241]}
   );
   gpc1_1 gpc2654 (
      {stage0_10[443]},
      {stage1_10[242]}
   );
   gpc1_1 gpc2655 (
      {stage0_10[444]},
      {stage1_10[243]}
   );
   gpc1_1 gpc2656 (
      {stage0_10[445]},
      {stage1_10[244]}
   );
   gpc1_1 gpc2657 (
      {stage0_10[446]},
      {stage1_10[245]}
   );
   gpc1_1 gpc2658 (
      {stage0_10[447]},
      {stage1_10[246]}
   );
   gpc1_1 gpc2659 (
      {stage0_10[448]},
      {stage1_10[247]}
   );
   gpc1_1 gpc2660 (
      {stage0_10[449]},
      {stage1_10[248]}
   );
   gpc1_1 gpc2661 (
      {stage0_10[450]},
      {stage1_10[249]}
   );
   gpc1_1 gpc2662 (
      {stage0_10[451]},
      {stage1_10[250]}
   );
   gpc1_1 gpc2663 (
      {stage0_10[452]},
      {stage1_10[251]}
   );
   gpc1_1 gpc2664 (
      {stage0_10[453]},
      {stage1_10[252]}
   );
   gpc1_1 gpc2665 (
      {stage0_10[454]},
      {stage1_10[253]}
   );
   gpc1_1 gpc2666 (
      {stage0_10[455]},
      {stage1_10[254]}
   );
   gpc1_1 gpc2667 (
      {stage0_10[456]},
      {stage1_10[255]}
   );
   gpc1_1 gpc2668 (
      {stage0_10[457]},
      {stage1_10[256]}
   );
   gpc1_1 gpc2669 (
      {stage0_10[458]},
      {stage1_10[257]}
   );
   gpc1_1 gpc2670 (
      {stage0_10[459]},
      {stage1_10[258]}
   );
   gpc1_1 gpc2671 (
      {stage0_10[460]},
      {stage1_10[259]}
   );
   gpc1_1 gpc2672 (
      {stage0_10[461]},
      {stage1_10[260]}
   );
   gpc1_1 gpc2673 (
      {stage0_10[462]},
      {stage1_10[261]}
   );
   gpc1_1 gpc2674 (
      {stage0_10[463]},
      {stage1_10[262]}
   );
   gpc1_1 gpc2675 (
      {stage0_10[464]},
      {stage1_10[263]}
   );
   gpc1_1 gpc2676 (
      {stage0_10[465]},
      {stage1_10[264]}
   );
   gpc1_1 gpc2677 (
      {stage0_10[466]},
      {stage1_10[265]}
   );
   gpc1_1 gpc2678 (
      {stage0_10[467]},
      {stage1_10[266]}
   );
   gpc1_1 gpc2679 (
      {stage0_10[468]},
      {stage1_10[267]}
   );
   gpc1_1 gpc2680 (
      {stage0_10[469]},
      {stage1_10[268]}
   );
   gpc1_1 gpc2681 (
      {stage0_10[470]},
      {stage1_10[269]}
   );
   gpc1_1 gpc2682 (
      {stage0_10[471]},
      {stage1_10[270]}
   );
   gpc1_1 gpc2683 (
      {stage0_10[472]},
      {stage1_10[271]}
   );
   gpc1_1 gpc2684 (
      {stage0_10[473]},
      {stage1_10[272]}
   );
   gpc1_1 gpc2685 (
      {stage0_10[474]},
      {stage1_10[273]}
   );
   gpc1_1 gpc2686 (
      {stage0_10[475]},
      {stage1_10[274]}
   );
   gpc1_1 gpc2687 (
      {stage0_10[476]},
      {stage1_10[275]}
   );
   gpc1_1 gpc2688 (
      {stage0_10[477]},
      {stage1_10[276]}
   );
   gpc1_1 gpc2689 (
      {stage0_10[478]},
      {stage1_10[277]}
   );
   gpc1_1 gpc2690 (
      {stage0_10[479]},
      {stage1_10[278]}
   );
   gpc1_1 gpc2691 (
      {stage0_10[480]},
      {stage1_10[279]}
   );
   gpc1_1 gpc2692 (
      {stage0_10[481]},
      {stage1_10[280]}
   );
   gpc1_1 gpc2693 (
      {stage0_10[482]},
      {stage1_10[281]}
   );
   gpc1_1 gpc2694 (
      {stage0_10[483]},
      {stage1_10[282]}
   );
   gpc1_1 gpc2695 (
      {stage0_10[484]},
      {stage1_10[283]}
   );
   gpc1_1 gpc2696 (
      {stage0_10[485]},
      {stage1_10[284]}
   );
   gpc1_1 gpc2697 (
      {stage0_11[367]},
      {stage1_11[158]}
   );
   gpc1_1 gpc2698 (
      {stage0_11[368]},
      {stage1_11[159]}
   );
   gpc1_1 gpc2699 (
      {stage0_11[369]},
      {stage1_11[160]}
   );
   gpc1_1 gpc2700 (
      {stage0_11[370]},
      {stage1_11[161]}
   );
   gpc1_1 gpc2701 (
      {stage0_11[371]},
      {stage1_11[162]}
   );
   gpc1_1 gpc2702 (
      {stage0_11[372]},
      {stage1_11[163]}
   );
   gpc1_1 gpc2703 (
      {stage0_11[373]},
      {stage1_11[164]}
   );
   gpc1_1 gpc2704 (
      {stage0_11[374]},
      {stage1_11[165]}
   );
   gpc1_1 gpc2705 (
      {stage0_11[375]},
      {stage1_11[166]}
   );
   gpc1_1 gpc2706 (
      {stage0_11[376]},
      {stage1_11[167]}
   );
   gpc1_1 gpc2707 (
      {stage0_11[377]},
      {stage1_11[168]}
   );
   gpc1_1 gpc2708 (
      {stage0_11[378]},
      {stage1_11[169]}
   );
   gpc1_1 gpc2709 (
      {stage0_11[379]},
      {stage1_11[170]}
   );
   gpc1_1 gpc2710 (
      {stage0_11[380]},
      {stage1_11[171]}
   );
   gpc1_1 gpc2711 (
      {stage0_11[381]},
      {stage1_11[172]}
   );
   gpc1_1 gpc2712 (
      {stage0_11[382]},
      {stage1_11[173]}
   );
   gpc1_1 gpc2713 (
      {stage0_11[383]},
      {stage1_11[174]}
   );
   gpc1_1 gpc2714 (
      {stage0_11[384]},
      {stage1_11[175]}
   );
   gpc1_1 gpc2715 (
      {stage0_11[385]},
      {stage1_11[176]}
   );
   gpc1_1 gpc2716 (
      {stage0_11[386]},
      {stage1_11[177]}
   );
   gpc1_1 gpc2717 (
      {stage0_11[387]},
      {stage1_11[178]}
   );
   gpc1_1 gpc2718 (
      {stage0_11[388]},
      {stage1_11[179]}
   );
   gpc1_1 gpc2719 (
      {stage0_11[389]},
      {stage1_11[180]}
   );
   gpc1_1 gpc2720 (
      {stage0_11[390]},
      {stage1_11[181]}
   );
   gpc1_1 gpc2721 (
      {stage0_11[391]},
      {stage1_11[182]}
   );
   gpc1_1 gpc2722 (
      {stage0_11[392]},
      {stage1_11[183]}
   );
   gpc1_1 gpc2723 (
      {stage0_11[393]},
      {stage1_11[184]}
   );
   gpc1_1 gpc2724 (
      {stage0_11[394]},
      {stage1_11[185]}
   );
   gpc1_1 gpc2725 (
      {stage0_11[395]},
      {stage1_11[186]}
   );
   gpc1_1 gpc2726 (
      {stage0_11[396]},
      {stage1_11[187]}
   );
   gpc1_1 gpc2727 (
      {stage0_11[397]},
      {stage1_11[188]}
   );
   gpc1_1 gpc2728 (
      {stage0_11[398]},
      {stage1_11[189]}
   );
   gpc1_1 gpc2729 (
      {stage0_11[399]},
      {stage1_11[190]}
   );
   gpc1_1 gpc2730 (
      {stage0_11[400]},
      {stage1_11[191]}
   );
   gpc1_1 gpc2731 (
      {stage0_11[401]},
      {stage1_11[192]}
   );
   gpc1_1 gpc2732 (
      {stage0_11[402]},
      {stage1_11[193]}
   );
   gpc1_1 gpc2733 (
      {stage0_11[403]},
      {stage1_11[194]}
   );
   gpc1_1 gpc2734 (
      {stage0_11[404]},
      {stage1_11[195]}
   );
   gpc1_1 gpc2735 (
      {stage0_11[405]},
      {stage1_11[196]}
   );
   gpc1_1 gpc2736 (
      {stage0_11[406]},
      {stage1_11[197]}
   );
   gpc1_1 gpc2737 (
      {stage0_11[407]},
      {stage1_11[198]}
   );
   gpc1_1 gpc2738 (
      {stage0_11[408]},
      {stage1_11[199]}
   );
   gpc1_1 gpc2739 (
      {stage0_11[409]},
      {stage1_11[200]}
   );
   gpc1_1 gpc2740 (
      {stage0_11[410]},
      {stage1_11[201]}
   );
   gpc1_1 gpc2741 (
      {stage0_11[411]},
      {stage1_11[202]}
   );
   gpc1_1 gpc2742 (
      {stage0_11[412]},
      {stage1_11[203]}
   );
   gpc1_1 gpc2743 (
      {stage0_11[413]},
      {stage1_11[204]}
   );
   gpc1_1 gpc2744 (
      {stage0_11[414]},
      {stage1_11[205]}
   );
   gpc1_1 gpc2745 (
      {stage0_11[415]},
      {stage1_11[206]}
   );
   gpc1_1 gpc2746 (
      {stage0_11[416]},
      {stage1_11[207]}
   );
   gpc1_1 gpc2747 (
      {stage0_11[417]},
      {stage1_11[208]}
   );
   gpc1_1 gpc2748 (
      {stage0_11[418]},
      {stage1_11[209]}
   );
   gpc1_1 gpc2749 (
      {stage0_11[419]},
      {stage1_11[210]}
   );
   gpc1_1 gpc2750 (
      {stage0_11[420]},
      {stage1_11[211]}
   );
   gpc1_1 gpc2751 (
      {stage0_11[421]},
      {stage1_11[212]}
   );
   gpc1_1 gpc2752 (
      {stage0_11[422]},
      {stage1_11[213]}
   );
   gpc1_1 gpc2753 (
      {stage0_11[423]},
      {stage1_11[214]}
   );
   gpc1_1 gpc2754 (
      {stage0_11[424]},
      {stage1_11[215]}
   );
   gpc1_1 gpc2755 (
      {stage0_11[425]},
      {stage1_11[216]}
   );
   gpc1_1 gpc2756 (
      {stage0_11[426]},
      {stage1_11[217]}
   );
   gpc1_1 gpc2757 (
      {stage0_11[427]},
      {stage1_11[218]}
   );
   gpc1_1 gpc2758 (
      {stage0_11[428]},
      {stage1_11[219]}
   );
   gpc1_1 gpc2759 (
      {stage0_11[429]},
      {stage1_11[220]}
   );
   gpc1_1 gpc2760 (
      {stage0_11[430]},
      {stage1_11[221]}
   );
   gpc1_1 gpc2761 (
      {stage0_11[431]},
      {stage1_11[222]}
   );
   gpc1_1 gpc2762 (
      {stage0_11[432]},
      {stage1_11[223]}
   );
   gpc1_1 gpc2763 (
      {stage0_11[433]},
      {stage1_11[224]}
   );
   gpc1_1 gpc2764 (
      {stage0_11[434]},
      {stage1_11[225]}
   );
   gpc1_1 gpc2765 (
      {stage0_11[435]},
      {stage1_11[226]}
   );
   gpc1_1 gpc2766 (
      {stage0_11[436]},
      {stage1_11[227]}
   );
   gpc1_1 gpc2767 (
      {stage0_11[437]},
      {stage1_11[228]}
   );
   gpc1_1 gpc2768 (
      {stage0_11[438]},
      {stage1_11[229]}
   );
   gpc1_1 gpc2769 (
      {stage0_11[439]},
      {stage1_11[230]}
   );
   gpc1_1 gpc2770 (
      {stage0_11[440]},
      {stage1_11[231]}
   );
   gpc1_1 gpc2771 (
      {stage0_11[441]},
      {stage1_11[232]}
   );
   gpc1_1 gpc2772 (
      {stage0_11[442]},
      {stage1_11[233]}
   );
   gpc1_1 gpc2773 (
      {stage0_11[443]},
      {stage1_11[234]}
   );
   gpc1_1 gpc2774 (
      {stage0_11[444]},
      {stage1_11[235]}
   );
   gpc1_1 gpc2775 (
      {stage0_11[445]},
      {stage1_11[236]}
   );
   gpc1_1 gpc2776 (
      {stage0_11[446]},
      {stage1_11[237]}
   );
   gpc1_1 gpc2777 (
      {stage0_11[447]},
      {stage1_11[238]}
   );
   gpc1_1 gpc2778 (
      {stage0_11[448]},
      {stage1_11[239]}
   );
   gpc1_1 gpc2779 (
      {stage0_11[449]},
      {stage1_11[240]}
   );
   gpc1_1 gpc2780 (
      {stage0_11[450]},
      {stage1_11[241]}
   );
   gpc1_1 gpc2781 (
      {stage0_11[451]},
      {stage1_11[242]}
   );
   gpc1_1 gpc2782 (
      {stage0_11[452]},
      {stage1_11[243]}
   );
   gpc1_1 gpc2783 (
      {stage0_11[453]},
      {stage1_11[244]}
   );
   gpc1_1 gpc2784 (
      {stage0_11[454]},
      {stage1_11[245]}
   );
   gpc1_1 gpc2785 (
      {stage0_11[455]},
      {stage1_11[246]}
   );
   gpc1_1 gpc2786 (
      {stage0_11[456]},
      {stage1_11[247]}
   );
   gpc1_1 gpc2787 (
      {stage0_11[457]},
      {stage1_11[248]}
   );
   gpc1_1 gpc2788 (
      {stage0_11[458]},
      {stage1_11[249]}
   );
   gpc1_1 gpc2789 (
      {stage0_11[459]},
      {stage1_11[250]}
   );
   gpc1_1 gpc2790 (
      {stage0_11[460]},
      {stage1_11[251]}
   );
   gpc1_1 gpc2791 (
      {stage0_11[461]},
      {stage1_11[252]}
   );
   gpc1_1 gpc2792 (
      {stage0_11[462]},
      {stage1_11[253]}
   );
   gpc1_1 gpc2793 (
      {stage0_11[463]},
      {stage1_11[254]}
   );
   gpc1_1 gpc2794 (
      {stage0_11[464]},
      {stage1_11[255]}
   );
   gpc1_1 gpc2795 (
      {stage0_11[465]},
      {stage1_11[256]}
   );
   gpc1_1 gpc2796 (
      {stage0_11[466]},
      {stage1_11[257]}
   );
   gpc1_1 gpc2797 (
      {stage0_11[467]},
      {stage1_11[258]}
   );
   gpc1_1 gpc2798 (
      {stage0_11[468]},
      {stage1_11[259]}
   );
   gpc1_1 gpc2799 (
      {stage0_11[469]},
      {stage1_11[260]}
   );
   gpc1_1 gpc2800 (
      {stage0_11[470]},
      {stage1_11[261]}
   );
   gpc1_1 gpc2801 (
      {stage0_11[471]},
      {stage1_11[262]}
   );
   gpc1_1 gpc2802 (
      {stage0_11[472]},
      {stage1_11[263]}
   );
   gpc1_1 gpc2803 (
      {stage0_11[473]},
      {stage1_11[264]}
   );
   gpc1_1 gpc2804 (
      {stage0_11[474]},
      {stage1_11[265]}
   );
   gpc1_1 gpc2805 (
      {stage0_11[475]},
      {stage1_11[266]}
   );
   gpc1_1 gpc2806 (
      {stage0_11[476]},
      {stage1_11[267]}
   );
   gpc1_1 gpc2807 (
      {stage0_11[477]},
      {stage1_11[268]}
   );
   gpc1_1 gpc2808 (
      {stage0_11[478]},
      {stage1_11[269]}
   );
   gpc1_1 gpc2809 (
      {stage0_11[479]},
      {stage1_11[270]}
   );
   gpc1_1 gpc2810 (
      {stage0_11[480]},
      {stage1_11[271]}
   );
   gpc1_1 gpc2811 (
      {stage0_11[481]},
      {stage1_11[272]}
   );
   gpc1_1 gpc2812 (
      {stage0_11[482]},
      {stage1_11[273]}
   );
   gpc1_1 gpc2813 (
      {stage0_11[483]},
      {stage1_11[274]}
   );
   gpc1_1 gpc2814 (
      {stage0_11[484]},
      {stage1_11[275]}
   );
   gpc1_1 gpc2815 (
      {stage0_11[485]},
      {stage1_11[276]}
   );
   gpc1_1 gpc2816 (
      {stage0_12[484]},
      {stage1_12[187]}
   );
   gpc1_1 gpc2817 (
      {stage0_12[485]},
      {stage1_12[188]}
   );
   gpc1_1 gpc2818 (
      {stage0_13[376]},
      {stage1_13[195]}
   );
   gpc1_1 gpc2819 (
      {stage0_13[377]},
      {stage1_13[196]}
   );
   gpc1_1 gpc2820 (
      {stage0_13[378]},
      {stage1_13[197]}
   );
   gpc1_1 gpc2821 (
      {stage0_13[379]},
      {stage1_13[198]}
   );
   gpc1_1 gpc2822 (
      {stage0_13[380]},
      {stage1_13[199]}
   );
   gpc1_1 gpc2823 (
      {stage0_13[381]},
      {stage1_13[200]}
   );
   gpc1_1 gpc2824 (
      {stage0_13[382]},
      {stage1_13[201]}
   );
   gpc1_1 gpc2825 (
      {stage0_13[383]},
      {stage1_13[202]}
   );
   gpc1_1 gpc2826 (
      {stage0_13[384]},
      {stage1_13[203]}
   );
   gpc1_1 gpc2827 (
      {stage0_13[385]},
      {stage1_13[204]}
   );
   gpc1_1 gpc2828 (
      {stage0_13[386]},
      {stage1_13[205]}
   );
   gpc1_1 gpc2829 (
      {stage0_13[387]},
      {stage1_13[206]}
   );
   gpc1_1 gpc2830 (
      {stage0_13[388]},
      {stage1_13[207]}
   );
   gpc1_1 gpc2831 (
      {stage0_13[389]},
      {stage1_13[208]}
   );
   gpc1_1 gpc2832 (
      {stage0_13[390]},
      {stage1_13[209]}
   );
   gpc1_1 gpc2833 (
      {stage0_13[391]},
      {stage1_13[210]}
   );
   gpc1_1 gpc2834 (
      {stage0_13[392]},
      {stage1_13[211]}
   );
   gpc1_1 gpc2835 (
      {stage0_13[393]},
      {stage1_13[212]}
   );
   gpc1_1 gpc2836 (
      {stage0_13[394]},
      {stage1_13[213]}
   );
   gpc1_1 gpc2837 (
      {stage0_13[395]},
      {stage1_13[214]}
   );
   gpc1_1 gpc2838 (
      {stage0_13[396]},
      {stage1_13[215]}
   );
   gpc1_1 gpc2839 (
      {stage0_13[397]},
      {stage1_13[216]}
   );
   gpc1_1 gpc2840 (
      {stage0_13[398]},
      {stage1_13[217]}
   );
   gpc1_1 gpc2841 (
      {stage0_13[399]},
      {stage1_13[218]}
   );
   gpc1_1 gpc2842 (
      {stage0_13[400]},
      {stage1_13[219]}
   );
   gpc1_1 gpc2843 (
      {stage0_13[401]},
      {stage1_13[220]}
   );
   gpc1_1 gpc2844 (
      {stage0_13[402]},
      {stage1_13[221]}
   );
   gpc1_1 gpc2845 (
      {stage0_13[403]},
      {stage1_13[222]}
   );
   gpc1_1 gpc2846 (
      {stage0_13[404]},
      {stage1_13[223]}
   );
   gpc1_1 gpc2847 (
      {stage0_13[405]},
      {stage1_13[224]}
   );
   gpc1_1 gpc2848 (
      {stage0_13[406]},
      {stage1_13[225]}
   );
   gpc1_1 gpc2849 (
      {stage0_13[407]},
      {stage1_13[226]}
   );
   gpc1_1 gpc2850 (
      {stage0_13[408]},
      {stage1_13[227]}
   );
   gpc1_1 gpc2851 (
      {stage0_13[409]},
      {stage1_13[228]}
   );
   gpc1_1 gpc2852 (
      {stage0_13[410]},
      {stage1_13[229]}
   );
   gpc1_1 gpc2853 (
      {stage0_13[411]},
      {stage1_13[230]}
   );
   gpc1_1 gpc2854 (
      {stage0_13[412]},
      {stage1_13[231]}
   );
   gpc1_1 gpc2855 (
      {stage0_13[413]},
      {stage1_13[232]}
   );
   gpc1_1 gpc2856 (
      {stage0_13[414]},
      {stage1_13[233]}
   );
   gpc1_1 gpc2857 (
      {stage0_13[415]},
      {stage1_13[234]}
   );
   gpc1_1 gpc2858 (
      {stage0_13[416]},
      {stage1_13[235]}
   );
   gpc1_1 gpc2859 (
      {stage0_13[417]},
      {stage1_13[236]}
   );
   gpc1_1 gpc2860 (
      {stage0_13[418]},
      {stage1_13[237]}
   );
   gpc1_1 gpc2861 (
      {stage0_13[419]},
      {stage1_13[238]}
   );
   gpc1_1 gpc2862 (
      {stage0_13[420]},
      {stage1_13[239]}
   );
   gpc1_1 gpc2863 (
      {stage0_13[421]},
      {stage1_13[240]}
   );
   gpc1_1 gpc2864 (
      {stage0_13[422]},
      {stage1_13[241]}
   );
   gpc1_1 gpc2865 (
      {stage0_13[423]},
      {stage1_13[242]}
   );
   gpc1_1 gpc2866 (
      {stage0_13[424]},
      {stage1_13[243]}
   );
   gpc1_1 gpc2867 (
      {stage0_13[425]},
      {stage1_13[244]}
   );
   gpc1_1 gpc2868 (
      {stage0_13[426]},
      {stage1_13[245]}
   );
   gpc1_1 gpc2869 (
      {stage0_13[427]},
      {stage1_13[246]}
   );
   gpc1_1 gpc2870 (
      {stage0_13[428]},
      {stage1_13[247]}
   );
   gpc1_1 gpc2871 (
      {stage0_13[429]},
      {stage1_13[248]}
   );
   gpc1_1 gpc2872 (
      {stage0_13[430]},
      {stage1_13[249]}
   );
   gpc1_1 gpc2873 (
      {stage0_13[431]},
      {stage1_13[250]}
   );
   gpc1_1 gpc2874 (
      {stage0_13[432]},
      {stage1_13[251]}
   );
   gpc1_1 gpc2875 (
      {stage0_13[433]},
      {stage1_13[252]}
   );
   gpc1_1 gpc2876 (
      {stage0_13[434]},
      {stage1_13[253]}
   );
   gpc1_1 gpc2877 (
      {stage0_13[435]},
      {stage1_13[254]}
   );
   gpc1_1 gpc2878 (
      {stage0_13[436]},
      {stage1_13[255]}
   );
   gpc1_1 gpc2879 (
      {stage0_13[437]},
      {stage1_13[256]}
   );
   gpc1_1 gpc2880 (
      {stage0_13[438]},
      {stage1_13[257]}
   );
   gpc1_1 gpc2881 (
      {stage0_13[439]},
      {stage1_13[258]}
   );
   gpc1_1 gpc2882 (
      {stage0_13[440]},
      {stage1_13[259]}
   );
   gpc1_1 gpc2883 (
      {stage0_13[441]},
      {stage1_13[260]}
   );
   gpc1_1 gpc2884 (
      {stage0_13[442]},
      {stage1_13[261]}
   );
   gpc1_1 gpc2885 (
      {stage0_13[443]},
      {stage1_13[262]}
   );
   gpc1_1 gpc2886 (
      {stage0_13[444]},
      {stage1_13[263]}
   );
   gpc1_1 gpc2887 (
      {stage0_13[445]},
      {stage1_13[264]}
   );
   gpc1_1 gpc2888 (
      {stage0_13[446]},
      {stage1_13[265]}
   );
   gpc1_1 gpc2889 (
      {stage0_13[447]},
      {stage1_13[266]}
   );
   gpc1_1 gpc2890 (
      {stage0_13[448]},
      {stage1_13[267]}
   );
   gpc1_1 gpc2891 (
      {stage0_13[449]},
      {stage1_13[268]}
   );
   gpc1_1 gpc2892 (
      {stage0_13[450]},
      {stage1_13[269]}
   );
   gpc1_1 gpc2893 (
      {stage0_13[451]},
      {stage1_13[270]}
   );
   gpc1_1 gpc2894 (
      {stage0_13[452]},
      {stage1_13[271]}
   );
   gpc1_1 gpc2895 (
      {stage0_13[453]},
      {stage1_13[272]}
   );
   gpc1_1 gpc2896 (
      {stage0_13[454]},
      {stage1_13[273]}
   );
   gpc1_1 gpc2897 (
      {stage0_13[455]},
      {stage1_13[274]}
   );
   gpc1_1 gpc2898 (
      {stage0_13[456]},
      {stage1_13[275]}
   );
   gpc1_1 gpc2899 (
      {stage0_13[457]},
      {stage1_13[276]}
   );
   gpc1_1 gpc2900 (
      {stage0_13[458]},
      {stage1_13[277]}
   );
   gpc1_1 gpc2901 (
      {stage0_13[459]},
      {stage1_13[278]}
   );
   gpc1_1 gpc2902 (
      {stage0_13[460]},
      {stage1_13[279]}
   );
   gpc1_1 gpc2903 (
      {stage0_13[461]},
      {stage1_13[280]}
   );
   gpc1_1 gpc2904 (
      {stage0_13[462]},
      {stage1_13[281]}
   );
   gpc1_1 gpc2905 (
      {stage0_13[463]},
      {stage1_13[282]}
   );
   gpc1_1 gpc2906 (
      {stage0_13[464]},
      {stage1_13[283]}
   );
   gpc1_1 gpc2907 (
      {stage0_13[465]},
      {stage1_13[284]}
   );
   gpc1_1 gpc2908 (
      {stage0_13[466]},
      {stage1_13[285]}
   );
   gpc1_1 gpc2909 (
      {stage0_13[467]},
      {stage1_13[286]}
   );
   gpc1_1 gpc2910 (
      {stage0_13[468]},
      {stage1_13[287]}
   );
   gpc1_1 gpc2911 (
      {stage0_13[469]},
      {stage1_13[288]}
   );
   gpc1_1 gpc2912 (
      {stage0_13[470]},
      {stage1_13[289]}
   );
   gpc1_1 gpc2913 (
      {stage0_13[471]},
      {stage1_13[290]}
   );
   gpc1_1 gpc2914 (
      {stage0_13[472]},
      {stage1_13[291]}
   );
   gpc1_1 gpc2915 (
      {stage0_13[473]},
      {stage1_13[292]}
   );
   gpc1_1 gpc2916 (
      {stage0_13[474]},
      {stage1_13[293]}
   );
   gpc1_1 gpc2917 (
      {stage0_13[475]},
      {stage1_13[294]}
   );
   gpc1_1 gpc2918 (
      {stage0_13[476]},
      {stage1_13[295]}
   );
   gpc1_1 gpc2919 (
      {stage0_13[477]},
      {stage1_13[296]}
   );
   gpc1_1 gpc2920 (
      {stage0_13[478]},
      {stage1_13[297]}
   );
   gpc1_1 gpc2921 (
      {stage0_13[479]},
      {stage1_13[298]}
   );
   gpc1_1 gpc2922 (
      {stage0_13[480]},
      {stage1_13[299]}
   );
   gpc1_1 gpc2923 (
      {stage0_13[481]},
      {stage1_13[300]}
   );
   gpc1_1 gpc2924 (
      {stage0_13[482]},
      {stage1_13[301]}
   );
   gpc1_1 gpc2925 (
      {stage0_13[483]},
      {stage1_13[302]}
   );
   gpc1_1 gpc2926 (
      {stage0_13[484]},
      {stage1_13[303]}
   );
   gpc1_1 gpc2927 (
      {stage0_13[485]},
      {stage1_13[304]}
   );
   gpc1_1 gpc2928 (
      {stage0_14[419]},
      {stage1_14[152]}
   );
   gpc1_1 gpc2929 (
      {stage0_14[420]},
      {stage1_14[153]}
   );
   gpc1_1 gpc2930 (
      {stage0_14[421]},
      {stage1_14[154]}
   );
   gpc1_1 gpc2931 (
      {stage0_14[422]},
      {stage1_14[155]}
   );
   gpc1_1 gpc2932 (
      {stage0_14[423]},
      {stage1_14[156]}
   );
   gpc1_1 gpc2933 (
      {stage0_14[424]},
      {stage1_14[157]}
   );
   gpc1_1 gpc2934 (
      {stage0_14[425]},
      {stage1_14[158]}
   );
   gpc1_1 gpc2935 (
      {stage0_14[426]},
      {stage1_14[159]}
   );
   gpc1_1 gpc2936 (
      {stage0_14[427]},
      {stage1_14[160]}
   );
   gpc1_1 gpc2937 (
      {stage0_14[428]},
      {stage1_14[161]}
   );
   gpc1_1 gpc2938 (
      {stage0_14[429]},
      {stage1_14[162]}
   );
   gpc1_1 gpc2939 (
      {stage0_14[430]},
      {stage1_14[163]}
   );
   gpc1_1 gpc2940 (
      {stage0_14[431]},
      {stage1_14[164]}
   );
   gpc1_1 gpc2941 (
      {stage0_14[432]},
      {stage1_14[165]}
   );
   gpc1_1 gpc2942 (
      {stage0_14[433]},
      {stage1_14[166]}
   );
   gpc1_1 gpc2943 (
      {stage0_14[434]},
      {stage1_14[167]}
   );
   gpc1_1 gpc2944 (
      {stage0_14[435]},
      {stage1_14[168]}
   );
   gpc1_1 gpc2945 (
      {stage0_14[436]},
      {stage1_14[169]}
   );
   gpc1_1 gpc2946 (
      {stage0_14[437]},
      {stage1_14[170]}
   );
   gpc1_1 gpc2947 (
      {stage0_14[438]},
      {stage1_14[171]}
   );
   gpc1_1 gpc2948 (
      {stage0_14[439]},
      {stage1_14[172]}
   );
   gpc1_1 gpc2949 (
      {stage0_14[440]},
      {stage1_14[173]}
   );
   gpc1_1 gpc2950 (
      {stage0_14[441]},
      {stage1_14[174]}
   );
   gpc1_1 gpc2951 (
      {stage0_14[442]},
      {stage1_14[175]}
   );
   gpc1_1 gpc2952 (
      {stage0_14[443]},
      {stage1_14[176]}
   );
   gpc1_1 gpc2953 (
      {stage0_14[444]},
      {stage1_14[177]}
   );
   gpc1_1 gpc2954 (
      {stage0_14[445]},
      {stage1_14[178]}
   );
   gpc1_1 gpc2955 (
      {stage0_14[446]},
      {stage1_14[179]}
   );
   gpc1_1 gpc2956 (
      {stage0_14[447]},
      {stage1_14[180]}
   );
   gpc1_1 gpc2957 (
      {stage0_14[448]},
      {stage1_14[181]}
   );
   gpc1_1 gpc2958 (
      {stage0_14[449]},
      {stage1_14[182]}
   );
   gpc1_1 gpc2959 (
      {stage0_14[450]},
      {stage1_14[183]}
   );
   gpc1_1 gpc2960 (
      {stage0_14[451]},
      {stage1_14[184]}
   );
   gpc1_1 gpc2961 (
      {stage0_14[452]},
      {stage1_14[185]}
   );
   gpc1_1 gpc2962 (
      {stage0_14[453]},
      {stage1_14[186]}
   );
   gpc1_1 gpc2963 (
      {stage0_14[454]},
      {stage1_14[187]}
   );
   gpc1_1 gpc2964 (
      {stage0_14[455]},
      {stage1_14[188]}
   );
   gpc1_1 gpc2965 (
      {stage0_14[456]},
      {stage1_14[189]}
   );
   gpc1_1 gpc2966 (
      {stage0_14[457]},
      {stage1_14[190]}
   );
   gpc1_1 gpc2967 (
      {stage0_14[458]},
      {stage1_14[191]}
   );
   gpc1_1 gpc2968 (
      {stage0_14[459]},
      {stage1_14[192]}
   );
   gpc1_1 gpc2969 (
      {stage0_14[460]},
      {stage1_14[193]}
   );
   gpc1_1 gpc2970 (
      {stage0_14[461]},
      {stage1_14[194]}
   );
   gpc1_1 gpc2971 (
      {stage0_14[462]},
      {stage1_14[195]}
   );
   gpc1_1 gpc2972 (
      {stage0_14[463]},
      {stage1_14[196]}
   );
   gpc1_1 gpc2973 (
      {stage0_14[464]},
      {stage1_14[197]}
   );
   gpc1_1 gpc2974 (
      {stage0_14[465]},
      {stage1_14[198]}
   );
   gpc1_1 gpc2975 (
      {stage0_14[466]},
      {stage1_14[199]}
   );
   gpc1_1 gpc2976 (
      {stage0_14[467]},
      {stage1_14[200]}
   );
   gpc1_1 gpc2977 (
      {stage0_14[468]},
      {stage1_14[201]}
   );
   gpc1_1 gpc2978 (
      {stage0_14[469]},
      {stage1_14[202]}
   );
   gpc1_1 gpc2979 (
      {stage0_14[470]},
      {stage1_14[203]}
   );
   gpc1_1 gpc2980 (
      {stage0_14[471]},
      {stage1_14[204]}
   );
   gpc1_1 gpc2981 (
      {stage0_14[472]},
      {stage1_14[205]}
   );
   gpc1_1 gpc2982 (
      {stage0_14[473]},
      {stage1_14[206]}
   );
   gpc1_1 gpc2983 (
      {stage0_14[474]},
      {stage1_14[207]}
   );
   gpc1_1 gpc2984 (
      {stage0_14[475]},
      {stage1_14[208]}
   );
   gpc1_1 gpc2985 (
      {stage0_14[476]},
      {stage1_14[209]}
   );
   gpc1_1 gpc2986 (
      {stage0_14[477]},
      {stage1_14[210]}
   );
   gpc1_1 gpc2987 (
      {stage0_14[478]},
      {stage1_14[211]}
   );
   gpc1_1 gpc2988 (
      {stage0_14[479]},
      {stage1_14[212]}
   );
   gpc1_1 gpc2989 (
      {stage0_14[480]},
      {stage1_14[213]}
   );
   gpc1_1 gpc2990 (
      {stage0_14[481]},
      {stage1_14[214]}
   );
   gpc1_1 gpc2991 (
      {stage0_14[482]},
      {stage1_14[215]}
   );
   gpc1_1 gpc2992 (
      {stage0_14[483]},
      {stage1_14[216]}
   );
   gpc1_1 gpc2993 (
      {stage0_14[484]},
      {stage1_14[217]}
   );
   gpc1_1 gpc2994 (
      {stage0_14[485]},
      {stage1_14[218]}
   );
   gpc1_1 gpc2995 (
      {stage0_15[479]},
      {stage1_15[164]}
   );
   gpc1_1 gpc2996 (
      {stage0_15[480]},
      {stage1_15[165]}
   );
   gpc1_1 gpc2997 (
      {stage0_15[481]},
      {stage1_15[166]}
   );
   gpc1_1 gpc2998 (
      {stage0_15[482]},
      {stage1_15[167]}
   );
   gpc1_1 gpc2999 (
      {stage0_15[483]},
      {stage1_15[168]}
   );
   gpc1_1 gpc3000 (
      {stage0_15[484]},
      {stage1_15[169]}
   );
   gpc1_1 gpc3001 (
      {stage0_15[485]},
      {stage1_15[170]}
   );
   gpc1_1 gpc3002 (
      {stage0_17[450]},
      {stage1_17[193]}
   );
   gpc1_1 gpc3003 (
      {stage0_17[451]},
      {stage1_17[194]}
   );
   gpc1_1 gpc3004 (
      {stage0_17[452]},
      {stage1_17[195]}
   );
   gpc1_1 gpc3005 (
      {stage0_17[453]},
      {stage1_17[196]}
   );
   gpc1_1 gpc3006 (
      {stage0_17[454]},
      {stage1_17[197]}
   );
   gpc1_1 gpc3007 (
      {stage0_17[455]},
      {stage1_17[198]}
   );
   gpc1_1 gpc3008 (
      {stage0_17[456]},
      {stage1_17[199]}
   );
   gpc1_1 gpc3009 (
      {stage0_17[457]},
      {stage1_17[200]}
   );
   gpc1_1 gpc3010 (
      {stage0_17[458]},
      {stage1_17[201]}
   );
   gpc1_1 gpc3011 (
      {stage0_17[459]},
      {stage1_17[202]}
   );
   gpc1_1 gpc3012 (
      {stage0_17[460]},
      {stage1_17[203]}
   );
   gpc1_1 gpc3013 (
      {stage0_17[461]},
      {stage1_17[204]}
   );
   gpc1_1 gpc3014 (
      {stage0_17[462]},
      {stage1_17[205]}
   );
   gpc1_1 gpc3015 (
      {stage0_17[463]},
      {stage1_17[206]}
   );
   gpc1_1 gpc3016 (
      {stage0_17[464]},
      {stage1_17[207]}
   );
   gpc1_1 gpc3017 (
      {stage0_17[465]},
      {stage1_17[208]}
   );
   gpc1_1 gpc3018 (
      {stage0_17[466]},
      {stage1_17[209]}
   );
   gpc1_1 gpc3019 (
      {stage0_17[467]},
      {stage1_17[210]}
   );
   gpc1_1 gpc3020 (
      {stage0_17[468]},
      {stage1_17[211]}
   );
   gpc1_1 gpc3021 (
      {stage0_17[469]},
      {stage1_17[212]}
   );
   gpc1_1 gpc3022 (
      {stage0_17[470]},
      {stage1_17[213]}
   );
   gpc1_1 gpc3023 (
      {stage0_17[471]},
      {stage1_17[214]}
   );
   gpc1_1 gpc3024 (
      {stage0_17[472]},
      {stage1_17[215]}
   );
   gpc1_1 gpc3025 (
      {stage0_17[473]},
      {stage1_17[216]}
   );
   gpc1_1 gpc3026 (
      {stage0_17[474]},
      {stage1_17[217]}
   );
   gpc1_1 gpc3027 (
      {stage0_17[475]},
      {stage1_17[218]}
   );
   gpc1_1 gpc3028 (
      {stage0_17[476]},
      {stage1_17[219]}
   );
   gpc1_1 gpc3029 (
      {stage0_17[477]},
      {stage1_17[220]}
   );
   gpc1_1 gpc3030 (
      {stage0_17[478]},
      {stage1_17[221]}
   );
   gpc1_1 gpc3031 (
      {stage0_17[479]},
      {stage1_17[222]}
   );
   gpc1_1 gpc3032 (
      {stage0_17[480]},
      {stage1_17[223]}
   );
   gpc1_1 gpc3033 (
      {stage0_17[481]},
      {stage1_17[224]}
   );
   gpc1_1 gpc3034 (
      {stage0_17[482]},
      {stage1_17[225]}
   );
   gpc1_1 gpc3035 (
      {stage0_17[483]},
      {stage1_17[226]}
   );
   gpc1_1 gpc3036 (
      {stage0_17[484]},
      {stage1_17[227]}
   );
   gpc1_1 gpc3037 (
      {stage0_17[485]},
      {stage1_17[228]}
   );
   gpc1_1 gpc3038 (
      {stage0_18[426]},
      {stage1_18[149]}
   );
   gpc1_1 gpc3039 (
      {stage0_18[427]},
      {stage1_18[150]}
   );
   gpc1_1 gpc3040 (
      {stage0_18[428]},
      {stage1_18[151]}
   );
   gpc1_1 gpc3041 (
      {stage0_18[429]},
      {stage1_18[152]}
   );
   gpc1_1 gpc3042 (
      {stage0_18[430]},
      {stage1_18[153]}
   );
   gpc1_1 gpc3043 (
      {stage0_18[431]},
      {stage1_18[154]}
   );
   gpc1_1 gpc3044 (
      {stage0_18[432]},
      {stage1_18[155]}
   );
   gpc1_1 gpc3045 (
      {stage0_18[433]},
      {stage1_18[156]}
   );
   gpc1_1 gpc3046 (
      {stage0_18[434]},
      {stage1_18[157]}
   );
   gpc1_1 gpc3047 (
      {stage0_18[435]},
      {stage1_18[158]}
   );
   gpc1_1 gpc3048 (
      {stage0_18[436]},
      {stage1_18[159]}
   );
   gpc1_1 gpc3049 (
      {stage0_18[437]},
      {stage1_18[160]}
   );
   gpc1_1 gpc3050 (
      {stage0_18[438]},
      {stage1_18[161]}
   );
   gpc1_1 gpc3051 (
      {stage0_18[439]},
      {stage1_18[162]}
   );
   gpc1_1 gpc3052 (
      {stage0_18[440]},
      {stage1_18[163]}
   );
   gpc1_1 gpc3053 (
      {stage0_18[441]},
      {stage1_18[164]}
   );
   gpc1_1 gpc3054 (
      {stage0_18[442]},
      {stage1_18[165]}
   );
   gpc1_1 gpc3055 (
      {stage0_18[443]},
      {stage1_18[166]}
   );
   gpc1_1 gpc3056 (
      {stage0_18[444]},
      {stage1_18[167]}
   );
   gpc1_1 gpc3057 (
      {stage0_18[445]},
      {stage1_18[168]}
   );
   gpc1_1 gpc3058 (
      {stage0_18[446]},
      {stage1_18[169]}
   );
   gpc1_1 gpc3059 (
      {stage0_18[447]},
      {stage1_18[170]}
   );
   gpc1_1 gpc3060 (
      {stage0_18[448]},
      {stage1_18[171]}
   );
   gpc1_1 gpc3061 (
      {stage0_18[449]},
      {stage1_18[172]}
   );
   gpc1_1 gpc3062 (
      {stage0_18[450]},
      {stage1_18[173]}
   );
   gpc1_1 gpc3063 (
      {stage0_18[451]},
      {stage1_18[174]}
   );
   gpc1_1 gpc3064 (
      {stage0_18[452]},
      {stage1_18[175]}
   );
   gpc1_1 gpc3065 (
      {stage0_18[453]},
      {stage1_18[176]}
   );
   gpc1_1 gpc3066 (
      {stage0_18[454]},
      {stage1_18[177]}
   );
   gpc1_1 gpc3067 (
      {stage0_18[455]},
      {stage1_18[178]}
   );
   gpc1_1 gpc3068 (
      {stage0_18[456]},
      {stage1_18[179]}
   );
   gpc1_1 gpc3069 (
      {stage0_18[457]},
      {stage1_18[180]}
   );
   gpc1_1 gpc3070 (
      {stage0_18[458]},
      {stage1_18[181]}
   );
   gpc1_1 gpc3071 (
      {stage0_18[459]},
      {stage1_18[182]}
   );
   gpc1_1 gpc3072 (
      {stage0_18[460]},
      {stage1_18[183]}
   );
   gpc1_1 gpc3073 (
      {stage0_18[461]},
      {stage1_18[184]}
   );
   gpc1_1 gpc3074 (
      {stage0_18[462]},
      {stage1_18[185]}
   );
   gpc1_1 gpc3075 (
      {stage0_18[463]},
      {stage1_18[186]}
   );
   gpc1_1 gpc3076 (
      {stage0_18[464]},
      {stage1_18[187]}
   );
   gpc1_1 gpc3077 (
      {stage0_18[465]},
      {stage1_18[188]}
   );
   gpc1_1 gpc3078 (
      {stage0_18[466]},
      {stage1_18[189]}
   );
   gpc1_1 gpc3079 (
      {stage0_18[467]},
      {stage1_18[190]}
   );
   gpc1_1 gpc3080 (
      {stage0_18[468]},
      {stage1_18[191]}
   );
   gpc1_1 gpc3081 (
      {stage0_18[469]},
      {stage1_18[192]}
   );
   gpc1_1 gpc3082 (
      {stage0_18[470]},
      {stage1_18[193]}
   );
   gpc1_1 gpc3083 (
      {stage0_18[471]},
      {stage1_18[194]}
   );
   gpc1_1 gpc3084 (
      {stage0_18[472]},
      {stage1_18[195]}
   );
   gpc1_1 gpc3085 (
      {stage0_18[473]},
      {stage1_18[196]}
   );
   gpc1_1 gpc3086 (
      {stage0_18[474]},
      {stage1_18[197]}
   );
   gpc1_1 gpc3087 (
      {stage0_18[475]},
      {stage1_18[198]}
   );
   gpc1_1 gpc3088 (
      {stage0_18[476]},
      {stage1_18[199]}
   );
   gpc1_1 gpc3089 (
      {stage0_18[477]},
      {stage1_18[200]}
   );
   gpc1_1 gpc3090 (
      {stage0_18[478]},
      {stage1_18[201]}
   );
   gpc1_1 gpc3091 (
      {stage0_18[479]},
      {stage1_18[202]}
   );
   gpc1_1 gpc3092 (
      {stage0_18[480]},
      {stage1_18[203]}
   );
   gpc1_1 gpc3093 (
      {stage0_18[481]},
      {stage1_18[204]}
   );
   gpc1_1 gpc3094 (
      {stage0_18[482]},
      {stage1_18[205]}
   );
   gpc1_1 gpc3095 (
      {stage0_18[483]},
      {stage1_18[206]}
   );
   gpc1_1 gpc3096 (
      {stage0_18[484]},
      {stage1_18[207]}
   );
   gpc1_1 gpc3097 (
      {stage0_18[485]},
      {stage1_18[208]}
   );
   gpc1_1 gpc3098 (
      {stage0_19[397]},
      {stage1_19[187]}
   );
   gpc1_1 gpc3099 (
      {stage0_19[398]},
      {stage1_19[188]}
   );
   gpc1_1 gpc3100 (
      {stage0_19[399]},
      {stage1_19[189]}
   );
   gpc1_1 gpc3101 (
      {stage0_19[400]},
      {stage1_19[190]}
   );
   gpc1_1 gpc3102 (
      {stage0_19[401]},
      {stage1_19[191]}
   );
   gpc1_1 gpc3103 (
      {stage0_19[402]},
      {stage1_19[192]}
   );
   gpc1_1 gpc3104 (
      {stage0_19[403]},
      {stage1_19[193]}
   );
   gpc1_1 gpc3105 (
      {stage0_19[404]},
      {stage1_19[194]}
   );
   gpc1_1 gpc3106 (
      {stage0_19[405]},
      {stage1_19[195]}
   );
   gpc1_1 gpc3107 (
      {stage0_19[406]},
      {stage1_19[196]}
   );
   gpc1_1 gpc3108 (
      {stage0_19[407]},
      {stage1_19[197]}
   );
   gpc1_1 gpc3109 (
      {stage0_19[408]},
      {stage1_19[198]}
   );
   gpc1_1 gpc3110 (
      {stage0_19[409]},
      {stage1_19[199]}
   );
   gpc1_1 gpc3111 (
      {stage0_19[410]},
      {stage1_19[200]}
   );
   gpc1_1 gpc3112 (
      {stage0_19[411]},
      {stage1_19[201]}
   );
   gpc1_1 gpc3113 (
      {stage0_19[412]},
      {stage1_19[202]}
   );
   gpc1_1 gpc3114 (
      {stage0_19[413]},
      {stage1_19[203]}
   );
   gpc1_1 gpc3115 (
      {stage0_19[414]},
      {stage1_19[204]}
   );
   gpc1_1 gpc3116 (
      {stage0_19[415]},
      {stage1_19[205]}
   );
   gpc1_1 gpc3117 (
      {stage0_19[416]},
      {stage1_19[206]}
   );
   gpc1_1 gpc3118 (
      {stage0_19[417]},
      {stage1_19[207]}
   );
   gpc1_1 gpc3119 (
      {stage0_19[418]},
      {stage1_19[208]}
   );
   gpc1_1 gpc3120 (
      {stage0_19[419]},
      {stage1_19[209]}
   );
   gpc1_1 gpc3121 (
      {stage0_19[420]},
      {stage1_19[210]}
   );
   gpc1_1 gpc3122 (
      {stage0_19[421]},
      {stage1_19[211]}
   );
   gpc1_1 gpc3123 (
      {stage0_19[422]},
      {stage1_19[212]}
   );
   gpc1_1 gpc3124 (
      {stage0_19[423]},
      {stage1_19[213]}
   );
   gpc1_1 gpc3125 (
      {stage0_19[424]},
      {stage1_19[214]}
   );
   gpc1_1 gpc3126 (
      {stage0_19[425]},
      {stage1_19[215]}
   );
   gpc1_1 gpc3127 (
      {stage0_19[426]},
      {stage1_19[216]}
   );
   gpc1_1 gpc3128 (
      {stage0_19[427]},
      {stage1_19[217]}
   );
   gpc1_1 gpc3129 (
      {stage0_19[428]},
      {stage1_19[218]}
   );
   gpc1_1 gpc3130 (
      {stage0_19[429]},
      {stage1_19[219]}
   );
   gpc1_1 gpc3131 (
      {stage0_19[430]},
      {stage1_19[220]}
   );
   gpc1_1 gpc3132 (
      {stage0_19[431]},
      {stage1_19[221]}
   );
   gpc1_1 gpc3133 (
      {stage0_19[432]},
      {stage1_19[222]}
   );
   gpc1_1 gpc3134 (
      {stage0_19[433]},
      {stage1_19[223]}
   );
   gpc1_1 gpc3135 (
      {stage0_19[434]},
      {stage1_19[224]}
   );
   gpc1_1 gpc3136 (
      {stage0_19[435]},
      {stage1_19[225]}
   );
   gpc1_1 gpc3137 (
      {stage0_19[436]},
      {stage1_19[226]}
   );
   gpc1_1 gpc3138 (
      {stage0_19[437]},
      {stage1_19[227]}
   );
   gpc1_1 gpc3139 (
      {stage0_19[438]},
      {stage1_19[228]}
   );
   gpc1_1 gpc3140 (
      {stage0_19[439]},
      {stage1_19[229]}
   );
   gpc1_1 gpc3141 (
      {stage0_19[440]},
      {stage1_19[230]}
   );
   gpc1_1 gpc3142 (
      {stage0_19[441]},
      {stage1_19[231]}
   );
   gpc1_1 gpc3143 (
      {stage0_19[442]},
      {stage1_19[232]}
   );
   gpc1_1 gpc3144 (
      {stage0_19[443]},
      {stage1_19[233]}
   );
   gpc1_1 gpc3145 (
      {stage0_19[444]},
      {stage1_19[234]}
   );
   gpc1_1 gpc3146 (
      {stage0_19[445]},
      {stage1_19[235]}
   );
   gpc1_1 gpc3147 (
      {stage0_19[446]},
      {stage1_19[236]}
   );
   gpc1_1 gpc3148 (
      {stage0_19[447]},
      {stage1_19[237]}
   );
   gpc1_1 gpc3149 (
      {stage0_19[448]},
      {stage1_19[238]}
   );
   gpc1_1 gpc3150 (
      {stage0_19[449]},
      {stage1_19[239]}
   );
   gpc1_1 gpc3151 (
      {stage0_19[450]},
      {stage1_19[240]}
   );
   gpc1_1 gpc3152 (
      {stage0_19[451]},
      {stage1_19[241]}
   );
   gpc1_1 gpc3153 (
      {stage0_19[452]},
      {stage1_19[242]}
   );
   gpc1_1 gpc3154 (
      {stage0_19[453]},
      {stage1_19[243]}
   );
   gpc1_1 gpc3155 (
      {stage0_19[454]},
      {stage1_19[244]}
   );
   gpc1_1 gpc3156 (
      {stage0_19[455]},
      {stage1_19[245]}
   );
   gpc1_1 gpc3157 (
      {stage0_19[456]},
      {stage1_19[246]}
   );
   gpc1_1 gpc3158 (
      {stage0_19[457]},
      {stage1_19[247]}
   );
   gpc1_1 gpc3159 (
      {stage0_19[458]},
      {stage1_19[248]}
   );
   gpc1_1 gpc3160 (
      {stage0_19[459]},
      {stage1_19[249]}
   );
   gpc1_1 gpc3161 (
      {stage0_19[460]},
      {stage1_19[250]}
   );
   gpc1_1 gpc3162 (
      {stage0_19[461]},
      {stage1_19[251]}
   );
   gpc1_1 gpc3163 (
      {stage0_19[462]},
      {stage1_19[252]}
   );
   gpc1_1 gpc3164 (
      {stage0_19[463]},
      {stage1_19[253]}
   );
   gpc1_1 gpc3165 (
      {stage0_19[464]},
      {stage1_19[254]}
   );
   gpc1_1 gpc3166 (
      {stage0_19[465]},
      {stage1_19[255]}
   );
   gpc1_1 gpc3167 (
      {stage0_19[466]},
      {stage1_19[256]}
   );
   gpc1_1 gpc3168 (
      {stage0_19[467]},
      {stage1_19[257]}
   );
   gpc1_1 gpc3169 (
      {stage0_19[468]},
      {stage1_19[258]}
   );
   gpc1_1 gpc3170 (
      {stage0_19[469]},
      {stage1_19[259]}
   );
   gpc1_1 gpc3171 (
      {stage0_19[470]},
      {stage1_19[260]}
   );
   gpc1_1 gpc3172 (
      {stage0_19[471]},
      {stage1_19[261]}
   );
   gpc1_1 gpc3173 (
      {stage0_19[472]},
      {stage1_19[262]}
   );
   gpc1_1 gpc3174 (
      {stage0_19[473]},
      {stage1_19[263]}
   );
   gpc1_1 gpc3175 (
      {stage0_19[474]},
      {stage1_19[264]}
   );
   gpc1_1 gpc3176 (
      {stage0_19[475]},
      {stage1_19[265]}
   );
   gpc1_1 gpc3177 (
      {stage0_19[476]},
      {stage1_19[266]}
   );
   gpc1_1 gpc3178 (
      {stage0_19[477]},
      {stage1_19[267]}
   );
   gpc1_1 gpc3179 (
      {stage0_19[478]},
      {stage1_19[268]}
   );
   gpc1_1 gpc3180 (
      {stage0_19[479]},
      {stage1_19[269]}
   );
   gpc1_1 gpc3181 (
      {stage0_19[480]},
      {stage1_19[270]}
   );
   gpc1_1 gpc3182 (
      {stage0_19[481]},
      {stage1_19[271]}
   );
   gpc1_1 gpc3183 (
      {stage0_19[482]},
      {stage1_19[272]}
   );
   gpc1_1 gpc3184 (
      {stage0_19[483]},
      {stage1_19[273]}
   );
   gpc1_1 gpc3185 (
      {stage0_19[484]},
      {stage1_19[274]}
   );
   gpc1_1 gpc3186 (
      {stage0_19[485]},
      {stage1_19[275]}
   );
   gpc1_1 gpc3187 (
      {stage0_20[432]},
      {stage1_20[214]}
   );
   gpc1_1 gpc3188 (
      {stage0_20[433]},
      {stage1_20[215]}
   );
   gpc1_1 gpc3189 (
      {stage0_20[434]},
      {stage1_20[216]}
   );
   gpc1_1 gpc3190 (
      {stage0_20[435]},
      {stage1_20[217]}
   );
   gpc1_1 gpc3191 (
      {stage0_20[436]},
      {stage1_20[218]}
   );
   gpc1_1 gpc3192 (
      {stage0_20[437]},
      {stage1_20[219]}
   );
   gpc1_1 gpc3193 (
      {stage0_20[438]},
      {stage1_20[220]}
   );
   gpc1_1 gpc3194 (
      {stage0_20[439]},
      {stage1_20[221]}
   );
   gpc1_1 gpc3195 (
      {stage0_20[440]},
      {stage1_20[222]}
   );
   gpc1_1 gpc3196 (
      {stage0_20[441]},
      {stage1_20[223]}
   );
   gpc1_1 gpc3197 (
      {stage0_20[442]},
      {stage1_20[224]}
   );
   gpc1_1 gpc3198 (
      {stage0_20[443]},
      {stage1_20[225]}
   );
   gpc1_1 gpc3199 (
      {stage0_20[444]},
      {stage1_20[226]}
   );
   gpc1_1 gpc3200 (
      {stage0_20[445]},
      {stage1_20[227]}
   );
   gpc1_1 gpc3201 (
      {stage0_20[446]},
      {stage1_20[228]}
   );
   gpc1_1 gpc3202 (
      {stage0_20[447]},
      {stage1_20[229]}
   );
   gpc1_1 gpc3203 (
      {stage0_20[448]},
      {stage1_20[230]}
   );
   gpc1_1 gpc3204 (
      {stage0_20[449]},
      {stage1_20[231]}
   );
   gpc1_1 gpc3205 (
      {stage0_20[450]},
      {stage1_20[232]}
   );
   gpc1_1 gpc3206 (
      {stage0_20[451]},
      {stage1_20[233]}
   );
   gpc1_1 gpc3207 (
      {stage0_20[452]},
      {stage1_20[234]}
   );
   gpc1_1 gpc3208 (
      {stage0_20[453]},
      {stage1_20[235]}
   );
   gpc1_1 gpc3209 (
      {stage0_20[454]},
      {stage1_20[236]}
   );
   gpc1_1 gpc3210 (
      {stage0_20[455]},
      {stage1_20[237]}
   );
   gpc1_1 gpc3211 (
      {stage0_20[456]},
      {stage1_20[238]}
   );
   gpc1_1 gpc3212 (
      {stage0_20[457]},
      {stage1_20[239]}
   );
   gpc1_1 gpc3213 (
      {stage0_20[458]},
      {stage1_20[240]}
   );
   gpc1_1 gpc3214 (
      {stage0_20[459]},
      {stage1_20[241]}
   );
   gpc1_1 gpc3215 (
      {stage0_20[460]},
      {stage1_20[242]}
   );
   gpc1_1 gpc3216 (
      {stage0_20[461]},
      {stage1_20[243]}
   );
   gpc1_1 gpc3217 (
      {stage0_20[462]},
      {stage1_20[244]}
   );
   gpc1_1 gpc3218 (
      {stage0_20[463]},
      {stage1_20[245]}
   );
   gpc1_1 gpc3219 (
      {stage0_20[464]},
      {stage1_20[246]}
   );
   gpc1_1 gpc3220 (
      {stage0_20[465]},
      {stage1_20[247]}
   );
   gpc1_1 gpc3221 (
      {stage0_20[466]},
      {stage1_20[248]}
   );
   gpc1_1 gpc3222 (
      {stage0_20[467]},
      {stage1_20[249]}
   );
   gpc1_1 gpc3223 (
      {stage0_20[468]},
      {stage1_20[250]}
   );
   gpc1_1 gpc3224 (
      {stage0_20[469]},
      {stage1_20[251]}
   );
   gpc1_1 gpc3225 (
      {stage0_20[470]},
      {stage1_20[252]}
   );
   gpc1_1 gpc3226 (
      {stage0_20[471]},
      {stage1_20[253]}
   );
   gpc1_1 gpc3227 (
      {stage0_20[472]},
      {stage1_20[254]}
   );
   gpc1_1 gpc3228 (
      {stage0_20[473]},
      {stage1_20[255]}
   );
   gpc1_1 gpc3229 (
      {stage0_20[474]},
      {stage1_20[256]}
   );
   gpc1_1 gpc3230 (
      {stage0_20[475]},
      {stage1_20[257]}
   );
   gpc1_1 gpc3231 (
      {stage0_20[476]},
      {stage1_20[258]}
   );
   gpc1_1 gpc3232 (
      {stage0_20[477]},
      {stage1_20[259]}
   );
   gpc1_1 gpc3233 (
      {stage0_20[478]},
      {stage1_20[260]}
   );
   gpc1_1 gpc3234 (
      {stage0_20[479]},
      {stage1_20[261]}
   );
   gpc1_1 gpc3235 (
      {stage0_20[480]},
      {stage1_20[262]}
   );
   gpc1_1 gpc3236 (
      {stage0_20[481]},
      {stage1_20[263]}
   );
   gpc1_1 gpc3237 (
      {stage0_20[482]},
      {stage1_20[264]}
   );
   gpc1_1 gpc3238 (
      {stage0_20[483]},
      {stage1_20[265]}
   );
   gpc1_1 gpc3239 (
      {stage0_20[484]},
      {stage1_20[266]}
   );
   gpc1_1 gpc3240 (
      {stage0_20[485]},
      {stage1_20[267]}
   );
   gpc1_1 gpc3241 (
      {stage0_21[468]},
      {stage1_21[172]}
   );
   gpc1_1 gpc3242 (
      {stage0_21[469]},
      {stage1_21[173]}
   );
   gpc1_1 gpc3243 (
      {stage0_21[470]},
      {stage1_21[174]}
   );
   gpc1_1 gpc3244 (
      {stage0_21[471]},
      {stage1_21[175]}
   );
   gpc1_1 gpc3245 (
      {stage0_21[472]},
      {stage1_21[176]}
   );
   gpc1_1 gpc3246 (
      {stage0_21[473]},
      {stage1_21[177]}
   );
   gpc1_1 gpc3247 (
      {stage0_21[474]},
      {stage1_21[178]}
   );
   gpc1_1 gpc3248 (
      {stage0_21[475]},
      {stage1_21[179]}
   );
   gpc1_1 gpc3249 (
      {stage0_21[476]},
      {stage1_21[180]}
   );
   gpc1_1 gpc3250 (
      {stage0_21[477]},
      {stage1_21[181]}
   );
   gpc1_1 gpc3251 (
      {stage0_21[478]},
      {stage1_21[182]}
   );
   gpc1_1 gpc3252 (
      {stage0_21[479]},
      {stage1_21[183]}
   );
   gpc1_1 gpc3253 (
      {stage0_21[480]},
      {stage1_21[184]}
   );
   gpc1_1 gpc3254 (
      {stage0_21[481]},
      {stage1_21[185]}
   );
   gpc1_1 gpc3255 (
      {stage0_21[482]},
      {stage1_21[186]}
   );
   gpc1_1 gpc3256 (
      {stage0_21[483]},
      {stage1_21[187]}
   );
   gpc1_1 gpc3257 (
      {stage0_21[484]},
      {stage1_21[188]}
   );
   gpc1_1 gpc3258 (
      {stage0_21[485]},
      {stage1_21[189]}
   );
   gpc1_1 gpc3259 (
      {stage0_22[472]},
      {stage1_22[157]}
   );
   gpc1_1 gpc3260 (
      {stage0_22[473]},
      {stage1_22[158]}
   );
   gpc1_1 gpc3261 (
      {stage0_22[474]},
      {stage1_22[159]}
   );
   gpc1_1 gpc3262 (
      {stage0_22[475]},
      {stage1_22[160]}
   );
   gpc1_1 gpc3263 (
      {stage0_22[476]},
      {stage1_22[161]}
   );
   gpc1_1 gpc3264 (
      {stage0_22[477]},
      {stage1_22[162]}
   );
   gpc1_1 gpc3265 (
      {stage0_22[478]},
      {stage1_22[163]}
   );
   gpc1_1 gpc3266 (
      {stage0_22[479]},
      {stage1_22[164]}
   );
   gpc1_1 gpc3267 (
      {stage0_22[480]},
      {stage1_22[165]}
   );
   gpc1_1 gpc3268 (
      {stage0_22[481]},
      {stage1_22[166]}
   );
   gpc1_1 gpc3269 (
      {stage0_22[482]},
      {stage1_22[167]}
   );
   gpc1_1 gpc3270 (
      {stage0_22[483]},
      {stage1_22[168]}
   );
   gpc1_1 gpc3271 (
      {stage0_22[484]},
      {stage1_22[169]}
   );
   gpc1_1 gpc3272 (
      {stage0_22[485]},
      {stage1_22[170]}
   );
   gpc1_1 gpc3273 (
      {stage0_23[396]},
      {stage1_23[197]}
   );
   gpc1_1 gpc3274 (
      {stage0_23[397]},
      {stage1_23[198]}
   );
   gpc1_1 gpc3275 (
      {stage0_23[398]},
      {stage1_23[199]}
   );
   gpc1_1 gpc3276 (
      {stage0_23[399]},
      {stage1_23[200]}
   );
   gpc1_1 gpc3277 (
      {stage0_23[400]},
      {stage1_23[201]}
   );
   gpc1_1 gpc3278 (
      {stage0_23[401]},
      {stage1_23[202]}
   );
   gpc1_1 gpc3279 (
      {stage0_23[402]},
      {stage1_23[203]}
   );
   gpc1_1 gpc3280 (
      {stage0_23[403]},
      {stage1_23[204]}
   );
   gpc1_1 gpc3281 (
      {stage0_23[404]},
      {stage1_23[205]}
   );
   gpc1_1 gpc3282 (
      {stage0_23[405]},
      {stage1_23[206]}
   );
   gpc1_1 gpc3283 (
      {stage0_23[406]},
      {stage1_23[207]}
   );
   gpc1_1 gpc3284 (
      {stage0_23[407]},
      {stage1_23[208]}
   );
   gpc1_1 gpc3285 (
      {stage0_23[408]},
      {stage1_23[209]}
   );
   gpc1_1 gpc3286 (
      {stage0_23[409]},
      {stage1_23[210]}
   );
   gpc1_1 gpc3287 (
      {stage0_23[410]},
      {stage1_23[211]}
   );
   gpc1_1 gpc3288 (
      {stage0_23[411]},
      {stage1_23[212]}
   );
   gpc1_1 gpc3289 (
      {stage0_23[412]},
      {stage1_23[213]}
   );
   gpc1_1 gpc3290 (
      {stage0_23[413]},
      {stage1_23[214]}
   );
   gpc1_1 gpc3291 (
      {stage0_23[414]},
      {stage1_23[215]}
   );
   gpc1_1 gpc3292 (
      {stage0_23[415]},
      {stage1_23[216]}
   );
   gpc1_1 gpc3293 (
      {stage0_23[416]},
      {stage1_23[217]}
   );
   gpc1_1 gpc3294 (
      {stage0_23[417]},
      {stage1_23[218]}
   );
   gpc1_1 gpc3295 (
      {stage0_23[418]},
      {stage1_23[219]}
   );
   gpc1_1 gpc3296 (
      {stage0_23[419]},
      {stage1_23[220]}
   );
   gpc1_1 gpc3297 (
      {stage0_23[420]},
      {stage1_23[221]}
   );
   gpc1_1 gpc3298 (
      {stage0_23[421]},
      {stage1_23[222]}
   );
   gpc1_1 gpc3299 (
      {stage0_23[422]},
      {stage1_23[223]}
   );
   gpc1_1 gpc3300 (
      {stage0_23[423]},
      {stage1_23[224]}
   );
   gpc1_1 gpc3301 (
      {stage0_23[424]},
      {stage1_23[225]}
   );
   gpc1_1 gpc3302 (
      {stage0_23[425]},
      {stage1_23[226]}
   );
   gpc1_1 gpc3303 (
      {stage0_23[426]},
      {stage1_23[227]}
   );
   gpc1_1 gpc3304 (
      {stage0_23[427]},
      {stage1_23[228]}
   );
   gpc1_1 gpc3305 (
      {stage0_23[428]},
      {stage1_23[229]}
   );
   gpc1_1 gpc3306 (
      {stage0_23[429]},
      {stage1_23[230]}
   );
   gpc1_1 gpc3307 (
      {stage0_23[430]},
      {stage1_23[231]}
   );
   gpc1_1 gpc3308 (
      {stage0_23[431]},
      {stage1_23[232]}
   );
   gpc1_1 gpc3309 (
      {stage0_23[432]},
      {stage1_23[233]}
   );
   gpc1_1 gpc3310 (
      {stage0_23[433]},
      {stage1_23[234]}
   );
   gpc1_1 gpc3311 (
      {stage0_23[434]},
      {stage1_23[235]}
   );
   gpc1_1 gpc3312 (
      {stage0_23[435]},
      {stage1_23[236]}
   );
   gpc1_1 gpc3313 (
      {stage0_23[436]},
      {stage1_23[237]}
   );
   gpc1_1 gpc3314 (
      {stage0_23[437]},
      {stage1_23[238]}
   );
   gpc1_1 gpc3315 (
      {stage0_23[438]},
      {stage1_23[239]}
   );
   gpc1_1 gpc3316 (
      {stage0_23[439]},
      {stage1_23[240]}
   );
   gpc1_1 gpc3317 (
      {stage0_23[440]},
      {stage1_23[241]}
   );
   gpc1_1 gpc3318 (
      {stage0_23[441]},
      {stage1_23[242]}
   );
   gpc1_1 gpc3319 (
      {stage0_23[442]},
      {stage1_23[243]}
   );
   gpc1_1 gpc3320 (
      {stage0_23[443]},
      {stage1_23[244]}
   );
   gpc1_1 gpc3321 (
      {stage0_23[444]},
      {stage1_23[245]}
   );
   gpc1_1 gpc3322 (
      {stage0_23[445]},
      {stage1_23[246]}
   );
   gpc1_1 gpc3323 (
      {stage0_23[446]},
      {stage1_23[247]}
   );
   gpc1_1 gpc3324 (
      {stage0_23[447]},
      {stage1_23[248]}
   );
   gpc1_1 gpc3325 (
      {stage0_23[448]},
      {stage1_23[249]}
   );
   gpc1_1 gpc3326 (
      {stage0_23[449]},
      {stage1_23[250]}
   );
   gpc1_1 gpc3327 (
      {stage0_23[450]},
      {stage1_23[251]}
   );
   gpc1_1 gpc3328 (
      {stage0_23[451]},
      {stage1_23[252]}
   );
   gpc1_1 gpc3329 (
      {stage0_23[452]},
      {stage1_23[253]}
   );
   gpc1_1 gpc3330 (
      {stage0_23[453]},
      {stage1_23[254]}
   );
   gpc1_1 gpc3331 (
      {stage0_23[454]},
      {stage1_23[255]}
   );
   gpc1_1 gpc3332 (
      {stage0_23[455]},
      {stage1_23[256]}
   );
   gpc1_1 gpc3333 (
      {stage0_23[456]},
      {stage1_23[257]}
   );
   gpc1_1 gpc3334 (
      {stage0_23[457]},
      {stage1_23[258]}
   );
   gpc1_1 gpc3335 (
      {stage0_23[458]},
      {stage1_23[259]}
   );
   gpc1_1 gpc3336 (
      {stage0_23[459]},
      {stage1_23[260]}
   );
   gpc1_1 gpc3337 (
      {stage0_23[460]},
      {stage1_23[261]}
   );
   gpc1_1 gpc3338 (
      {stage0_23[461]},
      {stage1_23[262]}
   );
   gpc1_1 gpc3339 (
      {stage0_23[462]},
      {stage1_23[263]}
   );
   gpc1_1 gpc3340 (
      {stage0_23[463]},
      {stage1_23[264]}
   );
   gpc1_1 gpc3341 (
      {stage0_23[464]},
      {stage1_23[265]}
   );
   gpc1_1 gpc3342 (
      {stage0_23[465]},
      {stage1_23[266]}
   );
   gpc1_1 gpc3343 (
      {stage0_23[466]},
      {stage1_23[267]}
   );
   gpc1_1 gpc3344 (
      {stage0_23[467]},
      {stage1_23[268]}
   );
   gpc1_1 gpc3345 (
      {stage0_23[468]},
      {stage1_23[269]}
   );
   gpc1_1 gpc3346 (
      {stage0_23[469]},
      {stage1_23[270]}
   );
   gpc1_1 gpc3347 (
      {stage0_23[470]},
      {stage1_23[271]}
   );
   gpc1_1 gpc3348 (
      {stage0_23[471]},
      {stage1_23[272]}
   );
   gpc1_1 gpc3349 (
      {stage0_23[472]},
      {stage1_23[273]}
   );
   gpc1_1 gpc3350 (
      {stage0_23[473]},
      {stage1_23[274]}
   );
   gpc1_1 gpc3351 (
      {stage0_23[474]},
      {stage1_23[275]}
   );
   gpc1_1 gpc3352 (
      {stage0_23[475]},
      {stage1_23[276]}
   );
   gpc1_1 gpc3353 (
      {stage0_23[476]},
      {stage1_23[277]}
   );
   gpc1_1 gpc3354 (
      {stage0_23[477]},
      {stage1_23[278]}
   );
   gpc1_1 gpc3355 (
      {stage0_23[478]},
      {stage1_23[279]}
   );
   gpc1_1 gpc3356 (
      {stage0_23[479]},
      {stage1_23[280]}
   );
   gpc1_1 gpc3357 (
      {stage0_23[480]},
      {stage1_23[281]}
   );
   gpc1_1 gpc3358 (
      {stage0_23[481]},
      {stage1_23[282]}
   );
   gpc1_1 gpc3359 (
      {stage0_23[482]},
      {stage1_23[283]}
   );
   gpc1_1 gpc3360 (
      {stage0_23[483]},
      {stage1_23[284]}
   );
   gpc1_1 gpc3361 (
      {stage0_23[484]},
      {stage1_23[285]}
   );
   gpc1_1 gpc3362 (
      {stage0_23[485]},
      {stage1_23[286]}
   );
   gpc1_1 gpc3363 (
      {stage0_24[485]},
      {stage1_24[213]}
   );
   gpc1_1 gpc3364 (
      {stage0_26[402]},
      {stage1_26[167]}
   );
   gpc1_1 gpc3365 (
      {stage0_26[403]},
      {stage1_26[168]}
   );
   gpc1_1 gpc3366 (
      {stage0_26[404]},
      {stage1_26[169]}
   );
   gpc1_1 gpc3367 (
      {stage0_26[405]},
      {stage1_26[170]}
   );
   gpc1_1 gpc3368 (
      {stage0_26[406]},
      {stage1_26[171]}
   );
   gpc1_1 gpc3369 (
      {stage0_26[407]},
      {stage1_26[172]}
   );
   gpc1_1 gpc3370 (
      {stage0_26[408]},
      {stage1_26[173]}
   );
   gpc1_1 gpc3371 (
      {stage0_26[409]},
      {stage1_26[174]}
   );
   gpc1_1 gpc3372 (
      {stage0_26[410]},
      {stage1_26[175]}
   );
   gpc1_1 gpc3373 (
      {stage0_26[411]},
      {stage1_26[176]}
   );
   gpc1_1 gpc3374 (
      {stage0_26[412]},
      {stage1_26[177]}
   );
   gpc1_1 gpc3375 (
      {stage0_26[413]},
      {stage1_26[178]}
   );
   gpc1_1 gpc3376 (
      {stage0_26[414]},
      {stage1_26[179]}
   );
   gpc1_1 gpc3377 (
      {stage0_26[415]},
      {stage1_26[180]}
   );
   gpc1_1 gpc3378 (
      {stage0_26[416]},
      {stage1_26[181]}
   );
   gpc1_1 gpc3379 (
      {stage0_26[417]},
      {stage1_26[182]}
   );
   gpc1_1 gpc3380 (
      {stage0_26[418]},
      {stage1_26[183]}
   );
   gpc1_1 gpc3381 (
      {stage0_26[419]},
      {stage1_26[184]}
   );
   gpc1_1 gpc3382 (
      {stage0_26[420]},
      {stage1_26[185]}
   );
   gpc1_1 gpc3383 (
      {stage0_26[421]},
      {stage1_26[186]}
   );
   gpc1_1 gpc3384 (
      {stage0_26[422]},
      {stage1_26[187]}
   );
   gpc1_1 gpc3385 (
      {stage0_26[423]},
      {stage1_26[188]}
   );
   gpc1_1 gpc3386 (
      {stage0_26[424]},
      {stage1_26[189]}
   );
   gpc1_1 gpc3387 (
      {stage0_26[425]},
      {stage1_26[190]}
   );
   gpc1_1 gpc3388 (
      {stage0_26[426]},
      {stage1_26[191]}
   );
   gpc1_1 gpc3389 (
      {stage0_26[427]},
      {stage1_26[192]}
   );
   gpc1_1 gpc3390 (
      {stage0_26[428]},
      {stage1_26[193]}
   );
   gpc1_1 gpc3391 (
      {stage0_26[429]},
      {stage1_26[194]}
   );
   gpc1_1 gpc3392 (
      {stage0_26[430]},
      {stage1_26[195]}
   );
   gpc1_1 gpc3393 (
      {stage0_26[431]},
      {stage1_26[196]}
   );
   gpc1_1 gpc3394 (
      {stage0_26[432]},
      {stage1_26[197]}
   );
   gpc1_1 gpc3395 (
      {stage0_26[433]},
      {stage1_26[198]}
   );
   gpc1_1 gpc3396 (
      {stage0_26[434]},
      {stage1_26[199]}
   );
   gpc1_1 gpc3397 (
      {stage0_26[435]},
      {stage1_26[200]}
   );
   gpc1_1 gpc3398 (
      {stage0_26[436]},
      {stage1_26[201]}
   );
   gpc1_1 gpc3399 (
      {stage0_26[437]},
      {stage1_26[202]}
   );
   gpc1_1 gpc3400 (
      {stage0_26[438]},
      {stage1_26[203]}
   );
   gpc1_1 gpc3401 (
      {stage0_26[439]},
      {stage1_26[204]}
   );
   gpc1_1 gpc3402 (
      {stage0_26[440]},
      {stage1_26[205]}
   );
   gpc1_1 gpc3403 (
      {stage0_26[441]},
      {stage1_26[206]}
   );
   gpc1_1 gpc3404 (
      {stage0_26[442]},
      {stage1_26[207]}
   );
   gpc1_1 gpc3405 (
      {stage0_26[443]},
      {stage1_26[208]}
   );
   gpc1_1 gpc3406 (
      {stage0_26[444]},
      {stage1_26[209]}
   );
   gpc1_1 gpc3407 (
      {stage0_26[445]},
      {stage1_26[210]}
   );
   gpc1_1 gpc3408 (
      {stage0_26[446]},
      {stage1_26[211]}
   );
   gpc1_1 gpc3409 (
      {stage0_26[447]},
      {stage1_26[212]}
   );
   gpc1_1 gpc3410 (
      {stage0_26[448]},
      {stage1_26[213]}
   );
   gpc1_1 gpc3411 (
      {stage0_26[449]},
      {stage1_26[214]}
   );
   gpc1_1 gpc3412 (
      {stage0_26[450]},
      {stage1_26[215]}
   );
   gpc1_1 gpc3413 (
      {stage0_26[451]},
      {stage1_26[216]}
   );
   gpc1_1 gpc3414 (
      {stage0_26[452]},
      {stage1_26[217]}
   );
   gpc1_1 gpc3415 (
      {stage0_26[453]},
      {stage1_26[218]}
   );
   gpc1_1 gpc3416 (
      {stage0_26[454]},
      {stage1_26[219]}
   );
   gpc1_1 gpc3417 (
      {stage0_26[455]},
      {stage1_26[220]}
   );
   gpc1_1 gpc3418 (
      {stage0_26[456]},
      {stage1_26[221]}
   );
   gpc1_1 gpc3419 (
      {stage0_26[457]},
      {stage1_26[222]}
   );
   gpc1_1 gpc3420 (
      {stage0_26[458]},
      {stage1_26[223]}
   );
   gpc1_1 gpc3421 (
      {stage0_26[459]},
      {stage1_26[224]}
   );
   gpc1_1 gpc3422 (
      {stage0_26[460]},
      {stage1_26[225]}
   );
   gpc1_1 gpc3423 (
      {stage0_26[461]},
      {stage1_26[226]}
   );
   gpc1_1 gpc3424 (
      {stage0_26[462]},
      {stage1_26[227]}
   );
   gpc1_1 gpc3425 (
      {stage0_26[463]},
      {stage1_26[228]}
   );
   gpc1_1 gpc3426 (
      {stage0_26[464]},
      {stage1_26[229]}
   );
   gpc1_1 gpc3427 (
      {stage0_26[465]},
      {stage1_26[230]}
   );
   gpc1_1 gpc3428 (
      {stage0_26[466]},
      {stage1_26[231]}
   );
   gpc1_1 gpc3429 (
      {stage0_26[467]},
      {stage1_26[232]}
   );
   gpc1_1 gpc3430 (
      {stage0_26[468]},
      {stage1_26[233]}
   );
   gpc1_1 gpc3431 (
      {stage0_26[469]},
      {stage1_26[234]}
   );
   gpc1_1 gpc3432 (
      {stage0_26[470]},
      {stage1_26[235]}
   );
   gpc1_1 gpc3433 (
      {stage0_26[471]},
      {stage1_26[236]}
   );
   gpc1_1 gpc3434 (
      {stage0_26[472]},
      {stage1_26[237]}
   );
   gpc1_1 gpc3435 (
      {stage0_26[473]},
      {stage1_26[238]}
   );
   gpc1_1 gpc3436 (
      {stage0_26[474]},
      {stage1_26[239]}
   );
   gpc1_1 gpc3437 (
      {stage0_26[475]},
      {stage1_26[240]}
   );
   gpc1_1 gpc3438 (
      {stage0_26[476]},
      {stage1_26[241]}
   );
   gpc1_1 gpc3439 (
      {stage0_26[477]},
      {stage1_26[242]}
   );
   gpc1_1 gpc3440 (
      {stage0_26[478]},
      {stage1_26[243]}
   );
   gpc1_1 gpc3441 (
      {stage0_26[479]},
      {stage1_26[244]}
   );
   gpc1_1 gpc3442 (
      {stage0_26[480]},
      {stage1_26[245]}
   );
   gpc1_1 gpc3443 (
      {stage0_26[481]},
      {stage1_26[246]}
   );
   gpc1_1 gpc3444 (
      {stage0_26[482]},
      {stage1_26[247]}
   );
   gpc1_1 gpc3445 (
      {stage0_26[483]},
      {stage1_26[248]}
   );
   gpc1_1 gpc3446 (
      {stage0_26[484]},
      {stage1_26[249]}
   );
   gpc1_1 gpc3447 (
      {stage0_26[485]},
      {stage1_26[250]}
   );
   gpc1_1 gpc3448 (
      {stage0_27[473]},
      {stage1_27[193]}
   );
   gpc1_1 gpc3449 (
      {stage0_27[474]},
      {stage1_27[194]}
   );
   gpc1_1 gpc3450 (
      {stage0_27[475]},
      {stage1_27[195]}
   );
   gpc1_1 gpc3451 (
      {stage0_27[476]},
      {stage1_27[196]}
   );
   gpc1_1 gpc3452 (
      {stage0_27[477]},
      {stage1_27[197]}
   );
   gpc1_1 gpc3453 (
      {stage0_27[478]},
      {stage1_27[198]}
   );
   gpc1_1 gpc3454 (
      {stage0_27[479]},
      {stage1_27[199]}
   );
   gpc1_1 gpc3455 (
      {stage0_27[480]},
      {stage1_27[200]}
   );
   gpc1_1 gpc3456 (
      {stage0_27[481]},
      {stage1_27[201]}
   );
   gpc1_1 gpc3457 (
      {stage0_27[482]},
      {stage1_27[202]}
   );
   gpc1_1 gpc3458 (
      {stage0_27[483]},
      {stage1_27[203]}
   );
   gpc1_1 gpc3459 (
      {stage0_27[484]},
      {stage1_27[204]}
   );
   gpc1_1 gpc3460 (
      {stage0_27[485]},
      {stage1_27[205]}
   );
   gpc1_1 gpc3461 (
      {stage0_28[475]},
      {stage1_28[213]}
   );
   gpc1_1 gpc3462 (
      {stage0_28[476]},
      {stage1_28[214]}
   );
   gpc1_1 gpc3463 (
      {stage0_28[477]},
      {stage1_28[215]}
   );
   gpc1_1 gpc3464 (
      {stage0_28[478]},
      {stage1_28[216]}
   );
   gpc1_1 gpc3465 (
      {stage0_28[479]},
      {stage1_28[217]}
   );
   gpc1_1 gpc3466 (
      {stage0_28[480]},
      {stage1_28[218]}
   );
   gpc1_1 gpc3467 (
      {stage0_28[481]},
      {stage1_28[219]}
   );
   gpc1_1 gpc3468 (
      {stage0_28[482]},
      {stage1_28[220]}
   );
   gpc1_1 gpc3469 (
      {stage0_28[483]},
      {stage1_28[221]}
   );
   gpc1_1 gpc3470 (
      {stage0_28[484]},
      {stage1_28[222]}
   );
   gpc1_1 gpc3471 (
      {stage0_28[485]},
      {stage1_28[223]}
   );
   gpc1_1 gpc3472 (
      {stage0_29[444]},
      {stage1_29[187]}
   );
   gpc1_1 gpc3473 (
      {stage0_29[445]},
      {stage1_29[188]}
   );
   gpc1_1 gpc3474 (
      {stage0_29[446]},
      {stage1_29[189]}
   );
   gpc1_1 gpc3475 (
      {stage0_29[447]},
      {stage1_29[190]}
   );
   gpc1_1 gpc3476 (
      {stage0_29[448]},
      {stage1_29[191]}
   );
   gpc1_1 gpc3477 (
      {stage0_29[449]},
      {stage1_29[192]}
   );
   gpc1_1 gpc3478 (
      {stage0_29[450]},
      {stage1_29[193]}
   );
   gpc1_1 gpc3479 (
      {stage0_29[451]},
      {stage1_29[194]}
   );
   gpc1_1 gpc3480 (
      {stage0_29[452]},
      {stage1_29[195]}
   );
   gpc1_1 gpc3481 (
      {stage0_29[453]},
      {stage1_29[196]}
   );
   gpc1_1 gpc3482 (
      {stage0_29[454]},
      {stage1_29[197]}
   );
   gpc1_1 gpc3483 (
      {stage0_29[455]},
      {stage1_29[198]}
   );
   gpc1_1 gpc3484 (
      {stage0_29[456]},
      {stage1_29[199]}
   );
   gpc1_1 gpc3485 (
      {stage0_29[457]},
      {stage1_29[200]}
   );
   gpc1_1 gpc3486 (
      {stage0_29[458]},
      {stage1_29[201]}
   );
   gpc1_1 gpc3487 (
      {stage0_29[459]},
      {stage1_29[202]}
   );
   gpc1_1 gpc3488 (
      {stage0_29[460]},
      {stage1_29[203]}
   );
   gpc1_1 gpc3489 (
      {stage0_29[461]},
      {stage1_29[204]}
   );
   gpc1_1 gpc3490 (
      {stage0_29[462]},
      {stage1_29[205]}
   );
   gpc1_1 gpc3491 (
      {stage0_29[463]},
      {stage1_29[206]}
   );
   gpc1_1 gpc3492 (
      {stage0_29[464]},
      {stage1_29[207]}
   );
   gpc1_1 gpc3493 (
      {stage0_29[465]},
      {stage1_29[208]}
   );
   gpc1_1 gpc3494 (
      {stage0_29[466]},
      {stage1_29[209]}
   );
   gpc1_1 gpc3495 (
      {stage0_29[467]},
      {stage1_29[210]}
   );
   gpc1_1 gpc3496 (
      {stage0_29[468]},
      {stage1_29[211]}
   );
   gpc1_1 gpc3497 (
      {stage0_29[469]},
      {stage1_29[212]}
   );
   gpc1_1 gpc3498 (
      {stage0_29[470]},
      {stage1_29[213]}
   );
   gpc1_1 gpc3499 (
      {stage0_29[471]},
      {stage1_29[214]}
   );
   gpc1_1 gpc3500 (
      {stage0_29[472]},
      {stage1_29[215]}
   );
   gpc1_1 gpc3501 (
      {stage0_29[473]},
      {stage1_29[216]}
   );
   gpc1_1 gpc3502 (
      {stage0_29[474]},
      {stage1_29[217]}
   );
   gpc1_1 gpc3503 (
      {stage0_29[475]},
      {stage1_29[218]}
   );
   gpc1_1 gpc3504 (
      {stage0_29[476]},
      {stage1_29[219]}
   );
   gpc1_1 gpc3505 (
      {stage0_29[477]},
      {stage1_29[220]}
   );
   gpc1_1 gpc3506 (
      {stage0_29[478]},
      {stage1_29[221]}
   );
   gpc1_1 gpc3507 (
      {stage0_29[479]},
      {stage1_29[222]}
   );
   gpc1_1 gpc3508 (
      {stage0_29[480]},
      {stage1_29[223]}
   );
   gpc1_1 gpc3509 (
      {stage0_29[481]},
      {stage1_29[224]}
   );
   gpc1_1 gpc3510 (
      {stage0_29[482]},
      {stage1_29[225]}
   );
   gpc1_1 gpc3511 (
      {stage0_29[483]},
      {stage1_29[226]}
   );
   gpc1_1 gpc3512 (
      {stage0_29[484]},
      {stage1_29[227]}
   );
   gpc1_1 gpc3513 (
      {stage0_29[485]},
      {stage1_29[228]}
   );
   gpc1_1 gpc3514 (
      {stage0_30[460]},
      {stage1_30[166]}
   );
   gpc1_1 gpc3515 (
      {stage0_30[461]},
      {stage1_30[167]}
   );
   gpc1_1 gpc3516 (
      {stage0_30[462]},
      {stage1_30[168]}
   );
   gpc1_1 gpc3517 (
      {stage0_30[463]},
      {stage1_30[169]}
   );
   gpc1_1 gpc3518 (
      {stage0_30[464]},
      {stage1_30[170]}
   );
   gpc1_1 gpc3519 (
      {stage0_30[465]},
      {stage1_30[171]}
   );
   gpc1_1 gpc3520 (
      {stage0_30[466]},
      {stage1_30[172]}
   );
   gpc1_1 gpc3521 (
      {stage0_30[467]},
      {stage1_30[173]}
   );
   gpc1_1 gpc3522 (
      {stage0_30[468]},
      {stage1_30[174]}
   );
   gpc1_1 gpc3523 (
      {stage0_30[469]},
      {stage1_30[175]}
   );
   gpc1_1 gpc3524 (
      {stage0_30[470]},
      {stage1_30[176]}
   );
   gpc1_1 gpc3525 (
      {stage0_30[471]},
      {stage1_30[177]}
   );
   gpc1_1 gpc3526 (
      {stage0_30[472]},
      {stage1_30[178]}
   );
   gpc1_1 gpc3527 (
      {stage0_30[473]},
      {stage1_30[179]}
   );
   gpc1_1 gpc3528 (
      {stage0_30[474]},
      {stage1_30[180]}
   );
   gpc1_1 gpc3529 (
      {stage0_30[475]},
      {stage1_30[181]}
   );
   gpc1_1 gpc3530 (
      {stage0_30[476]},
      {stage1_30[182]}
   );
   gpc1_1 gpc3531 (
      {stage0_30[477]},
      {stage1_30[183]}
   );
   gpc1_1 gpc3532 (
      {stage0_30[478]},
      {stage1_30[184]}
   );
   gpc1_1 gpc3533 (
      {stage0_30[479]},
      {stage1_30[185]}
   );
   gpc1_1 gpc3534 (
      {stage0_30[480]},
      {stage1_30[186]}
   );
   gpc1_1 gpc3535 (
      {stage0_30[481]},
      {stage1_30[187]}
   );
   gpc1_1 gpc3536 (
      {stage0_30[482]},
      {stage1_30[188]}
   );
   gpc1_1 gpc3537 (
      {stage0_30[483]},
      {stage1_30[189]}
   );
   gpc1_1 gpc3538 (
      {stage0_30[484]},
      {stage1_30[190]}
   );
   gpc1_1 gpc3539 (
      {stage0_30[485]},
      {stage1_30[191]}
   );
   gpc1_1 gpc3540 (
      {stage0_31[476]},
      {stage1_31[208]}
   );
   gpc1_1 gpc3541 (
      {stage0_31[477]},
      {stage1_31[209]}
   );
   gpc1_1 gpc3542 (
      {stage0_31[478]},
      {stage1_31[210]}
   );
   gpc1_1 gpc3543 (
      {stage0_31[479]},
      {stage1_31[211]}
   );
   gpc1_1 gpc3544 (
      {stage0_31[480]},
      {stage1_31[212]}
   );
   gpc1_1 gpc3545 (
      {stage0_31[481]},
      {stage1_31[213]}
   );
   gpc1_1 gpc3546 (
      {stage0_31[482]},
      {stage1_31[214]}
   );
   gpc1_1 gpc3547 (
      {stage0_31[483]},
      {stage1_31[215]}
   );
   gpc1_1 gpc3548 (
      {stage0_31[484]},
      {stage1_31[216]}
   );
   gpc1_1 gpc3549 (
      {stage0_31[485]},
      {stage1_31[217]}
   );
   gpc1_1 gpc3550 (
      {stage0_33[396]},
      {stage1_33[169]}
   );
   gpc1_1 gpc3551 (
      {stage0_33[397]},
      {stage1_33[170]}
   );
   gpc1_1 gpc3552 (
      {stage0_33[398]},
      {stage1_33[171]}
   );
   gpc1_1 gpc3553 (
      {stage0_33[399]},
      {stage1_33[172]}
   );
   gpc1_1 gpc3554 (
      {stage0_33[400]},
      {stage1_33[173]}
   );
   gpc1_1 gpc3555 (
      {stage0_33[401]},
      {stage1_33[174]}
   );
   gpc1_1 gpc3556 (
      {stage0_33[402]},
      {stage1_33[175]}
   );
   gpc1_1 gpc3557 (
      {stage0_33[403]},
      {stage1_33[176]}
   );
   gpc1_1 gpc3558 (
      {stage0_33[404]},
      {stage1_33[177]}
   );
   gpc1_1 gpc3559 (
      {stage0_33[405]},
      {stage1_33[178]}
   );
   gpc1_1 gpc3560 (
      {stage0_33[406]},
      {stage1_33[179]}
   );
   gpc1_1 gpc3561 (
      {stage0_33[407]},
      {stage1_33[180]}
   );
   gpc1_1 gpc3562 (
      {stage0_33[408]},
      {stage1_33[181]}
   );
   gpc1_1 gpc3563 (
      {stage0_33[409]},
      {stage1_33[182]}
   );
   gpc1_1 gpc3564 (
      {stage0_33[410]},
      {stage1_33[183]}
   );
   gpc1_1 gpc3565 (
      {stage0_33[411]},
      {stage1_33[184]}
   );
   gpc1_1 gpc3566 (
      {stage0_33[412]},
      {stage1_33[185]}
   );
   gpc1_1 gpc3567 (
      {stage0_33[413]},
      {stage1_33[186]}
   );
   gpc1_1 gpc3568 (
      {stage0_33[414]},
      {stage1_33[187]}
   );
   gpc1_1 gpc3569 (
      {stage0_33[415]},
      {stage1_33[188]}
   );
   gpc1_1 gpc3570 (
      {stage0_33[416]},
      {stage1_33[189]}
   );
   gpc1_1 gpc3571 (
      {stage0_33[417]},
      {stage1_33[190]}
   );
   gpc1_1 gpc3572 (
      {stage0_33[418]},
      {stage1_33[191]}
   );
   gpc1_1 gpc3573 (
      {stage0_33[419]},
      {stage1_33[192]}
   );
   gpc1_1 gpc3574 (
      {stage0_33[420]},
      {stage1_33[193]}
   );
   gpc1_1 gpc3575 (
      {stage0_33[421]},
      {stage1_33[194]}
   );
   gpc1_1 gpc3576 (
      {stage0_33[422]},
      {stage1_33[195]}
   );
   gpc1_1 gpc3577 (
      {stage0_33[423]},
      {stage1_33[196]}
   );
   gpc1_1 gpc3578 (
      {stage0_33[424]},
      {stage1_33[197]}
   );
   gpc1_1 gpc3579 (
      {stage0_33[425]},
      {stage1_33[198]}
   );
   gpc1_1 gpc3580 (
      {stage0_33[426]},
      {stage1_33[199]}
   );
   gpc1_1 gpc3581 (
      {stage0_33[427]},
      {stage1_33[200]}
   );
   gpc1_1 gpc3582 (
      {stage0_33[428]},
      {stage1_33[201]}
   );
   gpc1_1 gpc3583 (
      {stage0_33[429]},
      {stage1_33[202]}
   );
   gpc1_1 gpc3584 (
      {stage0_33[430]},
      {stage1_33[203]}
   );
   gpc1_1 gpc3585 (
      {stage0_33[431]},
      {stage1_33[204]}
   );
   gpc1_1 gpc3586 (
      {stage0_33[432]},
      {stage1_33[205]}
   );
   gpc1_1 gpc3587 (
      {stage0_33[433]},
      {stage1_33[206]}
   );
   gpc1_1 gpc3588 (
      {stage0_33[434]},
      {stage1_33[207]}
   );
   gpc1_1 gpc3589 (
      {stage0_33[435]},
      {stage1_33[208]}
   );
   gpc1_1 gpc3590 (
      {stage0_33[436]},
      {stage1_33[209]}
   );
   gpc1_1 gpc3591 (
      {stage0_33[437]},
      {stage1_33[210]}
   );
   gpc1_1 gpc3592 (
      {stage0_33[438]},
      {stage1_33[211]}
   );
   gpc1_1 gpc3593 (
      {stage0_33[439]},
      {stage1_33[212]}
   );
   gpc1_1 gpc3594 (
      {stage0_33[440]},
      {stage1_33[213]}
   );
   gpc1_1 gpc3595 (
      {stage0_33[441]},
      {stage1_33[214]}
   );
   gpc1_1 gpc3596 (
      {stage0_33[442]},
      {stage1_33[215]}
   );
   gpc1_1 gpc3597 (
      {stage0_33[443]},
      {stage1_33[216]}
   );
   gpc1_1 gpc3598 (
      {stage0_33[444]},
      {stage1_33[217]}
   );
   gpc1_1 gpc3599 (
      {stage0_33[445]},
      {stage1_33[218]}
   );
   gpc1_1 gpc3600 (
      {stage0_33[446]},
      {stage1_33[219]}
   );
   gpc1_1 gpc3601 (
      {stage0_33[447]},
      {stage1_33[220]}
   );
   gpc1_1 gpc3602 (
      {stage0_33[448]},
      {stage1_33[221]}
   );
   gpc1_1 gpc3603 (
      {stage0_33[449]},
      {stage1_33[222]}
   );
   gpc1_1 gpc3604 (
      {stage0_33[450]},
      {stage1_33[223]}
   );
   gpc1_1 gpc3605 (
      {stage0_33[451]},
      {stage1_33[224]}
   );
   gpc1_1 gpc3606 (
      {stage0_33[452]},
      {stage1_33[225]}
   );
   gpc1_1 gpc3607 (
      {stage0_33[453]},
      {stage1_33[226]}
   );
   gpc1_1 gpc3608 (
      {stage0_33[454]},
      {stage1_33[227]}
   );
   gpc1_1 gpc3609 (
      {stage0_33[455]},
      {stage1_33[228]}
   );
   gpc1_1 gpc3610 (
      {stage0_33[456]},
      {stage1_33[229]}
   );
   gpc1_1 gpc3611 (
      {stage0_33[457]},
      {stage1_33[230]}
   );
   gpc1_1 gpc3612 (
      {stage0_33[458]},
      {stage1_33[231]}
   );
   gpc1_1 gpc3613 (
      {stage0_33[459]},
      {stage1_33[232]}
   );
   gpc1_1 gpc3614 (
      {stage0_33[460]},
      {stage1_33[233]}
   );
   gpc1_1 gpc3615 (
      {stage0_33[461]},
      {stage1_33[234]}
   );
   gpc1_1 gpc3616 (
      {stage0_33[462]},
      {stage1_33[235]}
   );
   gpc1_1 gpc3617 (
      {stage0_33[463]},
      {stage1_33[236]}
   );
   gpc1_1 gpc3618 (
      {stage0_33[464]},
      {stage1_33[237]}
   );
   gpc1_1 gpc3619 (
      {stage0_33[465]},
      {stage1_33[238]}
   );
   gpc1_1 gpc3620 (
      {stage0_33[466]},
      {stage1_33[239]}
   );
   gpc1_1 gpc3621 (
      {stage0_33[467]},
      {stage1_33[240]}
   );
   gpc1_1 gpc3622 (
      {stage0_33[468]},
      {stage1_33[241]}
   );
   gpc1_1 gpc3623 (
      {stage0_33[469]},
      {stage1_33[242]}
   );
   gpc1_1 gpc3624 (
      {stage0_33[470]},
      {stage1_33[243]}
   );
   gpc1_1 gpc3625 (
      {stage0_33[471]},
      {stage1_33[244]}
   );
   gpc1_1 gpc3626 (
      {stage0_33[472]},
      {stage1_33[245]}
   );
   gpc1_1 gpc3627 (
      {stage0_33[473]},
      {stage1_33[246]}
   );
   gpc1_1 gpc3628 (
      {stage0_33[474]},
      {stage1_33[247]}
   );
   gpc1_1 gpc3629 (
      {stage0_33[475]},
      {stage1_33[248]}
   );
   gpc1_1 gpc3630 (
      {stage0_33[476]},
      {stage1_33[249]}
   );
   gpc1_1 gpc3631 (
      {stage0_33[477]},
      {stage1_33[250]}
   );
   gpc1_1 gpc3632 (
      {stage0_33[478]},
      {stage1_33[251]}
   );
   gpc1_1 gpc3633 (
      {stage0_33[479]},
      {stage1_33[252]}
   );
   gpc1_1 gpc3634 (
      {stage0_33[480]},
      {stage1_33[253]}
   );
   gpc1_1 gpc3635 (
      {stage0_33[481]},
      {stage1_33[254]}
   );
   gpc1_1 gpc3636 (
      {stage0_33[482]},
      {stage1_33[255]}
   );
   gpc1_1 gpc3637 (
      {stage0_33[483]},
      {stage1_33[256]}
   );
   gpc1_1 gpc3638 (
      {stage0_33[484]},
      {stage1_33[257]}
   );
   gpc1_1 gpc3639 (
      {stage0_33[485]},
      {stage1_33[258]}
   );
   gpc1_1 gpc3640 (
      {stage0_35[464]},
      {stage1_35[195]}
   );
   gpc1_1 gpc3641 (
      {stage0_35[465]},
      {stage1_35[196]}
   );
   gpc1_1 gpc3642 (
      {stage0_35[466]},
      {stage1_35[197]}
   );
   gpc1_1 gpc3643 (
      {stage0_35[467]},
      {stage1_35[198]}
   );
   gpc1_1 gpc3644 (
      {stage0_35[468]},
      {stage1_35[199]}
   );
   gpc1_1 gpc3645 (
      {stage0_35[469]},
      {stage1_35[200]}
   );
   gpc1_1 gpc3646 (
      {stage0_35[470]},
      {stage1_35[201]}
   );
   gpc1_1 gpc3647 (
      {stage0_35[471]},
      {stage1_35[202]}
   );
   gpc1_1 gpc3648 (
      {stage0_35[472]},
      {stage1_35[203]}
   );
   gpc1_1 gpc3649 (
      {stage0_35[473]},
      {stage1_35[204]}
   );
   gpc1_1 gpc3650 (
      {stage0_35[474]},
      {stage1_35[205]}
   );
   gpc1_1 gpc3651 (
      {stage0_35[475]},
      {stage1_35[206]}
   );
   gpc1_1 gpc3652 (
      {stage0_35[476]},
      {stage1_35[207]}
   );
   gpc1_1 gpc3653 (
      {stage0_35[477]},
      {stage1_35[208]}
   );
   gpc1_1 gpc3654 (
      {stage0_35[478]},
      {stage1_35[209]}
   );
   gpc1_1 gpc3655 (
      {stage0_35[479]},
      {stage1_35[210]}
   );
   gpc1_1 gpc3656 (
      {stage0_35[480]},
      {stage1_35[211]}
   );
   gpc1_1 gpc3657 (
      {stage0_35[481]},
      {stage1_35[212]}
   );
   gpc1_1 gpc3658 (
      {stage0_35[482]},
      {stage1_35[213]}
   );
   gpc1_1 gpc3659 (
      {stage0_35[483]},
      {stage1_35[214]}
   );
   gpc1_1 gpc3660 (
      {stage0_35[484]},
      {stage1_35[215]}
   );
   gpc1_1 gpc3661 (
      {stage0_35[485]},
      {stage1_35[216]}
   );
   gpc1_1 gpc3662 (
      {stage0_37[355]},
      {stage1_37[177]}
   );
   gpc1_1 gpc3663 (
      {stage0_37[356]},
      {stage1_37[178]}
   );
   gpc1_1 gpc3664 (
      {stage0_37[357]},
      {stage1_37[179]}
   );
   gpc1_1 gpc3665 (
      {stage0_37[358]},
      {stage1_37[180]}
   );
   gpc1_1 gpc3666 (
      {stage0_37[359]},
      {stage1_37[181]}
   );
   gpc1_1 gpc3667 (
      {stage0_37[360]},
      {stage1_37[182]}
   );
   gpc1_1 gpc3668 (
      {stage0_37[361]},
      {stage1_37[183]}
   );
   gpc1_1 gpc3669 (
      {stage0_37[362]},
      {stage1_37[184]}
   );
   gpc1_1 gpc3670 (
      {stage0_37[363]},
      {stage1_37[185]}
   );
   gpc1_1 gpc3671 (
      {stage0_37[364]},
      {stage1_37[186]}
   );
   gpc1_1 gpc3672 (
      {stage0_37[365]},
      {stage1_37[187]}
   );
   gpc1_1 gpc3673 (
      {stage0_37[366]},
      {stage1_37[188]}
   );
   gpc1_1 gpc3674 (
      {stage0_37[367]},
      {stage1_37[189]}
   );
   gpc1_1 gpc3675 (
      {stage0_37[368]},
      {stage1_37[190]}
   );
   gpc1_1 gpc3676 (
      {stage0_37[369]},
      {stage1_37[191]}
   );
   gpc1_1 gpc3677 (
      {stage0_37[370]},
      {stage1_37[192]}
   );
   gpc1_1 gpc3678 (
      {stage0_37[371]},
      {stage1_37[193]}
   );
   gpc1_1 gpc3679 (
      {stage0_37[372]},
      {stage1_37[194]}
   );
   gpc1_1 gpc3680 (
      {stage0_37[373]},
      {stage1_37[195]}
   );
   gpc1_1 gpc3681 (
      {stage0_37[374]},
      {stage1_37[196]}
   );
   gpc1_1 gpc3682 (
      {stage0_37[375]},
      {stage1_37[197]}
   );
   gpc1_1 gpc3683 (
      {stage0_37[376]},
      {stage1_37[198]}
   );
   gpc1_1 gpc3684 (
      {stage0_37[377]},
      {stage1_37[199]}
   );
   gpc1_1 gpc3685 (
      {stage0_37[378]},
      {stage1_37[200]}
   );
   gpc1_1 gpc3686 (
      {stage0_37[379]},
      {stage1_37[201]}
   );
   gpc1_1 gpc3687 (
      {stage0_37[380]},
      {stage1_37[202]}
   );
   gpc1_1 gpc3688 (
      {stage0_37[381]},
      {stage1_37[203]}
   );
   gpc1_1 gpc3689 (
      {stage0_37[382]},
      {stage1_37[204]}
   );
   gpc1_1 gpc3690 (
      {stage0_37[383]},
      {stage1_37[205]}
   );
   gpc1_1 gpc3691 (
      {stage0_37[384]},
      {stage1_37[206]}
   );
   gpc1_1 gpc3692 (
      {stage0_37[385]},
      {stage1_37[207]}
   );
   gpc1_1 gpc3693 (
      {stage0_37[386]},
      {stage1_37[208]}
   );
   gpc1_1 gpc3694 (
      {stage0_37[387]},
      {stage1_37[209]}
   );
   gpc1_1 gpc3695 (
      {stage0_37[388]},
      {stage1_37[210]}
   );
   gpc1_1 gpc3696 (
      {stage0_37[389]},
      {stage1_37[211]}
   );
   gpc1_1 gpc3697 (
      {stage0_37[390]},
      {stage1_37[212]}
   );
   gpc1_1 gpc3698 (
      {stage0_37[391]},
      {stage1_37[213]}
   );
   gpc1_1 gpc3699 (
      {stage0_37[392]},
      {stage1_37[214]}
   );
   gpc1_1 gpc3700 (
      {stage0_37[393]},
      {stage1_37[215]}
   );
   gpc1_1 gpc3701 (
      {stage0_37[394]},
      {stage1_37[216]}
   );
   gpc1_1 gpc3702 (
      {stage0_37[395]},
      {stage1_37[217]}
   );
   gpc1_1 gpc3703 (
      {stage0_37[396]},
      {stage1_37[218]}
   );
   gpc1_1 gpc3704 (
      {stage0_37[397]},
      {stage1_37[219]}
   );
   gpc1_1 gpc3705 (
      {stage0_37[398]},
      {stage1_37[220]}
   );
   gpc1_1 gpc3706 (
      {stage0_37[399]},
      {stage1_37[221]}
   );
   gpc1_1 gpc3707 (
      {stage0_37[400]},
      {stage1_37[222]}
   );
   gpc1_1 gpc3708 (
      {stage0_37[401]},
      {stage1_37[223]}
   );
   gpc1_1 gpc3709 (
      {stage0_37[402]},
      {stage1_37[224]}
   );
   gpc1_1 gpc3710 (
      {stage0_37[403]},
      {stage1_37[225]}
   );
   gpc1_1 gpc3711 (
      {stage0_37[404]},
      {stage1_37[226]}
   );
   gpc1_1 gpc3712 (
      {stage0_37[405]},
      {stage1_37[227]}
   );
   gpc1_1 gpc3713 (
      {stage0_37[406]},
      {stage1_37[228]}
   );
   gpc1_1 gpc3714 (
      {stage0_37[407]},
      {stage1_37[229]}
   );
   gpc1_1 gpc3715 (
      {stage0_37[408]},
      {stage1_37[230]}
   );
   gpc1_1 gpc3716 (
      {stage0_37[409]},
      {stage1_37[231]}
   );
   gpc1_1 gpc3717 (
      {stage0_37[410]},
      {stage1_37[232]}
   );
   gpc1_1 gpc3718 (
      {stage0_37[411]},
      {stage1_37[233]}
   );
   gpc1_1 gpc3719 (
      {stage0_37[412]},
      {stage1_37[234]}
   );
   gpc1_1 gpc3720 (
      {stage0_37[413]},
      {stage1_37[235]}
   );
   gpc1_1 gpc3721 (
      {stage0_37[414]},
      {stage1_37[236]}
   );
   gpc1_1 gpc3722 (
      {stage0_37[415]},
      {stage1_37[237]}
   );
   gpc1_1 gpc3723 (
      {stage0_37[416]},
      {stage1_37[238]}
   );
   gpc1_1 gpc3724 (
      {stage0_37[417]},
      {stage1_37[239]}
   );
   gpc1_1 gpc3725 (
      {stage0_37[418]},
      {stage1_37[240]}
   );
   gpc1_1 gpc3726 (
      {stage0_37[419]},
      {stage1_37[241]}
   );
   gpc1_1 gpc3727 (
      {stage0_37[420]},
      {stage1_37[242]}
   );
   gpc1_1 gpc3728 (
      {stage0_37[421]},
      {stage1_37[243]}
   );
   gpc1_1 gpc3729 (
      {stage0_37[422]},
      {stage1_37[244]}
   );
   gpc1_1 gpc3730 (
      {stage0_37[423]},
      {stage1_37[245]}
   );
   gpc1_1 gpc3731 (
      {stage0_37[424]},
      {stage1_37[246]}
   );
   gpc1_1 gpc3732 (
      {stage0_37[425]},
      {stage1_37[247]}
   );
   gpc1_1 gpc3733 (
      {stage0_37[426]},
      {stage1_37[248]}
   );
   gpc1_1 gpc3734 (
      {stage0_37[427]},
      {stage1_37[249]}
   );
   gpc1_1 gpc3735 (
      {stage0_37[428]},
      {stage1_37[250]}
   );
   gpc1_1 gpc3736 (
      {stage0_37[429]},
      {stage1_37[251]}
   );
   gpc1_1 gpc3737 (
      {stage0_37[430]},
      {stage1_37[252]}
   );
   gpc1_1 gpc3738 (
      {stage0_37[431]},
      {stage1_37[253]}
   );
   gpc1_1 gpc3739 (
      {stage0_37[432]},
      {stage1_37[254]}
   );
   gpc1_1 gpc3740 (
      {stage0_37[433]},
      {stage1_37[255]}
   );
   gpc1_1 gpc3741 (
      {stage0_37[434]},
      {stage1_37[256]}
   );
   gpc1_1 gpc3742 (
      {stage0_37[435]},
      {stage1_37[257]}
   );
   gpc1_1 gpc3743 (
      {stage0_37[436]},
      {stage1_37[258]}
   );
   gpc1_1 gpc3744 (
      {stage0_37[437]},
      {stage1_37[259]}
   );
   gpc1_1 gpc3745 (
      {stage0_37[438]},
      {stage1_37[260]}
   );
   gpc1_1 gpc3746 (
      {stage0_37[439]},
      {stage1_37[261]}
   );
   gpc1_1 gpc3747 (
      {stage0_37[440]},
      {stage1_37[262]}
   );
   gpc1_1 gpc3748 (
      {stage0_37[441]},
      {stage1_37[263]}
   );
   gpc1_1 gpc3749 (
      {stage0_37[442]},
      {stage1_37[264]}
   );
   gpc1_1 gpc3750 (
      {stage0_37[443]},
      {stage1_37[265]}
   );
   gpc1_1 gpc3751 (
      {stage0_37[444]},
      {stage1_37[266]}
   );
   gpc1_1 gpc3752 (
      {stage0_37[445]},
      {stage1_37[267]}
   );
   gpc1_1 gpc3753 (
      {stage0_37[446]},
      {stage1_37[268]}
   );
   gpc1_1 gpc3754 (
      {stage0_37[447]},
      {stage1_37[269]}
   );
   gpc1_1 gpc3755 (
      {stage0_37[448]},
      {stage1_37[270]}
   );
   gpc1_1 gpc3756 (
      {stage0_37[449]},
      {stage1_37[271]}
   );
   gpc1_1 gpc3757 (
      {stage0_37[450]},
      {stage1_37[272]}
   );
   gpc1_1 gpc3758 (
      {stage0_37[451]},
      {stage1_37[273]}
   );
   gpc1_1 gpc3759 (
      {stage0_37[452]},
      {stage1_37[274]}
   );
   gpc1_1 gpc3760 (
      {stage0_37[453]},
      {stage1_37[275]}
   );
   gpc1_1 gpc3761 (
      {stage0_37[454]},
      {stage1_37[276]}
   );
   gpc1_1 gpc3762 (
      {stage0_37[455]},
      {stage1_37[277]}
   );
   gpc1_1 gpc3763 (
      {stage0_37[456]},
      {stage1_37[278]}
   );
   gpc1_1 gpc3764 (
      {stage0_37[457]},
      {stage1_37[279]}
   );
   gpc1_1 gpc3765 (
      {stage0_37[458]},
      {stage1_37[280]}
   );
   gpc1_1 gpc3766 (
      {stage0_37[459]},
      {stage1_37[281]}
   );
   gpc1_1 gpc3767 (
      {stage0_37[460]},
      {stage1_37[282]}
   );
   gpc1_1 gpc3768 (
      {stage0_37[461]},
      {stage1_37[283]}
   );
   gpc1_1 gpc3769 (
      {stage0_37[462]},
      {stage1_37[284]}
   );
   gpc1_1 gpc3770 (
      {stage0_37[463]},
      {stage1_37[285]}
   );
   gpc1_1 gpc3771 (
      {stage0_37[464]},
      {stage1_37[286]}
   );
   gpc1_1 gpc3772 (
      {stage0_37[465]},
      {stage1_37[287]}
   );
   gpc1_1 gpc3773 (
      {stage0_37[466]},
      {stage1_37[288]}
   );
   gpc1_1 gpc3774 (
      {stage0_37[467]},
      {stage1_37[289]}
   );
   gpc1_1 gpc3775 (
      {stage0_37[468]},
      {stage1_37[290]}
   );
   gpc1_1 gpc3776 (
      {stage0_37[469]},
      {stage1_37[291]}
   );
   gpc1_1 gpc3777 (
      {stage0_37[470]},
      {stage1_37[292]}
   );
   gpc1_1 gpc3778 (
      {stage0_37[471]},
      {stage1_37[293]}
   );
   gpc1_1 gpc3779 (
      {stage0_37[472]},
      {stage1_37[294]}
   );
   gpc1_1 gpc3780 (
      {stage0_37[473]},
      {stage1_37[295]}
   );
   gpc1_1 gpc3781 (
      {stage0_37[474]},
      {stage1_37[296]}
   );
   gpc1_1 gpc3782 (
      {stage0_37[475]},
      {stage1_37[297]}
   );
   gpc1_1 gpc3783 (
      {stage0_37[476]},
      {stage1_37[298]}
   );
   gpc1_1 gpc3784 (
      {stage0_37[477]},
      {stage1_37[299]}
   );
   gpc1_1 gpc3785 (
      {stage0_37[478]},
      {stage1_37[300]}
   );
   gpc1_1 gpc3786 (
      {stage0_37[479]},
      {stage1_37[301]}
   );
   gpc1_1 gpc3787 (
      {stage0_37[480]},
      {stage1_37[302]}
   );
   gpc1_1 gpc3788 (
      {stage0_37[481]},
      {stage1_37[303]}
   );
   gpc1_1 gpc3789 (
      {stage0_37[482]},
      {stage1_37[304]}
   );
   gpc1_1 gpc3790 (
      {stage0_37[483]},
      {stage1_37[305]}
   );
   gpc1_1 gpc3791 (
      {stage0_37[484]},
      {stage1_37[306]}
   );
   gpc1_1 gpc3792 (
      {stage0_37[485]},
      {stage1_37[307]}
   );
   gpc1_1 gpc3793 (
      {stage0_38[391]},
      {stage1_38[170]}
   );
   gpc1_1 gpc3794 (
      {stage0_38[392]},
      {stage1_38[171]}
   );
   gpc1_1 gpc3795 (
      {stage0_38[393]},
      {stage1_38[172]}
   );
   gpc1_1 gpc3796 (
      {stage0_38[394]},
      {stage1_38[173]}
   );
   gpc1_1 gpc3797 (
      {stage0_38[395]},
      {stage1_38[174]}
   );
   gpc1_1 gpc3798 (
      {stage0_38[396]},
      {stage1_38[175]}
   );
   gpc1_1 gpc3799 (
      {stage0_38[397]},
      {stage1_38[176]}
   );
   gpc1_1 gpc3800 (
      {stage0_38[398]},
      {stage1_38[177]}
   );
   gpc1_1 gpc3801 (
      {stage0_38[399]},
      {stage1_38[178]}
   );
   gpc1_1 gpc3802 (
      {stage0_38[400]},
      {stage1_38[179]}
   );
   gpc1_1 gpc3803 (
      {stage0_38[401]},
      {stage1_38[180]}
   );
   gpc1_1 gpc3804 (
      {stage0_38[402]},
      {stage1_38[181]}
   );
   gpc1_1 gpc3805 (
      {stage0_38[403]},
      {stage1_38[182]}
   );
   gpc1_1 gpc3806 (
      {stage0_38[404]},
      {stage1_38[183]}
   );
   gpc1_1 gpc3807 (
      {stage0_38[405]},
      {stage1_38[184]}
   );
   gpc1_1 gpc3808 (
      {stage0_38[406]},
      {stage1_38[185]}
   );
   gpc1_1 gpc3809 (
      {stage0_38[407]},
      {stage1_38[186]}
   );
   gpc1_1 gpc3810 (
      {stage0_38[408]},
      {stage1_38[187]}
   );
   gpc1_1 gpc3811 (
      {stage0_38[409]},
      {stage1_38[188]}
   );
   gpc1_1 gpc3812 (
      {stage0_38[410]},
      {stage1_38[189]}
   );
   gpc1_1 gpc3813 (
      {stage0_38[411]},
      {stage1_38[190]}
   );
   gpc1_1 gpc3814 (
      {stage0_38[412]},
      {stage1_38[191]}
   );
   gpc1_1 gpc3815 (
      {stage0_38[413]},
      {stage1_38[192]}
   );
   gpc1_1 gpc3816 (
      {stage0_38[414]},
      {stage1_38[193]}
   );
   gpc1_1 gpc3817 (
      {stage0_38[415]},
      {stage1_38[194]}
   );
   gpc1_1 gpc3818 (
      {stage0_38[416]},
      {stage1_38[195]}
   );
   gpc1_1 gpc3819 (
      {stage0_38[417]},
      {stage1_38[196]}
   );
   gpc1_1 gpc3820 (
      {stage0_38[418]},
      {stage1_38[197]}
   );
   gpc1_1 gpc3821 (
      {stage0_38[419]},
      {stage1_38[198]}
   );
   gpc1_1 gpc3822 (
      {stage0_38[420]},
      {stage1_38[199]}
   );
   gpc1_1 gpc3823 (
      {stage0_38[421]},
      {stage1_38[200]}
   );
   gpc1_1 gpc3824 (
      {stage0_38[422]},
      {stage1_38[201]}
   );
   gpc1_1 gpc3825 (
      {stage0_38[423]},
      {stage1_38[202]}
   );
   gpc1_1 gpc3826 (
      {stage0_38[424]},
      {stage1_38[203]}
   );
   gpc1_1 gpc3827 (
      {stage0_38[425]},
      {stage1_38[204]}
   );
   gpc1_1 gpc3828 (
      {stage0_38[426]},
      {stage1_38[205]}
   );
   gpc1_1 gpc3829 (
      {stage0_38[427]},
      {stage1_38[206]}
   );
   gpc1_1 gpc3830 (
      {stage0_38[428]},
      {stage1_38[207]}
   );
   gpc1_1 gpc3831 (
      {stage0_38[429]},
      {stage1_38[208]}
   );
   gpc1_1 gpc3832 (
      {stage0_38[430]},
      {stage1_38[209]}
   );
   gpc1_1 gpc3833 (
      {stage0_38[431]},
      {stage1_38[210]}
   );
   gpc1_1 gpc3834 (
      {stage0_38[432]},
      {stage1_38[211]}
   );
   gpc1_1 gpc3835 (
      {stage0_38[433]},
      {stage1_38[212]}
   );
   gpc1_1 gpc3836 (
      {stage0_38[434]},
      {stage1_38[213]}
   );
   gpc1_1 gpc3837 (
      {stage0_38[435]},
      {stage1_38[214]}
   );
   gpc1_1 gpc3838 (
      {stage0_38[436]},
      {stage1_38[215]}
   );
   gpc1_1 gpc3839 (
      {stage0_38[437]},
      {stage1_38[216]}
   );
   gpc1_1 gpc3840 (
      {stage0_38[438]},
      {stage1_38[217]}
   );
   gpc1_1 gpc3841 (
      {stage0_38[439]},
      {stage1_38[218]}
   );
   gpc1_1 gpc3842 (
      {stage0_38[440]},
      {stage1_38[219]}
   );
   gpc1_1 gpc3843 (
      {stage0_38[441]},
      {stage1_38[220]}
   );
   gpc1_1 gpc3844 (
      {stage0_38[442]},
      {stage1_38[221]}
   );
   gpc1_1 gpc3845 (
      {stage0_38[443]},
      {stage1_38[222]}
   );
   gpc1_1 gpc3846 (
      {stage0_38[444]},
      {stage1_38[223]}
   );
   gpc1_1 gpc3847 (
      {stage0_38[445]},
      {stage1_38[224]}
   );
   gpc1_1 gpc3848 (
      {stage0_38[446]},
      {stage1_38[225]}
   );
   gpc1_1 gpc3849 (
      {stage0_38[447]},
      {stage1_38[226]}
   );
   gpc1_1 gpc3850 (
      {stage0_38[448]},
      {stage1_38[227]}
   );
   gpc1_1 gpc3851 (
      {stage0_38[449]},
      {stage1_38[228]}
   );
   gpc1_1 gpc3852 (
      {stage0_38[450]},
      {stage1_38[229]}
   );
   gpc1_1 gpc3853 (
      {stage0_38[451]},
      {stage1_38[230]}
   );
   gpc1_1 gpc3854 (
      {stage0_38[452]},
      {stage1_38[231]}
   );
   gpc1_1 gpc3855 (
      {stage0_38[453]},
      {stage1_38[232]}
   );
   gpc1_1 gpc3856 (
      {stage0_38[454]},
      {stage1_38[233]}
   );
   gpc1_1 gpc3857 (
      {stage0_38[455]},
      {stage1_38[234]}
   );
   gpc1_1 gpc3858 (
      {stage0_38[456]},
      {stage1_38[235]}
   );
   gpc1_1 gpc3859 (
      {stage0_38[457]},
      {stage1_38[236]}
   );
   gpc1_1 gpc3860 (
      {stage0_38[458]},
      {stage1_38[237]}
   );
   gpc1_1 gpc3861 (
      {stage0_38[459]},
      {stage1_38[238]}
   );
   gpc1_1 gpc3862 (
      {stage0_38[460]},
      {stage1_38[239]}
   );
   gpc1_1 gpc3863 (
      {stage0_38[461]},
      {stage1_38[240]}
   );
   gpc1_1 gpc3864 (
      {stage0_38[462]},
      {stage1_38[241]}
   );
   gpc1_1 gpc3865 (
      {stage0_38[463]},
      {stage1_38[242]}
   );
   gpc1_1 gpc3866 (
      {stage0_38[464]},
      {stage1_38[243]}
   );
   gpc1_1 gpc3867 (
      {stage0_38[465]},
      {stage1_38[244]}
   );
   gpc1_1 gpc3868 (
      {stage0_38[466]},
      {stage1_38[245]}
   );
   gpc1_1 gpc3869 (
      {stage0_38[467]},
      {stage1_38[246]}
   );
   gpc1_1 gpc3870 (
      {stage0_38[468]},
      {stage1_38[247]}
   );
   gpc1_1 gpc3871 (
      {stage0_38[469]},
      {stage1_38[248]}
   );
   gpc1_1 gpc3872 (
      {stage0_38[470]},
      {stage1_38[249]}
   );
   gpc1_1 gpc3873 (
      {stage0_38[471]},
      {stage1_38[250]}
   );
   gpc1_1 gpc3874 (
      {stage0_38[472]},
      {stage1_38[251]}
   );
   gpc1_1 gpc3875 (
      {stage0_38[473]},
      {stage1_38[252]}
   );
   gpc1_1 gpc3876 (
      {stage0_38[474]},
      {stage1_38[253]}
   );
   gpc1_1 gpc3877 (
      {stage0_38[475]},
      {stage1_38[254]}
   );
   gpc1_1 gpc3878 (
      {stage0_38[476]},
      {stage1_38[255]}
   );
   gpc1_1 gpc3879 (
      {stage0_38[477]},
      {stage1_38[256]}
   );
   gpc1_1 gpc3880 (
      {stage0_38[478]},
      {stage1_38[257]}
   );
   gpc1_1 gpc3881 (
      {stage0_38[479]},
      {stage1_38[258]}
   );
   gpc1_1 gpc3882 (
      {stage0_38[480]},
      {stage1_38[259]}
   );
   gpc1_1 gpc3883 (
      {stage0_38[481]},
      {stage1_38[260]}
   );
   gpc1_1 gpc3884 (
      {stage0_38[482]},
      {stage1_38[261]}
   );
   gpc1_1 gpc3885 (
      {stage0_38[483]},
      {stage1_38[262]}
   );
   gpc1_1 gpc3886 (
      {stage0_38[484]},
      {stage1_38[263]}
   );
   gpc1_1 gpc3887 (
      {stage0_38[485]},
      {stage1_38[264]}
   );
   gpc1_1 gpc3888 (
      {stage0_39[447]},
      {stage1_39[174]}
   );
   gpc1_1 gpc3889 (
      {stage0_39[448]},
      {stage1_39[175]}
   );
   gpc1_1 gpc3890 (
      {stage0_39[449]},
      {stage1_39[176]}
   );
   gpc1_1 gpc3891 (
      {stage0_39[450]},
      {stage1_39[177]}
   );
   gpc1_1 gpc3892 (
      {stage0_39[451]},
      {stage1_39[178]}
   );
   gpc1_1 gpc3893 (
      {stage0_39[452]},
      {stage1_39[179]}
   );
   gpc1_1 gpc3894 (
      {stage0_39[453]},
      {stage1_39[180]}
   );
   gpc1_1 gpc3895 (
      {stage0_39[454]},
      {stage1_39[181]}
   );
   gpc1_1 gpc3896 (
      {stage0_39[455]},
      {stage1_39[182]}
   );
   gpc1_1 gpc3897 (
      {stage0_39[456]},
      {stage1_39[183]}
   );
   gpc1_1 gpc3898 (
      {stage0_39[457]},
      {stage1_39[184]}
   );
   gpc1_1 gpc3899 (
      {stage0_39[458]},
      {stage1_39[185]}
   );
   gpc1_1 gpc3900 (
      {stage0_39[459]},
      {stage1_39[186]}
   );
   gpc1_1 gpc3901 (
      {stage0_39[460]},
      {stage1_39[187]}
   );
   gpc1_1 gpc3902 (
      {stage0_39[461]},
      {stage1_39[188]}
   );
   gpc1_1 gpc3903 (
      {stage0_39[462]},
      {stage1_39[189]}
   );
   gpc1_1 gpc3904 (
      {stage0_39[463]},
      {stage1_39[190]}
   );
   gpc1_1 gpc3905 (
      {stage0_39[464]},
      {stage1_39[191]}
   );
   gpc1_1 gpc3906 (
      {stage0_39[465]},
      {stage1_39[192]}
   );
   gpc1_1 gpc3907 (
      {stage0_39[466]},
      {stage1_39[193]}
   );
   gpc1_1 gpc3908 (
      {stage0_39[467]},
      {stage1_39[194]}
   );
   gpc1_1 gpc3909 (
      {stage0_39[468]},
      {stage1_39[195]}
   );
   gpc1_1 gpc3910 (
      {stage0_39[469]},
      {stage1_39[196]}
   );
   gpc1_1 gpc3911 (
      {stage0_39[470]},
      {stage1_39[197]}
   );
   gpc1_1 gpc3912 (
      {stage0_39[471]},
      {stage1_39[198]}
   );
   gpc1_1 gpc3913 (
      {stage0_39[472]},
      {stage1_39[199]}
   );
   gpc1_1 gpc3914 (
      {stage0_39[473]},
      {stage1_39[200]}
   );
   gpc1_1 gpc3915 (
      {stage0_39[474]},
      {stage1_39[201]}
   );
   gpc1_1 gpc3916 (
      {stage0_39[475]},
      {stage1_39[202]}
   );
   gpc1_1 gpc3917 (
      {stage0_39[476]},
      {stage1_39[203]}
   );
   gpc1_1 gpc3918 (
      {stage0_39[477]},
      {stage1_39[204]}
   );
   gpc1_1 gpc3919 (
      {stage0_39[478]},
      {stage1_39[205]}
   );
   gpc1_1 gpc3920 (
      {stage0_39[479]},
      {stage1_39[206]}
   );
   gpc1_1 gpc3921 (
      {stage0_39[480]},
      {stage1_39[207]}
   );
   gpc1_1 gpc3922 (
      {stage0_39[481]},
      {stage1_39[208]}
   );
   gpc1_1 gpc3923 (
      {stage0_39[482]},
      {stage1_39[209]}
   );
   gpc1_1 gpc3924 (
      {stage0_39[483]},
      {stage1_39[210]}
   );
   gpc1_1 gpc3925 (
      {stage0_39[484]},
      {stage1_39[211]}
   );
   gpc1_1 gpc3926 (
      {stage0_39[485]},
      {stage1_39[212]}
   );
   gpc1_1 gpc3927 (
      {stage0_40[380]},
      {stage1_40[198]}
   );
   gpc1_1 gpc3928 (
      {stage0_40[381]},
      {stage1_40[199]}
   );
   gpc1_1 gpc3929 (
      {stage0_40[382]},
      {stage1_40[200]}
   );
   gpc1_1 gpc3930 (
      {stage0_40[383]},
      {stage1_40[201]}
   );
   gpc1_1 gpc3931 (
      {stage0_40[384]},
      {stage1_40[202]}
   );
   gpc1_1 gpc3932 (
      {stage0_40[385]},
      {stage1_40[203]}
   );
   gpc1_1 gpc3933 (
      {stage0_40[386]},
      {stage1_40[204]}
   );
   gpc1_1 gpc3934 (
      {stage0_40[387]},
      {stage1_40[205]}
   );
   gpc1_1 gpc3935 (
      {stage0_40[388]},
      {stage1_40[206]}
   );
   gpc1_1 gpc3936 (
      {stage0_40[389]},
      {stage1_40[207]}
   );
   gpc1_1 gpc3937 (
      {stage0_40[390]},
      {stage1_40[208]}
   );
   gpc1_1 gpc3938 (
      {stage0_40[391]},
      {stage1_40[209]}
   );
   gpc1_1 gpc3939 (
      {stage0_40[392]},
      {stage1_40[210]}
   );
   gpc1_1 gpc3940 (
      {stage0_40[393]},
      {stage1_40[211]}
   );
   gpc1_1 gpc3941 (
      {stage0_40[394]},
      {stage1_40[212]}
   );
   gpc1_1 gpc3942 (
      {stage0_40[395]},
      {stage1_40[213]}
   );
   gpc1_1 gpc3943 (
      {stage0_40[396]},
      {stage1_40[214]}
   );
   gpc1_1 gpc3944 (
      {stage0_40[397]},
      {stage1_40[215]}
   );
   gpc1_1 gpc3945 (
      {stage0_40[398]},
      {stage1_40[216]}
   );
   gpc1_1 gpc3946 (
      {stage0_40[399]},
      {stage1_40[217]}
   );
   gpc1_1 gpc3947 (
      {stage0_40[400]},
      {stage1_40[218]}
   );
   gpc1_1 gpc3948 (
      {stage0_40[401]},
      {stage1_40[219]}
   );
   gpc1_1 gpc3949 (
      {stage0_40[402]},
      {stage1_40[220]}
   );
   gpc1_1 gpc3950 (
      {stage0_40[403]},
      {stage1_40[221]}
   );
   gpc1_1 gpc3951 (
      {stage0_40[404]},
      {stage1_40[222]}
   );
   gpc1_1 gpc3952 (
      {stage0_40[405]},
      {stage1_40[223]}
   );
   gpc1_1 gpc3953 (
      {stage0_40[406]},
      {stage1_40[224]}
   );
   gpc1_1 gpc3954 (
      {stage0_40[407]},
      {stage1_40[225]}
   );
   gpc1_1 gpc3955 (
      {stage0_40[408]},
      {stage1_40[226]}
   );
   gpc1_1 gpc3956 (
      {stage0_40[409]},
      {stage1_40[227]}
   );
   gpc1_1 gpc3957 (
      {stage0_40[410]},
      {stage1_40[228]}
   );
   gpc1_1 gpc3958 (
      {stage0_40[411]},
      {stage1_40[229]}
   );
   gpc1_1 gpc3959 (
      {stage0_40[412]},
      {stage1_40[230]}
   );
   gpc1_1 gpc3960 (
      {stage0_40[413]},
      {stage1_40[231]}
   );
   gpc1_1 gpc3961 (
      {stage0_40[414]},
      {stage1_40[232]}
   );
   gpc1_1 gpc3962 (
      {stage0_40[415]},
      {stage1_40[233]}
   );
   gpc1_1 gpc3963 (
      {stage0_40[416]},
      {stage1_40[234]}
   );
   gpc1_1 gpc3964 (
      {stage0_40[417]},
      {stage1_40[235]}
   );
   gpc1_1 gpc3965 (
      {stage0_40[418]},
      {stage1_40[236]}
   );
   gpc1_1 gpc3966 (
      {stage0_40[419]},
      {stage1_40[237]}
   );
   gpc1_1 gpc3967 (
      {stage0_40[420]},
      {stage1_40[238]}
   );
   gpc1_1 gpc3968 (
      {stage0_40[421]},
      {stage1_40[239]}
   );
   gpc1_1 gpc3969 (
      {stage0_40[422]},
      {stage1_40[240]}
   );
   gpc1_1 gpc3970 (
      {stage0_40[423]},
      {stage1_40[241]}
   );
   gpc1_1 gpc3971 (
      {stage0_40[424]},
      {stage1_40[242]}
   );
   gpc1_1 gpc3972 (
      {stage0_40[425]},
      {stage1_40[243]}
   );
   gpc1_1 gpc3973 (
      {stage0_40[426]},
      {stage1_40[244]}
   );
   gpc1_1 gpc3974 (
      {stage0_40[427]},
      {stage1_40[245]}
   );
   gpc1_1 gpc3975 (
      {stage0_40[428]},
      {stage1_40[246]}
   );
   gpc1_1 gpc3976 (
      {stage0_40[429]},
      {stage1_40[247]}
   );
   gpc1_1 gpc3977 (
      {stage0_40[430]},
      {stage1_40[248]}
   );
   gpc1_1 gpc3978 (
      {stage0_40[431]},
      {stage1_40[249]}
   );
   gpc1_1 gpc3979 (
      {stage0_40[432]},
      {stage1_40[250]}
   );
   gpc1_1 gpc3980 (
      {stage0_40[433]},
      {stage1_40[251]}
   );
   gpc1_1 gpc3981 (
      {stage0_40[434]},
      {stage1_40[252]}
   );
   gpc1_1 gpc3982 (
      {stage0_40[435]},
      {stage1_40[253]}
   );
   gpc1_1 gpc3983 (
      {stage0_40[436]},
      {stage1_40[254]}
   );
   gpc1_1 gpc3984 (
      {stage0_40[437]},
      {stage1_40[255]}
   );
   gpc1_1 gpc3985 (
      {stage0_40[438]},
      {stage1_40[256]}
   );
   gpc1_1 gpc3986 (
      {stage0_40[439]},
      {stage1_40[257]}
   );
   gpc1_1 gpc3987 (
      {stage0_40[440]},
      {stage1_40[258]}
   );
   gpc1_1 gpc3988 (
      {stage0_40[441]},
      {stage1_40[259]}
   );
   gpc1_1 gpc3989 (
      {stage0_40[442]},
      {stage1_40[260]}
   );
   gpc1_1 gpc3990 (
      {stage0_40[443]},
      {stage1_40[261]}
   );
   gpc1_1 gpc3991 (
      {stage0_40[444]},
      {stage1_40[262]}
   );
   gpc1_1 gpc3992 (
      {stage0_40[445]},
      {stage1_40[263]}
   );
   gpc1_1 gpc3993 (
      {stage0_40[446]},
      {stage1_40[264]}
   );
   gpc1_1 gpc3994 (
      {stage0_40[447]},
      {stage1_40[265]}
   );
   gpc1_1 gpc3995 (
      {stage0_40[448]},
      {stage1_40[266]}
   );
   gpc1_1 gpc3996 (
      {stage0_40[449]},
      {stage1_40[267]}
   );
   gpc1_1 gpc3997 (
      {stage0_40[450]},
      {stage1_40[268]}
   );
   gpc1_1 gpc3998 (
      {stage0_40[451]},
      {stage1_40[269]}
   );
   gpc1_1 gpc3999 (
      {stage0_40[452]},
      {stage1_40[270]}
   );
   gpc1_1 gpc4000 (
      {stage0_40[453]},
      {stage1_40[271]}
   );
   gpc1_1 gpc4001 (
      {stage0_40[454]},
      {stage1_40[272]}
   );
   gpc1_1 gpc4002 (
      {stage0_40[455]},
      {stage1_40[273]}
   );
   gpc1_1 gpc4003 (
      {stage0_40[456]},
      {stage1_40[274]}
   );
   gpc1_1 gpc4004 (
      {stage0_40[457]},
      {stage1_40[275]}
   );
   gpc1_1 gpc4005 (
      {stage0_40[458]},
      {stage1_40[276]}
   );
   gpc1_1 gpc4006 (
      {stage0_40[459]},
      {stage1_40[277]}
   );
   gpc1_1 gpc4007 (
      {stage0_40[460]},
      {stage1_40[278]}
   );
   gpc1_1 gpc4008 (
      {stage0_40[461]},
      {stage1_40[279]}
   );
   gpc1_1 gpc4009 (
      {stage0_40[462]},
      {stage1_40[280]}
   );
   gpc1_1 gpc4010 (
      {stage0_40[463]},
      {stage1_40[281]}
   );
   gpc1_1 gpc4011 (
      {stage0_40[464]},
      {stage1_40[282]}
   );
   gpc1_1 gpc4012 (
      {stage0_40[465]},
      {stage1_40[283]}
   );
   gpc1_1 gpc4013 (
      {stage0_40[466]},
      {stage1_40[284]}
   );
   gpc1_1 gpc4014 (
      {stage0_40[467]},
      {stage1_40[285]}
   );
   gpc1_1 gpc4015 (
      {stage0_40[468]},
      {stage1_40[286]}
   );
   gpc1_1 gpc4016 (
      {stage0_40[469]},
      {stage1_40[287]}
   );
   gpc1_1 gpc4017 (
      {stage0_40[470]},
      {stage1_40[288]}
   );
   gpc1_1 gpc4018 (
      {stage0_40[471]},
      {stage1_40[289]}
   );
   gpc1_1 gpc4019 (
      {stage0_40[472]},
      {stage1_40[290]}
   );
   gpc1_1 gpc4020 (
      {stage0_40[473]},
      {stage1_40[291]}
   );
   gpc1_1 gpc4021 (
      {stage0_40[474]},
      {stage1_40[292]}
   );
   gpc1_1 gpc4022 (
      {stage0_40[475]},
      {stage1_40[293]}
   );
   gpc1_1 gpc4023 (
      {stage0_40[476]},
      {stage1_40[294]}
   );
   gpc1_1 gpc4024 (
      {stage0_40[477]},
      {stage1_40[295]}
   );
   gpc1_1 gpc4025 (
      {stage0_40[478]},
      {stage1_40[296]}
   );
   gpc1_1 gpc4026 (
      {stage0_40[479]},
      {stage1_40[297]}
   );
   gpc1_1 gpc4027 (
      {stage0_40[480]},
      {stage1_40[298]}
   );
   gpc1_1 gpc4028 (
      {stage0_40[481]},
      {stage1_40[299]}
   );
   gpc1_1 gpc4029 (
      {stage0_40[482]},
      {stage1_40[300]}
   );
   gpc1_1 gpc4030 (
      {stage0_40[483]},
      {stage1_40[301]}
   );
   gpc1_1 gpc4031 (
      {stage0_40[484]},
      {stage1_40[302]}
   );
   gpc1_1 gpc4032 (
      {stage0_40[485]},
      {stage1_40[303]}
   );
   gpc1_1 gpc4033 (
      {stage0_41[477]},
      {stage1_41[162]}
   );
   gpc1_1 gpc4034 (
      {stage0_41[478]},
      {stage1_41[163]}
   );
   gpc1_1 gpc4035 (
      {stage0_41[479]},
      {stage1_41[164]}
   );
   gpc1_1 gpc4036 (
      {stage0_41[480]},
      {stage1_41[165]}
   );
   gpc1_1 gpc4037 (
      {stage0_41[481]},
      {stage1_41[166]}
   );
   gpc1_1 gpc4038 (
      {stage0_41[482]},
      {stage1_41[167]}
   );
   gpc1_1 gpc4039 (
      {stage0_41[483]},
      {stage1_41[168]}
   );
   gpc1_1 gpc4040 (
      {stage0_41[484]},
      {stage1_41[169]}
   );
   gpc1_1 gpc4041 (
      {stage0_41[485]},
      {stage1_41[170]}
   );
   gpc1_1 gpc4042 (
      {stage0_42[483]},
      {stage1_42[171]}
   );
   gpc1_1 gpc4043 (
      {stage0_42[484]},
      {stage1_42[172]}
   );
   gpc1_1 gpc4044 (
      {stage0_42[485]},
      {stage1_42[173]}
   );
   gpc1_1 gpc4045 (
      {stage0_43[451]},
      {stage1_43[219]}
   );
   gpc1_1 gpc4046 (
      {stage0_43[452]},
      {stage1_43[220]}
   );
   gpc1_1 gpc4047 (
      {stage0_43[453]},
      {stage1_43[221]}
   );
   gpc1_1 gpc4048 (
      {stage0_43[454]},
      {stage1_43[222]}
   );
   gpc1_1 gpc4049 (
      {stage0_43[455]},
      {stage1_43[223]}
   );
   gpc1_1 gpc4050 (
      {stage0_43[456]},
      {stage1_43[224]}
   );
   gpc1_1 gpc4051 (
      {stage0_43[457]},
      {stage1_43[225]}
   );
   gpc1_1 gpc4052 (
      {stage0_43[458]},
      {stage1_43[226]}
   );
   gpc1_1 gpc4053 (
      {stage0_43[459]},
      {stage1_43[227]}
   );
   gpc1_1 gpc4054 (
      {stage0_43[460]},
      {stage1_43[228]}
   );
   gpc1_1 gpc4055 (
      {stage0_43[461]},
      {stage1_43[229]}
   );
   gpc1_1 gpc4056 (
      {stage0_43[462]},
      {stage1_43[230]}
   );
   gpc1_1 gpc4057 (
      {stage0_43[463]},
      {stage1_43[231]}
   );
   gpc1_1 gpc4058 (
      {stage0_43[464]},
      {stage1_43[232]}
   );
   gpc1_1 gpc4059 (
      {stage0_43[465]},
      {stage1_43[233]}
   );
   gpc1_1 gpc4060 (
      {stage0_43[466]},
      {stage1_43[234]}
   );
   gpc1_1 gpc4061 (
      {stage0_43[467]},
      {stage1_43[235]}
   );
   gpc1_1 gpc4062 (
      {stage0_43[468]},
      {stage1_43[236]}
   );
   gpc1_1 gpc4063 (
      {stage0_43[469]},
      {stage1_43[237]}
   );
   gpc1_1 gpc4064 (
      {stage0_43[470]},
      {stage1_43[238]}
   );
   gpc1_1 gpc4065 (
      {stage0_43[471]},
      {stage1_43[239]}
   );
   gpc1_1 gpc4066 (
      {stage0_43[472]},
      {stage1_43[240]}
   );
   gpc1_1 gpc4067 (
      {stage0_43[473]},
      {stage1_43[241]}
   );
   gpc1_1 gpc4068 (
      {stage0_43[474]},
      {stage1_43[242]}
   );
   gpc1_1 gpc4069 (
      {stage0_43[475]},
      {stage1_43[243]}
   );
   gpc1_1 gpc4070 (
      {stage0_43[476]},
      {stage1_43[244]}
   );
   gpc1_1 gpc4071 (
      {stage0_43[477]},
      {stage1_43[245]}
   );
   gpc1_1 gpc4072 (
      {stage0_43[478]},
      {stage1_43[246]}
   );
   gpc1_1 gpc4073 (
      {stage0_43[479]},
      {stage1_43[247]}
   );
   gpc1_1 gpc4074 (
      {stage0_43[480]},
      {stage1_43[248]}
   );
   gpc1_1 gpc4075 (
      {stage0_43[481]},
      {stage1_43[249]}
   );
   gpc1_1 gpc4076 (
      {stage0_43[482]},
      {stage1_43[250]}
   );
   gpc1_1 gpc4077 (
      {stage0_43[483]},
      {stage1_43[251]}
   );
   gpc1_1 gpc4078 (
      {stage0_43[484]},
      {stage1_43[252]}
   );
   gpc1_1 gpc4079 (
      {stage0_43[485]},
      {stage1_43[253]}
   );
   gpc1_1 gpc4080 (
      {stage0_44[424]},
      {stage1_44[194]}
   );
   gpc1_1 gpc4081 (
      {stage0_44[425]},
      {stage1_44[195]}
   );
   gpc1_1 gpc4082 (
      {stage0_44[426]},
      {stage1_44[196]}
   );
   gpc1_1 gpc4083 (
      {stage0_44[427]},
      {stage1_44[197]}
   );
   gpc1_1 gpc4084 (
      {stage0_44[428]},
      {stage1_44[198]}
   );
   gpc1_1 gpc4085 (
      {stage0_44[429]},
      {stage1_44[199]}
   );
   gpc1_1 gpc4086 (
      {stage0_44[430]},
      {stage1_44[200]}
   );
   gpc1_1 gpc4087 (
      {stage0_44[431]},
      {stage1_44[201]}
   );
   gpc1_1 gpc4088 (
      {stage0_44[432]},
      {stage1_44[202]}
   );
   gpc1_1 gpc4089 (
      {stage0_44[433]},
      {stage1_44[203]}
   );
   gpc1_1 gpc4090 (
      {stage0_44[434]},
      {stage1_44[204]}
   );
   gpc1_1 gpc4091 (
      {stage0_44[435]},
      {stage1_44[205]}
   );
   gpc1_1 gpc4092 (
      {stage0_44[436]},
      {stage1_44[206]}
   );
   gpc1_1 gpc4093 (
      {stage0_44[437]},
      {stage1_44[207]}
   );
   gpc1_1 gpc4094 (
      {stage0_44[438]},
      {stage1_44[208]}
   );
   gpc1_1 gpc4095 (
      {stage0_44[439]},
      {stage1_44[209]}
   );
   gpc1_1 gpc4096 (
      {stage0_44[440]},
      {stage1_44[210]}
   );
   gpc1_1 gpc4097 (
      {stage0_44[441]},
      {stage1_44[211]}
   );
   gpc1_1 gpc4098 (
      {stage0_44[442]},
      {stage1_44[212]}
   );
   gpc1_1 gpc4099 (
      {stage0_44[443]},
      {stage1_44[213]}
   );
   gpc1_1 gpc4100 (
      {stage0_44[444]},
      {stage1_44[214]}
   );
   gpc1_1 gpc4101 (
      {stage0_44[445]},
      {stage1_44[215]}
   );
   gpc1_1 gpc4102 (
      {stage0_44[446]},
      {stage1_44[216]}
   );
   gpc1_1 gpc4103 (
      {stage0_44[447]},
      {stage1_44[217]}
   );
   gpc1_1 gpc4104 (
      {stage0_44[448]},
      {stage1_44[218]}
   );
   gpc1_1 gpc4105 (
      {stage0_44[449]},
      {stage1_44[219]}
   );
   gpc1_1 gpc4106 (
      {stage0_44[450]},
      {stage1_44[220]}
   );
   gpc1_1 gpc4107 (
      {stage0_44[451]},
      {stage1_44[221]}
   );
   gpc1_1 gpc4108 (
      {stage0_44[452]},
      {stage1_44[222]}
   );
   gpc1_1 gpc4109 (
      {stage0_44[453]},
      {stage1_44[223]}
   );
   gpc1_1 gpc4110 (
      {stage0_44[454]},
      {stage1_44[224]}
   );
   gpc1_1 gpc4111 (
      {stage0_44[455]},
      {stage1_44[225]}
   );
   gpc1_1 gpc4112 (
      {stage0_44[456]},
      {stage1_44[226]}
   );
   gpc1_1 gpc4113 (
      {stage0_44[457]},
      {stage1_44[227]}
   );
   gpc1_1 gpc4114 (
      {stage0_44[458]},
      {stage1_44[228]}
   );
   gpc1_1 gpc4115 (
      {stage0_44[459]},
      {stage1_44[229]}
   );
   gpc1_1 gpc4116 (
      {stage0_44[460]},
      {stage1_44[230]}
   );
   gpc1_1 gpc4117 (
      {stage0_44[461]},
      {stage1_44[231]}
   );
   gpc1_1 gpc4118 (
      {stage0_44[462]},
      {stage1_44[232]}
   );
   gpc1_1 gpc4119 (
      {stage0_44[463]},
      {stage1_44[233]}
   );
   gpc1_1 gpc4120 (
      {stage0_44[464]},
      {stage1_44[234]}
   );
   gpc1_1 gpc4121 (
      {stage0_44[465]},
      {stage1_44[235]}
   );
   gpc1_1 gpc4122 (
      {stage0_44[466]},
      {stage1_44[236]}
   );
   gpc1_1 gpc4123 (
      {stage0_44[467]},
      {stage1_44[237]}
   );
   gpc1_1 gpc4124 (
      {stage0_44[468]},
      {stage1_44[238]}
   );
   gpc1_1 gpc4125 (
      {stage0_44[469]},
      {stage1_44[239]}
   );
   gpc1_1 gpc4126 (
      {stage0_44[470]},
      {stage1_44[240]}
   );
   gpc1_1 gpc4127 (
      {stage0_44[471]},
      {stage1_44[241]}
   );
   gpc1_1 gpc4128 (
      {stage0_44[472]},
      {stage1_44[242]}
   );
   gpc1_1 gpc4129 (
      {stage0_44[473]},
      {stage1_44[243]}
   );
   gpc1_1 gpc4130 (
      {stage0_44[474]},
      {stage1_44[244]}
   );
   gpc1_1 gpc4131 (
      {stage0_44[475]},
      {stage1_44[245]}
   );
   gpc1_1 gpc4132 (
      {stage0_44[476]},
      {stage1_44[246]}
   );
   gpc1_1 gpc4133 (
      {stage0_44[477]},
      {stage1_44[247]}
   );
   gpc1_1 gpc4134 (
      {stage0_44[478]},
      {stage1_44[248]}
   );
   gpc1_1 gpc4135 (
      {stage0_44[479]},
      {stage1_44[249]}
   );
   gpc1_1 gpc4136 (
      {stage0_44[480]},
      {stage1_44[250]}
   );
   gpc1_1 gpc4137 (
      {stage0_44[481]},
      {stage1_44[251]}
   );
   gpc1_1 gpc4138 (
      {stage0_44[482]},
      {stage1_44[252]}
   );
   gpc1_1 gpc4139 (
      {stage0_44[483]},
      {stage1_44[253]}
   );
   gpc1_1 gpc4140 (
      {stage0_44[484]},
      {stage1_44[254]}
   );
   gpc1_1 gpc4141 (
      {stage0_44[485]},
      {stage1_44[255]}
   );
   gpc1_1 gpc4142 (
      {stage0_45[433]},
      {stage1_45[159]}
   );
   gpc1_1 gpc4143 (
      {stage0_45[434]},
      {stage1_45[160]}
   );
   gpc1_1 gpc4144 (
      {stage0_45[435]},
      {stage1_45[161]}
   );
   gpc1_1 gpc4145 (
      {stage0_45[436]},
      {stage1_45[162]}
   );
   gpc1_1 gpc4146 (
      {stage0_45[437]},
      {stage1_45[163]}
   );
   gpc1_1 gpc4147 (
      {stage0_45[438]},
      {stage1_45[164]}
   );
   gpc1_1 gpc4148 (
      {stage0_45[439]},
      {stage1_45[165]}
   );
   gpc1_1 gpc4149 (
      {stage0_45[440]},
      {stage1_45[166]}
   );
   gpc1_1 gpc4150 (
      {stage0_45[441]},
      {stage1_45[167]}
   );
   gpc1_1 gpc4151 (
      {stage0_45[442]},
      {stage1_45[168]}
   );
   gpc1_1 gpc4152 (
      {stage0_45[443]},
      {stage1_45[169]}
   );
   gpc1_1 gpc4153 (
      {stage0_45[444]},
      {stage1_45[170]}
   );
   gpc1_1 gpc4154 (
      {stage0_45[445]},
      {stage1_45[171]}
   );
   gpc1_1 gpc4155 (
      {stage0_45[446]},
      {stage1_45[172]}
   );
   gpc1_1 gpc4156 (
      {stage0_45[447]},
      {stage1_45[173]}
   );
   gpc1_1 gpc4157 (
      {stage0_45[448]},
      {stage1_45[174]}
   );
   gpc1_1 gpc4158 (
      {stage0_45[449]},
      {stage1_45[175]}
   );
   gpc1_1 gpc4159 (
      {stage0_45[450]},
      {stage1_45[176]}
   );
   gpc1_1 gpc4160 (
      {stage0_45[451]},
      {stage1_45[177]}
   );
   gpc1_1 gpc4161 (
      {stage0_45[452]},
      {stage1_45[178]}
   );
   gpc1_1 gpc4162 (
      {stage0_45[453]},
      {stage1_45[179]}
   );
   gpc1_1 gpc4163 (
      {stage0_45[454]},
      {stage1_45[180]}
   );
   gpc1_1 gpc4164 (
      {stage0_45[455]},
      {stage1_45[181]}
   );
   gpc1_1 gpc4165 (
      {stage0_45[456]},
      {stage1_45[182]}
   );
   gpc1_1 gpc4166 (
      {stage0_45[457]},
      {stage1_45[183]}
   );
   gpc1_1 gpc4167 (
      {stage0_45[458]},
      {stage1_45[184]}
   );
   gpc1_1 gpc4168 (
      {stage0_45[459]},
      {stage1_45[185]}
   );
   gpc1_1 gpc4169 (
      {stage0_45[460]},
      {stage1_45[186]}
   );
   gpc1_1 gpc4170 (
      {stage0_45[461]},
      {stage1_45[187]}
   );
   gpc1_1 gpc4171 (
      {stage0_45[462]},
      {stage1_45[188]}
   );
   gpc1_1 gpc4172 (
      {stage0_45[463]},
      {stage1_45[189]}
   );
   gpc1_1 gpc4173 (
      {stage0_45[464]},
      {stage1_45[190]}
   );
   gpc1_1 gpc4174 (
      {stage0_45[465]},
      {stage1_45[191]}
   );
   gpc1_1 gpc4175 (
      {stage0_45[466]},
      {stage1_45[192]}
   );
   gpc1_1 gpc4176 (
      {stage0_45[467]},
      {stage1_45[193]}
   );
   gpc1_1 gpc4177 (
      {stage0_45[468]},
      {stage1_45[194]}
   );
   gpc1_1 gpc4178 (
      {stage0_45[469]},
      {stage1_45[195]}
   );
   gpc1_1 gpc4179 (
      {stage0_45[470]},
      {stage1_45[196]}
   );
   gpc1_1 gpc4180 (
      {stage0_45[471]},
      {stage1_45[197]}
   );
   gpc1_1 gpc4181 (
      {stage0_45[472]},
      {stage1_45[198]}
   );
   gpc1_1 gpc4182 (
      {stage0_45[473]},
      {stage1_45[199]}
   );
   gpc1_1 gpc4183 (
      {stage0_45[474]},
      {stage1_45[200]}
   );
   gpc1_1 gpc4184 (
      {stage0_45[475]},
      {stage1_45[201]}
   );
   gpc1_1 gpc4185 (
      {stage0_45[476]},
      {stage1_45[202]}
   );
   gpc1_1 gpc4186 (
      {stage0_45[477]},
      {stage1_45[203]}
   );
   gpc1_1 gpc4187 (
      {stage0_45[478]},
      {stage1_45[204]}
   );
   gpc1_1 gpc4188 (
      {stage0_45[479]},
      {stage1_45[205]}
   );
   gpc1_1 gpc4189 (
      {stage0_45[480]},
      {stage1_45[206]}
   );
   gpc1_1 gpc4190 (
      {stage0_45[481]},
      {stage1_45[207]}
   );
   gpc1_1 gpc4191 (
      {stage0_45[482]},
      {stage1_45[208]}
   );
   gpc1_1 gpc4192 (
      {stage0_45[483]},
      {stage1_45[209]}
   );
   gpc1_1 gpc4193 (
      {stage0_45[484]},
      {stage1_45[210]}
   );
   gpc1_1 gpc4194 (
      {stage0_45[485]},
      {stage1_45[211]}
   );
   gpc1_1 gpc4195 (
      {stage0_46[356]},
      {stage1_46[168]}
   );
   gpc1_1 gpc4196 (
      {stage0_46[357]},
      {stage1_46[169]}
   );
   gpc1_1 gpc4197 (
      {stage0_46[358]},
      {stage1_46[170]}
   );
   gpc1_1 gpc4198 (
      {stage0_46[359]},
      {stage1_46[171]}
   );
   gpc1_1 gpc4199 (
      {stage0_46[360]},
      {stage1_46[172]}
   );
   gpc1_1 gpc4200 (
      {stage0_46[361]},
      {stage1_46[173]}
   );
   gpc1_1 gpc4201 (
      {stage0_46[362]},
      {stage1_46[174]}
   );
   gpc1_1 gpc4202 (
      {stage0_46[363]},
      {stage1_46[175]}
   );
   gpc1_1 gpc4203 (
      {stage0_46[364]},
      {stage1_46[176]}
   );
   gpc1_1 gpc4204 (
      {stage0_46[365]},
      {stage1_46[177]}
   );
   gpc1_1 gpc4205 (
      {stage0_46[366]},
      {stage1_46[178]}
   );
   gpc1_1 gpc4206 (
      {stage0_46[367]},
      {stage1_46[179]}
   );
   gpc1_1 gpc4207 (
      {stage0_46[368]},
      {stage1_46[180]}
   );
   gpc1_1 gpc4208 (
      {stage0_46[369]},
      {stage1_46[181]}
   );
   gpc1_1 gpc4209 (
      {stage0_46[370]},
      {stage1_46[182]}
   );
   gpc1_1 gpc4210 (
      {stage0_46[371]},
      {stage1_46[183]}
   );
   gpc1_1 gpc4211 (
      {stage0_46[372]},
      {stage1_46[184]}
   );
   gpc1_1 gpc4212 (
      {stage0_46[373]},
      {stage1_46[185]}
   );
   gpc1_1 gpc4213 (
      {stage0_46[374]},
      {stage1_46[186]}
   );
   gpc1_1 gpc4214 (
      {stage0_46[375]},
      {stage1_46[187]}
   );
   gpc1_1 gpc4215 (
      {stage0_46[376]},
      {stage1_46[188]}
   );
   gpc1_1 gpc4216 (
      {stage0_46[377]},
      {stage1_46[189]}
   );
   gpc1_1 gpc4217 (
      {stage0_46[378]},
      {stage1_46[190]}
   );
   gpc1_1 gpc4218 (
      {stage0_46[379]},
      {stage1_46[191]}
   );
   gpc1_1 gpc4219 (
      {stage0_46[380]},
      {stage1_46[192]}
   );
   gpc1_1 gpc4220 (
      {stage0_46[381]},
      {stage1_46[193]}
   );
   gpc1_1 gpc4221 (
      {stage0_46[382]},
      {stage1_46[194]}
   );
   gpc1_1 gpc4222 (
      {stage0_46[383]},
      {stage1_46[195]}
   );
   gpc1_1 gpc4223 (
      {stage0_46[384]},
      {stage1_46[196]}
   );
   gpc1_1 gpc4224 (
      {stage0_46[385]},
      {stage1_46[197]}
   );
   gpc1_1 gpc4225 (
      {stage0_46[386]},
      {stage1_46[198]}
   );
   gpc1_1 gpc4226 (
      {stage0_46[387]},
      {stage1_46[199]}
   );
   gpc1_1 gpc4227 (
      {stage0_46[388]},
      {stage1_46[200]}
   );
   gpc1_1 gpc4228 (
      {stage0_46[389]},
      {stage1_46[201]}
   );
   gpc1_1 gpc4229 (
      {stage0_46[390]},
      {stage1_46[202]}
   );
   gpc1_1 gpc4230 (
      {stage0_46[391]},
      {stage1_46[203]}
   );
   gpc1_1 gpc4231 (
      {stage0_46[392]},
      {stage1_46[204]}
   );
   gpc1_1 gpc4232 (
      {stage0_46[393]},
      {stage1_46[205]}
   );
   gpc1_1 gpc4233 (
      {stage0_46[394]},
      {stage1_46[206]}
   );
   gpc1_1 gpc4234 (
      {stage0_46[395]},
      {stage1_46[207]}
   );
   gpc1_1 gpc4235 (
      {stage0_46[396]},
      {stage1_46[208]}
   );
   gpc1_1 gpc4236 (
      {stage0_46[397]},
      {stage1_46[209]}
   );
   gpc1_1 gpc4237 (
      {stage0_46[398]},
      {stage1_46[210]}
   );
   gpc1_1 gpc4238 (
      {stage0_46[399]},
      {stage1_46[211]}
   );
   gpc1_1 gpc4239 (
      {stage0_46[400]},
      {stage1_46[212]}
   );
   gpc1_1 gpc4240 (
      {stage0_46[401]},
      {stage1_46[213]}
   );
   gpc1_1 gpc4241 (
      {stage0_46[402]},
      {stage1_46[214]}
   );
   gpc1_1 gpc4242 (
      {stage0_46[403]},
      {stage1_46[215]}
   );
   gpc1_1 gpc4243 (
      {stage0_46[404]},
      {stage1_46[216]}
   );
   gpc1_1 gpc4244 (
      {stage0_46[405]},
      {stage1_46[217]}
   );
   gpc1_1 gpc4245 (
      {stage0_46[406]},
      {stage1_46[218]}
   );
   gpc1_1 gpc4246 (
      {stage0_46[407]},
      {stage1_46[219]}
   );
   gpc1_1 gpc4247 (
      {stage0_46[408]},
      {stage1_46[220]}
   );
   gpc1_1 gpc4248 (
      {stage0_46[409]},
      {stage1_46[221]}
   );
   gpc1_1 gpc4249 (
      {stage0_46[410]},
      {stage1_46[222]}
   );
   gpc1_1 gpc4250 (
      {stage0_46[411]},
      {stage1_46[223]}
   );
   gpc1_1 gpc4251 (
      {stage0_46[412]},
      {stage1_46[224]}
   );
   gpc1_1 gpc4252 (
      {stage0_46[413]},
      {stage1_46[225]}
   );
   gpc1_1 gpc4253 (
      {stage0_46[414]},
      {stage1_46[226]}
   );
   gpc1_1 gpc4254 (
      {stage0_46[415]},
      {stage1_46[227]}
   );
   gpc1_1 gpc4255 (
      {stage0_46[416]},
      {stage1_46[228]}
   );
   gpc1_1 gpc4256 (
      {stage0_46[417]},
      {stage1_46[229]}
   );
   gpc1_1 gpc4257 (
      {stage0_46[418]},
      {stage1_46[230]}
   );
   gpc1_1 gpc4258 (
      {stage0_46[419]},
      {stage1_46[231]}
   );
   gpc1_1 gpc4259 (
      {stage0_46[420]},
      {stage1_46[232]}
   );
   gpc1_1 gpc4260 (
      {stage0_46[421]},
      {stage1_46[233]}
   );
   gpc1_1 gpc4261 (
      {stage0_46[422]},
      {stage1_46[234]}
   );
   gpc1_1 gpc4262 (
      {stage0_46[423]},
      {stage1_46[235]}
   );
   gpc1_1 gpc4263 (
      {stage0_46[424]},
      {stage1_46[236]}
   );
   gpc1_1 gpc4264 (
      {stage0_46[425]},
      {stage1_46[237]}
   );
   gpc1_1 gpc4265 (
      {stage0_46[426]},
      {stage1_46[238]}
   );
   gpc1_1 gpc4266 (
      {stage0_46[427]},
      {stage1_46[239]}
   );
   gpc1_1 gpc4267 (
      {stage0_46[428]},
      {stage1_46[240]}
   );
   gpc1_1 gpc4268 (
      {stage0_46[429]},
      {stage1_46[241]}
   );
   gpc1_1 gpc4269 (
      {stage0_46[430]},
      {stage1_46[242]}
   );
   gpc1_1 gpc4270 (
      {stage0_46[431]},
      {stage1_46[243]}
   );
   gpc1_1 gpc4271 (
      {stage0_46[432]},
      {stage1_46[244]}
   );
   gpc1_1 gpc4272 (
      {stage0_46[433]},
      {stage1_46[245]}
   );
   gpc1_1 gpc4273 (
      {stage0_46[434]},
      {stage1_46[246]}
   );
   gpc1_1 gpc4274 (
      {stage0_46[435]},
      {stage1_46[247]}
   );
   gpc1_1 gpc4275 (
      {stage0_46[436]},
      {stage1_46[248]}
   );
   gpc1_1 gpc4276 (
      {stage0_46[437]},
      {stage1_46[249]}
   );
   gpc1_1 gpc4277 (
      {stage0_46[438]},
      {stage1_46[250]}
   );
   gpc1_1 gpc4278 (
      {stage0_46[439]},
      {stage1_46[251]}
   );
   gpc1_1 gpc4279 (
      {stage0_46[440]},
      {stage1_46[252]}
   );
   gpc1_1 gpc4280 (
      {stage0_46[441]},
      {stage1_46[253]}
   );
   gpc1_1 gpc4281 (
      {stage0_46[442]},
      {stage1_46[254]}
   );
   gpc1_1 gpc4282 (
      {stage0_46[443]},
      {stage1_46[255]}
   );
   gpc1_1 gpc4283 (
      {stage0_46[444]},
      {stage1_46[256]}
   );
   gpc1_1 gpc4284 (
      {stage0_46[445]},
      {stage1_46[257]}
   );
   gpc1_1 gpc4285 (
      {stage0_46[446]},
      {stage1_46[258]}
   );
   gpc1_1 gpc4286 (
      {stage0_46[447]},
      {stage1_46[259]}
   );
   gpc1_1 gpc4287 (
      {stage0_46[448]},
      {stage1_46[260]}
   );
   gpc1_1 gpc4288 (
      {stage0_46[449]},
      {stage1_46[261]}
   );
   gpc1_1 gpc4289 (
      {stage0_46[450]},
      {stage1_46[262]}
   );
   gpc1_1 gpc4290 (
      {stage0_46[451]},
      {stage1_46[263]}
   );
   gpc1_1 gpc4291 (
      {stage0_46[452]},
      {stage1_46[264]}
   );
   gpc1_1 gpc4292 (
      {stage0_46[453]},
      {stage1_46[265]}
   );
   gpc1_1 gpc4293 (
      {stage0_46[454]},
      {stage1_46[266]}
   );
   gpc1_1 gpc4294 (
      {stage0_46[455]},
      {stage1_46[267]}
   );
   gpc1_1 gpc4295 (
      {stage0_46[456]},
      {stage1_46[268]}
   );
   gpc1_1 gpc4296 (
      {stage0_46[457]},
      {stage1_46[269]}
   );
   gpc1_1 gpc4297 (
      {stage0_46[458]},
      {stage1_46[270]}
   );
   gpc1_1 gpc4298 (
      {stage0_46[459]},
      {stage1_46[271]}
   );
   gpc1_1 gpc4299 (
      {stage0_46[460]},
      {stage1_46[272]}
   );
   gpc1_1 gpc4300 (
      {stage0_46[461]},
      {stage1_46[273]}
   );
   gpc1_1 gpc4301 (
      {stage0_46[462]},
      {stage1_46[274]}
   );
   gpc1_1 gpc4302 (
      {stage0_46[463]},
      {stage1_46[275]}
   );
   gpc1_1 gpc4303 (
      {stage0_46[464]},
      {stage1_46[276]}
   );
   gpc1_1 gpc4304 (
      {stage0_46[465]},
      {stage1_46[277]}
   );
   gpc1_1 gpc4305 (
      {stage0_46[466]},
      {stage1_46[278]}
   );
   gpc1_1 gpc4306 (
      {stage0_46[467]},
      {stage1_46[279]}
   );
   gpc1_1 gpc4307 (
      {stage0_46[468]},
      {stage1_46[280]}
   );
   gpc1_1 gpc4308 (
      {stage0_46[469]},
      {stage1_46[281]}
   );
   gpc1_1 gpc4309 (
      {stage0_46[470]},
      {stage1_46[282]}
   );
   gpc1_1 gpc4310 (
      {stage0_46[471]},
      {stage1_46[283]}
   );
   gpc1_1 gpc4311 (
      {stage0_46[472]},
      {stage1_46[284]}
   );
   gpc1_1 gpc4312 (
      {stage0_46[473]},
      {stage1_46[285]}
   );
   gpc1_1 gpc4313 (
      {stage0_46[474]},
      {stage1_46[286]}
   );
   gpc1_1 gpc4314 (
      {stage0_46[475]},
      {stage1_46[287]}
   );
   gpc1_1 gpc4315 (
      {stage0_46[476]},
      {stage1_46[288]}
   );
   gpc1_1 gpc4316 (
      {stage0_46[477]},
      {stage1_46[289]}
   );
   gpc1_1 gpc4317 (
      {stage0_46[478]},
      {stage1_46[290]}
   );
   gpc1_1 gpc4318 (
      {stage0_46[479]},
      {stage1_46[291]}
   );
   gpc1_1 gpc4319 (
      {stage0_46[480]},
      {stage1_46[292]}
   );
   gpc1_1 gpc4320 (
      {stage0_46[481]},
      {stage1_46[293]}
   );
   gpc1_1 gpc4321 (
      {stage0_46[482]},
      {stage1_46[294]}
   );
   gpc1_1 gpc4322 (
      {stage0_46[483]},
      {stage1_46[295]}
   );
   gpc1_1 gpc4323 (
      {stage0_46[484]},
      {stage1_46[296]}
   );
   gpc1_1 gpc4324 (
      {stage0_46[485]},
      {stage1_46[297]}
   );
   gpc1_1 gpc4325 (
      {stage0_47[443]},
      {stage1_47[193]}
   );
   gpc1_1 gpc4326 (
      {stage0_47[444]},
      {stage1_47[194]}
   );
   gpc1_1 gpc4327 (
      {stage0_47[445]},
      {stage1_47[195]}
   );
   gpc1_1 gpc4328 (
      {stage0_47[446]},
      {stage1_47[196]}
   );
   gpc1_1 gpc4329 (
      {stage0_47[447]},
      {stage1_47[197]}
   );
   gpc1_1 gpc4330 (
      {stage0_47[448]},
      {stage1_47[198]}
   );
   gpc1_1 gpc4331 (
      {stage0_47[449]},
      {stage1_47[199]}
   );
   gpc1_1 gpc4332 (
      {stage0_47[450]},
      {stage1_47[200]}
   );
   gpc1_1 gpc4333 (
      {stage0_47[451]},
      {stage1_47[201]}
   );
   gpc1_1 gpc4334 (
      {stage0_47[452]},
      {stage1_47[202]}
   );
   gpc1_1 gpc4335 (
      {stage0_47[453]},
      {stage1_47[203]}
   );
   gpc1_1 gpc4336 (
      {stage0_47[454]},
      {stage1_47[204]}
   );
   gpc1_1 gpc4337 (
      {stage0_47[455]},
      {stage1_47[205]}
   );
   gpc1_1 gpc4338 (
      {stage0_47[456]},
      {stage1_47[206]}
   );
   gpc1_1 gpc4339 (
      {stage0_47[457]},
      {stage1_47[207]}
   );
   gpc1_1 gpc4340 (
      {stage0_47[458]},
      {stage1_47[208]}
   );
   gpc1_1 gpc4341 (
      {stage0_47[459]},
      {stage1_47[209]}
   );
   gpc1_1 gpc4342 (
      {stage0_47[460]},
      {stage1_47[210]}
   );
   gpc1_1 gpc4343 (
      {stage0_47[461]},
      {stage1_47[211]}
   );
   gpc1_1 gpc4344 (
      {stage0_47[462]},
      {stage1_47[212]}
   );
   gpc1_1 gpc4345 (
      {stage0_47[463]},
      {stage1_47[213]}
   );
   gpc1_1 gpc4346 (
      {stage0_47[464]},
      {stage1_47[214]}
   );
   gpc1_1 gpc4347 (
      {stage0_47[465]},
      {stage1_47[215]}
   );
   gpc1_1 gpc4348 (
      {stage0_47[466]},
      {stage1_47[216]}
   );
   gpc1_1 gpc4349 (
      {stage0_47[467]},
      {stage1_47[217]}
   );
   gpc1_1 gpc4350 (
      {stage0_47[468]},
      {stage1_47[218]}
   );
   gpc1_1 gpc4351 (
      {stage0_47[469]},
      {stage1_47[219]}
   );
   gpc1_1 gpc4352 (
      {stage0_47[470]},
      {stage1_47[220]}
   );
   gpc1_1 gpc4353 (
      {stage0_47[471]},
      {stage1_47[221]}
   );
   gpc1_1 gpc4354 (
      {stage0_47[472]},
      {stage1_47[222]}
   );
   gpc1_1 gpc4355 (
      {stage0_47[473]},
      {stage1_47[223]}
   );
   gpc1_1 gpc4356 (
      {stage0_47[474]},
      {stage1_47[224]}
   );
   gpc1_1 gpc4357 (
      {stage0_47[475]},
      {stage1_47[225]}
   );
   gpc1_1 gpc4358 (
      {stage0_47[476]},
      {stage1_47[226]}
   );
   gpc1_1 gpc4359 (
      {stage0_47[477]},
      {stage1_47[227]}
   );
   gpc1_1 gpc4360 (
      {stage0_47[478]},
      {stage1_47[228]}
   );
   gpc1_1 gpc4361 (
      {stage0_47[479]},
      {stage1_47[229]}
   );
   gpc1_1 gpc4362 (
      {stage0_47[480]},
      {stage1_47[230]}
   );
   gpc1_1 gpc4363 (
      {stage0_47[481]},
      {stage1_47[231]}
   );
   gpc1_1 gpc4364 (
      {stage0_47[482]},
      {stage1_47[232]}
   );
   gpc1_1 gpc4365 (
      {stage0_47[483]},
      {stage1_47[233]}
   );
   gpc1_1 gpc4366 (
      {stage0_47[484]},
      {stage1_47[234]}
   );
   gpc1_1 gpc4367 (
      {stage0_47[485]},
      {stage1_47[235]}
   );
   gpc1_1 gpc4368 (
      {stage0_48[478]},
      {stage1_48[190]}
   );
   gpc1_1 gpc4369 (
      {stage0_48[479]},
      {stage1_48[191]}
   );
   gpc1_1 gpc4370 (
      {stage0_48[480]},
      {stage1_48[192]}
   );
   gpc1_1 gpc4371 (
      {stage0_48[481]},
      {stage1_48[193]}
   );
   gpc1_1 gpc4372 (
      {stage0_48[482]},
      {stage1_48[194]}
   );
   gpc1_1 gpc4373 (
      {stage0_48[483]},
      {stage1_48[195]}
   );
   gpc1_1 gpc4374 (
      {stage0_48[484]},
      {stage1_48[196]}
   );
   gpc1_1 gpc4375 (
      {stage0_48[485]},
      {stage1_48[197]}
   );
   gpc1_1 gpc4376 (
      {stage0_50[481]},
      {stage1_50[185]}
   );
   gpc1_1 gpc4377 (
      {stage0_50[482]},
      {stage1_50[186]}
   );
   gpc1_1 gpc4378 (
      {stage0_50[483]},
      {stage1_50[187]}
   );
   gpc1_1 gpc4379 (
      {stage0_50[484]},
      {stage1_50[188]}
   );
   gpc1_1 gpc4380 (
      {stage0_50[485]},
      {stage1_50[189]}
   );
   gpc1_1 gpc4381 (
      {stage0_51[435]},
      {stage1_51[224]}
   );
   gpc1_1 gpc4382 (
      {stage0_51[436]},
      {stage1_51[225]}
   );
   gpc1_1 gpc4383 (
      {stage0_51[437]},
      {stage1_51[226]}
   );
   gpc1_1 gpc4384 (
      {stage0_51[438]},
      {stage1_51[227]}
   );
   gpc1_1 gpc4385 (
      {stage0_51[439]},
      {stage1_51[228]}
   );
   gpc1_1 gpc4386 (
      {stage0_51[440]},
      {stage1_51[229]}
   );
   gpc1_1 gpc4387 (
      {stage0_51[441]},
      {stage1_51[230]}
   );
   gpc1_1 gpc4388 (
      {stage0_51[442]},
      {stage1_51[231]}
   );
   gpc1_1 gpc4389 (
      {stage0_51[443]},
      {stage1_51[232]}
   );
   gpc1_1 gpc4390 (
      {stage0_51[444]},
      {stage1_51[233]}
   );
   gpc1_1 gpc4391 (
      {stage0_51[445]},
      {stage1_51[234]}
   );
   gpc1_1 gpc4392 (
      {stage0_51[446]},
      {stage1_51[235]}
   );
   gpc1_1 gpc4393 (
      {stage0_51[447]},
      {stage1_51[236]}
   );
   gpc1_1 gpc4394 (
      {stage0_51[448]},
      {stage1_51[237]}
   );
   gpc1_1 gpc4395 (
      {stage0_51[449]},
      {stage1_51[238]}
   );
   gpc1_1 gpc4396 (
      {stage0_51[450]},
      {stage1_51[239]}
   );
   gpc1_1 gpc4397 (
      {stage0_51[451]},
      {stage1_51[240]}
   );
   gpc1_1 gpc4398 (
      {stage0_51[452]},
      {stage1_51[241]}
   );
   gpc1_1 gpc4399 (
      {stage0_51[453]},
      {stage1_51[242]}
   );
   gpc1_1 gpc4400 (
      {stage0_51[454]},
      {stage1_51[243]}
   );
   gpc1_1 gpc4401 (
      {stage0_51[455]},
      {stage1_51[244]}
   );
   gpc1_1 gpc4402 (
      {stage0_51[456]},
      {stage1_51[245]}
   );
   gpc1_1 gpc4403 (
      {stage0_51[457]},
      {stage1_51[246]}
   );
   gpc1_1 gpc4404 (
      {stage0_51[458]},
      {stage1_51[247]}
   );
   gpc1_1 gpc4405 (
      {stage0_51[459]},
      {stage1_51[248]}
   );
   gpc1_1 gpc4406 (
      {stage0_51[460]},
      {stage1_51[249]}
   );
   gpc1_1 gpc4407 (
      {stage0_51[461]},
      {stage1_51[250]}
   );
   gpc1_1 gpc4408 (
      {stage0_51[462]},
      {stage1_51[251]}
   );
   gpc1_1 gpc4409 (
      {stage0_51[463]},
      {stage1_51[252]}
   );
   gpc1_1 gpc4410 (
      {stage0_51[464]},
      {stage1_51[253]}
   );
   gpc1_1 gpc4411 (
      {stage0_51[465]},
      {stage1_51[254]}
   );
   gpc1_1 gpc4412 (
      {stage0_51[466]},
      {stage1_51[255]}
   );
   gpc1_1 gpc4413 (
      {stage0_51[467]},
      {stage1_51[256]}
   );
   gpc1_1 gpc4414 (
      {stage0_51[468]},
      {stage1_51[257]}
   );
   gpc1_1 gpc4415 (
      {stage0_51[469]},
      {stage1_51[258]}
   );
   gpc1_1 gpc4416 (
      {stage0_51[470]},
      {stage1_51[259]}
   );
   gpc1_1 gpc4417 (
      {stage0_51[471]},
      {stage1_51[260]}
   );
   gpc1_1 gpc4418 (
      {stage0_51[472]},
      {stage1_51[261]}
   );
   gpc1_1 gpc4419 (
      {stage0_51[473]},
      {stage1_51[262]}
   );
   gpc1_1 gpc4420 (
      {stage0_51[474]},
      {stage1_51[263]}
   );
   gpc1_1 gpc4421 (
      {stage0_51[475]},
      {stage1_51[264]}
   );
   gpc1_1 gpc4422 (
      {stage0_51[476]},
      {stage1_51[265]}
   );
   gpc1_1 gpc4423 (
      {stage0_51[477]},
      {stage1_51[266]}
   );
   gpc1_1 gpc4424 (
      {stage0_51[478]},
      {stage1_51[267]}
   );
   gpc1_1 gpc4425 (
      {stage0_51[479]},
      {stage1_51[268]}
   );
   gpc1_1 gpc4426 (
      {stage0_51[480]},
      {stage1_51[269]}
   );
   gpc1_1 gpc4427 (
      {stage0_51[481]},
      {stage1_51[270]}
   );
   gpc1_1 gpc4428 (
      {stage0_51[482]},
      {stage1_51[271]}
   );
   gpc1_1 gpc4429 (
      {stage0_51[483]},
      {stage1_51[272]}
   );
   gpc1_1 gpc4430 (
      {stage0_51[484]},
      {stage1_51[273]}
   );
   gpc1_1 gpc4431 (
      {stage0_51[485]},
      {stage1_51[274]}
   );
   gpc1_1 gpc4432 (
      {stage0_54[453]},
      {stage1_54[198]}
   );
   gpc1_1 gpc4433 (
      {stage0_54[454]},
      {stage1_54[199]}
   );
   gpc1_1 gpc4434 (
      {stage0_54[455]},
      {stage1_54[200]}
   );
   gpc1_1 gpc4435 (
      {stage0_54[456]},
      {stage1_54[201]}
   );
   gpc1_1 gpc4436 (
      {stage0_54[457]},
      {stage1_54[202]}
   );
   gpc1_1 gpc4437 (
      {stage0_54[458]},
      {stage1_54[203]}
   );
   gpc1_1 gpc4438 (
      {stage0_54[459]},
      {stage1_54[204]}
   );
   gpc1_1 gpc4439 (
      {stage0_54[460]},
      {stage1_54[205]}
   );
   gpc1_1 gpc4440 (
      {stage0_54[461]},
      {stage1_54[206]}
   );
   gpc1_1 gpc4441 (
      {stage0_54[462]},
      {stage1_54[207]}
   );
   gpc1_1 gpc4442 (
      {stage0_54[463]},
      {stage1_54[208]}
   );
   gpc1_1 gpc4443 (
      {stage0_54[464]},
      {stage1_54[209]}
   );
   gpc1_1 gpc4444 (
      {stage0_54[465]},
      {stage1_54[210]}
   );
   gpc1_1 gpc4445 (
      {stage0_54[466]},
      {stage1_54[211]}
   );
   gpc1_1 gpc4446 (
      {stage0_54[467]},
      {stage1_54[212]}
   );
   gpc1_1 gpc4447 (
      {stage0_54[468]},
      {stage1_54[213]}
   );
   gpc1_1 gpc4448 (
      {stage0_54[469]},
      {stage1_54[214]}
   );
   gpc1_1 gpc4449 (
      {stage0_54[470]},
      {stage1_54[215]}
   );
   gpc1_1 gpc4450 (
      {stage0_54[471]},
      {stage1_54[216]}
   );
   gpc1_1 gpc4451 (
      {stage0_54[472]},
      {stage1_54[217]}
   );
   gpc1_1 gpc4452 (
      {stage0_54[473]},
      {stage1_54[218]}
   );
   gpc1_1 gpc4453 (
      {stage0_54[474]},
      {stage1_54[219]}
   );
   gpc1_1 gpc4454 (
      {stage0_54[475]},
      {stage1_54[220]}
   );
   gpc1_1 gpc4455 (
      {stage0_54[476]},
      {stage1_54[221]}
   );
   gpc1_1 gpc4456 (
      {stage0_54[477]},
      {stage1_54[222]}
   );
   gpc1_1 gpc4457 (
      {stage0_54[478]},
      {stage1_54[223]}
   );
   gpc1_1 gpc4458 (
      {stage0_54[479]},
      {stage1_54[224]}
   );
   gpc1_1 gpc4459 (
      {stage0_54[480]},
      {stage1_54[225]}
   );
   gpc1_1 gpc4460 (
      {stage0_54[481]},
      {stage1_54[226]}
   );
   gpc1_1 gpc4461 (
      {stage0_54[482]},
      {stage1_54[227]}
   );
   gpc1_1 gpc4462 (
      {stage0_54[483]},
      {stage1_54[228]}
   );
   gpc1_1 gpc4463 (
      {stage0_54[484]},
      {stage1_54[229]}
   );
   gpc1_1 gpc4464 (
      {stage0_54[485]},
      {stage1_54[230]}
   );
   gpc1_1 gpc4465 (
      {stage0_55[425]},
      {stage1_55[206]}
   );
   gpc1_1 gpc4466 (
      {stage0_55[426]},
      {stage1_55[207]}
   );
   gpc1_1 gpc4467 (
      {stage0_55[427]},
      {stage1_55[208]}
   );
   gpc1_1 gpc4468 (
      {stage0_55[428]},
      {stage1_55[209]}
   );
   gpc1_1 gpc4469 (
      {stage0_55[429]},
      {stage1_55[210]}
   );
   gpc1_1 gpc4470 (
      {stage0_55[430]},
      {stage1_55[211]}
   );
   gpc1_1 gpc4471 (
      {stage0_55[431]},
      {stage1_55[212]}
   );
   gpc1_1 gpc4472 (
      {stage0_55[432]},
      {stage1_55[213]}
   );
   gpc1_1 gpc4473 (
      {stage0_55[433]},
      {stage1_55[214]}
   );
   gpc1_1 gpc4474 (
      {stage0_55[434]},
      {stage1_55[215]}
   );
   gpc1_1 gpc4475 (
      {stage0_55[435]},
      {stage1_55[216]}
   );
   gpc1_1 gpc4476 (
      {stage0_55[436]},
      {stage1_55[217]}
   );
   gpc1_1 gpc4477 (
      {stage0_55[437]},
      {stage1_55[218]}
   );
   gpc1_1 gpc4478 (
      {stage0_55[438]},
      {stage1_55[219]}
   );
   gpc1_1 gpc4479 (
      {stage0_55[439]},
      {stage1_55[220]}
   );
   gpc1_1 gpc4480 (
      {stage0_55[440]},
      {stage1_55[221]}
   );
   gpc1_1 gpc4481 (
      {stage0_55[441]},
      {stage1_55[222]}
   );
   gpc1_1 gpc4482 (
      {stage0_55[442]},
      {stage1_55[223]}
   );
   gpc1_1 gpc4483 (
      {stage0_55[443]},
      {stage1_55[224]}
   );
   gpc1_1 gpc4484 (
      {stage0_55[444]},
      {stage1_55[225]}
   );
   gpc1_1 gpc4485 (
      {stage0_55[445]},
      {stage1_55[226]}
   );
   gpc1_1 gpc4486 (
      {stage0_55[446]},
      {stage1_55[227]}
   );
   gpc1_1 gpc4487 (
      {stage0_55[447]},
      {stage1_55[228]}
   );
   gpc1_1 gpc4488 (
      {stage0_55[448]},
      {stage1_55[229]}
   );
   gpc1_1 gpc4489 (
      {stage0_55[449]},
      {stage1_55[230]}
   );
   gpc1_1 gpc4490 (
      {stage0_55[450]},
      {stage1_55[231]}
   );
   gpc1_1 gpc4491 (
      {stage0_55[451]},
      {stage1_55[232]}
   );
   gpc1_1 gpc4492 (
      {stage0_55[452]},
      {stage1_55[233]}
   );
   gpc1_1 gpc4493 (
      {stage0_55[453]},
      {stage1_55[234]}
   );
   gpc1_1 gpc4494 (
      {stage0_55[454]},
      {stage1_55[235]}
   );
   gpc1_1 gpc4495 (
      {stage0_55[455]},
      {stage1_55[236]}
   );
   gpc1_1 gpc4496 (
      {stage0_55[456]},
      {stage1_55[237]}
   );
   gpc1_1 gpc4497 (
      {stage0_55[457]},
      {stage1_55[238]}
   );
   gpc1_1 gpc4498 (
      {stage0_55[458]},
      {stage1_55[239]}
   );
   gpc1_1 gpc4499 (
      {stage0_55[459]},
      {stage1_55[240]}
   );
   gpc1_1 gpc4500 (
      {stage0_55[460]},
      {stage1_55[241]}
   );
   gpc1_1 gpc4501 (
      {stage0_55[461]},
      {stage1_55[242]}
   );
   gpc1_1 gpc4502 (
      {stage0_55[462]},
      {stage1_55[243]}
   );
   gpc1_1 gpc4503 (
      {stage0_55[463]},
      {stage1_55[244]}
   );
   gpc1_1 gpc4504 (
      {stage0_55[464]},
      {stage1_55[245]}
   );
   gpc1_1 gpc4505 (
      {stage0_55[465]},
      {stage1_55[246]}
   );
   gpc1_1 gpc4506 (
      {stage0_55[466]},
      {stage1_55[247]}
   );
   gpc1_1 gpc4507 (
      {stage0_55[467]},
      {stage1_55[248]}
   );
   gpc1_1 gpc4508 (
      {stage0_55[468]},
      {stage1_55[249]}
   );
   gpc1_1 gpc4509 (
      {stage0_55[469]},
      {stage1_55[250]}
   );
   gpc1_1 gpc4510 (
      {stage0_55[470]},
      {stage1_55[251]}
   );
   gpc1_1 gpc4511 (
      {stage0_55[471]},
      {stage1_55[252]}
   );
   gpc1_1 gpc4512 (
      {stage0_55[472]},
      {stage1_55[253]}
   );
   gpc1_1 gpc4513 (
      {stage0_55[473]},
      {stage1_55[254]}
   );
   gpc1_1 gpc4514 (
      {stage0_55[474]},
      {stage1_55[255]}
   );
   gpc1_1 gpc4515 (
      {stage0_55[475]},
      {stage1_55[256]}
   );
   gpc1_1 gpc4516 (
      {stage0_55[476]},
      {stage1_55[257]}
   );
   gpc1_1 gpc4517 (
      {stage0_55[477]},
      {stage1_55[258]}
   );
   gpc1_1 gpc4518 (
      {stage0_55[478]},
      {stage1_55[259]}
   );
   gpc1_1 gpc4519 (
      {stage0_55[479]},
      {stage1_55[260]}
   );
   gpc1_1 gpc4520 (
      {stage0_55[480]},
      {stage1_55[261]}
   );
   gpc1_1 gpc4521 (
      {stage0_55[481]},
      {stage1_55[262]}
   );
   gpc1_1 gpc4522 (
      {stage0_55[482]},
      {stage1_55[263]}
   );
   gpc1_1 gpc4523 (
      {stage0_55[483]},
      {stage1_55[264]}
   );
   gpc1_1 gpc4524 (
      {stage0_55[484]},
      {stage1_55[265]}
   );
   gpc1_1 gpc4525 (
      {stage0_55[485]},
      {stage1_55[266]}
   );
   gpc1_1 gpc4526 (
      {stage0_58[460]},
      {stage1_58[194]}
   );
   gpc1_1 gpc4527 (
      {stage0_58[461]},
      {stage1_58[195]}
   );
   gpc1_1 gpc4528 (
      {stage0_58[462]},
      {stage1_58[196]}
   );
   gpc1_1 gpc4529 (
      {stage0_58[463]},
      {stage1_58[197]}
   );
   gpc1_1 gpc4530 (
      {stage0_58[464]},
      {stage1_58[198]}
   );
   gpc1_1 gpc4531 (
      {stage0_58[465]},
      {stage1_58[199]}
   );
   gpc1_1 gpc4532 (
      {stage0_58[466]},
      {stage1_58[200]}
   );
   gpc1_1 gpc4533 (
      {stage0_58[467]},
      {stage1_58[201]}
   );
   gpc1_1 gpc4534 (
      {stage0_58[468]},
      {stage1_58[202]}
   );
   gpc1_1 gpc4535 (
      {stage0_58[469]},
      {stage1_58[203]}
   );
   gpc1_1 gpc4536 (
      {stage0_58[470]},
      {stage1_58[204]}
   );
   gpc1_1 gpc4537 (
      {stage0_58[471]},
      {stage1_58[205]}
   );
   gpc1_1 gpc4538 (
      {stage0_58[472]},
      {stage1_58[206]}
   );
   gpc1_1 gpc4539 (
      {stage0_58[473]},
      {stage1_58[207]}
   );
   gpc1_1 gpc4540 (
      {stage0_58[474]},
      {stage1_58[208]}
   );
   gpc1_1 gpc4541 (
      {stage0_58[475]},
      {stage1_58[209]}
   );
   gpc1_1 gpc4542 (
      {stage0_58[476]},
      {stage1_58[210]}
   );
   gpc1_1 gpc4543 (
      {stage0_58[477]},
      {stage1_58[211]}
   );
   gpc1_1 gpc4544 (
      {stage0_58[478]},
      {stage1_58[212]}
   );
   gpc1_1 gpc4545 (
      {stage0_58[479]},
      {stage1_58[213]}
   );
   gpc1_1 gpc4546 (
      {stage0_58[480]},
      {stage1_58[214]}
   );
   gpc1_1 gpc4547 (
      {stage0_58[481]},
      {stage1_58[215]}
   );
   gpc1_1 gpc4548 (
      {stage0_58[482]},
      {stage1_58[216]}
   );
   gpc1_1 gpc4549 (
      {stage0_58[483]},
      {stage1_58[217]}
   );
   gpc1_1 gpc4550 (
      {stage0_58[484]},
      {stage1_58[218]}
   );
   gpc1_1 gpc4551 (
      {stage0_58[485]},
      {stage1_58[219]}
   );
   gpc1_1 gpc4552 (
      {stage0_59[469]},
      {stage1_59[189]}
   );
   gpc1_1 gpc4553 (
      {stage0_59[470]},
      {stage1_59[190]}
   );
   gpc1_1 gpc4554 (
      {stage0_59[471]},
      {stage1_59[191]}
   );
   gpc1_1 gpc4555 (
      {stage0_59[472]},
      {stage1_59[192]}
   );
   gpc1_1 gpc4556 (
      {stage0_59[473]},
      {stage1_59[193]}
   );
   gpc1_1 gpc4557 (
      {stage0_59[474]},
      {stage1_59[194]}
   );
   gpc1_1 gpc4558 (
      {stage0_59[475]},
      {stage1_59[195]}
   );
   gpc1_1 gpc4559 (
      {stage0_59[476]},
      {stage1_59[196]}
   );
   gpc1_1 gpc4560 (
      {stage0_59[477]},
      {stage1_59[197]}
   );
   gpc1_1 gpc4561 (
      {stage0_59[478]},
      {stage1_59[198]}
   );
   gpc1_1 gpc4562 (
      {stage0_59[479]},
      {stage1_59[199]}
   );
   gpc1_1 gpc4563 (
      {stage0_59[480]},
      {stage1_59[200]}
   );
   gpc1_1 gpc4564 (
      {stage0_59[481]},
      {stage1_59[201]}
   );
   gpc1_1 gpc4565 (
      {stage0_59[482]},
      {stage1_59[202]}
   );
   gpc1_1 gpc4566 (
      {stage0_59[483]},
      {stage1_59[203]}
   );
   gpc1_1 gpc4567 (
      {stage0_59[484]},
      {stage1_59[204]}
   );
   gpc1_1 gpc4568 (
      {stage0_59[485]},
      {stage1_59[205]}
   );
   gpc1_1 gpc4569 (
      {stage0_62[474]},
      {stage1_62[181]}
   );
   gpc1_1 gpc4570 (
      {stage0_62[475]},
      {stage1_62[182]}
   );
   gpc1_1 gpc4571 (
      {stage0_62[476]},
      {stage1_62[183]}
   );
   gpc1_1 gpc4572 (
      {stage0_62[477]},
      {stage1_62[184]}
   );
   gpc1_1 gpc4573 (
      {stage0_62[478]},
      {stage1_62[185]}
   );
   gpc1_1 gpc4574 (
      {stage0_62[479]},
      {stage1_62[186]}
   );
   gpc1_1 gpc4575 (
      {stage0_62[480]},
      {stage1_62[187]}
   );
   gpc1_1 gpc4576 (
      {stage0_62[481]},
      {stage1_62[188]}
   );
   gpc1_1 gpc4577 (
      {stage0_62[482]},
      {stage1_62[189]}
   );
   gpc1_1 gpc4578 (
      {stage0_62[483]},
      {stage1_62[190]}
   );
   gpc1_1 gpc4579 (
      {stage0_62[484]},
      {stage1_62[191]}
   );
   gpc1_1 gpc4580 (
      {stage0_62[485]},
      {stage1_62[192]}
   );
   gpc1_1 gpc4581 (
      {stage0_63[324]},
      {stage1_63[146]}
   );
   gpc1_1 gpc4582 (
      {stage0_63[325]},
      {stage1_63[147]}
   );
   gpc1_1 gpc4583 (
      {stage0_63[326]},
      {stage1_63[148]}
   );
   gpc1_1 gpc4584 (
      {stage0_63[327]},
      {stage1_63[149]}
   );
   gpc1_1 gpc4585 (
      {stage0_63[328]},
      {stage1_63[150]}
   );
   gpc1_1 gpc4586 (
      {stage0_63[329]},
      {stage1_63[151]}
   );
   gpc1_1 gpc4587 (
      {stage0_63[330]},
      {stage1_63[152]}
   );
   gpc1_1 gpc4588 (
      {stage0_63[331]},
      {stage1_63[153]}
   );
   gpc1_1 gpc4589 (
      {stage0_63[332]},
      {stage1_63[154]}
   );
   gpc1_1 gpc4590 (
      {stage0_63[333]},
      {stage1_63[155]}
   );
   gpc1_1 gpc4591 (
      {stage0_63[334]},
      {stage1_63[156]}
   );
   gpc1_1 gpc4592 (
      {stage0_63[335]},
      {stage1_63[157]}
   );
   gpc1_1 gpc4593 (
      {stage0_63[336]},
      {stage1_63[158]}
   );
   gpc1_1 gpc4594 (
      {stage0_63[337]},
      {stage1_63[159]}
   );
   gpc1_1 gpc4595 (
      {stage0_63[338]},
      {stage1_63[160]}
   );
   gpc1_1 gpc4596 (
      {stage0_63[339]},
      {stage1_63[161]}
   );
   gpc1_1 gpc4597 (
      {stage0_63[340]},
      {stage1_63[162]}
   );
   gpc1_1 gpc4598 (
      {stage0_63[341]},
      {stage1_63[163]}
   );
   gpc1_1 gpc4599 (
      {stage0_63[342]},
      {stage1_63[164]}
   );
   gpc1_1 gpc4600 (
      {stage0_63[343]},
      {stage1_63[165]}
   );
   gpc1_1 gpc4601 (
      {stage0_63[344]},
      {stage1_63[166]}
   );
   gpc1_1 gpc4602 (
      {stage0_63[345]},
      {stage1_63[167]}
   );
   gpc1_1 gpc4603 (
      {stage0_63[346]},
      {stage1_63[168]}
   );
   gpc1_1 gpc4604 (
      {stage0_63[347]},
      {stage1_63[169]}
   );
   gpc1_1 gpc4605 (
      {stage0_63[348]},
      {stage1_63[170]}
   );
   gpc1_1 gpc4606 (
      {stage0_63[349]},
      {stage1_63[171]}
   );
   gpc1_1 gpc4607 (
      {stage0_63[350]},
      {stage1_63[172]}
   );
   gpc1_1 gpc4608 (
      {stage0_63[351]},
      {stage1_63[173]}
   );
   gpc1_1 gpc4609 (
      {stage0_63[352]},
      {stage1_63[174]}
   );
   gpc1_1 gpc4610 (
      {stage0_63[353]},
      {stage1_63[175]}
   );
   gpc1_1 gpc4611 (
      {stage0_63[354]},
      {stage1_63[176]}
   );
   gpc1_1 gpc4612 (
      {stage0_63[355]},
      {stage1_63[177]}
   );
   gpc1_1 gpc4613 (
      {stage0_63[356]},
      {stage1_63[178]}
   );
   gpc1_1 gpc4614 (
      {stage0_63[357]},
      {stage1_63[179]}
   );
   gpc1_1 gpc4615 (
      {stage0_63[358]},
      {stage1_63[180]}
   );
   gpc1_1 gpc4616 (
      {stage0_63[359]},
      {stage1_63[181]}
   );
   gpc1_1 gpc4617 (
      {stage0_63[360]},
      {stage1_63[182]}
   );
   gpc1_1 gpc4618 (
      {stage0_63[361]},
      {stage1_63[183]}
   );
   gpc1_1 gpc4619 (
      {stage0_63[362]},
      {stage1_63[184]}
   );
   gpc1_1 gpc4620 (
      {stage0_63[363]},
      {stage1_63[185]}
   );
   gpc1_1 gpc4621 (
      {stage0_63[364]},
      {stage1_63[186]}
   );
   gpc1_1 gpc4622 (
      {stage0_63[365]},
      {stage1_63[187]}
   );
   gpc1_1 gpc4623 (
      {stage0_63[366]},
      {stage1_63[188]}
   );
   gpc1_1 gpc4624 (
      {stage0_63[367]},
      {stage1_63[189]}
   );
   gpc1_1 gpc4625 (
      {stage0_63[368]},
      {stage1_63[190]}
   );
   gpc1_1 gpc4626 (
      {stage0_63[369]},
      {stage1_63[191]}
   );
   gpc1_1 gpc4627 (
      {stage0_63[370]},
      {stage1_63[192]}
   );
   gpc1_1 gpc4628 (
      {stage0_63[371]},
      {stage1_63[193]}
   );
   gpc1_1 gpc4629 (
      {stage0_63[372]},
      {stage1_63[194]}
   );
   gpc1_1 gpc4630 (
      {stage0_63[373]},
      {stage1_63[195]}
   );
   gpc1_1 gpc4631 (
      {stage0_63[374]},
      {stage1_63[196]}
   );
   gpc1_1 gpc4632 (
      {stage0_63[375]},
      {stage1_63[197]}
   );
   gpc1_1 gpc4633 (
      {stage0_63[376]},
      {stage1_63[198]}
   );
   gpc1_1 gpc4634 (
      {stage0_63[377]},
      {stage1_63[199]}
   );
   gpc1_1 gpc4635 (
      {stage0_63[378]},
      {stage1_63[200]}
   );
   gpc1_1 gpc4636 (
      {stage0_63[379]},
      {stage1_63[201]}
   );
   gpc1_1 gpc4637 (
      {stage0_63[380]},
      {stage1_63[202]}
   );
   gpc1_1 gpc4638 (
      {stage0_63[381]},
      {stage1_63[203]}
   );
   gpc1_1 gpc4639 (
      {stage0_63[382]},
      {stage1_63[204]}
   );
   gpc1_1 gpc4640 (
      {stage0_63[383]},
      {stage1_63[205]}
   );
   gpc1_1 gpc4641 (
      {stage0_63[384]},
      {stage1_63[206]}
   );
   gpc1_1 gpc4642 (
      {stage0_63[385]},
      {stage1_63[207]}
   );
   gpc1_1 gpc4643 (
      {stage0_63[386]},
      {stage1_63[208]}
   );
   gpc1_1 gpc4644 (
      {stage0_63[387]},
      {stage1_63[209]}
   );
   gpc1_1 gpc4645 (
      {stage0_63[388]},
      {stage1_63[210]}
   );
   gpc1_1 gpc4646 (
      {stage0_63[389]},
      {stage1_63[211]}
   );
   gpc1_1 gpc4647 (
      {stage0_63[390]},
      {stage1_63[212]}
   );
   gpc1_1 gpc4648 (
      {stage0_63[391]},
      {stage1_63[213]}
   );
   gpc1_1 gpc4649 (
      {stage0_63[392]},
      {stage1_63[214]}
   );
   gpc1_1 gpc4650 (
      {stage0_63[393]},
      {stage1_63[215]}
   );
   gpc1_1 gpc4651 (
      {stage0_63[394]},
      {stage1_63[216]}
   );
   gpc1_1 gpc4652 (
      {stage0_63[395]},
      {stage1_63[217]}
   );
   gpc1_1 gpc4653 (
      {stage0_63[396]},
      {stage1_63[218]}
   );
   gpc1_1 gpc4654 (
      {stage0_63[397]},
      {stage1_63[219]}
   );
   gpc1_1 gpc4655 (
      {stage0_63[398]},
      {stage1_63[220]}
   );
   gpc1_1 gpc4656 (
      {stage0_63[399]},
      {stage1_63[221]}
   );
   gpc1_1 gpc4657 (
      {stage0_63[400]},
      {stage1_63[222]}
   );
   gpc1_1 gpc4658 (
      {stage0_63[401]},
      {stage1_63[223]}
   );
   gpc1_1 gpc4659 (
      {stage0_63[402]},
      {stage1_63[224]}
   );
   gpc1_1 gpc4660 (
      {stage0_63[403]},
      {stage1_63[225]}
   );
   gpc1_1 gpc4661 (
      {stage0_63[404]},
      {stage1_63[226]}
   );
   gpc1_1 gpc4662 (
      {stage0_63[405]},
      {stage1_63[227]}
   );
   gpc1_1 gpc4663 (
      {stage0_63[406]},
      {stage1_63[228]}
   );
   gpc1_1 gpc4664 (
      {stage0_63[407]},
      {stage1_63[229]}
   );
   gpc1_1 gpc4665 (
      {stage0_63[408]},
      {stage1_63[230]}
   );
   gpc1_1 gpc4666 (
      {stage0_63[409]},
      {stage1_63[231]}
   );
   gpc1_1 gpc4667 (
      {stage0_63[410]},
      {stage1_63[232]}
   );
   gpc1_1 gpc4668 (
      {stage0_63[411]},
      {stage1_63[233]}
   );
   gpc1_1 gpc4669 (
      {stage0_63[412]},
      {stage1_63[234]}
   );
   gpc1_1 gpc4670 (
      {stage0_63[413]},
      {stage1_63[235]}
   );
   gpc1_1 gpc4671 (
      {stage0_63[414]},
      {stage1_63[236]}
   );
   gpc1_1 gpc4672 (
      {stage0_63[415]},
      {stage1_63[237]}
   );
   gpc1_1 gpc4673 (
      {stage0_63[416]},
      {stage1_63[238]}
   );
   gpc1_1 gpc4674 (
      {stage0_63[417]},
      {stage1_63[239]}
   );
   gpc1_1 gpc4675 (
      {stage0_63[418]},
      {stage1_63[240]}
   );
   gpc1_1 gpc4676 (
      {stage0_63[419]},
      {stage1_63[241]}
   );
   gpc1_1 gpc4677 (
      {stage0_63[420]},
      {stage1_63[242]}
   );
   gpc1_1 gpc4678 (
      {stage0_63[421]},
      {stage1_63[243]}
   );
   gpc1_1 gpc4679 (
      {stage0_63[422]},
      {stage1_63[244]}
   );
   gpc1_1 gpc4680 (
      {stage0_63[423]},
      {stage1_63[245]}
   );
   gpc1_1 gpc4681 (
      {stage0_63[424]},
      {stage1_63[246]}
   );
   gpc1_1 gpc4682 (
      {stage0_63[425]},
      {stage1_63[247]}
   );
   gpc1_1 gpc4683 (
      {stage0_63[426]},
      {stage1_63[248]}
   );
   gpc1_1 gpc4684 (
      {stage0_63[427]},
      {stage1_63[249]}
   );
   gpc1_1 gpc4685 (
      {stage0_63[428]},
      {stage1_63[250]}
   );
   gpc1_1 gpc4686 (
      {stage0_63[429]},
      {stage1_63[251]}
   );
   gpc1_1 gpc4687 (
      {stage0_63[430]},
      {stage1_63[252]}
   );
   gpc1_1 gpc4688 (
      {stage0_63[431]},
      {stage1_63[253]}
   );
   gpc1_1 gpc4689 (
      {stage0_63[432]},
      {stage1_63[254]}
   );
   gpc1_1 gpc4690 (
      {stage0_63[433]},
      {stage1_63[255]}
   );
   gpc1_1 gpc4691 (
      {stage0_63[434]},
      {stage1_63[256]}
   );
   gpc1_1 gpc4692 (
      {stage0_63[435]},
      {stage1_63[257]}
   );
   gpc1_1 gpc4693 (
      {stage0_63[436]},
      {stage1_63[258]}
   );
   gpc1_1 gpc4694 (
      {stage0_63[437]},
      {stage1_63[259]}
   );
   gpc1_1 gpc4695 (
      {stage0_63[438]},
      {stage1_63[260]}
   );
   gpc1_1 gpc4696 (
      {stage0_63[439]},
      {stage1_63[261]}
   );
   gpc1_1 gpc4697 (
      {stage0_63[440]},
      {stage1_63[262]}
   );
   gpc1_1 gpc4698 (
      {stage0_63[441]},
      {stage1_63[263]}
   );
   gpc1_1 gpc4699 (
      {stage0_63[442]},
      {stage1_63[264]}
   );
   gpc1_1 gpc4700 (
      {stage0_63[443]},
      {stage1_63[265]}
   );
   gpc1_1 gpc4701 (
      {stage0_63[444]},
      {stage1_63[266]}
   );
   gpc1_1 gpc4702 (
      {stage0_63[445]},
      {stage1_63[267]}
   );
   gpc1_1 gpc4703 (
      {stage0_63[446]},
      {stage1_63[268]}
   );
   gpc1_1 gpc4704 (
      {stage0_63[447]},
      {stage1_63[269]}
   );
   gpc1_1 gpc4705 (
      {stage0_63[448]},
      {stage1_63[270]}
   );
   gpc1_1 gpc4706 (
      {stage0_63[449]},
      {stage1_63[271]}
   );
   gpc1_1 gpc4707 (
      {stage0_63[450]},
      {stage1_63[272]}
   );
   gpc1_1 gpc4708 (
      {stage0_63[451]},
      {stage1_63[273]}
   );
   gpc1_1 gpc4709 (
      {stage0_63[452]},
      {stage1_63[274]}
   );
   gpc1_1 gpc4710 (
      {stage0_63[453]},
      {stage1_63[275]}
   );
   gpc1_1 gpc4711 (
      {stage0_63[454]},
      {stage1_63[276]}
   );
   gpc1_1 gpc4712 (
      {stage0_63[455]},
      {stage1_63[277]}
   );
   gpc1_1 gpc4713 (
      {stage0_63[456]},
      {stage1_63[278]}
   );
   gpc1_1 gpc4714 (
      {stage0_63[457]},
      {stage1_63[279]}
   );
   gpc1_1 gpc4715 (
      {stage0_63[458]},
      {stage1_63[280]}
   );
   gpc1_1 gpc4716 (
      {stage0_63[459]},
      {stage1_63[281]}
   );
   gpc1_1 gpc4717 (
      {stage0_63[460]},
      {stage1_63[282]}
   );
   gpc1_1 gpc4718 (
      {stage0_63[461]},
      {stage1_63[283]}
   );
   gpc1_1 gpc4719 (
      {stage0_63[462]},
      {stage1_63[284]}
   );
   gpc1_1 gpc4720 (
      {stage0_63[463]},
      {stage1_63[285]}
   );
   gpc1_1 gpc4721 (
      {stage0_63[464]},
      {stage1_63[286]}
   );
   gpc1_1 gpc4722 (
      {stage0_63[465]},
      {stage1_63[287]}
   );
   gpc1_1 gpc4723 (
      {stage0_63[466]},
      {stage1_63[288]}
   );
   gpc1_1 gpc4724 (
      {stage0_63[467]},
      {stage1_63[289]}
   );
   gpc1_1 gpc4725 (
      {stage0_63[468]},
      {stage1_63[290]}
   );
   gpc1_1 gpc4726 (
      {stage0_63[469]},
      {stage1_63[291]}
   );
   gpc1_1 gpc4727 (
      {stage0_63[470]},
      {stage1_63[292]}
   );
   gpc1_1 gpc4728 (
      {stage0_63[471]},
      {stage1_63[293]}
   );
   gpc1_1 gpc4729 (
      {stage0_63[472]},
      {stage1_63[294]}
   );
   gpc1_1 gpc4730 (
      {stage0_63[473]},
      {stage1_63[295]}
   );
   gpc1_1 gpc4731 (
      {stage0_63[474]},
      {stage1_63[296]}
   );
   gpc1_1 gpc4732 (
      {stage0_63[475]},
      {stage1_63[297]}
   );
   gpc1_1 gpc4733 (
      {stage0_63[476]},
      {stage1_63[298]}
   );
   gpc1_1 gpc4734 (
      {stage0_63[477]},
      {stage1_63[299]}
   );
   gpc1_1 gpc4735 (
      {stage0_63[478]},
      {stage1_63[300]}
   );
   gpc1_1 gpc4736 (
      {stage0_63[479]},
      {stage1_63[301]}
   );
   gpc1_1 gpc4737 (
      {stage0_63[480]},
      {stage1_63[302]}
   );
   gpc1_1 gpc4738 (
      {stage0_63[481]},
      {stage1_63[303]}
   );
   gpc1_1 gpc4739 (
      {stage0_63[482]},
      {stage1_63[304]}
   );
   gpc1_1 gpc4740 (
      {stage0_63[483]},
      {stage1_63[305]}
   );
   gpc1_1 gpc4741 (
      {stage0_63[484]},
      {stage1_63[306]}
   );
   gpc1_1 gpc4742 (
      {stage0_63[485]},
      {stage1_63[307]}
   );
   gpc606_5 gpc4743 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc4744 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc4745 (
      {stage1_0[12], stage1_0[13], stage1_0[14], stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc615_5 gpc4746 (
      {stage1_0[18], stage1_0[19], stage1_0[20], stage1_0[21], stage1_0[22]},
      {stage1_1[0]},
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc4747 (
      {stage1_0[23], stage1_0[24], stage1_0[25], stage1_0[26], stage1_0[27]},
      {stage1_1[1]},
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc615_5 gpc4748 (
      {stage1_0[28], stage1_0[29], stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[2]},
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc615_5 gpc4749 (
      {stage1_0[33], stage1_0[34], stage1_0[35], stage1_0[36], stage1_0[37]},
      {stage1_1[3]},
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc615_5 gpc4750 (
      {stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41], stage1_0[42]},
      {stage1_1[4]},
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc615_5 gpc4751 (
      {stage1_0[43], stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_1[5]},
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc615_5 gpc4752 (
      {stage1_0[48], stage1_0[49], stage1_0[50], stage1_0[51], stage1_0[52]},
      {stage1_1[6]},
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc615_5 gpc4753 (
      {stage1_0[53], stage1_0[54], stage1_0[55], stage1_0[56], stage1_0[57]},
      {stage1_1[7]},
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc615_5 gpc4754 (
      {stage1_0[58], stage1_0[59], stage1_0[60], stage1_0[61], stage1_0[62]},
      {stage1_1[8]},
      {stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc615_5 gpc4755 (
      {stage1_0[63], stage1_0[64], stage1_0[65], stage1_0[66], stage1_0[67]},
      {stage1_1[9]},
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc615_5 gpc4756 (
      {stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71], stage1_0[72]},
      {stage1_1[10]},
      {stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82], stage1_2[83]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc615_5 gpc4757 (
      {stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_1[11]},
      {stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87], stage1_2[88], stage1_2[89]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc615_5 gpc4758 (
      {stage1_0[78], stage1_0[79], stage1_0[80], stage1_0[81], stage1_0[82]},
      {stage1_1[12]},
      {stage1_2[90], stage1_2[91], stage1_2[92], stage1_2[93], stage1_2[94], stage1_2[95]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc615_5 gpc4759 (
      {stage1_0[83], stage1_0[84], stage1_0[85], stage1_0[86], stage1_0[87]},
      {stage1_1[13]},
      {stage1_2[96], stage1_2[97], stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc615_5 gpc4760 (
      {stage1_0[88], stage1_0[89], stage1_0[90], stage1_0[91], stage1_0[92]},
      {stage1_1[14]},
      {stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106], stage1_2[107]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc615_5 gpc4761 (
      {stage1_0[93], stage1_0[94], stage1_0[95], stage1_0[96], stage1_0[97]},
      {stage1_1[15]},
      {stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111], stage1_2[112], stage1_2[113]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc615_5 gpc4762 (
      {stage1_0[98], stage1_0[99], stage1_0[100], stage1_0[101], stage1_0[102]},
      {stage1_1[16]},
      {stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117], stage1_2[118], stage1_2[119]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc615_5 gpc4763 (
      {stage1_0[103], stage1_0[104], stage1_0[105], stage1_0[106], stage1_0[107]},
      {stage1_1[17]},
      {stage1_2[120], stage1_2[121], stage1_2[122], stage1_2[123], stage1_2[124], stage1_2[125]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc4764 (
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21]}
   );
   gpc606_5 gpc4765 (
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22]}
   );
   gpc606_5 gpc4766 (
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc4767 (
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[3],stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24]}
   );
   gpc606_5 gpc4768 (
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29]},
      {stage2_5[4],stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25]}
   );
   gpc606_5 gpc4769 (
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35]},
      {stage2_5[5],stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26]}
   );
   gpc606_5 gpc4770 (
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage2_5[6],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc4771 (
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47]},
      {stage2_5[7],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc4772 (
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage2_5[8],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc4773 (
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59]},
      {stage2_5[9],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc4774 (
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage2_5[10],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc4775 (
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage2_5[11],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc4776 (
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77]},
      {stage2_5[12],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc4777 (
      {stage1_1[96], stage1_1[97], stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101]},
      {stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83]},
      {stage2_5[13],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc4778 (
      {stage1_1[102], stage1_1[103], stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107]},
      {stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89]},
      {stage2_5[14],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc606_5 gpc4779 (
      {stage1_1[108], stage1_1[109], stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113]},
      {stage1_3[90], stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage2_5[15],stage2_4[36],stage2_3[36],stage2_2[36],stage2_1[36]}
   );
   gpc606_5 gpc4780 (
      {stage1_1[114], stage1_1[115], stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119]},
      {stage1_3[96], stage1_3[97], stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101]},
      {stage2_5[16],stage2_4[37],stage2_3[37],stage2_2[37],stage2_1[37]}
   );
   gpc606_5 gpc4781 (
      {stage1_1[120], stage1_1[121], stage1_1[122], stage1_1[123], stage1_1[124], stage1_1[125]},
      {stage1_3[102], stage1_3[103], stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107]},
      {stage2_5[17],stage2_4[38],stage2_3[38],stage2_2[38],stage2_1[38]}
   );
   gpc606_5 gpc4782 (
      {stage1_1[126], stage1_1[127], stage1_1[128], stage1_1[129], stage1_1[130], stage1_1[131]},
      {stage1_3[108], stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112], stage1_3[113]},
      {stage2_5[18],stage2_4[39],stage2_3[39],stage2_2[39],stage2_1[39]}
   );
   gpc606_5 gpc4783 (
      {stage1_1[132], stage1_1[133], stage1_1[134], stage1_1[135], stage1_1[136], stage1_1[137]},
      {stage1_3[114], stage1_3[115], stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119]},
      {stage2_5[19],stage2_4[40],stage2_3[40],stage2_2[40],stage2_1[40]}
   );
   gpc606_5 gpc4784 (
      {stage1_1[138], stage1_1[139], stage1_1[140], stage1_1[141], stage1_1[142], stage1_1[143]},
      {stage1_3[120], stage1_3[121], stage1_3[122], stage1_3[123], stage1_3[124], stage1_3[125]},
      {stage2_5[20],stage2_4[41],stage2_3[41],stage2_2[41],stage2_1[41]}
   );
   gpc606_5 gpc4785 (
      {stage1_1[144], stage1_1[145], stage1_1[146], stage1_1[147], stage1_1[148], stage1_1[149]},
      {stage1_3[126], stage1_3[127], stage1_3[128], stage1_3[129], stage1_3[130], stage1_3[131]},
      {stage2_5[21],stage2_4[42],stage2_3[42],stage2_2[42],stage2_1[42]}
   );
   gpc606_5 gpc4786 (
      {stage1_1[150], stage1_1[151], stage1_1[152], stage1_1[153], stage1_1[154], stage1_1[155]},
      {stage1_3[132], stage1_3[133], stage1_3[134], stage1_3[135], stage1_3[136], stage1_3[137]},
      {stage2_5[22],stage2_4[43],stage2_3[43],stage2_2[43],stage2_1[43]}
   );
   gpc606_5 gpc4787 (
      {stage1_1[156], stage1_1[157], stage1_1[158], stage1_1[159], stage1_1[160], stage1_1[161]},
      {stage1_3[138], stage1_3[139], stage1_3[140], stage1_3[141], stage1_3[142], stage1_3[143]},
      {stage2_5[23],stage2_4[44],stage2_3[44],stage2_2[44],stage2_1[44]}
   );
   gpc606_5 gpc4788 (
      {stage1_1[162], stage1_1[163], stage1_1[164], stage1_1[165], stage1_1[166], stage1_1[167]},
      {stage1_3[144], stage1_3[145], stage1_3[146], stage1_3[147], stage1_3[148], stage1_3[149]},
      {stage2_5[24],stage2_4[45],stage2_3[45],stage2_2[45],stage2_1[45]}
   );
   gpc606_5 gpc4789 (
      {stage1_2[126], stage1_2[127], stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[25],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc606_5 gpc4790 (
      {stage1_2[132], stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[26],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc606_5 gpc4791 (
      {stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142], stage1_2[143]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[27],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc1343_5 gpc4792 (
      {stage1_4[18], stage1_4[19], stage1_4[20]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3]},
      {stage1_6[0], stage1_6[1], stage1_6[2]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[0],stage2_6[3],stage2_5[28],stage2_4[49]}
   );
   gpc1406_5 gpc4793 (
      {stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage1_7[1]},
      {stage2_8[1],stage2_7[1],stage2_6[4],stage2_5[29],stage2_4[50]}
   );
   gpc606_5 gpc4794 (
      {stage1_4[27], stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31], stage1_4[32]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[2],stage2_7[2],stage2_6[5],stage2_5[30],stage2_4[51]}
   );
   gpc606_5 gpc4795 (
      {stage1_4[33], stage1_4[34], stage1_4[35], stage1_4[36], stage1_4[37], stage1_4[38]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[3],stage2_7[3],stage2_6[6],stage2_5[31],stage2_4[52]}
   );
   gpc606_5 gpc4796 (
      {stage1_4[39], stage1_4[40], stage1_4[41], stage1_4[42], stage1_4[43], stage1_4[44]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[4],stage2_7[4],stage2_6[7],stage2_5[32],stage2_4[53]}
   );
   gpc606_5 gpc4797 (
      {stage1_4[45], stage1_4[46], stage1_4[47], stage1_4[48], stage1_4[49], stage1_4[50]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[5],stage2_7[5],stage2_6[8],stage2_5[33],stage2_4[54]}
   );
   gpc606_5 gpc4798 (
      {stage1_4[51], stage1_4[52], stage1_4[53], stage1_4[54], stage1_4[55], stage1_4[56]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[6],stage2_7[6],stage2_6[9],stage2_5[34],stage2_4[55]}
   );
   gpc606_5 gpc4799 (
      {stage1_4[57], stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61], stage1_4[62]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[7],stage2_7[7],stage2_6[10],stage2_5[35],stage2_4[56]}
   );
   gpc606_5 gpc4800 (
      {stage1_4[63], stage1_4[64], stage1_4[65], stage1_4[66], stage1_4[67], stage1_4[68]},
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage2_8[8],stage2_7[8],stage2_6[11],stage2_5[36],stage2_4[57]}
   );
   gpc606_5 gpc4801 (
      {stage1_4[69], stage1_4[70], stage1_4[71], stage1_4[72], stage1_4[73], stage1_4[74]},
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54]},
      {stage2_8[9],stage2_7[9],stage2_6[12],stage2_5[37],stage2_4[58]}
   );
   gpc606_5 gpc4802 (
      {stage1_4[75], stage1_4[76], stage1_4[77], stage1_4[78], stage1_4[79], stage1_4[80]},
      {stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage2_8[10],stage2_7[10],stage2_6[13],stage2_5[38],stage2_4[59]}
   );
   gpc606_5 gpc4803 (
      {stage1_4[81], stage1_4[82], stage1_4[83], stage1_4[84], stage1_4[85], stage1_4[86]},
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66]},
      {stage2_8[11],stage2_7[11],stage2_6[14],stage2_5[39],stage2_4[60]}
   );
   gpc606_5 gpc4804 (
      {stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91], stage1_4[92]},
      {stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71], stage1_6[72]},
      {stage2_8[12],stage2_7[12],stage2_6[15],stage2_5[40],stage2_4[61]}
   );
   gpc606_5 gpc4805 (
      {stage1_4[93], stage1_4[94], stage1_4[95], stage1_4[96], stage1_4[97], stage1_4[98]},
      {stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78]},
      {stage2_8[13],stage2_7[13],stage2_6[16],stage2_5[41],stage2_4[62]}
   );
   gpc606_5 gpc4806 (
      {stage1_4[99], stage1_4[100], stage1_4[101], stage1_4[102], stage1_4[103], stage1_4[104]},
      {stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84]},
      {stage2_8[14],stage2_7[14],stage2_6[17],stage2_5[42],stage2_4[63]}
   );
   gpc606_5 gpc4807 (
      {stage1_4[105], stage1_4[106], stage1_4[107], stage1_4[108], stage1_4[109], stage1_4[110]},
      {stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage2_8[15],stage2_7[15],stage2_6[18],stage2_5[43],stage2_4[64]}
   );
   gpc606_5 gpc4808 (
      {stage1_4[111], stage1_4[112], stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116]},
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96]},
      {stage2_8[16],stage2_7[16],stage2_6[19],stage2_5[44],stage2_4[65]}
   );
   gpc606_5 gpc4809 (
      {stage1_4[117], stage1_4[118], stage1_4[119], stage1_4[120], stage1_4[121], stage1_4[122]},
      {stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101], stage1_6[102]},
      {stage2_8[17],stage2_7[17],stage2_6[20],stage2_5[45],stage2_4[66]}
   );
   gpc606_5 gpc4810 (
      {stage1_4[123], stage1_4[124], stage1_4[125], stage1_4[126], stage1_4[127], stage1_4[128]},
      {stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107], stage1_6[108]},
      {stage2_8[18],stage2_7[18],stage2_6[21],stage2_5[46],stage2_4[67]}
   );
   gpc606_5 gpc4811 (
      {stage1_4[129], stage1_4[130], stage1_4[131], stage1_4[132], stage1_4[133], stage1_4[134]},
      {stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114]},
      {stage2_8[19],stage2_7[19],stage2_6[22],stage2_5[47],stage2_4[68]}
   );
   gpc606_5 gpc4812 (
      {stage1_4[135], stage1_4[136], stage1_4[137], stage1_4[138], stage1_4[139], stage1_4[140]},
      {stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119], stage1_6[120]},
      {stage2_8[20],stage2_7[20],stage2_6[23],stage2_5[48],stage2_4[69]}
   );
   gpc606_5 gpc4813 (
      {stage1_4[141], stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145], stage1_4[146]},
      {stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125], stage1_6[126]},
      {stage2_8[21],stage2_7[21],stage2_6[24],stage2_5[49],stage2_4[70]}
   );
   gpc606_5 gpc4814 (
      {stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150], stage1_4[151], stage1_4[152]},
      {stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131], stage1_6[132]},
      {stage2_8[22],stage2_7[22],stage2_6[25],stage2_5[50],stage2_4[71]}
   );
   gpc606_5 gpc4815 (
      {stage1_4[153], stage1_4[154], stage1_4[155], stage1_4[156], stage1_4[157], stage1_4[158]},
      {stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137], stage1_6[138]},
      {stage2_8[23],stage2_7[23],stage2_6[26],stage2_5[51],stage2_4[72]}
   );
   gpc606_5 gpc4816 (
      {stage1_4[159], stage1_4[160], stage1_4[161], stage1_4[162], stage1_4[163], stage1_4[164]},
      {stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143], stage1_6[144]},
      {stage2_8[24],stage2_7[24],stage2_6[27],stage2_5[52],stage2_4[73]}
   );
   gpc606_5 gpc4817 (
      {stage1_4[165], stage1_4[166], stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170]},
      {stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149], stage1_6[150]},
      {stage2_8[25],stage2_7[25],stage2_6[28],stage2_5[53],stage2_4[74]}
   );
   gpc606_5 gpc4818 (
      {stage1_4[171], stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175], stage1_4[176]},
      {stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155], stage1_6[156]},
      {stage2_8[26],stage2_7[26],stage2_6[29],stage2_5[54],stage2_4[75]}
   );
   gpc606_5 gpc4819 (
      {stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180], stage1_4[181], stage1_4[182]},
      {stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161], stage1_6[162]},
      {stage2_8[27],stage2_7[27],stage2_6[30],stage2_5[55],stage2_4[76]}
   );
   gpc606_5 gpc4820 (
      {stage1_4[183], stage1_4[184], stage1_4[185], stage1_4[186], stage1_4[187], stage1_4[188]},
      {stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166], stage1_6[167], stage1_6[168]},
      {stage2_8[28],stage2_7[28],stage2_6[31],stage2_5[56],stage2_4[77]}
   );
   gpc606_5 gpc4821 (
      {stage1_4[189], stage1_4[190], stage1_4[191], stage1_4[192], stage1_4[193], stage1_4[194]},
      {stage1_6[169], stage1_6[170], stage1_6[171], stage1_6[172], stage1_6[173], stage1_6[174]},
      {stage2_8[29],stage2_7[29],stage2_6[32],stage2_5[57],stage2_4[78]}
   );
   gpc606_5 gpc4822 (
      {stage1_5[4], stage1_5[5], stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9]},
      {stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7]},
      {stage2_9[0],stage2_8[30],stage2_7[30],stage2_6[33],stage2_5[58]}
   );
   gpc606_5 gpc4823 (
      {stage1_5[10], stage1_5[11], stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15]},
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13]},
      {stage2_9[1],stage2_8[31],stage2_7[31],stage2_6[34],stage2_5[59]}
   );
   gpc606_5 gpc4824 (
      {stage1_5[16], stage1_5[17], stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21]},
      {stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18], stage1_7[19]},
      {stage2_9[2],stage2_8[32],stage2_7[32],stage2_6[35],stage2_5[60]}
   );
   gpc606_5 gpc4825 (
      {stage1_5[22], stage1_5[23], stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27]},
      {stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24], stage1_7[25]},
      {stage2_9[3],stage2_8[33],stage2_7[33],stage2_6[36],stage2_5[61]}
   );
   gpc606_5 gpc4826 (
      {stage1_5[28], stage1_5[29], stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33]},
      {stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30], stage1_7[31]},
      {stage2_9[4],stage2_8[34],stage2_7[34],stage2_6[37],stage2_5[62]}
   );
   gpc606_5 gpc4827 (
      {stage1_5[34], stage1_5[35], stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39]},
      {stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37]},
      {stage2_9[5],stage2_8[35],stage2_7[35],stage2_6[38],stage2_5[63]}
   );
   gpc606_5 gpc4828 (
      {stage1_5[40], stage1_5[41], stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45]},
      {stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage2_9[6],stage2_8[36],stage2_7[36],stage2_6[39],stage2_5[64]}
   );
   gpc606_5 gpc4829 (
      {stage1_5[46], stage1_5[47], stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51]},
      {stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48], stage1_7[49]},
      {stage2_9[7],stage2_8[37],stage2_7[37],stage2_6[40],stage2_5[65]}
   );
   gpc606_5 gpc4830 (
      {stage1_5[52], stage1_5[53], stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57]},
      {stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53], stage1_7[54], stage1_7[55]},
      {stage2_9[8],stage2_8[38],stage2_7[38],stage2_6[41],stage2_5[66]}
   );
   gpc606_5 gpc4831 (
      {stage1_5[58], stage1_5[59], stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63]},
      {stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60], stage1_7[61]},
      {stage2_9[9],stage2_8[39],stage2_7[39],stage2_6[42],stage2_5[67]}
   );
   gpc606_5 gpc4832 (
      {stage1_5[64], stage1_5[65], stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69]},
      {stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66], stage1_7[67]},
      {stage2_9[10],stage2_8[40],stage2_7[40],stage2_6[43],stage2_5[68]}
   );
   gpc606_5 gpc4833 (
      {stage1_5[70], stage1_5[71], stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75]},
      {stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71], stage1_7[72], stage1_7[73]},
      {stage2_9[11],stage2_8[41],stage2_7[41],stage2_6[44],stage2_5[69]}
   );
   gpc606_5 gpc4834 (
      {stage1_5[76], stage1_5[77], stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81]},
      {stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77], stage1_7[78], stage1_7[79]},
      {stage2_9[12],stage2_8[42],stage2_7[42],stage2_6[45],stage2_5[70]}
   );
   gpc606_5 gpc4835 (
      {stage1_5[82], stage1_5[83], stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87]},
      {stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85]},
      {stage2_9[13],stage2_8[43],stage2_7[43],stage2_6[46],stage2_5[71]}
   );
   gpc606_5 gpc4836 (
      {stage1_5[88], stage1_5[89], stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93]},
      {stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], stage1_7[91]},
      {stage2_9[14],stage2_8[44],stage2_7[44],stage2_6[47],stage2_5[72]}
   );
   gpc606_5 gpc4837 (
      {stage1_5[94], stage1_5[95], stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99]},
      {stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95], stage1_7[96], stage1_7[97]},
      {stage2_9[15],stage2_8[45],stage2_7[45],stage2_6[48],stage2_5[73]}
   );
   gpc606_5 gpc4838 (
      {stage1_5[100], stage1_5[101], stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105]},
      {stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101], stage1_7[102], stage1_7[103]},
      {stage2_9[16],stage2_8[46],stage2_7[46],stage2_6[49],stage2_5[74]}
   );
   gpc606_5 gpc4839 (
      {stage1_5[106], stage1_5[107], stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111]},
      {stage1_7[104], stage1_7[105], stage1_7[106], stage1_7[107], stage1_7[108], stage1_7[109]},
      {stage2_9[17],stage2_8[47],stage2_7[47],stage2_6[50],stage2_5[75]}
   );
   gpc606_5 gpc4840 (
      {stage1_5[112], stage1_5[113], stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117]},
      {stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113], stage1_7[114], stage1_7[115]},
      {stage2_9[18],stage2_8[48],stage2_7[48],stage2_6[51],stage2_5[76]}
   );
   gpc606_5 gpc4841 (
      {stage1_5[118], stage1_5[119], stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123]},
      {stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120], stage1_7[121]},
      {stage2_9[19],stage2_8[49],stage2_7[49],stage2_6[52],stage2_5[77]}
   );
   gpc615_5 gpc4842 (
      {stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125], stage1_7[126]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[20],stage2_8[50],stage2_7[50]}
   );
   gpc615_5 gpc4843 (
      {stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130], stage1_7[131]},
      {stage1_8[1]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[1],stage2_9[21],stage2_8[51],stage2_7[51]}
   );
   gpc615_5 gpc4844 (
      {stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135], stage1_7[136]},
      {stage1_8[2]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[2],stage2_9[22],stage2_8[52],stage2_7[52]}
   );
   gpc615_5 gpc4845 (
      {stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140], stage1_7[141]},
      {stage1_8[3]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[3],stage2_9[23],stage2_8[53],stage2_7[53]}
   );
   gpc615_5 gpc4846 (
      {stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145], stage1_7[146]},
      {stage1_8[4]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[4],stage2_9[24],stage2_8[54],stage2_7[54]}
   );
   gpc615_5 gpc4847 (
      {stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150], stage1_7[151]},
      {stage1_8[5]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[5],stage2_9[25],stage2_8[55],stage2_7[55]}
   );
   gpc615_5 gpc4848 (
      {stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155], stage1_7[156]},
      {stage1_8[6]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[6],stage2_9[26],stage2_8[56],stage2_7[56]}
   );
   gpc615_5 gpc4849 (
      {stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160], stage1_7[161]},
      {stage1_8[7]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[7],stage2_9[27],stage2_8[57],stage2_7[57]}
   );
   gpc615_5 gpc4850 (
      {stage1_7[162], stage1_7[163], stage1_7[164], stage1_7[165], stage1_7[166]},
      {stage1_8[8]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[8],stage2_9[28],stage2_8[58],stage2_7[58]}
   );
   gpc615_5 gpc4851 (
      {stage1_7[167], stage1_7[168], stage1_7[169], stage1_7[170], stage1_7[171]},
      {stage1_8[9]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[9],stage2_9[29],stage2_8[59],stage2_7[59]}
   );
   gpc615_5 gpc4852 (
      {stage1_7[172], stage1_7[173], stage1_7[174], stage1_7[175], stage1_7[176]},
      {stage1_8[10]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[10],stage2_9[30],stage2_8[60],stage2_7[60]}
   );
   gpc615_5 gpc4853 (
      {stage1_7[177], stage1_7[178], stage1_7[179], stage1_7[180], stage1_7[181]},
      {stage1_8[11]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[11],stage2_9[31],stage2_8[61],stage2_7[61]}
   );
   gpc615_5 gpc4854 (
      {stage1_7[182], stage1_7[183], stage1_7[184], stage1_7[185], stage1_7[186]},
      {stage1_8[12]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[12],stage2_9[32],stage2_8[62],stage2_7[62]}
   );
   gpc615_5 gpc4855 (
      {stage1_7[187], stage1_7[188], stage1_7[189], stage1_7[190], stage1_7[191]},
      {stage1_8[13]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[13],stage2_9[33],stage2_8[63],stage2_7[63]}
   );
   gpc615_5 gpc4856 (
      {stage1_7[192], stage1_7[193], stage1_7[194], stage1_7[195], stage1_7[196]},
      {stage1_8[14]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[14],stage2_9[34],stage2_8[64],stage2_7[64]}
   );
   gpc615_5 gpc4857 (
      {stage1_7[197], stage1_7[198], stage1_7[199], stage1_7[200], stage1_7[201]},
      {stage1_8[15]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[15],stage2_9[35],stage2_8[65],stage2_7[65]}
   );
   gpc615_5 gpc4858 (
      {stage1_7[202], stage1_7[203], stage1_7[204], stage1_7[205], stage1_7[206]},
      {stage1_8[16]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[16],stage2_9[36],stage2_8[66],stage2_7[66]}
   );
   gpc615_5 gpc4859 (
      {stage1_7[207], stage1_7[208], stage1_7[209], stage1_7[210], stage1_7[211]},
      {stage1_8[17]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[17],stage2_9[37],stage2_8[67],stage2_7[67]}
   );
   gpc615_5 gpc4860 (
      {stage1_7[212], stage1_7[213], stage1_7[214], stage1_7[215], stage1_7[216]},
      {stage1_8[18]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[18],stage2_9[38],stage2_8[68],stage2_7[68]}
   );
   gpc207_4 gpc4861 (
      {stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25]},
      {stage1_10[0], stage1_10[1]},
      {stage2_11[19],stage2_10[19],stage2_9[39],stage2_8[69]}
   );
   gpc606_5 gpc4862 (
      {stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29], stage1_8[30], stage1_8[31]},
      {stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6], stage1_10[7]},
      {stage2_12[0],stage2_11[20],stage2_10[20],stage2_9[40],stage2_8[70]}
   );
   gpc606_5 gpc4863 (
      {stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35], stage1_8[36], stage1_8[37]},
      {stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12], stage1_10[13]},
      {stage2_12[1],stage2_11[21],stage2_10[21],stage2_9[41],stage2_8[71]}
   );
   gpc606_5 gpc4864 (
      {stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41], stage1_8[42], stage1_8[43]},
      {stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19]},
      {stage2_12[2],stage2_11[22],stage2_10[22],stage2_9[42],stage2_8[72]}
   );
   gpc606_5 gpc4865 (
      {stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48], stage1_8[49]},
      {stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23], stage1_10[24], stage1_10[25]},
      {stage2_12[3],stage2_11[23],stage2_10[23],stage2_9[43],stage2_8[73]}
   );
   gpc606_5 gpc4866 (
      {stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53], stage1_8[54], stage1_8[55]},
      {stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29], stage1_10[30], stage1_10[31]},
      {stage2_12[4],stage2_11[24],stage2_10[24],stage2_9[44],stage2_8[74]}
   );
   gpc606_5 gpc4867 (
      {stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59], stage1_8[60], stage1_8[61]},
      {stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36], stage1_10[37]},
      {stage2_12[5],stage2_11[25],stage2_10[25],stage2_9[45],stage2_8[75]}
   );
   gpc606_5 gpc4868 (
      {stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65], stage1_8[66], stage1_8[67]},
      {stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41], stage1_10[42], stage1_10[43]},
      {stage2_12[6],stage2_11[26],stage2_10[26],stage2_9[46],stage2_8[76]}
   );
   gpc606_5 gpc4869 (
      {stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71], stage1_8[72], stage1_8[73]},
      {stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47], stage1_10[48], stage1_10[49]},
      {stage2_12[7],stage2_11[27],stage2_10[27],stage2_9[47],stage2_8[77]}
   );
   gpc606_5 gpc4870 (
      {stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77], stage1_8[78], stage1_8[79]},
      {stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55]},
      {stage2_12[8],stage2_11[28],stage2_10[28],stage2_9[48],stage2_8[78]}
   );
   gpc606_5 gpc4871 (
      {stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83], stage1_8[84], stage1_8[85]},
      {stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59], stage1_10[60], stage1_10[61]},
      {stage2_12[9],stage2_11[29],stage2_10[29],stage2_9[49],stage2_8[79]}
   );
   gpc606_5 gpc4872 (
      {stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89], stage1_8[90], stage1_8[91]},
      {stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65], stage1_10[66], stage1_10[67]},
      {stage2_12[10],stage2_11[30],stage2_10[30],stage2_9[50],stage2_8[80]}
   );
   gpc606_5 gpc4873 (
      {stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95], stage1_8[96], stage1_8[97]},
      {stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71], stage1_10[72], stage1_10[73]},
      {stage2_12[11],stage2_11[31],stage2_10[31],stage2_9[51],stage2_8[81]}
   );
   gpc606_5 gpc4874 (
      {stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101], stage1_8[102], stage1_8[103]},
      {stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77], stage1_10[78], stage1_10[79]},
      {stage2_12[12],stage2_11[32],stage2_10[32],stage2_9[52],stage2_8[82]}
   );
   gpc606_5 gpc4875 (
      {stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107], stage1_8[108], stage1_8[109]},
      {stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83], stage1_10[84], stage1_10[85]},
      {stage2_12[13],stage2_11[33],stage2_10[33],stage2_9[53],stage2_8[83]}
   );
   gpc606_5 gpc4876 (
      {stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113], stage1_8[114], stage1_8[115]},
      {stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89], stage1_10[90], stage1_10[91]},
      {stage2_12[14],stage2_11[34],stage2_10[34],stage2_9[54],stage2_8[84]}
   );
   gpc606_5 gpc4877 (
      {stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119], stage1_8[120], stage1_8[121]},
      {stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95], stage1_10[96], stage1_10[97]},
      {stage2_12[15],stage2_11[35],stage2_10[35],stage2_9[55],stage2_8[85]}
   );
   gpc606_5 gpc4878 (
      {stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125], stage1_8[126], stage1_8[127]},
      {stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101], stage1_10[102], stage1_10[103]},
      {stage2_12[16],stage2_11[36],stage2_10[36],stage2_9[56],stage2_8[86]}
   );
   gpc606_5 gpc4879 (
      {stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131], stage1_8[132], stage1_8[133]},
      {stage1_10[104], stage1_10[105], stage1_10[106], stage1_10[107], stage1_10[108], stage1_10[109]},
      {stage2_12[17],stage2_11[37],stage2_10[37],stage2_9[57],stage2_8[87]}
   );
   gpc606_5 gpc4880 (
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[18],stage2_11[38],stage2_10[38],stage2_9[58]}
   );
   gpc606_5 gpc4881 (
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[19],stage2_11[39],stage2_10[39],stage2_9[59]}
   );
   gpc606_5 gpc4882 (
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[20],stage2_11[40],stage2_10[40],stage2_9[60]}
   );
   gpc615_5 gpc4883 (
      {stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113], stage1_10[114]},
      {stage1_11[18]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[3],stage2_12[21],stage2_11[41],stage2_10[41]}
   );
   gpc615_5 gpc4884 (
      {stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119]},
      {stage1_11[19]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[4],stage2_12[22],stage2_11[42],stage2_10[42]}
   );
   gpc615_5 gpc4885 (
      {stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124]},
      {stage1_11[20]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[5],stage2_12[23],stage2_11[43],stage2_10[43]}
   );
   gpc615_5 gpc4886 (
      {stage1_10[125], stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129]},
      {stage1_11[21]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[6],stage2_12[24],stage2_11[44],stage2_10[44]}
   );
   gpc615_5 gpc4887 (
      {stage1_10[130], stage1_10[131], stage1_10[132], stage1_10[133], stage1_10[134]},
      {stage1_11[22]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[7],stage2_12[25],stage2_11[45],stage2_10[45]}
   );
   gpc615_5 gpc4888 (
      {stage1_10[135], stage1_10[136], stage1_10[137], stage1_10[138], stage1_10[139]},
      {stage1_11[23]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[8],stage2_12[26],stage2_11[46],stage2_10[46]}
   );
   gpc615_5 gpc4889 (
      {stage1_10[140], stage1_10[141], stage1_10[142], stage1_10[143], stage1_10[144]},
      {stage1_11[24]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[9],stage2_12[27],stage2_11[47],stage2_10[47]}
   );
   gpc615_5 gpc4890 (
      {stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148], stage1_10[149]},
      {stage1_11[25]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[10],stage2_12[28],stage2_11[48],stage2_10[48]}
   );
   gpc615_5 gpc4891 (
      {stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154]},
      {stage1_11[26]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[11],stage2_12[29],stage2_11[49],stage2_10[49]}
   );
   gpc615_5 gpc4892 (
      {stage1_10[155], stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159]},
      {stage1_11[27]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[12],stage2_12[30],stage2_11[50],stage2_10[50]}
   );
   gpc615_5 gpc4893 (
      {stage1_10[160], stage1_10[161], stage1_10[162], stage1_10[163], stage1_10[164]},
      {stage1_11[28]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[13],stage2_12[31],stage2_11[51],stage2_10[51]}
   );
   gpc615_5 gpc4894 (
      {stage1_10[165], stage1_10[166], stage1_10[167], stage1_10[168], stage1_10[169]},
      {stage1_11[29]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[14],stage2_12[32],stage2_11[52],stage2_10[52]}
   );
   gpc615_5 gpc4895 (
      {stage1_10[170], stage1_10[171], stage1_10[172], stage1_10[173], stage1_10[174]},
      {stage1_11[30]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[15],stage2_12[33],stage2_11[53],stage2_10[53]}
   );
   gpc606_5 gpc4896 (
      {stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35], stage1_11[36]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[13],stage2_13[16],stage2_12[34],stage2_11[54]}
   );
   gpc606_5 gpc4897 (
      {stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[14],stage2_13[17],stage2_12[35],stage2_11[55]}
   );
   gpc606_5 gpc4898 (
      {stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[15],stage2_13[18],stage2_12[36],stage2_11[56]}
   );
   gpc606_5 gpc4899 (
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53], stage1_11[54]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[16],stage2_13[19],stage2_12[37],stage2_11[57]}
   );
   gpc606_5 gpc4900 (
      {stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59], stage1_11[60]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[17],stage2_13[20],stage2_12[38],stage2_11[58]}
   );
   gpc606_5 gpc4901 (
      {stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65], stage1_11[66]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[18],stage2_13[21],stage2_12[39],stage2_11[59]}
   );
   gpc606_5 gpc4902 (
      {stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71], stage1_11[72]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[19],stage2_13[22],stage2_12[40],stage2_11[60]}
   );
   gpc606_5 gpc4903 (
      {stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77], stage1_11[78]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[20],stage2_13[23],stage2_12[41],stage2_11[61]}
   );
   gpc606_5 gpc4904 (
      {stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83], stage1_11[84]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[21],stage2_13[24],stage2_12[42],stage2_11[62]}
   );
   gpc606_5 gpc4905 (
      {stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89], stage1_11[90]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[22],stage2_13[25],stage2_12[43],stage2_11[63]}
   );
   gpc606_5 gpc4906 (
      {stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95], stage1_11[96]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[23],stage2_13[26],stage2_12[44],stage2_11[64]}
   );
   gpc606_5 gpc4907 (
      {stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101], stage1_11[102]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[24],stage2_13[27],stage2_12[45],stage2_11[65]}
   );
   gpc606_5 gpc4908 (
      {stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108]},
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage2_15[12],stage2_14[25],stage2_13[28],stage2_12[46],stage2_11[66]}
   );
   gpc606_5 gpc4909 (
      {stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage2_15[13],stage2_14[26],stage2_13[29],stage2_12[47],stage2_11[67]}
   );
   gpc606_5 gpc4910 (
      {stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119], stage1_11[120]},
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage2_15[14],stage2_14[27],stage2_13[30],stage2_12[48],stage2_11[68]}
   );
   gpc606_5 gpc4911 (
      {stage1_11[121], stage1_11[122], stage1_11[123], stage1_11[124], stage1_11[125], stage1_11[126]},
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage2_15[15],stage2_14[28],stage2_13[31],stage2_12[49],stage2_11[69]}
   );
   gpc606_5 gpc4912 (
      {stage1_11[127], stage1_11[128], stage1_11[129], stage1_11[130], stage1_11[131], stage1_11[132]},
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage2_15[16],stage2_14[29],stage2_13[32],stage2_12[50],stage2_11[70]}
   );
   gpc615_5 gpc4913 (
      {stage1_11[133], stage1_11[134], stage1_11[135], stage1_11[136], stage1_11[137]},
      {stage1_12[78]},
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage2_15[17],stage2_14[30],stage2_13[33],stage2_12[51],stage2_11[71]}
   );
   gpc615_5 gpc4914 (
      {stage1_11[138], stage1_11[139], stage1_11[140], stage1_11[141], stage1_11[142]},
      {stage1_12[79]},
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage2_15[18],stage2_14[31],stage2_13[34],stage2_12[52],stage2_11[72]}
   );
   gpc615_5 gpc4915 (
      {stage1_11[143], stage1_11[144], stage1_11[145], stage1_11[146], stage1_11[147]},
      {stage1_12[80]},
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage2_15[19],stage2_14[32],stage2_13[35],stage2_12[53],stage2_11[73]}
   );
   gpc615_5 gpc4916 (
      {stage1_11[148], stage1_11[149], stage1_11[150], stage1_11[151], stage1_11[152]},
      {stage1_12[81]},
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage2_15[20],stage2_14[33],stage2_13[36],stage2_12[54],stage2_11[74]}
   );
   gpc615_5 gpc4917 (
      {stage1_11[153], stage1_11[154], stage1_11[155], stage1_11[156], stage1_11[157]},
      {stage1_12[82]},
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage2_15[21],stage2_14[34],stage2_13[37],stage2_12[55],stage2_11[75]}
   );
   gpc615_5 gpc4918 (
      {stage1_11[158], stage1_11[159], stage1_11[160], stage1_11[161], stage1_11[162]},
      {stage1_12[83]},
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136], stage1_13[137]},
      {stage2_15[22],stage2_14[35],stage2_13[38],stage2_12[56],stage2_11[76]}
   );
   gpc615_5 gpc4919 (
      {stage1_11[163], stage1_11[164], stage1_11[165], stage1_11[166], stage1_11[167]},
      {stage1_12[84]},
      {stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141], stage1_13[142], stage1_13[143]},
      {stage2_15[23],stage2_14[36],stage2_13[39],stage2_12[57],stage2_11[77]}
   );
   gpc615_5 gpc4920 (
      {stage1_11[168], stage1_11[169], stage1_11[170], stage1_11[171], stage1_11[172]},
      {stage1_12[85]},
      {stage1_13[144], stage1_13[145], stage1_13[146], stage1_13[147], stage1_13[148], stage1_13[149]},
      {stage2_15[24],stage2_14[37],stage2_13[40],stage2_12[58],stage2_11[78]}
   );
   gpc615_5 gpc4921 (
      {stage1_11[173], stage1_11[174], stage1_11[175], stage1_11[176], stage1_11[177]},
      {stage1_12[86]},
      {stage1_13[150], stage1_13[151], stage1_13[152], stage1_13[153], stage1_13[154], stage1_13[155]},
      {stage2_15[25],stage2_14[38],stage2_13[41],stage2_12[59],stage2_11[79]}
   );
   gpc615_5 gpc4922 (
      {stage1_11[178], stage1_11[179], stage1_11[180], stage1_11[181], stage1_11[182]},
      {stage1_12[87]},
      {stage1_13[156], stage1_13[157], stage1_13[158], stage1_13[159], stage1_13[160], stage1_13[161]},
      {stage2_15[26],stage2_14[39],stage2_13[42],stage2_12[60],stage2_11[80]}
   );
   gpc615_5 gpc4923 (
      {stage1_11[183], stage1_11[184], stage1_11[185], stage1_11[186], stage1_11[187]},
      {stage1_12[88]},
      {stage1_13[162], stage1_13[163], stage1_13[164], stage1_13[165], stage1_13[166], stage1_13[167]},
      {stage2_15[27],stage2_14[40],stage2_13[43],stage2_12[61],stage2_11[81]}
   );
   gpc615_5 gpc4924 (
      {stage1_11[188], stage1_11[189], stage1_11[190], stage1_11[191], stage1_11[192]},
      {stage1_12[89]},
      {stage1_13[168], stage1_13[169], stage1_13[170], stage1_13[171], stage1_13[172], stage1_13[173]},
      {stage2_15[28],stage2_14[41],stage2_13[44],stage2_12[62],stage2_11[82]}
   );
   gpc615_5 gpc4925 (
      {stage1_11[193], stage1_11[194], stage1_11[195], stage1_11[196], stage1_11[197]},
      {stage1_12[90]},
      {stage1_13[174], stage1_13[175], stage1_13[176], stage1_13[177], stage1_13[178], stage1_13[179]},
      {stage2_15[29],stage2_14[42],stage2_13[45],stage2_12[63],stage2_11[83]}
   );
   gpc615_5 gpc4926 (
      {stage1_11[198], stage1_11[199], stage1_11[200], stage1_11[201], stage1_11[202]},
      {stage1_12[91]},
      {stage1_13[180], stage1_13[181], stage1_13[182], stage1_13[183], stage1_13[184], stage1_13[185]},
      {stage2_15[30],stage2_14[43],stage2_13[46],stage2_12[64],stage2_11[84]}
   );
   gpc615_5 gpc4927 (
      {stage1_11[203], stage1_11[204], stage1_11[205], stage1_11[206], stage1_11[207]},
      {stage1_12[92]},
      {stage1_13[186], stage1_13[187], stage1_13[188], stage1_13[189], stage1_13[190], stage1_13[191]},
      {stage2_15[31],stage2_14[44],stage2_13[47],stage2_12[65],stage2_11[85]}
   );
   gpc615_5 gpc4928 (
      {stage1_11[208], stage1_11[209], stage1_11[210], stage1_11[211], stage1_11[212]},
      {stage1_12[93]},
      {stage1_13[192], stage1_13[193], stage1_13[194], stage1_13[195], stage1_13[196], stage1_13[197]},
      {stage2_15[32],stage2_14[45],stage2_13[48],stage2_12[66],stage2_11[86]}
   );
   gpc615_5 gpc4929 (
      {stage1_11[213], stage1_11[214], stage1_11[215], stage1_11[216], stage1_11[217]},
      {stage1_12[94]},
      {stage1_13[198], stage1_13[199], stage1_13[200], stage1_13[201], stage1_13[202], stage1_13[203]},
      {stage2_15[33],stage2_14[46],stage2_13[49],stage2_12[67],stage2_11[87]}
   );
   gpc615_5 gpc4930 (
      {stage1_11[218], stage1_11[219], stage1_11[220], stage1_11[221], stage1_11[222]},
      {stage1_12[95]},
      {stage1_13[204], stage1_13[205], stage1_13[206], stage1_13[207], stage1_13[208], stage1_13[209]},
      {stage2_15[34],stage2_14[47],stage2_13[50],stage2_12[68],stage2_11[88]}
   );
   gpc1325_5 gpc4931 (
      {stage1_11[223], stage1_11[224], stage1_11[225], stage1_11[226], stage1_11[227]},
      {stage1_12[96], stage1_12[97]},
      {stage1_13[210], stage1_13[211], stage1_13[212]},
      {stage1_14[0]},
      {stage2_15[35],stage2_14[48],stage2_13[51],stage2_12[69],stage2_11[89]}
   );
   gpc2135_5 gpc4932 (
      {stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101], stage1_12[102]},
      {stage1_13[213], stage1_13[214], stage1_13[215]},
      {stage1_14[1]},
      {stage1_15[0], stage1_15[1]},
      {stage2_16[0],stage2_15[36],stage2_14[49],stage2_13[52],stage2_12[70]}
   );
   gpc606_5 gpc4933 (
      {stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107], stage1_12[108]},
      {stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6], stage1_14[7]},
      {stage2_16[1],stage2_15[37],stage2_14[50],stage2_13[53],stage2_12[71]}
   );
   gpc606_5 gpc4934 (
      {stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113], stage1_12[114]},
      {stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12], stage1_14[13]},
      {stage2_16[2],stage2_15[38],stage2_14[51],stage2_13[54],stage2_12[72]}
   );
   gpc606_5 gpc4935 (
      {stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119], stage1_12[120]},
      {stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18], stage1_14[19]},
      {stage2_16[3],stage2_15[39],stage2_14[52],stage2_13[55],stage2_12[73]}
   );
   gpc606_5 gpc4936 (
      {stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125], stage1_12[126]},
      {stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25]},
      {stage2_16[4],stage2_15[40],stage2_14[53],stage2_13[56],stage2_12[74]}
   );
   gpc606_5 gpc4937 (
      {stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131], stage1_12[132]},
      {stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31]},
      {stage2_16[5],stage2_15[41],stage2_14[54],stage2_13[57],stage2_12[75]}
   );
   gpc606_5 gpc4938 (
      {stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136], stage1_12[137], stage1_12[138]},
      {stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36], stage1_14[37]},
      {stage2_16[6],stage2_15[42],stage2_14[55],stage2_13[58],stage2_12[76]}
   );
   gpc606_5 gpc4939 (
      {stage1_12[139], stage1_12[140], stage1_12[141], stage1_12[142], stage1_12[143], stage1_12[144]},
      {stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42], stage1_14[43]},
      {stage2_16[7],stage2_15[43],stage2_14[56],stage2_13[59],stage2_12[77]}
   );
   gpc606_5 gpc4940 (
      {stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148], stage1_12[149], stage1_12[150]},
      {stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47], stage1_14[48], stage1_14[49]},
      {stage2_16[8],stage2_15[44],stage2_14[57],stage2_13[60],stage2_12[78]}
   );
   gpc606_5 gpc4941 (
      {stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154], stage1_12[155], stage1_12[156]},
      {stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53], stage1_14[54], stage1_14[55]},
      {stage2_16[9],stage2_15[45],stage2_14[58],stage2_13[61],stage2_12[79]}
   );
   gpc606_5 gpc4942 (
      {stage1_12[157], stage1_12[158], stage1_12[159], stage1_12[160], stage1_12[161], stage1_12[162]},
      {stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59], stage1_14[60], stage1_14[61]},
      {stage2_16[10],stage2_15[46],stage2_14[59],stage2_13[62],stage2_12[80]}
   );
   gpc606_5 gpc4943 (
      {stage1_13[216], stage1_13[217], stage1_13[218], stage1_13[219], stage1_13[220], stage1_13[221]},
      {stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5], stage1_15[6], stage1_15[7]},
      {stage2_17[0],stage2_16[11],stage2_15[47],stage2_14[60],stage2_13[63]}
   );
   gpc606_5 gpc4944 (
      {stage1_13[222], stage1_13[223], stage1_13[224], stage1_13[225], stage1_13[226], stage1_13[227]},
      {stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11], stage1_15[12], stage1_15[13]},
      {stage2_17[1],stage2_16[12],stage2_15[48],stage2_14[61],stage2_13[64]}
   );
   gpc606_5 gpc4945 (
      {stage1_13[228], stage1_13[229], stage1_13[230], stage1_13[231], stage1_13[232], stage1_13[233]},
      {stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19]},
      {stage2_17[2],stage2_16[13],stage2_15[49],stage2_14[62],stage2_13[65]}
   );
   gpc606_5 gpc4946 (
      {stage1_13[234], stage1_13[235], stage1_13[236], stage1_13[237], stage1_13[238], stage1_13[239]},
      {stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23], stage1_15[24], stage1_15[25]},
      {stage2_17[3],stage2_16[14],stage2_15[50],stage2_14[63],stage2_13[66]}
   );
   gpc606_5 gpc4947 (
      {stage1_13[240], stage1_13[241], stage1_13[242], stage1_13[243], stage1_13[244], stage1_13[245]},
      {stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31]},
      {stage2_17[4],stage2_16[15],stage2_15[51],stage2_14[64],stage2_13[67]}
   );
   gpc606_5 gpc4948 (
      {stage1_13[246], stage1_13[247], stage1_13[248], stage1_13[249], stage1_13[250], stage1_13[251]},
      {stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37]},
      {stage2_17[5],stage2_16[16],stage2_15[52],stage2_14[65],stage2_13[68]}
   );
   gpc606_5 gpc4949 (
      {stage1_13[252], stage1_13[253], stage1_13[254], stage1_13[255], stage1_13[256], stage1_13[257]},
      {stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43]},
      {stage2_17[6],stage2_16[17],stage2_15[53],stage2_14[66],stage2_13[69]}
   );
   gpc606_5 gpc4950 (
      {stage1_13[258], stage1_13[259], stage1_13[260], stage1_13[261], stage1_13[262], stage1_13[263]},
      {stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47], stage1_15[48], stage1_15[49]},
      {stage2_17[7],stage2_16[18],stage2_15[54],stage2_14[67],stage2_13[70]}
   );
   gpc606_5 gpc4951 (
      {stage1_13[264], stage1_13[265], stage1_13[266], stage1_13[267], stage1_13[268], stage1_13[269]},
      {stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53], stage1_15[54], stage1_15[55]},
      {stage2_17[8],stage2_16[19],stage2_15[55],stage2_14[68],stage2_13[71]}
   );
   gpc606_5 gpc4952 (
      {stage1_13[270], stage1_13[271], stage1_13[272], stage1_13[273], stage1_13[274], stage1_13[275]},
      {stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59], stage1_15[60], stage1_15[61]},
      {stage2_17[9],stage2_16[20],stage2_15[56],stage2_14[69],stage2_13[72]}
   );
   gpc606_5 gpc4953 (
      {stage1_13[276], stage1_13[277], stage1_13[278], stage1_13[279], stage1_13[280], stage1_13[281]},
      {stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65], stage1_15[66], stage1_15[67]},
      {stage2_17[10],stage2_16[21],stage2_15[57],stage2_14[70],stage2_13[73]}
   );
   gpc606_5 gpc4954 (
      {stage1_13[282], stage1_13[283], stage1_13[284], stage1_13[285], stage1_13[286], stage1_13[287]},
      {stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71], stage1_15[72], stage1_15[73]},
      {stage2_17[11],stage2_16[22],stage2_15[58],stage2_14[71],stage2_13[74]}
   );
   gpc606_5 gpc4955 (
      {stage1_13[288], stage1_13[289], stage1_13[290], stage1_13[291], stage1_13[292], stage1_13[293]},
      {stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77], stage1_15[78], stage1_15[79]},
      {stage2_17[12],stage2_16[23],stage2_15[59],stage2_14[72],stage2_13[75]}
   );
   gpc606_5 gpc4956 (
      {stage1_13[294], stage1_13[295], stage1_13[296], stage1_13[297], stage1_13[298], stage1_13[299]},
      {stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83], stage1_15[84], stage1_15[85]},
      {stage2_17[13],stage2_16[24],stage2_15[60],stage2_14[73],stage2_13[76]}
   );
   gpc606_5 gpc4957 (
      {stage1_13[300], stage1_13[301], stage1_13[302], stage1_13[303], stage1_13[304], 1'b0},
      {stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89], stage1_15[90], stage1_15[91]},
      {stage2_17[14],stage2_16[25],stage2_15[61],stage2_14[74],stage2_13[77]}
   );
   gpc615_5 gpc4958 (
      {stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65], stage1_14[66]},
      {stage1_15[92]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[15],stage2_16[26],stage2_15[62],stage2_14[75]}
   );
   gpc615_5 gpc4959 (
      {stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage1_15[93]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[16],stage2_16[27],stage2_15[63],stage2_14[76]}
   );
   gpc615_5 gpc4960 (
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76]},
      {stage1_15[94]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[17],stage2_16[28],stage2_15[64],stage2_14[77]}
   );
   gpc615_5 gpc4961 (
      {stage1_14[77], stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81]},
      {stage1_15[95]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[18],stage2_16[29],stage2_15[65],stage2_14[78]}
   );
   gpc615_5 gpc4962 (
      {stage1_14[82], stage1_14[83], stage1_14[84], stage1_14[85], stage1_14[86]},
      {stage1_15[96]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[19],stage2_16[30],stage2_15[66],stage2_14[79]}
   );
   gpc615_5 gpc4963 (
      {stage1_14[87], stage1_14[88], stage1_14[89], stage1_14[90], stage1_14[91]},
      {stage1_15[97]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[20],stage2_16[31],stage2_15[67],stage2_14[80]}
   );
   gpc615_5 gpc4964 (
      {stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95], stage1_14[96]},
      {stage1_15[98]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[21],stage2_16[32],stage2_15[68],stage2_14[81]}
   );
   gpc615_5 gpc4965 (
      {stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage1_15[99]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[22],stage2_16[33],stage2_15[69],stage2_14[82]}
   );
   gpc615_5 gpc4966 (
      {stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106]},
      {stage1_15[100]},
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage2_18[8],stage2_17[23],stage2_16[34],stage2_15[70],stage2_14[83]}
   );
   gpc615_5 gpc4967 (
      {stage1_14[107], stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111]},
      {stage1_15[101]},
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage2_18[9],stage2_17[24],stage2_16[35],stage2_15[71],stage2_14[84]}
   );
   gpc615_5 gpc4968 (
      {stage1_14[112], stage1_14[113], stage1_14[114], stage1_14[115], stage1_14[116]},
      {stage1_15[102]},
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65]},
      {stage2_18[10],stage2_17[25],stage2_16[36],stage2_15[72],stage2_14[85]}
   );
   gpc615_5 gpc4969 (
      {stage1_14[117], stage1_14[118], stage1_14[119], stage1_14[120], stage1_14[121]},
      {stage1_15[103]},
      {stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71]},
      {stage2_18[11],stage2_17[26],stage2_16[37],stage2_15[73],stage2_14[86]}
   );
   gpc615_5 gpc4970 (
      {stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125], stage1_14[126]},
      {stage1_15[104]},
      {stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77]},
      {stage2_18[12],stage2_17[27],stage2_16[38],stage2_15[74],stage2_14[87]}
   );
   gpc615_5 gpc4971 (
      {stage1_14[127], stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage1_15[105]},
      {stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83]},
      {stage2_18[13],stage2_17[28],stage2_16[39],stage2_15[75],stage2_14[88]}
   );
   gpc615_5 gpc4972 (
      {stage1_14[132], stage1_14[133], stage1_14[134], stage1_14[135], stage1_14[136]},
      {stage1_15[106]},
      {stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage2_18[14],stage2_17[29],stage2_16[40],stage2_15[76],stage2_14[89]}
   );
   gpc615_5 gpc4973 (
      {stage1_14[137], stage1_14[138], stage1_14[139], stage1_14[140], stage1_14[141]},
      {stage1_15[107]},
      {stage1_16[90], stage1_16[91], stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95]},
      {stage2_18[15],stage2_17[30],stage2_16[41],stage2_15[77],stage2_14[90]}
   );
   gpc615_5 gpc4974 (
      {stage1_14[142], stage1_14[143], stage1_14[144], stage1_14[145], stage1_14[146]},
      {stage1_15[108]},
      {stage1_16[96], stage1_16[97], stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101]},
      {stage2_18[16],stage2_17[31],stage2_16[42],stage2_15[78],stage2_14[91]}
   );
   gpc615_5 gpc4975 (
      {stage1_14[147], stage1_14[148], stage1_14[149], stage1_14[150], stage1_14[151]},
      {stage1_15[109]},
      {stage1_16[102], stage1_16[103], stage1_16[104], stage1_16[105], stage1_16[106], stage1_16[107]},
      {stage2_18[17],stage2_17[32],stage2_16[43],stage2_15[79],stage2_14[92]}
   );
   gpc615_5 gpc4976 (
      {stage1_14[152], stage1_14[153], stage1_14[154], stage1_14[155], stage1_14[156]},
      {stage1_15[110]},
      {stage1_16[108], stage1_16[109], stage1_16[110], stage1_16[111], stage1_16[112], stage1_16[113]},
      {stage2_18[18],stage2_17[33],stage2_16[44],stage2_15[80],stage2_14[93]}
   );
   gpc615_5 gpc4977 (
      {stage1_14[157], stage1_14[158], stage1_14[159], stage1_14[160], stage1_14[161]},
      {stage1_15[111]},
      {stage1_16[114], stage1_16[115], stage1_16[116], stage1_16[117], stage1_16[118], stage1_16[119]},
      {stage2_18[19],stage2_17[34],stage2_16[45],stage2_15[81],stage2_14[94]}
   );
   gpc615_5 gpc4978 (
      {stage1_14[162], stage1_14[163], stage1_14[164], stage1_14[165], stage1_14[166]},
      {stage1_15[112]},
      {stage1_16[120], stage1_16[121], stage1_16[122], stage1_16[123], stage1_16[124], stage1_16[125]},
      {stage2_18[20],stage2_17[35],stage2_16[46],stage2_15[82],stage2_14[95]}
   );
   gpc615_5 gpc4979 (
      {stage1_14[167], stage1_14[168], stage1_14[169], stage1_14[170], stage1_14[171]},
      {stage1_15[113]},
      {stage1_16[126], stage1_16[127], stage1_16[128], stage1_16[129], stage1_16[130], stage1_16[131]},
      {stage2_18[21],stage2_17[36],stage2_16[47],stage2_15[83],stage2_14[96]}
   );
   gpc615_5 gpc4980 (
      {stage1_14[172], stage1_14[173], stage1_14[174], stage1_14[175], stage1_14[176]},
      {stage1_15[114]},
      {stage1_16[132], stage1_16[133], stage1_16[134], stage1_16[135], stage1_16[136], stage1_16[137]},
      {stage2_18[22],stage2_17[37],stage2_16[48],stage2_15[84],stage2_14[97]}
   );
   gpc615_5 gpc4981 (
      {stage1_14[177], stage1_14[178], stage1_14[179], stage1_14[180], stage1_14[181]},
      {stage1_15[115]},
      {stage1_16[138], stage1_16[139], stage1_16[140], stage1_16[141], stage1_16[142], stage1_16[143]},
      {stage2_18[23],stage2_17[38],stage2_16[49],stage2_15[85],stage2_14[98]}
   );
   gpc615_5 gpc4982 (
      {stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185], stage1_14[186]},
      {stage1_15[116]},
      {stage1_16[144], stage1_16[145], stage1_16[146], stage1_16[147], stage1_16[148], stage1_16[149]},
      {stage2_18[24],stage2_17[39],stage2_16[50],stage2_15[86],stage2_14[99]}
   );
   gpc615_5 gpc4983 (
      {stage1_14[187], stage1_14[188], stage1_14[189], stage1_14[190], stage1_14[191]},
      {stage1_15[117]},
      {stage1_16[150], stage1_16[151], stage1_16[152], stage1_16[153], stage1_16[154], stage1_16[155]},
      {stage2_18[25],stage2_17[40],stage2_16[51],stage2_15[87],stage2_14[100]}
   );
   gpc615_5 gpc4984 (
      {stage1_14[192], stage1_14[193], stage1_14[194], stage1_14[195], stage1_14[196]},
      {stage1_15[118]},
      {stage1_16[156], stage1_16[157], stage1_16[158], stage1_16[159], stage1_16[160], stage1_16[161]},
      {stage2_18[26],stage2_17[41],stage2_16[52],stage2_15[88],stage2_14[101]}
   );
   gpc615_5 gpc4985 (
      {stage1_14[197], stage1_14[198], stage1_14[199], stage1_14[200], stage1_14[201]},
      {stage1_15[119]},
      {stage1_16[162], stage1_16[163], stage1_16[164], stage1_16[165], stage1_16[166], stage1_16[167]},
      {stage2_18[27],stage2_17[42],stage2_16[53],stage2_15[89],stage2_14[102]}
   );
   gpc615_5 gpc4986 (
      {stage1_14[202], stage1_14[203], stage1_14[204], stage1_14[205], stage1_14[206]},
      {stage1_15[120]},
      {stage1_16[168], stage1_16[169], stage1_16[170], stage1_16[171], stage1_16[172], stage1_16[173]},
      {stage2_18[28],stage2_17[43],stage2_16[54],stage2_15[90],stage2_14[103]}
   );
   gpc615_5 gpc4987 (
      {stage1_14[207], stage1_14[208], stage1_14[209], stage1_14[210], stage1_14[211]},
      {stage1_15[121]},
      {stage1_16[174], stage1_16[175], stage1_16[176], stage1_16[177], stage1_16[178], stage1_16[179]},
      {stage2_18[29],stage2_17[44],stage2_16[55],stage2_15[91],stage2_14[104]}
   );
   gpc615_5 gpc4988 (
      {stage1_14[212], stage1_14[213], stage1_14[214], stage1_14[215], stage1_14[216]},
      {stage1_15[122]},
      {stage1_16[180], stage1_16[181], stage1_16[182], stage1_16[183], stage1_16[184], stage1_16[185]},
      {stage2_18[30],stage2_17[45],stage2_16[56],stage2_15[92],stage2_14[105]}
   );
   gpc606_5 gpc4989 (
      {stage1_16[186], stage1_16[187], stage1_16[188], stage1_16[189], stage1_16[190], stage1_16[191]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[0],stage2_18[31],stage2_17[46],stage2_16[57]}
   );
   gpc606_5 gpc4990 (
      {stage1_16[192], stage1_16[193], stage1_16[194], stage1_16[195], stage1_16[196], stage1_16[197]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[1],stage2_18[32],stage2_17[47],stage2_16[58]}
   );
   gpc606_5 gpc4991 (
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[2],stage2_18[33],stage2_17[48]}
   );
   gpc606_5 gpc4992 (
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[3],stage2_19[3],stage2_18[34],stage2_17[49]}
   );
   gpc606_5 gpc4993 (
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[4],stage2_19[4],stage2_18[35],stage2_17[50]}
   );
   gpc606_5 gpc4994 (
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[5],stage2_19[5],stage2_18[36],stage2_17[51]}
   );
   gpc606_5 gpc4995 (
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[6],stage2_19[6],stage2_18[37],stage2_17[52]}
   );
   gpc606_5 gpc4996 (
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[7],stage2_19[7],stage2_18[38],stage2_17[53]}
   );
   gpc606_5 gpc4997 (
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[8],stage2_19[8],stage2_18[39],stage2_17[54]}
   );
   gpc606_5 gpc4998 (
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[9],stage2_19[9],stage2_18[40],stage2_17[55]}
   );
   gpc606_5 gpc4999 (
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[10],stage2_19[10],stage2_18[41],stage2_17[56]}
   );
   gpc606_5 gpc5000 (
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[11],stage2_19[11],stage2_18[42],stage2_17[57]}
   );
   gpc606_5 gpc5001 (
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[12],stage2_19[12],stage2_18[43],stage2_17[58]}
   );
   gpc606_5 gpc5002 (
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[13],stage2_19[13],stage2_18[44],stage2_17[59]}
   );
   gpc606_5 gpc5003 (
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage1_19[72], stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage2_21[12],stage2_20[14],stage2_19[14],stage2_18[45],stage2_17[60]}
   );
   gpc606_5 gpc5004 (
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82], stage1_19[83]},
      {stage2_21[13],stage2_20[15],stage2_19[15],stage2_18[46],stage2_17[61]}
   );
   gpc606_5 gpc5005 (
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87], stage1_19[88], stage1_19[89]},
      {stage2_21[14],stage2_20[16],stage2_19[16],stage2_18[47],stage2_17[62]}
   );
   gpc606_5 gpc5006 (
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93], stage1_19[94], stage1_19[95]},
      {stage2_21[15],stage2_20[17],stage2_19[17],stage2_18[48],stage2_17[63]}
   );
   gpc606_5 gpc5007 (
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage1_19[96], stage1_19[97], stage1_19[98], stage1_19[99], stage1_19[100], stage1_19[101]},
      {stage2_21[16],stage2_20[18],stage2_19[18],stage2_18[49],stage2_17[64]}
   );
   gpc606_5 gpc5008 (
      {stage1_17[102], stage1_17[103], stage1_17[104], stage1_17[105], stage1_17[106], stage1_17[107]},
      {stage1_19[102], stage1_19[103], stage1_19[104], stage1_19[105], stage1_19[106], stage1_19[107]},
      {stage2_21[17],stage2_20[19],stage2_19[19],stage2_18[50],stage2_17[65]}
   );
   gpc606_5 gpc5009 (
      {stage1_17[108], stage1_17[109], stage1_17[110], stage1_17[111], stage1_17[112], stage1_17[113]},
      {stage1_19[108], stage1_19[109], stage1_19[110], stage1_19[111], stage1_19[112], stage1_19[113]},
      {stage2_21[18],stage2_20[20],stage2_19[20],stage2_18[51],stage2_17[66]}
   );
   gpc606_5 gpc5010 (
      {stage1_17[114], stage1_17[115], stage1_17[116], stage1_17[117], stage1_17[118], stage1_17[119]},
      {stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117], stage1_19[118], stage1_19[119]},
      {stage2_21[19],stage2_20[21],stage2_19[21],stage2_18[52],stage2_17[67]}
   );
   gpc606_5 gpc5011 (
      {stage1_17[120], stage1_17[121], stage1_17[122], stage1_17[123], stage1_17[124], stage1_17[125]},
      {stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123], stage1_19[124], stage1_19[125]},
      {stage2_21[20],stage2_20[22],stage2_19[22],stage2_18[53],stage2_17[68]}
   );
   gpc606_5 gpc5012 (
      {stage1_17[126], stage1_17[127], stage1_17[128], stage1_17[129], stage1_17[130], stage1_17[131]},
      {stage1_19[126], stage1_19[127], stage1_19[128], stage1_19[129], stage1_19[130], stage1_19[131]},
      {stage2_21[21],stage2_20[23],stage2_19[23],stage2_18[54],stage2_17[69]}
   );
   gpc606_5 gpc5013 (
      {stage1_17[132], stage1_17[133], stage1_17[134], stage1_17[135], stage1_17[136], stage1_17[137]},
      {stage1_19[132], stage1_19[133], stage1_19[134], stage1_19[135], stage1_19[136], stage1_19[137]},
      {stage2_21[22],stage2_20[24],stage2_19[24],stage2_18[55],stage2_17[70]}
   );
   gpc606_5 gpc5014 (
      {stage1_17[138], stage1_17[139], stage1_17[140], stage1_17[141], stage1_17[142], stage1_17[143]},
      {stage1_19[138], stage1_19[139], stage1_19[140], stage1_19[141], stage1_19[142], stage1_19[143]},
      {stage2_21[23],stage2_20[25],stage2_19[25],stage2_18[56],stage2_17[71]}
   );
   gpc606_5 gpc5015 (
      {stage1_17[144], stage1_17[145], stage1_17[146], stage1_17[147], stage1_17[148], stage1_17[149]},
      {stage1_19[144], stage1_19[145], stage1_19[146], stage1_19[147], stage1_19[148], stage1_19[149]},
      {stage2_21[24],stage2_20[26],stage2_19[26],stage2_18[57],stage2_17[72]}
   );
   gpc606_5 gpc5016 (
      {stage1_17[150], stage1_17[151], stage1_17[152], stage1_17[153], stage1_17[154], stage1_17[155]},
      {stage1_19[150], stage1_19[151], stage1_19[152], stage1_19[153], stage1_19[154], stage1_19[155]},
      {stage2_21[25],stage2_20[27],stage2_19[27],stage2_18[58],stage2_17[73]}
   );
   gpc606_5 gpc5017 (
      {stage1_17[156], stage1_17[157], stage1_17[158], stage1_17[159], stage1_17[160], stage1_17[161]},
      {stage1_19[156], stage1_19[157], stage1_19[158], stage1_19[159], stage1_19[160], stage1_19[161]},
      {stage2_21[26],stage2_20[28],stage2_19[28],stage2_18[59],stage2_17[74]}
   );
   gpc606_5 gpc5018 (
      {stage1_17[162], stage1_17[163], stage1_17[164], stage1_17[165], stage1_17[166], stage1_17[167]},
      {stage1_19[162], stage1_19[163], stage1_19[164], stage1_19[165], stage1_19[166], stage1_19[167]},
      {stage2_21[27],stage2_20[29],stage2_19[29],stage2_18[60],stage2_17[75]}
   );
   gpc606_5 gpc5019 (
      {stage1_17[168], stage1_17[169], stage1_17[170], stage1_17[171], stage1_17[172], stage1_17[173]},
      {stage1_19[168], stage1_19[169], stage1_19[170], stage1_19[171], stage1_19[172], stage1_19[173]},
      {stage2_21[28],stage2_20[30],stage2_19[30],stage2_18[61],stage2_17[76]}
   );
   gpc606_5 gpc5020 (
      {stage1_17[174], stage1_17[175], stage1_17[176], stage1_17[177], stage1_17[178], stage1_17[179]},
      {stage1_19[174], stage1_19[175], stage1_19[176], stage1_19[177], stage1_19[178], stage1_19[179]},
      {stage2_21[29],stage2_20[31],stage2_19[31],stage2_18[62],stage2_17[77]}
   );
   gpc606_5 gpc5021 (
      {stage1_17[180], stage1_17[181], stage1_17[182], stage1_17[183], stage1_17[184], stage1_17[185]},
      {stage1_19[180], stage1_19[181], stage1_19[182], stage1_19[183], stage1_19[184], stage1_19[185]},
      {stage2_21[30],stage2_20[32],stage2_19[32],stage2_18[63],stage2_17[78]}
   );
   gpc606_5 gpc5022 (
      {stage1_17[186], stage1_17[187], stage1_17[188], stage1_17[189], stage1_17[190], stage1_17[191]},
      {stage1_19[186], stage1_19[187], stage1_19[188], stage1_19[189], stage1_19[190], stage1_19[191]},
      {stage2_21[31],stage2_20[33],stage2_19[33],stage2_18[64],stage2_17[79]}
   );
   gpc606_5 gpc5023 (
      {stage1_17[192], stage1_17[193], stage1_17[194], stage1_17[195], stage1_17[196], stage1_17[197]},
      {stage1_19[192], stage1_19[193], stage1_19[194], stage1_19[195], stage1_19[196], stage1_19[197]},
      {stage2_21[32],stage2_20[34],stage2_19[34],stage2_18[65],stage2_17[80]}
   );
   gpc606_5 gpc5024 (
      {stage1_17[198], stage1_17[199], stage1_17[200], stage1_17[201], stage1_17[202], stage1_17[203]},
      {stage1_19[198], stage1_19[199], stage1_19[200], stage1_19[201], stage1_19[202], stage1_19[203]},
      {stage2_21[33],stage2_20[35],stage2_19[35],stage2_18[66],stage2_17[81]}
   );
   gpc606_5 gpc5025 (
      {stage1_17[204], stage1_17[205], stage1_17[206], stage1_17[207], stage1_17[208], stage1_17[209]},
      {stage1_19[204], stage1_19[205], stage1_19[206], stage1_19[207], stage1_19[208], stage1_19[209]},
      {stage2_21[34],stage2_20[36],stage2_19[36],stage2_18[67],stage2_17[82]}
   );
   gpc606_5 gpc5026 (
      {stage1_17[210], stage1_17[211], stage1_17[212], stage1_17[213], stage1_17[214], stage1_17[215]},
      {stage1_19[210], stage1_19[211], stage1_19[212], stage1_19[213], stage1_19[214], stage1_19[215]},
      {stage2_21[35],stage2_20[37],stage2_19[37],stage2_18[68],stage2_17[83]}
   );
   gpc606_5 gpc5027 (
      {stage1_17[216], stage1_17[217], stage1_17[218], stage1_17[219], stage1_17[220], stage1_17[221]},
      {stage1_19[216], stage1_19[217], stage1_19[218], stage1_19[219], stage1_19[220], stage1_19[221]},
      {stage2_21[36],stage2_20[38],stage2_19[38],stage2_18[69],stage2_17[84]}
   );
   gpc606_5 gpc5028 (
      {stage1_17[222], stage1_17[223], stage1_17[224], stage1_17[225], stage1_17[226], stage1_17[227]},
      {stage1_19[222], stage1_19[223], stage1_19[224], stage1_19[225], stage1_19[226], stage1_19[227]},
      {stage2_21[37],stage2_20[39],stage2_19[39],stage2_18[70],stage2_17[85]}
   );
   gpc606_5 gpc5029 (
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[38],stage2_20[40],stage2_19[40],stage2_18[71]}
   );
   gpc606_5 gpc5030 (
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[39],stage2_20[41],stage2_19[41],stage2_18[72]}
   );
   gpc606_5 gpc5031 (
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[40],stage2_20[42],stage2_19[42],stage2_18[73]}
   );
   gpc606_5 gpc5032 (
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage2_22[3],stage2_21[41],stage2_20[43],stage2_19[43],stage2_18[74]}
   );
   gpc606_5 gpc5033 (
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27], stage1_20[28], stage1_20[29]},
      {stage2_22[4],stage2_21[42],stage2_20[44],stage2_19[44],stage2_18[75]}
   );
   gpc606_5 gpc5034 (
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage1_20[30], stage1_20[31], stage1_20[32], stage1_20[33], stage1_20[34], stage1_20[35]},
      {stage2_22[5],stage2_21[43],stage2_20[45],stage2_19[45],stage2_18[76]}
   );
   gpc606_5 gpc5035 (
      {stage1_18[48], stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53]},
      {stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39], stage1_20[40], stage1_20[41]},
      {stage2_22[6],stage2_21[44],stage2_20[46],stage2_19[46],stage2_18[77]}
   );
   gpc606_5 gpc5036 (
      {stage1_18[54], stage1_18[55], stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59]},
      {stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46], stage1_20[47]},
      {stage2_22[7],stage2_21[45],stage2_20[47],stage2_19[47],stage2_18[78]}
   );
   gpc606_5 gpc5037 (
      {stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51], stage1_20[52], stage1_20[53]},
      {stage2_22[8],stage2_21[46],stage2_20[48],stage2_19[48],stage2_18[79]}
   );
   gpc606_5 gpc5038 (
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71]},
      {stage1_20[54], stage1_20[55], stage1_20[56], stage1_20[57], stage1_20[58], stage1_20[59]},
      {stage2_22[9],stage2_21[47],stage2_20[49],stage2_19[49],stage2_18[80]}
   );
   gpc606_5 gpc5039 (
      {stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77]},
      {stage1_20[60], stage1_20[61], stage1_20[62], stage1_20[63], stage1_20[64], stage1_20[65]},
      {stage2_22[10],stage2_21[48],stage2_20[50],stage2_19[50],stage2_18[81]}
   );
   gpc606_5 gpc5040 (
      {stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage1_20[66], stage1_20[67], stage1_20[68], stage1_20[69], stage1_20[70], stage1_20[71]},
      {stage2_22[11],stage2_21[49],stage2_20[51],stage2_19[51],stage2_18[82]}
   );
   gpc606_5 gpc5041 (
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88], stage1_18[89]},
      {stage1_20[72], stage1_20[73], stage1_20[74], stage1_20[75], stage1_20[76], stage1_20[77]},
      {stage2_22[12],stage2_21[50],stage2_20[52],stage2_19[52],stage2_18[83]}
   );
   gpc606_5 gpc5042 (
      {stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93], stage1_18[94], stage1_18[95]},
      {stage1_20[78], stage1_20[79], stage1_20[80], stage1_20[81], stage1_20[82], stage1_20[83]},
      {stage2_22[13],stage2_21[51],stage2_20[53],stage2_19[53],stage2_18[84]}
   );
   gpc606_5 gpc5043 (
      {stage1_18[96], stage1_18[97], stage1_18[98], stage1_18[99], stage1_18[100], stage1_18[101]},
      {stage1_20[84], stage1_20[85], stage1_20[86], stage1_20[87], stage1_20[88], stage1_20[89]},
      {stage2_22[14],stage2_21[52],stage2_20[54],stage2_19[54],stage2_18[85]}
   );
   gpc606_5 gpc5044 (
      {stage1_18[102], stage1_18[103], stage1_18[104], stage1_18[105], stage1_18[106], stage1_18[107]},
      {stage1_20[90], stage1_20[91], stage1_20[92], stage1_20[93], stage1_20[94], stage1_20[95]},
      {stage2_22[15],stage2_21[53],stage2_20[55],stage2_19[55],stage2_18[86]}
   );
   gpc606_5 gpc5045 (
      {stage1_18[108], stage1_18[109], stage1_18[110], stage1_18[111], stage1_18[112], stage1_18[113]},
      {stage1_20[96], stage1_20[97], stage1_20[98], stage1_20[99], stage1_20[100], stage1_20[101]},
      {stage2_22[16],stage2_21[54],stage2_20[56],stage2_19[56],stage2_18[87]}
   );
   gpc606_5 gpc5046 (
      {stage1_18[114], stage1_18[115], stage1_18[116], stage1_18[117], stage1_18[118], stage1_18[119]},
      {stage1_20[102], stage1_20[103], stage1_20[104], stage1_20[105], stage1_20[106], stage1_20[107]},
      {stage2_22[17],stage2_21[55],stage2_20[57],stage2_19[57],stage2_18[88]}
   );
   gpc606_5 gpc5047 (
      {stage1_18[120], stage1_18[121], stage1_18[122], stage1_18[123], stage1_18[124], stage1_18[125]},
      {stage1_20[108], stage1_20[109], stage1_20[110], stage1_20[111], stage1_20[112], stage1_20[113]},
      {stage2_22[18],stage2_21[56],stage2_20[58],stage2_19[58],stage2_18[89]}
   );
   gpc606_5 gpc5048 (
      {stage1_18[126], stage1_18[127], stage1_18[128], stage1_18[129], stage1_18[130], stage1_18[131]},
      {stage1_20[114], stage1_20[115], stage1_20[116], stage1_20[117], stage1_20[118], stage1_20[119]},
      {stage2_22[19],stage2_21[57],stage2_20[59],stage2_19[59],stage2_18[90]}
   );
   gpc606_5 gpc5049 (
      {stage1_18[132], stage1_18[133], stage1_18[134], stage1_18[135], stage1_18[136], stage1_18[137]},
      {stage1_20[120], stage1_20[121], stage1_20[122], stage1_20[123], stage1_20[124], stage1_20[125]},
      {stage2_22[20],stage2_21[58],stage2_20[60],stage2_19[60],stage2_18[91]}
   );
   gpc606_5 gpc5050 (
      {stage1_18[138], stage1_18[139], stage1_18[140], stage1_18[141], stage1_18[142], stage1_18[143]},
      {stage1_20[126], stage1_20[127], stage1_20[128], stage1_20[129], stage1_20[130], stage1_20[131]},
      {stage2_22[21],stage2_21[59],stage2_20[61],stage2_19[61],stage2_18[92]}
   );
   gpc606_5 gpc5051 (
      {stage1_18[144], stage1_18[145], stage1_18[146], stage1_18[147], stage1_18[148], stage1_18[149]},
      {stage1_20[132], stage1_20[133], stage1_20[134], stage1_20[135], stage1_20[136], stage1_20[137]},
      {stage2_22[22],stage2_21[60],stage2_20[62],stage2_19[62],stage2_18[93]}
   );
   gpc606_5 gpc5052 (
      {stage1_18[150], stage1_18[151], stage1_18[152], stage1_18[153], stage1_18[154], stage1_18[155]},
      {stage1_20[138], stage1_20[139], stage1_20[140], stage1_20[141], stage1_20[142], stage1_20[143]},
      {stage2_22[23],stage2_21[61],stage2_20[63],stage2_19[63],stage2_18[94]}
   );
   gpc606_5 gpc5053 (
      {stage1_18[156], stage1_18[157], stage1_18[158], stage1_18[159], stage1_18[160], stage1_18[161]},
      {stage1_20[144], stage1_20[145], stage1_20[146], stage1_20[147], stage1_20[148], stage1_20[149]},
      {stage2_22[24],stage2_21[62],stage2_20[64],stage2_19[64],stage2_18[95]}
   );
   gpc606_5 gpc5054 (
      {stage1_18[162], stage1_18[163], stage1_18[164], stage1_18[165], stage1_18[166], stage1_18[167]},
      {stage1_20[150], stage1_20[151], stage1_20[152], stage1_20[153], stage1_20[154], stage1_20[155]},
      {stage2_22[25],stage2_21[63],stage2_20[65],stage2_19[65],stage2_18[96]}
   );
   gpc606_5 gpc5055 (
      {stage1_18[168], stage1_18[169], stage1_18[170], stage1_18[171], stage1_18[172], stage1_18[173]},
      {stage1_20[156], stage1_20[157], stage1_20[158], stage1_20[159], stage1_20[160], stage1_20[161]},
      {stage2_22[26],stage2_21[64],stage2_20[66],stage2_19[66],stage2_18[97]}
   );
   gpc606_5 gpc5056 (
      {stage1_18[174], stage1_18[175], stage1_18[176], stage1_18[177], stage1_18[178], stage1_18[179]},
      {stage1_20[162], stage1_20[163], stage1_20[164], stage1_20[165], stage1_20[166], stage1_20[167]},
      {stage2_22[27],stage2_21[65],stage2_20[67],stage2_19[67],stage2_18[98]}
   );
   gpc606_5 gpc5057 (
      {stage1_18[180], stage1_18[181], stage1_18[182], stage1_18[183], stage1_18[184], stage1_18[185]},
      {stage1_20[168], stage1_20[169], stage1_20[170], stage1_20[171], stage1_20[172], stage1_20[173]},
      {stage2_22[28],stage2_21[66],stage2_20[68],stage2_19[68],stage2_18[99]}
   );
   gpc615_5 gpc5058 (
      {stage1_18[186], stage1_18[187], stage1_18[188], stage1_18[189], stage1_18[190]},
      {stage1_19[228]},
      {stage1_20[174], stage1_20[175], stage1_20[176], stage1_20[177], stage1_20[178], stage1_20[179]},
      {stage2_22[29],stage2_21[67],stage2_20[69],stage2_19[69],stage2_18[100]}
   );
   gpc615_5 gpc5059 (
      {stage1_19[229], stage1_19[230], stage1_19[231], stage1_19[232], stage1_19[233]},
      {stage1_20[180]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[30],stage2_21[68],stage2_20[70],stage2_19[70]}
   );
   gpc606_5 gpc5060 (
      {stage1_20[181], stage1_20[182], stage1_20[183], stage1_20[184], stage1_20[185], stage1_20[186]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[1],stage2_22[31],stage2_21[69],stage2_20[71]}
   );
   gpc615_5 gpc5061 (
      {stage1_20[187], stage1_20[188], stage1_20[189], stage1_20[190], stage1_20[191]},
      {stage1_21[6]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[2],stage2_22[32],stage2_21[70],stage2_20[72]}
   );
   gpc615_5 gpc5062 (
      {stage1_20[192], stage1_20[193], stage1_20[194], stage1_20[195], stage1_20[196]},
      {stage1_21[7]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[3],stage2_22[33],stage2_21[71],stage2_20[73]}
   );
   gpc615_5 gpc5063 (
      {stage1_20[197], stage1_20[198], stage1_20[199], stage1_20[200], stage1_20[201]},
      {stage1_21[8]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[4],stage2_22[34],stage2_21[72],stage2_20[74]}
   );
   gpc615_5 gpc5064 (
      {stage1_20[202], stage1_20[203], stage1_20[204], stage1_20[205], stage1_20[206]},
      {stage1_21[9]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[5],stage2_22[35],stage2_21[73],stage2_20[75]}
   );
   gpc615_5 gpc5065 (
      {stage1_20[207], stage1_20[208], stage1_20[209], stage1_20[210], stage1_20[211]},
      {stage1_21[10]},
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage2_24[5],stage2_23[6],stage2_22[36],stage2_21[74],stage2_20[76]}
   );
   gpc615_5 gpc5066 (
      {stage1_20[212], stage1_20[213], stage1_20[214], stage1_20[215], stage1_20[216]},
      {stage1_21[11]},
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage2_24[6],stage2_23[7],stage2_22[37],stage2_21[75],stage2_20[77]}
   );
   gpc615_5 gpc5067 (
      {stage1_20[217], stage1_20[218], stage1_20[219], stage1_20[220], stage1_20[221]},
      {stage1_21[12]},
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage2_24[7],stage2_23[8],stage2_22[38],stage2_21[76],stage2_20[78]}
   );
   gpc615_5 gpc5068 (
      {stage1_20[222], stage1_20[223], stage1_20[224], stage1_20[225], stage1_20[226]},
      {stage1_21[13]},
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage2_24[8],stage2_23[9],stage2_22[39],stage2_21[77],stage2_20[79]}
   );
   gpc615_5 gpc5069 (
      {stage1_20[227], stage1_20[228], stage1_20[229], stage1_20[230], stage1_20[231]},
      {stage1_21[14]},
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage2_24[9],stage2_23[10],stage2_22[40],stage2_21[78],stage2_20[80]}
   );
   gpc615_5 gpc5070 (
      {stage1_20[232], stage1_20[233], stage1_20[234], stage1_20[235], stage1_20[236]},
      {stage1_21[15]},
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage2_24[10],stage2_23[11],stage2_22[41],stage2_21[79],stage2_20[81]}
   );
   gpc615_5 gpc5071 (
      {stage1_20[237], stage1_20[238], stage1_20[239], stage1_20[240], stage1_20[241]},
      {stage1_21[16]},
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage2_24[11],stage2_23[12],stage2_22[42],stage2_21[80],stage2_20[82]}
   );
   gpc615_5 gpc5072 (
      {stage1_20[242], stage1_20[243], stage1_20[244], stage1_20[245], stage1_20[246]},
      {stage1_21[17]},
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77]},
      {stage2_24[12],stage2_23[13],stage2_22[43],stage2_21[81],stage2_20[83]}
   );
   gpc615_5 gpc5073 (
      {stage1_20[247], stage1_20[248], stage1_20[249], stage1_20[250], stage1_20[251]},
      {stage1_21[18]},
      {stage1_22[78], stage1_22[79], stage1_22[80], stage1_22[81], stage1_22[82], stage1_22[83]},
      {stage2_24[13],stage2_23[14],stage2_22[44],stage2_21[82],stage2_20[84]}
   );
   gpc615_5 gpc5074 (
      {stage1_20[252], stage1_20[253], stage1_20[254], stage1_20[255], stage1_20[256]},
      {stage1_21[19]},
      {stage1_22[84], stage1_22[85], stage1_22[86], stage1_22[87], stage1_22[88], stage1_22[89]},
      {stage2_24[14],stage2_23[15],stage2_22[45],stage2_21[83],stage2_20[85]}
   );
   gpc615_5 gpc5075 (
      {stage1_20[257], stage1_20[258], stage1_20[259], stage1_20[260], stage1_20[261]},
      {stage1_21[20]},
      {stage1_22[90], stage1_22[91], stage1_22[92], stage1_22[93], stage1_22[94], stage1_22[95]},
      {stage2_24[15],stage2_23[16],stage2_22[46],stage2_21[84],stage2_20[86]}
   );
   gpc606_5 gpc5076 (
      {stage1_21[21], stage1_21[22], stage1_21[23], stage1_21[24], stage1_21[25], stage1_21[26]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[16],stage2_23[17],stage2_22[47],stage2_21[85]}
   );
   gpc606_5 gpc5077 (
      {stage1_21[27], stage1_21[28], stage1_21[29], stage1_21[30], stage1_21[31], stage1_21[32]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[17],stage2_23[18],stage2_22[48],stage2_21[86]}
   );
   gpc606_5 gpc5078 (
      {stage1_21[33], stage1_21[34], stage1_21[35], stage1_21[36], stage1_21[37], stage1_21[38]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[18],stage2_23[19],stage2_22[49],stage2_21[87]}
   );
   gpc606_5 gpc5079 (
      {stage1_21[39], stage1_21[40], stage1_21[41], stage1_21[42], stage1_21[43], stage1_21[44]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[19],stage2_23[20],stage2_22[50],stage2_21[88]}
   );
   gpc606_5 gpc5080 (
      {stage1_21[45], stage1_21[46], stage1_21[47], stage1_21[48], stage1_21[49], stage1_21[50]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[20],stage2_23[21],stage2_22[51],stage2_21[89]}
   );
   gpc606_5 gpc5081 (
      {stage1_21[51], stage1_21[52], stage1_21[53], stage1_21[54], stage1_21[55], stage1_21[56]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage2_25[5],stage2_24[21],stage2_23[22],stage2_22[52],stage2_21[90]}
   );
   gpc606_5 gpc5082 (
      {stage1_21[57], stage1_21[58], stage1_21[59], stage1_21[60], stage1_21[61], stage1_21[62]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage2_25[6],stage2_24[22],stage2_23[23],stage2_22[53],stage2_21[91]}
   );
   gpc606_5 gpc5083 (
      {stage1_21[63], stage1_21[64], stage1_21[65], stage1_21[66], stage1_21[67], stage1_21[68]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage2_25[7],stage2_24[23],stage2_23[24],stage2_22[54],stage2_21[92]}
   );
   gpc606_5 gpc5084 (
      {stage1_21[69], stage1_21[70], stage1_21[71], stage1_21[72], stage1_21[73], stage1_21[74]},
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage2_25[8],stage2_24[24],stage2_23[25],stage2_22[55],stage2_21[93]}
   );
   gpc606_5 gpc5085 (
      {stage1_21[75], stage1_21[76], stage1_21[77], stage1_21[78], stage1_21[79], stage1_21[80]},
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage2_25[9],stage2_24[25],stage2_23[26],stage2_22[56],stage2_21[94]}
   );
   gpc606_5 gpc5086 (
      {stage1_21[81], stage1_21[82], stage1_21[83], stage1_21[84], stage1_21[85], stage1_21[86]},
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage2_25[10],stage2_24[26],stage2_23[27],stage2_22[57],stage2_21[95]}
   );
   gpc606_5 gpc5087 (
      {stage1_21[87], stage1_21[88], stage1_21[89], stage1_21[90], stage1_21[91], stage1_21[92]},
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage2_25[11],stage2_24[27],stage2_23[28],stage2_22[58],stage2_21[96]}
   );
   gpc606_5 gpc5088 (
      {stage1_21[93], stage1_21[94], stage1_21[95], stage1_21[96], stage1_21[97], stage1_21[98]},
      {stage1_23[72], stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage2_25[12],stage2_24[28],stage2_23[29],stage2_22[59],stage2_21[97]}
   );
   gpc606_5 gpc5089 (
      {stage1_21[99], stage1_21[100], stage1_21[101], stage1_21[102], stage1_21[103], stage1_21[104]},
      {stage1_23[78], stage1_23[79], stage1_23[80], stage1_23[81], stage1_23[82], stage1_23[83]},
      {stage2_25[13],stage2_24[29],stage2_23[30],stage2_22[60],stage2_21[98]}
   );
   gpc606_5 gpc5090 (
      {stage1_21[105], stage1_21[106], stage1_21[107], stage1_21[108], stage1_21[109], stage1_21[110]},
      {stage1_23[84], stage1_23[85], stage1_23[86], stage1_23[87], stage1_23[88], stage1_23[89]},
      {stage2_25[14],stage2_24[30],stage2_23[31],stage2_22[61],stage2_21[99]}
   );
   gpc606_5 gpc5091 (
      {stage1_21[111], stage1_21[112], stage1_21[113], stage1_21[114], stage1_21[115], stage1_21[116]},
      {stage1_23[90], stage1_23[91], stage1_23[92], stage1_23[93], stage1_23[94], stage1_23[95]},
      {stage2_25[15],stage2_24[31],stage2_23[32],stage2_22[62],stage2_21[100]}
   );
   gpc606_5 gpc5092 (
      {stage1_21[117], stage1_21[118], stage1_21[119], stage1_21[120], stage1_21[121], stage1_21[122]},
      {stage1_23[96], stage1_23[97], stage1_23[98], stage1_23[99], stage1_23[100], stage1_23[101]},
      {stage2_25[16],stage2_24[32],stage2_23[33],stage2_22[63],stage2_21[101]}
   );
   gpc606_5 gpc5093 (
      {stage1_21[123], stage1_21[124], stage1_21[125], stage1_21[126], stage1_21[127], stage1_21[128]},
      {stage1_23[102], stage1_23[103], stage1_23[104], stage1_23[105], stage1_23[106], stage1_23[107]},
      {stage2_25[17],stage2_24[33],stage2_23[34],stage2_22[64],stage2_21[102]}
   );
   gpc615_5 gpc5094 (
      {stage1_21[129], stage1_21[130], stage1_21[131], stage1_21[132], stage1_21[133]},
      {stage1_22[96]},
      {stage1_23[108], stage1_23[109], stage1_23[110], stage1_23[111], stage1_23[112], stage1_23[113]},
      {stage2_25[18],stage2_24[34],stage2_23[35],stage2_22[65],stage2_21[103]}
   );
   gpc615_5 gpc5095 (
      {stage1_21[134], stage1_21[135], stage1_21[136], stage1_21[137], stage1_21[138]},
      {stage1_22[97]},
      {stage1_23[114], stage1_23[115], stage1_23[116], stage1_23[117], stage1_23[118], stage1_23[119]},
      {stage2_25[19],stage2_24[35],stage2_23[36],stage2_22[66],stage2_21[104]}
   );
   gpc615_5 gpc5096 (
      {stage1_21[139], stage1_21[140], stage1_21[141], stage1_21[142], stage1_21[143]},
      {stage1_22[98]},
      {stage1_23[120], stage1_23[121], stage1_23[122], stage1_23[123], stage1_23[124], stage1_23[125]},
      {stage2_25[20],stage2_24[36],stage2_23[37],stage2_22[67],stage2_21[105]}
   );
   gpc615_5 gpc5097 (
      {stage1_21[144], stage1_21[145], stage1_21[146], stage1_21[147], stage1_21[148]},
      {stage1_22[99]},
      {stage1_23[126], stage1_23[127], stage1_23[128], stage1_23[129], stage1_23[130], stage1_23[131]},
      {stage2_25[21],stage2_24[37],stage2_23[38],stage2_22[68],stage2_21[106]}
   );
   gpc615_5 gpc5098 (
      {stage1_21[149], stage1_21[150], stage1_21[151], stage1_21[152], stage1_21[153]},
      {stage1_22[100]},
      {stage1_23[132], stage1_23[133], stage1_23[134], stage1_23[135], stage1_23[136], stage1_23[137]},
      {stage2_25[22],stage2_24[38],stage2_23[39],stage2_22[69],stage2_21[107]}
   );
   gpc615_5 gpc5099 (
      {stage1_21[154], stage1_21[155], stage1_21[156], stage1_21[157], stage1_21[158]},
      {stage1_22[101]},
      {stage1_23[138], stage1_23[139], stage1_23[140], stage1_23[141], stage1_23[142], stage1_23[143]},
      {stage2_25[23],stage2_24[39],stage2_23[40],stage2_22[70],stage2_21[108]}
   );
   gpc615_5 gpc5100 (
      {stage1_21[159], stage1_21[160], stage1_21[161], stage1_21[162], stage1_21[163]},
      {stage1_22[102]},
      {stage1_23[144], stage1_23[145], stage1_23[146], stage1_23[147], stage1_23[148], stage1_23[149]},
      {stage2_25[24],stage2_24[40],stage2_23[41],stage2_22[71],stage2_21[109]}
   );
   gpc615_5 gpc5101 (
      {stage1_21[164], stage1_21[165], stage1_21[166], stage1_21[167], stage1_21[168]},
      {stage1_22[103]},
      {stage1_23[150], stage1_23[151], stage1_23[152], stage1_23[153], stage1_23[154], stage1_23[155]},
      {stage2_25[25],stage2_24[41],stage2_23[42],stage2_22[72],stage2_21[110]}
   );
   gpc615_5 gpc5102 (
      {stage1_21[169], stage1_21[170], stage1_21[171], stage1_21[172], stage1_21[173]},
      {stage1_22[104]},
      {stage1_23[156], stage1_23[157], stage1_23[158], stage1_23[159], stage1_23[160], stage1_23[161]},
      {stage2_25[26],stage2_24[42],stage2_23[43],stage2_22[73],stage2_21[111]}
   );
   gpc615_5 gpc5103 (
      {stage1_22[105], stage1_22[106], stage1_22[107], stage1_22[108], stage1_22[109]},
      {stage1_23[162]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[27],stage2_24[43],stage2_23[44],stage2_22[74]}
   );
   gpc615_5 gpc5104 (
      {stage1_22[110], stage1_22[111], stage1_22[112], stage1_22[113], stage1_22[114]},
      {stage1_23[163]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[28],stage2_24[44],stage2_23[45],stage2_22[75]}
   );
   gpc615_5 gpc5105 (
      {stage1_22[115], stage1_22[116], stage1_22[117], stage1_22[118], stage1_22[119]},
      {stage1_23[164]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[29],stage2_24[45],stage2_23[46],stage2_22[76]}
   );
   gpc615_5 gpc5106 (
      {stage1_22[120], stage1_22[121], stage1_22[122], stage1_22[123], stage1_22[124]},
      {stage1_23[165]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[30],stage2_24[46],stage2_23[47],stage2_22[77]}
   );
   gpc615_5 gpc5107 (
      {stage1_22[125], stage1_22[126], stage1_22[127], stage1_22[128], stage1_22[129]},
      {stage1_23[166]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[31],stage2_24[47],stage2_23[48],stage2_22[78]}
   );
   gpc615_5 gpc5108 (
      {stage1_22[130], stage1_22[131], stage1_22[132], stage1_22[133], stage1_22[134]},
      {stage1_23[167]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[32],stage2_24[48],stage2_23[49],stage2_22[79]}
   );
   gpc615_5 gpc5109 (
      {stage1_22[135], stage1_22[136], stage1_22[137], stage1_22[138], stage1_22[139]},
      {stage1_23[168]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[33],stage2_24[49],stage2_23[50],stage2_22[80]}
   );
   gpc615_5 gpc5110 (
      {stage1_22[140], stage1_22[141], stage1_22[142], stage1_22[143], stage1_22[144]},
      {stage1_23[169]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[34],stage2_24[50],stage2_23[51],stage2_22[81]}
   );
   gpc615_5 gpc5111 (
      {stage1_23[170], stage1_23[171], stage1_23[172], stage1_23[173], stage1_23[174]},
      {stage1_24[48]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[8],stage2_25[35],stage2_24[51],stage2_23[52]}
   );
   gpc615_5 gpc5112 (
      {stage1_23[175], stage1_23[176], stage1_23[177], stage1_23[178], stage1_23[179]},
      {stage1_24[49]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[9],stage2_25[36],stage2_24[52],stage2_23[53]}
   );
   gpc615_5 gpc5113 (
      {stage1_23[180], stage1_23[181], stage1_23[182], stage1_23[183], stage1_23[184]},
      {stage1_24[50]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[10],stage2_25[37],stage2_24[53],stage2_23[54]}
   );
   gpc615_5 gpc5114 (
      {stage1_23[185], stage1_23[186], stage1_23[187], stage1_23[188], stage1_23[189]},
      {stage1_24[51]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[11],stage2_25[38],stage2_24[54],stage2_23[55]}
   );
   gpc615_5 gpc5115 (
      {stage1_23[190], stage1_23[191], stage1_23[192], stage1_23[193], stage1_23[194]},
      {stage1_24[52]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[12],stage2_25[39],stage2_24[55],stage2_23[56]}
   );
   gpc615_5 gpc5116 (
      {stage1_23[195], stage1_23[196], stage1_23[197], stage1_23[198], stage1_23[199]},
      {stage1_24[53]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[13],stage2_25[40],stage2_24[56],stage2_23[57]}
   );
   gpc615_5 gpc5117 (
      {stage1_23[200], stage1_23[201], stage1_23[202], stage1_23[203], stage1_23[204]},
      {stage1_24[54]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[14],stage2_25[41],stage2_24[57],stage2_23[58]}
   );
   gpc615_5 gpc5118 (
      {stage1_23[205], stage1_23[206], stage1_23[207], stage1_23[208], stage1_23[209]},
      {stage1_24[55]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[15],stage2_25[42],stage2_24[58],stage2_23[59]}
   );
   gpc615_5 gpc5119 (
      {stage1_23[210], stage1_23[211], stage1_23[212], stage1_23[213], stage1_23[214]},
      {stage1_24[56]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage2_27[8],stage2_26[16],stage2_25[43],stage2_24[59],stage2_23[60]}
   );
   gpc615_5 gpc5120 (
      {stage1_23[215], stage1_23[216], stage1_23[217], stage1_23[218], stage1_23[219]},
      {stage1_24[57]},
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage2_27[9],stage2_26[17],stage2_25[44],stage2_24[60],stage2_23[61]}
   );
   gpc615_5 gpc5121 (
      {stage1_23[220], stage1_23[221], stage1_23[222], stage1_23[223], stage1_23[224]},
      {stage1_24[58]},
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage2_27[10],stage2_26[18],stage2_25[45],stage2_24[61],stage2_23[62]}
   );
   gpc615_5 gpc5122 (
      {stage1_23[225], stage1_23[226], stage1_23[227], stage1_23[228], stage1_23[229]},
      {stage1_24[59]},
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage2_27[11],stage2_26[19],stage2_25[46],stage2_24[62],stage2_23[63]}
   );
   gpc615_5 gpc5123 (
      {stage1_23[230], stage1_23[231], stage1_23[232], stage1_23[233], stage1_23[234]},
      {stage1_24[60]},
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage2_27[12],stage2_26[20],stage2_25[47],stage2_24[63],stage2_23[64]}
   );
   gpc615_5 gpc5124 (
      {stage1_23[235], stage1_23[236], stage1_23[237], stage1_23[238], stage1_23[239]},
      {stage1_24[61]},
      {stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82], stage1_25[83]},
      {stage2_27[13],stage2_26[21],stage2_25[48],stage2_24[64],stage2_23[65]}
   );
   gpc615_5 gpc5125 (
      {stage1_23[240], stage1_23[241], stage1_23[242], stage1_23[243], stage1_23[244]},
      {stage1_24[62]},
      {stage1_25[84], stage1_25[85], stage1_25[86], stage1_25[87], stage1_25[88], stage1_25[89]},
      {stage2_27[14],stage2_26[22],stage2_25[49],stage2_24[65],stage2_23[66]}
   );
   gpc615_5 gpc5126 (
      {stage1_23[245], stage1_23[246], stage1_23[247], stage1_23[248], stage1_23[249]},
      {stage1_24[63]},
      {stage1_25[90], stage1_25[91], stage1_25[92], stage1_25[93], stage1_25[94], stage1_25[95]},
      {stage2_27[15],stage2_26[23],stage2_25[50],stage2_24[66],stage2_23[67]}
   );
   gpc615_5 gpc5127 (
      {stage1_23[250], stage1_23[251], stage1_23[252], stage1_23[253], stage1_23[254]},
      {stage1_24[64]},
      {stage1_25[96], stage1_25[97], stage1_25[98], stage1_25[99], stage1_25[100], stage1_25[101]},
      {stage2_27[16],stage2_26[24],stage2_25[51],stage2_24[67],stage2_23[68]}
   );
   gpc615_5 gpc5128 (
      {stage1_23[255], stage1_23[256], stage1_23[257], stage1_23[258], stage1_23[259]},
      {stage1_24[65]},
      {stage1_25[102], stage1_25[103], stage1_25[104], stage1_25[105], stage1_25[106], stage1_25[107]},
      {stage2_27[17],stage2_26[25],stage2_25[52],stage2_24[68],stage2_23[69]}
   );
   gpc615_5 gpc5129 (
      {stage1_23[260], stage1_23[261], stage1_23[262], stage1_23[263], stage1_23[264]},
      {stage1_24[66]},
      {stage1_25[108], stage1_25[109], stage1_25[110], stage1_25[111], stage1_25[112], stage1_25[113]},
      {stage2_27[18],stage2_26[26],stage2_25[53],stage2_24[69],stage2_23[70]}
   );
   gpc615_5 gpc5130 (
      {stage1_23[265], stage1_23[266], stage1_23[267], stage1_23[268], stage1_23[269]},
      {stage1_24[67]},
      {stage1_25[114], stage1_25[115], stage1_25[116], stage1_25[117], stage1_25[118], stage1_25[119]},
      {stage2_27[19],stage2_26[27],stage2_25[54],stage2_24[70],stage2_23[71]}
   );
   gpc615_5 gpc5131 (
      {stage1_23[270], stage1_23[271], stage1_23[272], stage1_23[273], stage1_23[274]},
      {stage1_24[68]},
      {stage1_25[120], stage1_25[121], stage1_25[122], stage1_25[123], stage1_25[124], stage1_25[125]},
      {stage2_27[20],stage2_26[28],stage2_25[55],stage2_24[71],stage2_23[72]}
   );
   gpc615_5 gpc5132 (
      {stage1_23[275], stage1_23[276], stage1_23[277], stage1_23[278], stage1_23[279]},
      {stage1_24[69]},
      {stage1_25[126], stage1_25[127], stage1_25[128], stage1_25[129], stage1_25[130], stage1_25[131]},
      {stage2_27[21],stage2_26[29],stage2_25[56],stage2_24[72],stage2_23[73]}
   );
   gpc615_5 gpc5133 (
      {stage1_23[280], stage1_23[281], stage1_23[282], stage1_23[283], stage1_23[284]},
      {stage1_24[70]},
      {stage1_25[132], stage1_25[133], stage1_25[134], stage1_25[135], stage1_25[136], stage1_25[137]},
      {stage2_27[22],stage2_26[30],stage2_25[57],stage2_24[73],stage2_23[74]}
   );
   gpc615_5 gpc5134 (
      {stage1_23[285], stage1_23[286], 1'b0, 1'b0, 1'b0},
      {stage1_24[71]},
      {stage1_25[138], stage1_25[139], stage1_25[140], stage1_25[141], stage1_25[142], stage1_25[143]},
      {stage2_27[23],stage2_26[31],stage2_25[58],stage2_24[74],stage2_23[75]}
   );
   gpc606_5 gpc5135 (
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[24],stage2_26[32],stage2_25[59],stage2_24[75]}
   );
   gpc606_5 gpc5136 (
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[25],stage2_26[33],stage2_25[60],stage2_24[76]}
   );
   gpc606_5 gpc5137 (
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[26],stage2_26[34],stage2_25[61],stage2_24[77]}
   );
   gpc606_5 gpc5138 (
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94], stage1_24[95]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[27],stage2_26[35],stage2_25[62],stage2_24[78]}
   );
   gpc606_5 gpc5139 (
      {stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99], stage1_24[100], stage1_24[101]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[28],stage2_26[36],stage2_25[63],stage2_24[79]}
   );
   gpc606_5 gpc5140 (
      {stage1_24[102], stage1_24[103], stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107]},
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage2_28[5],stage2_27[29],stage2_26[37],stage2_25[64],stage2_24[80]}
   );
   gpc606_5 gpc5141 (
      {stage1_24[108], stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage2_28[6],stage2_27[30],stage2_26[38],stage2_25[65],stage2_24[81]}
   );
   gpc606_5 gpc5142 (
      {stage1_24[114], stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118], stage1_24[119]},
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage2_28[7],stage2_27[31],stage2_26[39],stage2_25[66],stage2_24[82]}
   );
   gpc606_5 gpc5143 (
      {stage1_24[120], stage1_24[121], stage1_24[122], stage1_24[123], stage1_24[124], stage1_24[125]},
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage2_28[8],stage2_27[32],stage2_26[40],stage2_25[67],stage2_24[83]}
   );
   gpc606_5 gpc5144 (
      {stage1_24[126], stage1_24[127], stage1_24[128], stage1_24[129], stage1_24[130], stage1_24[131]},
      {stage1_26[54], stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59]},
      {stage2_28[9],stage2_27[33],stage2_26[41],stage2_25[68],stage2_24[84]}
   );
   gpc606_5 gpc5145 (
      {stage1_24[132], stage1_24[133], stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137]},
      {stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64], stage1_26[65]},
      {stage2_28[10],stage2_27[34],stage2_26[42],stage2_25[69],stage2_24[85]}
   );
   gpc606_5 gpc5146 (
      {stage1_24[138], stage1_24[139], stage1_24[140], stage1_24[141], stage1_24[142], stage1_24[143]},
      {stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69], stage1_26[70], stage1_26[71]},
      {stage2_28[11],stage2_27[35],stage2_26[43],stage2_25[70],stage2_24[86]}
   );
   gpc606_5 gpc5147 (
      {stage1_24[144], stage1_24[145], stage1_24[146], stage1_24[147], stage1_24[148], stage1_24[149]},
      {stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75], stage1_26[76], stage1_26[77]},
      {stage2_28[12],stage2_27[36],stage2_26[44],stage2_25[71],stage2_24[87]}
   );
   gpc606_5 gpc5148 (
      {stage1_24[150], stage1_24[151], stage1_24[152], stage1_24[153], stage1_24[154], stage1_24[155]},
      {stage1_26[78], stage1_26[79], stage1_26[80], stage1_26[81], stage1_26[82], stage1_26[83]},
      {stage2_28[13],stage2_27[37],stage2_26[45],stage2_25[72],stage2_24[88]}
   );
   gpc606_5 gpc5149 (
      {stage1_24[156], stage1_24[157], stage1_24[158], stage1_24[159], stage1_24[160], stage1_24[161]},
      {stage1_26[84], stage1_26[85], stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89]},
      {stage2_28[14],stage2_27[38],stage2_26[46],stage2_25[73],stage2_24[89]}
   );
   gpc606_5 gpc5150 (
      {stage1_24[162], stage1_24[163], stage1_24[164], stage1_24[165], stage1_24[166], stage1_24[167]},
      {stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94], stage1_26[95]},
      {stage2_28[15],stage2_27[39],stage2_26[47],stage2_25[74],stage2_24[90]}
   );
   gpc606_5 gpc5151 (
      {stage1_24[168], stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173]},
      {stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99], stage1_26[100], stage1_26[101]},
      {stage2_28[16],stage2_27[40],stage2_26[48],stage2_25[75],stage2_24[91]}
   );
   gpc606_5 gpc5152 (
      {stage1_24[174], stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178], stage1_24[179]},
      {stage1_26[102], stage1_26[103], stage1_26[104], stage1_26[105], stage1_26[106], stage1_26[107]},
      {stage2_28[17],stage2_27[41],stage2_26[49],stage2_25[76],stage2_24[92]}
   );
   gpc606_5 gpc5153 (
      {stage1_24[180], stage1_24[181], stage1_24[182], stage1_24[183], stage1_24[184], stage1_24[185]},
      {stage1_26[108], stage1_26[109], stage1_26[110], stage1_26[111], stage1_26[112], stage1_26[113]},
      {stage2_28[18],stage2_27[42],stage2_26[50],stage2_25[77],stage2_24[93]}
   );
   gpc606_5 gpc5154 (
      {stage1_24[186], stage1_24[187], stage1_24[188], stage1_24[189], stage1_24[190], stage1_24[191]},
      {stage1_26[114], stage1_26[115], stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119]},
      {stage2_28[19],stage2_27[43],stage2_26[51],stage2_25[78],stage2_24[94]}
   );
   gpc606_5 gpc5155 (
      {stage1_24[192], stage1_24[193], stage1_24[194], stage1_24[195], stage1_24[196], stage1_24[197]},
      {stage1_26[120], stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124], stage1_26[125]},
      {stage2_28[20],stage2_27[44],stage2_26[52],stage2_25[79],stage2_24[95]}
   );
   gpc606_5 gpc5156 (
      {stage1_24[198], stage1_24[199], stage1_24[200], stage1_24[201], stage1_24[202], stage1_24[203]},
      {stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129], stage1_26[130], stage1_26[131]},
      {stage2_28[21],stage2_27[45],stage2_26[53],stage2_25[80],stage2_24[96]}
   );
   gpc606_5 gpc5157 (
      {stage1_24[204], stage1_24[205], stage1_24[206], stage1_24[207], stage1_24[208], stage1_24[209]},
      {stage1_26[132], stage1_26[133], stage1_26[134], stage1_26[135], stage1_26[136], stage1_26[137]},
      {stage2_28[22],stage2_27[46],stage2_26[54],stage2_25[81],stage2_24[97]}
   );
   gpc207_4 gpc5158 (
      {stage1_25[144], stage1_25[145], stage1_25[146], stage1_25[147], stage1_25[148], stage1_25[149], stage1_25[150]},
      {stage1_27[0], stage1_27[1]},
      {stage2_28[23],stage2_27[47],stage2_26[55],stage2_25[82]}
   );
   gpc606_5 gpc5159 (
      {stage1_25[151], stage1_25[152], stage1_25[153], stage1_25[154], stage1_25[155], stage1_25[156]},
      {stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5], stage1_27[6], stage1_27[7]},
      {stage2_29[0],stage2_28[24],stage2_27[48],stage2_26[56],stage2_25[83]}
   );
   gpc606_5 gpc5160 (
      {stage1_25[157], stage1_25[158], stage1_25[159], stage1_25[160], stage1_25[161], stage1_25[162]},
      {stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11], stage1_27[12], stage1_27[13]},
      {stage2_29[1],stage2_28[25],stage2_27[49],stage2_26[57],stage2_25[84]}
   );
   gpc606_5 gpc5161 (
      {stage1_25[163], stage1_25[164], stage1_25[165], stage1_25[166], stage1_25[167], stage1_25[168]},
      {stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17], stage1_27[18], stage1_27[19]},
      {stage2_29[2],stage2_28[26],stage2_27[50],stage2_26[58],stage2_25[85]}
   );
   gpc606_5 gpc5162 (
      {stage1_25[169], stage1_25[170], stage1_25[171], stage1_25[172], stage1_25[173], stage1_25[174]},
      {stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23], stage1_27[24], stage1_27[25]},
      {stage2_29[3],stage2_28[27],stage2_27[51],stage2_26[59],stage2_25[86]}
   );
   gpc615_5 gpc5163 (
      {stage1_26[138], stage1_26[139], stage1_26[140], stage1_26[141], stage1_26[142]},
      {stage1_27[26]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[4],stage2_28[28],stage2_27[52],stage2_26[60]}
   );
   gpc615_5 gpc5164 (
      {stage1_26[143], stage1_26[144], stage1_26[145], stage1_26[146], stage1_26[147]},
      {stage1_27[27]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[5],stage2_28[29],stage2_27[53],stage2_26[61]}
   );
   gpc615_5 gpc5165 (
      {stage1_26[148], stage1_26[149], stage1_26[150], stage1_26[151], stage1_26[152]},
      {stage1_27[28]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[6],stage2_28[30],stage2_27[54],stage2_26[62]}
   );
   gpc615_5 gpc5166 (
      {stage1_26[153], stage1_26[154], stage1_26[155], stage1_26[156], stage1_26[157]},
      {stage1_27[29]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[7],stage2_28[31],stage2_27[55],stage2_26[63]}
   );
   gpc615_5 gpc5167 (
      {stage1_26[158], stage1_26[159], stage1_26[160], stage1_26[161], stage1_26[162]},
      {stage1_27[30]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[8],stage2_28[32],stage2_27[56],stage2_26[64]}
   );
   gpc615_5 gpc5168 (
      {stage1_26[163], stage1_26[164], stage1_26[165], stage1_26[166], stage1_26[167]},
      {stage1_27[31]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[9],stage2_28[33],stage2_27[57],stage2_26[65]}
   );
   gpc615_5 gpc5169 (
      {stage1_26[168], stage1_26[169], stage1_26[170], stage1_26[171], stage1_26[172]},
      {stage1_27[32]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[10],stage2_28[34],stage2_27[58],stage2_26[66]}
   );
   gpc615_5 gpc5170 (
      {stage1_26[173], stage1_26[174], stage1_26[175], stage1_26[176], stage1_26[177]},
      {stage1_27[33]},
      {stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47]},
      {stage2_30[7],stage2_29[11],stage2_28[35],stage2_27[59],stage2_26[67]}
   );
   gpc615_5 gpc5171 (
      {stage1_26[178], stage1_26[179], stage1_26[180], stage1_26[181], stage1_26[182]},
      {stage1_27[34]},
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage2_30[8],stage2_29[12],stage2_28[36],stage2_27[60],stage2_26[68]}
   );
   gpc615_5 gpc5172 (
      {stage1_26[183], stage1_26[184], stage1_26[185], stage1_26[186], stage1_26[187]},
      {stage1_27[35]},
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage2_30[9],stage2_29[13],stage2_28[37],stage2_27[61],stage2_26[69]}
   );
   gpc615_5 gpc5173 (
      {stage1_26[188], stage1_26[189], stage1_26[190], stage1_26[191], stage1_26[192]},
      {stage1_27[36]},
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage2_30[10],stage2_29[14],stage2_28[38],stage2_27[62],stage2_26[70]}
   );
   gpc615_5 gpc5174 (
      {stage1_26[193], stage1_26[194], stage1_26[195], stage1_26[196], stage1_26[197]},
      {stage1_27[37]},
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage2_30[11],stage2_29[15],stage2_28[39],stage2_27[63],stage2_26[71]}
   );
   gpc615_5 gpc5175 (
      {stage1_26[198], stage1_26[199], stage1_26[200], stage1_26[201], stage1_26[202]},
      {stage1_27[38]},
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage2_30[12],stage2_29[16],stage2_28[40],stage2_27[64],stage2_26[72]}
   );
   gpc615_5 gpc5176 (
      {stage1_26[203], stage1_26[204], stage1_26[205], stage1_26[206], stage1_26[207]},
      {stage1_27[39]},
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage2_30[13],stage2_29[17],stage2_28[41],stage2_27[65],stage2_26[73]}
   );
   gpc615_5 gpc5177 (
      {stage1_26[208], stage1_26[209], stage1_26[210], stage1_26[211], stage1_26[212]},
      {stage1_27[40]},
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage2_30[14],stage2_29[18],stage2_28[42],stage2_27[66],stage2_26[74]}
   );
   gpc615_5 gpc5178 (
      {stage1_26[213], stage1_26[214], stage1_26[215], stage1_26[216], stage1_26[217]},
      {stage1_27[41]},
      {stage1_28[90], stage1_28[91], stage1_28[92], stage1_28[93], stage1_28[94], stage1_28[95]},
      {stage2_30[15],stage2_29[19],stage2_28[43],stage2_27[67],stage2_26[75]}
   );
   gpc615_5 gpc5179 (
      {stage1_26[218], stage1_26[219], stage1_26[220], stage1_26[221], stage1_26[222]},
      {stage1_27[42]},
      {stage1_28[96], stage1_28[97], stage1_28[98], stage1_28[99], stage1_28[100], stage1_28[101]},
      {stage2_30[16],stage2_29[20],stage2_28[44],stage2_27[68],stage2_26[76]}
   );
   gpc615_5 gpc5180 (
      {stage1_26[223], stage1_26[224], stage1_26[225], stage1_26[226], stage1_26[227]},
      {stage1_27[43]},
      {stage1_28[102], stage1_28[103], stage1_28[104], stage1_28[105], stage1_28[106], stage1_28[107]},
      {stage2_30[17],stage2_29[21],stage2_28[45],stage2_27[69],stage2_26[77]}
   );
   gpc615_5 gpc5181 (
      {stage1_26[228], stage1_26[229], stage1_26[230], stage1_26[231], stage1_26[232]},
      {stage1_27[44]},
      {stage1_28[108], stage1_28[109], stage1_28[110], stage1_28[111], stage1_28[112], stage1_28[113]},
      {stage2_30[18],stage2_29[22],stage2_28[46],stage2_27[70],stage2_26[78]}
   );
   gpc615_5 gpc5182 (
      {stage1_26[233], stage1_26[234], stage1_26[235], stage1_26[236], stage1_26[237]},
      {stage1_27[45]},
      {stage1_28[114], stage1_28[115], stage1_28[116], stage1_28[117], stage1_28[118], stage1_28[119]},
      {stage2_30[19],stage2_29[23],stage2_28[47],stage2_27[71],stage2_26[79]}
   );
   gpc615_5 gpc5183 (
      {stage1_26[238], stage1_26[239], stage1_26[240], stage1_26[241], stage1_26[242]},
      {stage1_27[46]},
      {stage1_28[120], stage1_28[121], stage1_28[122], stage1_28[123], stage1_28[124], stage1_28[125]},
      {stage2_30[20],stage2_29[24],stage2_28[48],stage2_27[72],stage2_26[80]}
   );
   gpc615_5 gpc5184 (
      {stage1_26[243], stage1_26[244], stage1_26[245], stage1_26[246], stage1_26[247]},
      {stage1_27[47]},
      {stage1_28[126], stage1_28[127], stage1_28[128], stage1_28[129], stage1_28[130], stage1_28[131]},
      {stage2_30[21],stage2_29[25],stage2_28[49],stage2_27[73],stage2_26[81]}
   );
   gpc615_5 gpc5185 (
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52]},
      {stage1_28[132]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[22],stage2_29[26],stage2_28[50],stage2_27[74]}
   );
   gpc615_5 gpc5186 (
      {stage1_27[53], stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57]},
      {stage1_28[133]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[23],stage2_29[27],stage2_28[51],stage2_27[75]}
   );
   gpc615_5 gpc5187 (
      {stage1_27[58], stage1_27[59], stage1_27[60], stage1_27[61], stage1_27[62]},
      {stage1_28[134]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[24],stage2_29[28],stage2_28[52],stage2_27[76]}
   );
   gpc615_5 gpc5188 (
      {stage1_27[63], stage1_27[64], stage1_27[65], stage1_27[66], stage1_27[67]},
      {stage1_28[135]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[25],stage2_29[29],stage2_28[53],stage2_27[77]}
   );
   gpc615_5 gpc5189 (
      {stage1_27[68], stage1_27[69], stage1_27[70], stage1_27[71], stage1_27[72]},
      {stage1_28[136]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[26],stage2_29[30],stage2_28[54],stage2_27[78]}
   );
   gpc615_5 gpc5190 (
      {stage1_27[73], stage1_27[74], stage1_27[75], stage1_27[76], stage1_27[77]},
      {stage1_28[137]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[27],stage2_29[31],stage2_28[55],stage2_27[79]}
   );
   gpc615_5 gpc5191 (
      {stage1_27[78], stage1_27[79], stage1_27[80], stage1_27[81], stage1_27[82]},
      {stage1_28[138]},
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage2_31[6],stage2_30[28],stage2_29[32],stage2_28[56],stage2_27[80]}
   );
   gpc615_5 gpc5192 (
      {stage1_27[83], stage1_27[84], stage1_27[85], stage1_27[86], stage1_27[87]},
      {stage1_28[139]},
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage2_31[7],stage2_30[29],stage2_29[33],stage2_28[57],stage2_27[81]}
   );
   gpc615_5 gpc5193 (
      {stage1_27[88], stage1_27[89], stage1_27[90], stage1_27[91], stage1_27[92]},
      {stage1_28[140]},
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage2_31[8],stage2_30[30],stage2_29[34],stage2_28[58],stage2_27[82]}
   );
   gpc615_5 gpc5194 (
      {stage1_27[93], stage1_27[94], stage1_27[95], stage1_27[96], stage1_27[97]},
      {stage1_28[141]},
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage2_31[9],stage2_30[31],stage2_29[35],stage2_28[59],stage2_27[83]}
   );
   gpc615_5 gpc5195 (
      {stage1_27[98], stage1_27[99], stage1_27[100], stage1_27[101], stage1_27[102]},
      {stage1_28[142]},
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage2_31[10],stage2_30[32],stage2_29[36],stage2_28[60],stage2_27[84]}
   );
   gpc615_5 gpc5196 (
      {stage1_27[103], stage1_27[104], stage1_27[105], stage1_27[106], stage1_27[107]},
      {stage1_28[143]},
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage2_31[11],stage2_30[33],stage2_29[37],stage2_28[61],stage2_27[85]}
   );
   gpc615_5 gpc5197 (
      {stage1_27[108], stage1_27[109], stage1_27[110], stage1_27[111], stage1_27[112]},
      {stage1_28[144]},
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage2_31[12],stage2_30[34],stage2_29[38],stage2_28[62],stage2_27[86]}
   );
   gpc615_5 gpc5198 (
      {stage1_27[113], stage1_27[114], stage1_27[115], stage1_27[116], stage1_27[117]},
      {stage1_28[145]},
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage2_31[13],stage2_30[35],stage2_29[39],stage2_28[63],stage2_27[87]}
   );
   gpc615_5 gpc5199 (
      {stage1_27[118], stage1_27[119], stage1_27[120], stage1_27[121], stage1_27[122]},
      {stage1_28[146]},
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage2_31[14],stage2_30[36],stage2_29[40],stage2_28[64],stage2_27[88]}
   );
   gpc615_5 gpc5200 (
      {stage1_27[123], stage1_27[124], stage1_27[125], stage1_27[126], stage1_27[127]},
      {stage1_28[147]},
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage2_31[15],stage2_30[37],stage2_29[41],stage2_28[65],stage2_27[89]}
   );
   gpc615_5 gpc5201 (
      {stage1_27[128], stage1_27[129], stage1_27[130], stage1_27[131], stage1_27[132]},
      {stage1_28[148]},
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage2_31[16],stage2_30[38],stage2_29[42],stage2_28[66],stage2_27[90]}
   );
   gpc615_5 gpc5202 (
      {stage1_27[133], stage1_27[134], stage1_27[135], stage1_27[136], stage1_27[137]},
      {stage1_28[149]},
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage2_31[17],stage2_30[39],stage2_29[43],stage2_28[67],stage2_27[91]}
   );
   gpc615_5 gpc5203 (
      {stage1_27[138], stage1_27[139], stage1_27[140], stage1_27[141], stage1_27[142]},
      {stage1_28[150]},
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage2_31[18],stage2_30[40],stage2_29[44],stage2_28[68],stage2_27[92]}
   );
   gpc615_5 gpc5204 (
      {stage1_27[143], stage1_27[144], stage1_27[145], stage1_27[146], stage1_27[147]},
      {stage1_28[151]},
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], stage1_29[118], stage1_29[119]},
      {stage2_31[19],stage2_30[41],stage2_29[45],stage2_28[69],stage2_27[93]}
   );
   gpc615_5 gpc5205 (
      {stage1_27[148], stage1_27[149], stage1_27[150], stage1_27[151], stage1_27[152]},
      {stage1_28[152]},
      {stage1_29[120], stage1_29[121], stage1_29[122], stage1_29[123], stage1_29[124], stage1_29[125]},
      {stage2_31[20],stage2_30[42],stage2_29[46],stage2_28[70],stage2_27[94]}
   );
   gpc615_5 gpc5206 (
      {stage1_27[153], stage1_27[154], stage1_27[155], stage1_27[156], stage1_27[157]},
      {stage1_28[153]},
      {stage1_29[126], stage1_29[127], stage1_29[128], stage1_29[129], stage1_29[130], stage1_29[131]},
      {stage2_31[21],stage2_30[43],stage2_29[47],stage2_28[71],stage2_27[95]}
   );
   gpc615_5 gpc5207 (
      {stage1_27[158], stage1_27[159], stage1_27[160], stage1_27[161], stage1_27[162]},
      {stage1_28[154]},
      {stage1_29[132], stage1_29[133], stage1_29[134], stage1_29[135], stage1_29[136], stage1_29[137]},
      {stage2_31[22],stage2_30[44],stage2_29[48],stage2_28[72],stage2_27[96]}
   );
   gpc615_5 gpc5208 (
      {stage1_27[163], stage1_27[164], stage1_27[165], stage1_27[166], stage1_27[167]},
      {stage1_28[155]},
      {stage1_29[138], stage1_29[139], stage1_29[140], stage1_29[141], stage1_29[142], stage1_29[143]},
      {stage2_31[23],stage2_30[45],stage2_29[49],stage2_28[73],stage2_27[97]}
   );
   gpc615_5 gpc5209 (
      {stage1_27[168], stage1_27[169], stage1_27[170], stage1_27[171], stage1_27[172]},
      {stage1_28[156]},
      {stage1_29[144], stage1_29[145], stage1_29[146], stage1_29[147], stage1_29[148], stage1_29[149]},
      {stage2_31[24],stage2_30[46],stage2_29[50],stage2_28[74],stage2_27[98]}
   );
   gpc615_5 gpc5210 (
      {stage1_27[173], stage1_27[174], stage1_27[175], stage1_27[176], stage1_27[177]},
      {stage1_28[157]},
      {stage1_29[150], stage1_29[151], stage1_29[152], stage1_29[153], stage1_29[154], stage1_29[155]},
      {stage2_31[25],stage2_30[47],stage2_29[51],stage2_28[75],stage2_27[99]}
   );
   gpc615_5 gpc5211 (
      {stage1_27[178], stage1_27[179], stage1_27[180], stage1_27[181], stage1_27[182]},
      {stage1_28[158]},
      {stage1_29[156], stage1_29[157], stage1_29[158], stage1_29[159], stage1_29[160], stage1_29[161]},
      {stage2_31[26],stage2_30[48],stage2_29[52],stage2_28[76],stage2_27[100]}
   );
   gpc615_5 gpc5212 (
      {stage1_27[183], stage1_27[184], stage1_27[185], stage1_27[186], stage1_27[187]},
      {stage1_28[159]},
      {stage1_29[162], stage1_29[163], stage1_29[164], stage1_29[165], stage1_29[166], stage1_29[167]},
      {stage2_31[27],stage2_30[49],stage2_29[53],stage2_28[77],stage2_27[101]}
   );
   gpc615_5 gpc5213 (
      {stage1_27[188], stage1_27[189], stage1_27[190], stage1_27[191], stage1_27[192]},
      {stage1_28[160]},
      {stage1_29[168], stage1_29[169], stage1_29[170], stage1_29[171], stage1_29[172], stage1_29[173]},
      {stage2_31[28],stage2_30[50],stage2_29[54],stage2_28[78],stage2_27[102]}
   );
   gpc615_5 gpc5214 (
      {stage1_27[193], stage1_27[194], stage1_27[195], stage1_27[196], stage1_27[197]},
      {stage1_28[161]},
      {stage1_29[174], stage1_29[175], stage1_29[176], stage1_29[177], stage1_29[178], stage1_29[179]},
      {stage2_31[29],stage2_30[51],stage2_29[55],stage2_28[79],stage2_27[103]}
   );
   gpc615_5 gpc5215 (
      {stage1_27[198], stage1_27[199], stage1_27[200], stage1_27[201], stage1_27[202]},
      {stage1_28[162]},
      {stage1_29[180], stage1_29[181], stage1_29[182], stage1_29[183], stage1_29[184], stage1_29[185]},
      {stage2_31[30],stage2_30[52],stage2_29[56],stage2_28[80],stage2_27[104]}
   );
   gpc615_5 gpc5216 (
      {stage1_27[203], stage1_27[204], stage1_27[205], 1'b0, 1'b0},
      {stage1_28[163]},
      {stage1_29[186], stage1_29[187], stage1_29[188], stage1_29[189], stage1_29[190], stage1_29[191]},
      {stage2_31[31],stage2_30[53],stage2_29[57],stage2_28[81],stage2_27[105]}
   );
   gpc606_5 gpc5217 (
      {stage1_28[164], stage1_28[165], stage1_28[166], stage1_28[167], stage1_28[168], stage1_28[169]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[32],stage2_30[54],stage2_29[58],stage2_28[82]}
   );
   gpc606_5 gpc5218 (
      {stage1_28[170], stage1_28[171], stage1_28[172], stage1_28[173], stage1_28[174], stage1_28[175]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[33],stage2_30[55],stage2_29[59],stage2_28[83]}
   );
   gpc606_5 gpc5219 (
      {stage1_28[176], stage1_28[177], stage1_28[178], stage1_28[179], stage1_28[180], stage1_28[181]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[34],stage2_30[56],stage2_29[60],stage2_28[84]}
   );
   gpc606_5 gpc5220 (
      {stage1_28[182], stage1_28[183], stage1_28[184], stage1_28[185], stage1_28[186], stage1_28[187]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[35],stage2_30[57],stage2_29[61],stage2_28[85]}
   );
   gpc606_5 gpc5221 (
      {stage1_28[188], stage1_28[189], stage1_28[190], stage1_28[191], stage1_28[192], stage1_28[193]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[36],stage2_30[58],stage2_29[62],stage2_28[86]}
   );
   gpc606_5 gpc5222 (
      {stage1_28[194], stage1_28[195], stage1_28[196], stage1_28[197], stage1_28[198], stage1_28[199]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[37],stage2_30[59],stage2_29[63],stage2_28[87]}
   );
   gpc606_5 gpc5223 (
      {stage1_28[200], stage1_28[201], stage1_28[202], stage1_28[203], stage1_28[204], stage1_28[205]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[38],stage2_30[60],stage2_29[64],stage2_28[88]}
   );
   gpc606_5 gpc5224 (
      {stage1_28[206], stage1_28[207], stage1_28[208], stage1_28[209], stage1_28[210], stage1_28[211]},
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage2_32[7],stage2_31[39],stage2_30[61],stage2_29[65],stage2_28[89]}
   );
   gpc606_5 gpc5225 (
      {stage1_28[212], stage1_28[213], stage1_28[214], stage1_28[215], stage1_28[216], stage1_28[217]},
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage2_32[8],stage2_31[40],stage2_30[62],stage2_29[66],stage2_28[90]}
   );
   gpc606_5 gpc5226 (
      {stage1_28[218], stage1_28[219], stage1_28[220], stage1_28[221], stage1_28[222], stage1_28[223]},
      {stage1_30[54], stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59]},
      {stage2_32[9],stage2_31[41],stage2_30[63],stage2_29[67],stage2_28[91]}
   );
   gpc1163_5 gpc5227 (
      {stage1_29[192], stage1_29[193], stage1_29[194]},
      {stage1_30[60], stage1_30[61], stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65]},
      {stage1_31[0]},
      {stage1_32[0]},
      {stage2_33[0],stage2_32[10],stage2_31[42],stage2_30[64],stage2_29[68]}
   );
   gpc1163_5 gpc5228 (
      {stage1_29[195], stage1_29[196], stage1_29[197]},
      {stage1_30[66], stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_31[1]},
      {stage1_32[1]},
      {stage2_33[1],stage2_32[11],stage2_31[43],stage2_30[65],stage2_29[69]}
   );
   gpc1163_5 gpc5229 (
      {stage1_29[198], stage1_29[199], stage1_29[200]},
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76], stage1_30[77]},
      {stage1_31[2]},
      {stage1_32[2]},
      {stage2_33[2],stage2_32[12],stage2_31[44],stage2_30[66],stage2_29[70]}
   );
   gpc1163_5 gpc5230 (
      {stage1_29[201], stage1_29[202], stage1_29[203]},
      {stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81], stage1_30[82], stage1_30[83]},
      {stage1_31[3]},
      {stage1_32[3]},
      {stage2_33[3],stage2_32[13],stage2_31[45],stage2_30[67],stage2_29[71]}
   );
   gpc606_5 gpc5231 (
      {stage1_29[204], stage1_29[205], stage1_29[206], stage1_29[207], stage1_29[208], stage1_29[209]},
      {stage1_31[4], stage1_31[5], stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9]},
      {stage2_33[4],stage2_32[14],stage2_31[46],stage2_30[68],stage2_29[72]}
   );
   gpc606_5 gpc5232 (
      {stage1_29[210], stage1_29[211], stage1_29[212], stage1_29[213], stage1_29[214], stage1_29[215]},
      {stage1_31[10], stage1_31[11], stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15]},
      {stage2_33[5],stage2_32[15],stage2_31[47],stage2_30[69],stage2_29[73]}
   );
   gpc606_5 gpc5233 (
      {stage1_30[84], stage1_30[85], stage1_30[86], stage1_30[87], stage1_30[88], stage1_30[89]},
      {stage1_32[4], stage1_32[5], stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9]},
      {stage2_34[0],stage2_33[6],stage2_32[16],stage2_31[48],stage2_30[70]}
   );
   gpc615_5 gpc5234 (
      {stage1_30[90], stage1_30[91], stage1_30[92], stage1_30[93], stage1_30[94]},
      {stage1_31[16]},
      {stage1_32[10], stage1_32[11], stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15]},
      {stage2_34[1],stage2_33[7],stage2_32[17],stage2_31[49],stage2_30[71]}
   );
   gpc615_5 gpc5235 (
      {stage1_30[95], stage1_30[96], stage1_30[97], stage1_30[98], stage1_30[99]},
      {stage1_31[17]},
      {stage1_32[16], stage1_32[17], stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21]},
      {stage2_34[2],stage2_33[8],stage2_32[18],stage2_31[50],stage2_30[72]}
   );
   gpc615_5 gpc5236 (
      {stage1_30[100], stage1_30[101], stage1_30[102], stage1_30[103], stage1_30[104]},
      {stage1_31[18]},
      {stage1_32[22], stage1_32[23], stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27]},
      {stage2_34[3],stage2_33[9],stage2_32[19],stage2_31[51],stage2_30[73]}
   );
   gpc615_5 gpc5237 (
      {stage1_30[105], stage1_30[106], stage1_30[107], stage1_30[108], stage1_30[109]},
      {stage1_31[19]},
      {stage1_32[28], stage1_32[29], stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33]},
      {stage2_34[4],stage2_33[10],stage2_32[20],stage2_31[52],stage2_30[74]}
   );
   gpc615_5 gpc5238 (
      {stage1_30[110], stage1_30[111], stage1_30[112], stage1_30[113], stage1_30[114]},
      {stage1_31[20]},
      {stage1_32[34], stage1_32[35], stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39]},
      {stage2_34[5],stage2_33[11],stage2_32[21],stage2_31[53],stage2_30[75]}
   );
   gpc615_5 gpc5239 (
      {stage1_30[115], stage1_30[116], stage1_30[117], stage1_30[118], stage1_30[119]},
      {stage1_31[21]},
      {stage1_32[40], stage1_32[41], stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45]},
      {stage2_34[6],stage2_33[12],stage2_32[22],stage2_31[54],stage2_30[76]}
   );
   gpc615_5 gpc5240 (
      {stage1_30[120], stage1_30[121], stage1_30[122], stage1_30[123], stage1_30[124]},
      {stage1_31[22]},
      {stage1_32[46], stage1_32[47], stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51]},
      {stage2_34[7],stage2_33[13],stage2_32[23],stage2_31[55],stage2_30[77]}
   );
   gpc615_5 gpc5241 (
      {stage1_30[125], stage1_30[126], stage1_30[127], stage1_30[128], stage1_30[129]},
      {stage1_31[23]},
      {stage1_32[52], stage1_32[53], stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57]},
      {stage2_34[8],stage2_33[14],stage2_32[24],stage2_31[56],stage2_30[78]}
   );
   gpc615_5 gpc5242 (
      {stage1_30[130], stage1_30[131], stage1_30[132], stage1_30[133], stage1_30[134]},
      {stage1_31[24]},
      {stage1_32[58], stage1_32[59], stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63]},
      {stage2_34[9],stage2_33[15],stage2_32[25],stage2_31[57],stage2_30[79]}
   );
   gpc615_5 gpc5243 (
      {stage1_30[135], stage1_30[136], stage1_30[137], stage1_30[138], stage1_30[139]},
      {stage1_31[25]},
      {stage1_32[64], stage1_32[65], stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69]},
      {stage2_34[10],stage2_33[16],stage2_32[26],stage2_31[58],stage2_30[80]}
   );
   gpc615_5 gpc5244 (
      {stage1_30[140], stage1_30[141], stage1_30[142], stage1_30[143], stage1_30[144]},
      {stage1_31[26]},
      {stage1_32[70], stage1_32[71], stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75]},
      {stage2_34[11],stage2_33[17],stage2_32[27],stage2_31[59],stage2_30[81]}
   );
   gpc615_5 gpc5245 (
      {stage1_30[145], stage1_30[146], stage1_30[147], stage1_30[148], stage1_30[149]},
      {stage1_31[27]},
      {stage1_32[76], stage1_32[77], stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81]},
      {stage2_34[12],stage2_33[18],stage2_32[28],stage2_31[60],stage2_30[82]}
   );
   gpc615_5 gpc5246 (
      {stage1_30[150], stage1_30[151], stage1_30[152], stage1_30[153], stage1_30[154]},
      {stage1_31[28]},
      {stage1_32[82], stage1_32[83], stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87]},
      {stage2_34[13],stage2_33[19],stage2_32[29],stage2_31[61],stage2_30[83]}
   );
   gpc615_5 gpc5247 (
      {stage1_30[155], stage1_30[156], stage1_30[157], stage1_30[158], stage1_30[159]},
      {stage1_31[29]},
      {stage1_32[88], stage1_32[89], stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93]},
      {stage2_34[14],stage2_33[20],stage2_32[30],stage2_31[62],stage2_30[84]}
   );
   gpc1163_5 gpc5248 (
      {stage1_31[30], stage1_31[31], stage1_31[32]},
      {stage1_32[94], stage1_32[95], stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99]},
      {stage1_33[0]},
      {stage1_34[0]},
      {stage2_35[0],stage2_34[15],stage2_33[21],stage2_32[31],stage2_31[63]}
   );
   gpc606_5 gpc5249 (
      {stage1_31[33], stage1_31[34], stage1_31[35], stage1_31[36], stage1_31[37], stage1_31[38]},
      {stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5], stage1_33[6]},
      {stage2_35[1],stage2_34[16],stage2_33[22],stage2_32[32],stage2_31[64]}
   );
   gpc606_5 gpc5250 (
      {stage1_31[39], stage1_31[40], stage1_31[41], stage1_31[42], stage1_31[43], stage1_31[44]},
      {stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11], stage1_33[12]},
      {stage2_35[2],stage2_34[17],stage2_33[23],stage2_32[33],stage2_31[65]}
   );
   gpc606_5 gpc5251 (
      {stage1_31[45], stage1_31[46], stage1_31[47], stage1_31[48], stage1_31[49], stage1_31[50]},
      {stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17], stage1_33[18]},
      {stage2_35[3],stage2_34[18],stage2_33[24],stage2_32[34],stage2_31[66]}
   );
   gpc606_5 gpc5252 (
      {stage1_31[51], stage1_31[52], stage1_31[53], stage1_31[54], stage1_31[55], stage1_31[56]},
      {stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23], stage1_33[24]},
      {stage2_35[4],stage2_34[19],stage2_33[25],stage2_32[35],stage2_31[67]}
   );
   gpc606_5 gpc5253 (
      {stage1_31[57], stage1_31[58], stage1_31[59], stage1_31[60], stage1_31[61], stage1_31[62]},
      {stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29], stage1_33[30]},
      {stage2_35[5],stage2_34[20],stage2_33[26],stage2_32[36],stage2_31[68]}
   );
   gpc606_5 gpc5254 (
      {stage1_31[63], stage1_31[64], stage1_31[65], stage1_31[66], stage1_31[67], stage1_31[68]},
      {stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35], stage1_33[36]},
      {stage2_35[6],stage2_34[21],stage2_33[27],stage2_32[37],stage2_31[69]}
   );
   gpc606_5 gpc5255 (
      {stage1_31[69], stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73], stage1_31[74]},
      {stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41], stage1_33[42]},
      {stage2_35[7],stage2_34[22],stage2_33[28],stage2_32[38],stage2_31[70]}
   );
   gpc606_5 gpc5256 (
      {stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78], stage1_31[79], stage1_31[80]},
      {stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47], stage1_33[48]},
      {stage2_35[8],stage2_34[23],stage2_33[29],stage2_32[39],stage2_31[71]}
   );
   gpc606_5 gpc5257 (
      {stage1_31[81], stage1_31[82], stage1_31[83], stage1_31[84], stage1_31[85], stage1_31[86]},
      {stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53], stage1_33[54]},
      {stage2_35[9],stage2_34[24],stage2_33[30],stage2_32[40],stage2_31[72]}
   );
   gpc606_5 gpc5258 (
      {stage1_31[87], stage1_31[88], stage1_31[89], stage1_31[90], stage1_31[91], stage1_31[92]},
      {stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59], stage1_33[60]},
      {stage2_35[10],stage2_34[25],stage2_33[31],stage2_32[41],stage2_31[73]}
   );
   gpc606_5 gpc5259 (
      {stage1_31[93], stage1_31[94], stage1_31[95], stage1_31[96], stage1_31[97], stage1_31[98]},
      {stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65], stage1_33[66]},
      {stage2_35[11],stage2_34[26],stage2_33[32],stage2_32[42],stage2_31[74]}
   );
   gpc606_5 gpc5260 (
      {stage1_31[99], stage1_31[100], stage1_31[101], stage1_31[102], stage1_31[103], stage1_31[104]},
      {stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71], stage1_33[72]},
      {stage2_35[12],stage2_34[27],stage2_33[33],stage2_32[43],stage2_31[75]}
   );
   gpc615_5 gpc5261 (
      {stage1_31[105], stage1_31[106], stage1_31[107], stage1_31[108], stage1_31[109]},
      {stage1_32[100]},
      {stage1_33[73], stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77], stage1_33[78]},
      {stage2_35[13],stage2_34[28],stage2_33[34],stage2_32[44],stage2_31[76]}
   );
   gpc615_5 gpc5262 (
      {stage1_31[110], stage1_31[111], stage1_31[112], stage1_31[113], stage1_31[114]},
      {stage1_32[101]},
      {stage1_33[79], stage1_33[80], stage1_33[81], stage1_33[82], stage1_33[83], stage1_33[84]},
      {stage2_35[14],stage2_34[29],stage2_33[35],stage2_32[45],stage2_31[77]}
   );
   gpc615_5 gpc5263 (
      {stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118], stage1_31[119]},
      {stage1_32[102]},
      {stage1_33[85], stage1_33[86], stage1_33[87], stage1_33[88], stage1_33[89], stage1_33[90]},
      {stage2_35[15],stage2_34[30],stage2_33[36],stage2_32[46],stage2_31[78]}
   );
   gpc615_5 gpc5264 (
      {stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123], stage1_31[124]},
      {stage1_32[103]},
      {stage1_33[91], stage1_33[92], stage1_33[93], stage1_33[94], stage1_33[95], stage1_33[96]},
      {stage2_35[16],stage2_34[31],stage2_33[37],stage2_32[47],stage2_31[79]}
   );
   gpc615_5 gpc5265 (
      {stage1_31[125], stage1_31[126], stage1_31[127], stage1_31[128], stage1_31[129]},
      {stage1_32[104]},
      {stage1_33[97], stage1_33[98], stage1_33[99], stage1_33[100], stage1_33[101], stage1_33[102]},
      {stage2_35[17],stage2_34[32],stage2_33[38],stage2_32[48],stage2_31[80]}
   );
   gpc615_5 gpc5266 (
      {stage1_31[130], stage1_31[131], stage1_31[132], stage1_31[133], stage1_31[134]},
      {stage1_32[105]},
      {stage1_33[103], stage1_33[104], stage1_33[105], stage1_33[106], stage1_33[107], stage1_33[108]},
      {stage2_35[18],stage2_34[33],stage2_33[39],stage2_32[49],stage2_31[81]}
   );
   gpc615_5 gpc5267 (
      {stage1_31[135], stage1_31[136], stage1_31[137], stage1_31[138], stage1_31[139]},
      {stage1_32[106]},
      {stage1_33[109], stage1_33[110], stage1_33[111], stage1_33[112], stage1_33[113], stage1_33[114]},
      {stage2_35[19],stage2_34[34],stage2_33[40],stage2_32[50],stage2_31[82]}
   );
   gpc615_5 gpc5268 (
      {stage1_31[140], stage1_31[141], stage1_31[142], stage1_31[143], stage1_31[144]},
      {stage1_32[107]},
      {stage1_33[115], stage1_33[116], stage1_33[117], stage1_33[118], stage1_33[119], stage1_33[120]},
      {stage2_35[20],stage2_34[35],stage2_33[41],stage2_32[51],stage2_31[83]}
   );
   gpc615_5 gpc5269 (
      {stage1_31[145], stage1_31[146], stage1_31[147], stage1_31[148], stage1_31[149]},
      {stage1_32[108]},
      {stage1_33[121], stage1_33[122], stage1_33[123], stage1_33[124], stage1_33[125], stage1_33[126]},
      {stage2_35[21],stage2_34[36],stage2_33[42],stage2_32[52],stage2_31[84]}
   );
   gpc615_5 gpc5270 (
      {stage1_31[150], stage1_31[151], stage1_31[152], stage1_31[153], stage1_31[154]},
      {stage1_32[109]},
      {stage1_33[127], stage1_33[128], stage1_33[129], stage1_33[130], stage1_33[131], stage1_33[132]},
      {stage2_35[22],stage2_34[37],stage2_33[43],stage2_32[53],stage2_31[85]}
   );
   gpc615_5 gpc5271 (
      {stage1_31[155], stage1_31[156], stage1_31[157], stage1_31[158], stage1_31[159]},
      {stage1_32[110]},
      {stage1_33[133], stage1_33[134], stage1_33[135], stage1_33[136], stage1_33[137], stage1_33[138]},
      {stage2_35[23],stage2_34[38],stage2_33[44],stage2_32[54],stage2_31[86]}
   );
   gpc615_5 gpc5272 (
      {stage1_31[160], stage1_31[161], stage1_31[162], stage1_31[163], stage1_31[164]},
      {stage1_32[111]},
      {stage1_33[139], stage1_33[140], stage1_33[141], stage1_33[142], stage1_33[143], stage1_33[144]},
      {stage2_35[24],stage2_34[39],stage2_33[45],stage2_32[55],stage2_31[87]}
   );
   gpc615_5 gpc5273 (
      {stage1_31[165], stage1_31[166], stage1_31[167], stage1_31[168], stage1_31[169]},
      {stage1_32[112]},
      {stage1_33[145], stage1_33[146], stage1_33[147], stage1_33[148], stage1_33[149], stage1_33[150]},
      {stage2_35[25],stage2_34[40],stage2_33[46],stage2_32[56],stage2_31[88]}
   );
   gpc615_5 gpc5274 (
      {stage1_31[170], stage1_31[171], stage1_31[172], stage1_31[173], stage1_31[174]},
      {stage1_32[113]},
      {stage1_33[151], stage1_33[152], stage1_33[153], stage1_33[154], stage1_33[155], stage1_33[156]},
      {stage2_35[26],stage2_34[41],stage2_33[47],stage2_32[57],stage2_31[89]}
   );
   gpc615_5 gpc5275 (
      {stage1_31[175], stage1_31[176], stage1_31[177], stage1_31[178], stage1_31[179]},
      {stage1_32[114]},
      {stage1_33[157], stage1_33[158], stage1_33[159], stage1_33[160], stage1_33[161], stage1_33[162]},
      {stage2_35[27],stage2_34[42],stage2_33[48],stage2_32[58],stage2_31[90]}
   );
   gpc615_5 gpc5276 (
      {stage1_31[180], stage1_31[181], stage1_31[182], stage1_31[183], stage1_31[184]},
      {stage1_32[115]},
      {stage1_33[163], stage1_33[164], stage1_33[165], stage1_33[166], stage1_33[167], stage1_33[168]},
      {stage2_35[28],stage2_34[43],stage2_33[49],stage2_32[59],stage2_31[91]}
   );
   gpc615_5 gpc5277 (
      {stage1_31[185], stage1_31[186], stage1_31[187], stage1_31[188], stage1_31[189]},
      {stage1_32[116]},
      {stage1_33[169], stage1_33[170], stage1_33[171], stage1_33[172], stage1_33[173], stage1_33[174]},
      {stage2_35[29],stage2_34[44],stage2_33[50],stage2_32[60],stage2_31[92]}
   );
   gpc615_5 gpc5278 (
      {stage1_31[190], stage1_31[191], stage1_31[192], stage1_31[193], stage1_31[194]},
      {stage1_32[117]},
      {stage1_33[175], stage1_33[176], stage1_33[177], stage1_33[178], stage1_33[179], stage1_33[180]},
      {stage2_35[30],stage2_34[45],stage2_33[51],stage2_32[61],stage2_31[93]}
   );
   gpc615_5 gpc5279 (
      {stage1_31[195], stage1_31[196], stage1_31[197], stage1_31[198], stage1_31[199]},
      {stage1_32[118]},
      {stage1_33[181], stage1_33[182], stage1_33[183], stage1_33[184], stage1_33[185], stage1_33[186]},
      {stage2_35[31],stage2_34[46],stage2_33[52],stage2_32[62],stage2_31[94]}
   );
   gpc615_5 gpc5280 (
      {stage1_31[200], stage1_31[201], stage1_31[202], stage1_31[203], stage1_31[204]},
      {stage1_32[119]},
      {stage1_33[187], stage1_33[188], stage1_33[189], stage1_33[190], stage1_33[191], stage1_33[192]},
      {stage2_35[32],stage2_34[47],stage2_33[53],stage2_32[63],stage2_31[95]}
   );
   gpc615_5 gpc5281 (
      {stage1_31[205], stage1_31[206], stage1_31[207], stage1_31[208], stage1_31[209]},
      {stage1_32[120]},
      {stage1_33[193], stage1_33[194], stage1_33[195], stage1_33[196], stage1_33[197], stage1_33[198]},
      {stage2_35[33],stage2_34[48],stage2_33[54],stage2_32[64],stage2_31[96]}
   );
   gpc615_5 gpc5282 (
      {stage1_31[210], stage1_31[211], stage1_31[212], stage1_31[213], stage1_31[214]},
      {stage1_32[121]},
      {stage1_33[199], stage1_33[200], stage1_33[201], stage1_33[202], stage1_33[203], stage1_33[204]},
      {stage2_35[34],stage2_34[49],stage2_33[55],stage2_32[65],stage2_31[97]}
   );
   gpc615_5 gpc5283 (
      {stage1_31[215], stage1_31[216], stage1_31[217], 1'b0, 1'b0},
      {stage1_32[122]},
      {stage1_33[205], stage1_33[206], stage1_33[207], stage1_33[208], stage1_33[209], stage1_33[210]},
      {stage2_35[35],stage2_34[50],stage2_33[56],stage2_32[66],stage2_31[98]}
   );
   gpc606_5 gpc5284 (
      {stage1_32[123], stage1_32[124], stage1_32[125], stage1_32[126], stage1_32[127], stage1_32[128]},
      {stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5], stage1_34[6]},
      {stage2_36[0],stage2_35[36],stage2_34[51],stage2_33[57],stage2_32[67]}
   );
   gpc606_5 gpc5285 (
      {stage1_32[129], stage1_32[130], stage1_32[131], stage1_32[132], stage1_32[133], stage1_32[134]},
      {stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11], stage1_34[12]},
      {stage2_36[1],stage2_35[37],stage2_34[52],stage2_33[58],stage2_32[68]}
   );
   gpc606_5 gpc5286 (
      {stage1_32[135], stage1_32[136], stage1_32[137], stage1_32[138], stage1_32[139], stage1_32[140]},
      {stage1_34[13], stage1_34[14], stage1_34[15], stage1_34[16], stage1_34[17], stage1_34[18]},
      {stage2_36[2],stage2_35[38],stage2_34[53],stage2_33[59],stage2_32[69]}
   );
   gpc606_5 gpc5287 (
      {stage1_32[141], stage1_32[142], stage1_32[143], stage1_32[144], stage1_32[145], stage1_32[146]},
      {stage1_34[19], stage1_34[20], stage1_34[21], stage1_34[22], stage1_34[23], stage1_34[24]},
      {stage2_36[3],stage2_35[39],stage2_34[54],stage2_33[60],stage2_32[70]}
   );
   gpc606_5 gpc5288 (
      {stage1_32[147], stage1_32[148], stage1_32[149], stage1_32[150], stage1_32[151], stage1_32[152]},
      {stage1_34[25], stage1_34[26], stage1_34[27], stage1_34[28], stage1_34[29], stage1_34[30]},
      {stage2_36[4],stage2_35[40],stage2_34[55],stage2_33[61],stage2_32[71]}
   );
   gpc606_5 gpc5289 (
      {stage1_32[153], stage1_32[154], stage1_32[155], stage1_32[156], stage1_32[157], stage1_32[158]},
      {stage1_34[31], stage1_34[32], stage1_34[33], stage1_34[34], stage1_34[35], stage1_34[36]},
      {stage2_36[5],stage2_35[41],stage2_34[56],stage2_33[62],stage2_32[72]}
   );
   gpc606_5 gpc5290 (
      {stage1_32[159], stage1_32[160], stage1_32[161], stage1_32[162], stage1_32[163], stage1_32[164]},
      {stage1_34[37], stage1_34[38], stage1_34[39], stage1_34[40], stage1_34[41], stage1_34[42]},
      {stage2_36[6],stage2_35[42],stage2_34[57],stage2_33[63],stage2_32[73]}
   );
   gpc606_5 gpc5291 (
      {stage1_32[165], stage1_32[166], stage1_32[167], stage1_32[168], stage1_32[169], stage1_32[170]},
      {stage1_34[43], stage1_34[44], stage1_34[45], stage1_34[46], stage1_34[47], stage1_34[48]},
      {stage2_36[7],stage2_35[43],stage2_34[58],stage2_33[64],stage2_32[74]}
   );
   gpc606_5 gpc5292 (
      {stage1_32[171], stage1_32[172], stage1_32[173], stage1_32[174], stage1_32[175], stage1_32[176]},
      {stage1_34[49], stage1_34[50], stage1_34[51], stage1_34[52], stage1_34[53], stage1_34[54]},
      {stage2_36[8],stage2_35[44],stage2_34[59],stage2_33[65],stage2_32[75]}
   );
   gpc606_5 gpc5293 (
      {stage1_32[177], stage1_32[178], stage1_32[179], stage1_32[180], stage1_32[181], stage1_32[182]},
      {stage1_34[55], stage1_34[56], stage1_34[57], stage1_34[58], stage1_34[59], stage1_34[60]},
      {stage2_36[9],stage2_35[45],stage2_34[60],stage2_33[66],stage2_32[76]}
   );
   gpc606_5 gpc5294 (
      {stage1_32[183], stage1_32[184], stage1_32[185], stage1_32[186], stage1_32[187], stage1_32[188]},
      {stage1_34[61], stage1_34[62], stage1_34[63], stage1_34[64], stage1_34[65], stage1_34[66]},
      {stage2_36[10],stage2_35[46],stage2_34[61],stage2_33[67],stage2_32[77]}
   );
   gpc2116_5 gpc5295 (
      {stage1_33[211], stage1_33[212], stage1_33[213], stage1_33[214], stage1_33[215], stage1_33[216]},
      {stage1_34[67]},
      {stage1_35[0]},
      {stage1_36[0], stage1_36[1]},
      {stage2_37[0],stage2_36[11],stage2_35[47],stage2_34[62],stage2_33[68]}
   );
   gpc606_5 gpc5296 (
      {stage1_33[217], stage1_33[218], stage1_33[219], stage1_33[220], stage1_33[221], stage1_33[222]},
      {stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5], stage1_35[6]},
      {stage2_37[1],stage2_36[12],stage2_35[48],stage2_34[63],stage2_33[69]}
   );
   gpc606_5 gpc5297 (
      {stage1_33[223], stage1_33[224], stage1_33[225], stage1_33[226], stage1_33[227], stage1_33[228]},
      {stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11], stage1_35[12]},
      {stage2_37[2],stage2_36[13],stage2_35[49],stage2_34[64],stage2_33[70]}
   );
   gpc606_5 gpc5298 (
      {stage1_33[229], stage1_33[230], stage1_33[231], stage1_33[232], stage1_33[233], stage1_33[234]},
      {stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17], stage1_35[18]},
      {stage2_37[3],stage2_36[14],stage2_35[50],stage2_34[65],stage2_33[71]}
   );
   gpc606_5 gpc5299 (
      {stage1_33[235], stage1_33[236], stage1_33[237], stage1_33[238], stage1_33[239], stage1_33[240]},
      {stage1_35[19], stage1_35[20], stage1_35[21], stage1_35[22], stage1_35[23], stage1_35[24]},
      {stage2_37[4],stage2_36[15],stage2_35[51],stage2_34[66],stage2_33[72]}
   );
   gpc606_5 gpc5300 (
      {stage1_33[241], stage1_33[242], stage1_33[243], stage1_33[244], stage1_33[245], stage1_33[246]},
      {stage1_35[25], stage1_35[26], stage1_35[27], stage1_35[28], stage1_35[29], stage1_35[30]},
      {stage2_37[5],stage2_36[16],stage2_35[52],stage2_34[67],stage2_33[73]}
   );
   gpc606_5 gpc5301 (
      {stage1_33[247], stage1_33[248], stage1_33[249], stage1_33[250], stage1_33[251], stage1_33[252]},
      {stage1_35[31], stage1_35[32], stage1_35[33], stage1_35[34], stage1_35[35], stage1_35[36]},
      {stage2_37[6],stage2_36[17],stage2_35[53],stage2_34[68],stage2_33[74]}
   );
   gpc606_5 gpc5302 (
      {stage1_33[253], stage1_33[254], stage1_33[255], stage1_33[256], stage1_33[257], stage1_33[258]},
      {stage1_35[37], stage1_35[38], stage1_35[39], stage1_35[40], stage1_35[41], stage1_35[42]},
      {stage2_37[7],stage2_36[18],stage2_35[54],stage2_34[69],stage2_33[75]}
   );
   gpc606_5 gpc5303 (
      {stage1_34[68], stage1_34[69], stage1_34[70], stage1_34[71], stage1_34[72], stage1_34[73]},
      {stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5], stage1_36[6], stage1_36[7]},
      {stage2_38[0],stage2_37[8],stage2_36[19],stage2_35[55],stage2_34[70]}
   );
   gpc606_5 gpc5304 (
      {stage1_34[74], stage1_34[75], stage1_34[76], stage1_34[77], stage1_34[78], stage1_34[79]},
      {stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11], stage1_36[12], stage1_36[13]},
      {stage2_38[1],stage2_37[9],stage2_36[20],stage2_35[56],stage2_34[71]}
   );
   gpc606_5 gpc5305 (
      {stage1_34[80], stage1_34[81], stage1_34[82], stage1_34[83], stage1_34[84], stage1_34[85]},
      {stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17], stage1_36[18], stage1_36[19]},
      {stage2_38[2],stage2_37[10],stage2_36[21],stage2_35[57],stage2_34[72]}
   );
   gpc606_5 gpc5306 (
      {stage1_34[86], stage1_34[87], stage1_34[88], stage1_34[89], stage1_34[90], stage1_34[91]},
      {stage1_36[20], stage1_36[21], stage1_36[22], stage1_36[23], stage1_36[24], stage1_36[25]},
      {stage2_38[3],stage2_37[11],stage2_36[22],stage2_35[58],stage2_34[73]}
   );
   gpc606_5 gpc5307 (
      {stage1_34[92], stage1_34[93], stage1_34[94], stage1_34[95], stage1_34[96], stage1_34[97]},
      {stage1_36[26], stage1_36[27], stage1_36[28], stage1_36[29], stage1_36[30], stage1_36[31]},
      {stage2_38[4],stage2_37[12],stage2_36[23],stage2_35[59],stage2_34[74]}
   );
   gpc606_5 gpc5308 (
      {stage1_34[98], stage1_34[99], stage1_34[100], stage1_34[101], stage1_34[102], stage1_34[103]},
      {stage1_36[32], stage1_36[33], stage1_36[34], stage1_36[35], stage1_36[36], stage1_36[37]},
      {stage2_38[5],stage2_37[13],stage2_36[24],stage2_35[60],stage2_34[75]}
   );
   gpc606_5 gpc5309 (
      {stage1_34[104], stage1_34[105], stage1_34[106], stage1_34[107], stage1_34[108], stage1_34[109]},
      {stage1_36[38], stage1_36[39], stage1_36[40], stage1_36[41], stage1_36[42], stage1_36[43]},
      {stage2_38[6],stage2_37[14],stage2_36[25],stage2_35[61],stage2_34[76]}
   );
   gpc606_5 gpc5310 (
      {stage1_34[110], stage1_34[111], stage1_34[112], stage1_34[113], stage1_34[114], stage1_34[115]},
      {stage1_36[44], stage1_36[45], stage1_36[46], stage1_36[47], stage1_36[48], stage1_36[49]},
      {stage2_38[7],stage2_37[15],stage2_36[26],stage2_35[62],stage2_34[77]}
   );
   gpc606_5 gpc5311 (
      {stage1_34[116], stage1_34[117], stage1_34[118], stage1_34[119], stage1_34[120], stage1_34[121]},
      {stage1_36[50], stage1_36[51], stage1_36[52], stage1_36[53], stage1_36[54], stage1_36[55]},
      {stage2_38[8],stage2_37[16],stage2_36[27],stage2_35[63],stage2_34[78]}
   );
   gpc606_5 gpc5312 (
      {stage1_34[122], stage1_34[123], stage1_34[124], stage1_34[125], stage1_34[126], stage1_34[127]},
      {stage1_36[56], stage1_36[57], stage1_36[58], stage1_36[59], stage1_36[60], stage1_36[61]},
      {stage2_38[9],stage2_37[17],stage2_36[28],stage2_35[64],stage2_34[79]}
   );
   gpc606_5 gpc5313 (
      {stage1_34[128], stage1_34[129], stage1_34[130], stage1_34[131], stage1_34[132], stage1_34[133]},
      {stage1_36[62], stage1_36[63], stage1_36[64], stage1_36[65], stage1_36[66], stage1_36[67]},
      {stage2_38[10],stage2_37[18],stage2_36[29],stage2_35[65],stage2_34[80]}
   );
   gpc606_5 gpc5314 (
      {stage1_34[134], stage1_34[135], stage1_34[136], stage1_34[137], stage1_34[138], stage1_34[139]},
      {stage1_36[68], stage1_36[69], stage1_36[70], stage1_36[71], stage1_36[72], stage1_36[73]},
      {stage2_38[11],stage2_37[19],stage2_36[30],stage2_35[66],stage2_34[81]}
   );
   gpc615_5 gpc5315 (
      {stage1_35[43], stage1_35[44], stage1_35[45], stage1_35[46], stage1_35[47]},
      {stage1_36[74]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[12],stage2_37[20],stage2_36[31],stage2_35[67]}
   );
   gpc615_5 gpc5316 (
      {stage1_35[48], stage1_35[49], stage1_35[50], stage1_35[51], stage1_35[52]},
      {stage1_36[75]},
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage2_39[1],stage2_38[13],stage2_37[21],stage2_36[32],stage2_35[68]}
   );
   gpc615_5 gpc5317 (
      {stage1_35[53], stage1_35[54], stage1_35[55], stage1_35[56], stage1_35[57]},
      {stage1_36[76]},
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage2_39[2],stage2_38[14],stage2_37[22],stage2_36[33],stage2_35[69]}
   );
   gpc615_5 gpc5318 (
      {stage1_35[58], stage1_35[59], stage1_35[60], stage1_35[61], stage1_35[62]},
      {stage1_36[77]},
      {stage1_37[18], stage1_37[19], stage1_37[20], stage1_37[21], stage1_37[22], stage1_37[23]},
      {stage2_39[3],stage2_38[15],stage2_37[23],stage2_36[34],stage2_35[70]}
   );
   gpc615_5 gpc5319 (
      {stage1_35[63], stage1_35[64], stage1_35[65], stage1_35[66], stage1_35[67]},
      {stage1_36[78]},
      {stage1_37[24], stage1_37[25], stage1_37[26], stage1_37[27], stage1_37[28], stage1_37[29]},
      {stage2_39[4],stage2_38[16],stage2_37[24],stage2_36[35],stage2_35[71]}
   );
   gpc615_5 gpc5320 (
      {stage1_35[68], stage1_35[69], stage1_35[70], stage1_35[71], stage1_35[72]},
      {stage1_36[79]},
      {stage1_37[30], stage1_37[31], stage1_37[32], stage1_37[33], stage1_37[34], stage1_37[35]},
      {stage2_39[5],stage2_38[17],stage2_37[25],stage2_36[36],stage2_35[72]}
   );
   gpc615_5 gpc5321 (
      {stage1_35[73], stage1_35[74], stage1_35[75], stage1_35[76], stage1_35[77]},
      {stage1_36[80]},
      {stage1_37[36], stage1_37[37], stage1_37[38], stage1_37[39], stage1_37[40], stage1_37[41]},
      {stage2_39[6],stage2_38[18],stage2_37[26],stage2_36[37],stage2_35[73]}
   );
   gpc615_5 gpc5322 (
      {stage1_35[78], stage1_35[79], stage1_35[80], stage1_35[81], stage1_35[82]},
      {stage1_36[81]},
      {stage1_37[42], stage1_37[43], stage1_37[44], stage1_37[45], stage1_37[46], stage1_37[47]},
      {stage2_39[7],stage2_38[19],stage2_37[27],stage2_36[38],stage2_35[74]}
   );
   gpc615_5 gpc5323 (
      {stage1_35[83], stage1_35[84], stage1_35[85], stage1_35[86], stage1_35[87]},
      {stage1_36[82]},
      {stage1_37[48], stage1_37[49], stage1_37[50], stage1_37[51], stage1_37[52], stage1_37[53]},
      {stage2_39[8],stage2_38[20],stage2_37[28],stage2_36[39],stage2_35[75]}
   );
   gpc615_5 gpc5324 (
      {stage1_35[88], stage1_35[89], stage1_35[90], stage1_35[91], stage1_35[92]},
      {stage1_36[83]},
      {stage1_37[54], stage1_37[55], stage1_37[56], stage1_37[57], stage1_37[58], stage1_37[59]},
      {stage2_39[9],stage2_38[21],stage2_37[29],stage2_36[40],stage2_35[76]}
   );
   gpc615_5 gpc5325 (
      {stage1_35[93], stage1_35[94], stage1_35[95], stage1_35[96], stage1_35[97]},
      {stage1_36[84]},
      {stage1_37[60], stage1_37[61], stage1_37[62], stage1_37[63], stage1_37[64], stage1_37[65]},
      {stage2_39[10],stage2_38[22],stage2_37[30],stage2_36[41],stage2_35[77]}
   );
   gpc615_5 gpc5326 (
      {stage1_35[98], stage1_35[99], stage1_35[100], stage1_35[101], stage1_35[102]},
      {stage1_36[85]},
      {stage1_37[66], stage1_37[67], stage1_37[68], stage1_37[69], stage1_37[70], stage1_37[71]},
      {stage2_39[11],stage2_38[23],stage2_37[31],stage2_36[42],stage2_35[78]}
   );
   gpc615_5 gpc5327 (
      {stage1_35[103], stage1_35[104], stage1_35[105], stage1_35[106], stage1_35[107]},
      {stage1_36[86]},
      {stage1_37[72], stage1_37[73], stage1_37[74], stage1_37[75], stage1_37[76], stage1_37[77]},
      {stage2_39[12],stage2_38[24],stage2_37[32],stage2_36[43],stage2_35[79]}
   );
   gpc615_5 gpc5328 (
      {stage1_35[108], stage1_35[109], stage1_35[110], stage1_35[111], stage1_35[112]},
      {stage1_36[87]},
      {stage1_37[78], stage1_37[79], stage1_37[80], stage1_37[81], stage1_37[82], stage1_37[83]},
      {stage2_39[13],stage2_38[25],stage2_37[33],stage2_36[44],stage2_35[80]}
   );
   gpc615_5 gpc5329 (
      {stage1_35[113], stage1_35[114], stage1_35[115], stage1_35[116], stage1_35[117]},
      {stage1_36[88]},
      {stage1_37[84], stage1_37[85], stage1_37[86], stage1_37[87], stage1_37[88], stage1_37[89]},
      {stage2_39[14],stage2_38[26],stage2_37[34],stage2_36[45],stage2_35[81]}
   );
   gpc615_5 gpc5330 (
      {stage1_35[118], stage1_35[119], stage1_35[120], stage1_35[121], stage1_35[122]},
      {stage1_36[89]},
      {stage1_37[90], stage1_37[91], stage1_37[92], stage1_37[93], stage1_37[94], stage1_37[95]},
      {stage2_39[15],stage2_38[27],stage2_37[35],stage2_36[46],stage2_35[82]}
   );
   gpc615_5 gpc5331 (
      {stage1_35[123], stage1_35[124], stage1_35[125], stage1_35[126], stage1_35[127]},
      {stage1_36[90]},
      {stage1_37[96], stage1_37[97], stage1_37[98], stage1_37[99], stage1_37[100], stage1_37[101]},
      {stage2_39[16],stage2_38[28],stage2_37[36],stage2_36[47],stage2_35[83]}
   );
   gpc615_5 gpc5332 (
      {stage1_35[128], stage1_35[129], stage1_35[130], stage1_35[131], stage1_35[132]},
      {stage1_36[91]},
      {stage1_37[102], stage1_37[103], stage1_37[104], stage1_37[105], stage1_37[106], stage1_37[107]},
      {stage2_39[17],stage2_38[29],stage2_37[37],stage2_36[48],stage2_35[84]}
   );
   gpc615_5 gpc5333 (
      {stage1_35[133], stage1_35[134], stage1_35[135], stage1_35[136], stage1_35[137]},
      {stage1_36[92]},
      {stage1_37[108], stage1_37[109], stage1_37[110], stage1_37[111], stage1_37[112], stage1_37[113]},
      {stage2_39[18],stage2_38[30],stage2_37[38],stage2_36[49],stage2_35[85]}
   );
   gpc615_5 gpc5334 (
      {stage1_35[138], stage1_35[139], stage1_35[140], stage1_35[141], stage1_35[142]},
      {stage1_36[93]},
      {stage1_37[114], stage1_37[115], stage1_37[116], stage1_37[117], stage1_37[118], stage1_37[119]},
      {stage2_39[19],stage2_38[31],stage2_37[39],stage2_36[50],stage2_35[86]}
   );
   gpc615_5 gpc5335 (
      {stage1_35[143], stage1_35[144], stage1_35[145], stage1_35[146], stage1_35[147]},
      {stage1_36[94]},
      {stage1_37[120], stage1_37[121], stage1_37[122], stage1_37[123], stage1_37[124], stage1_37[125]},
      {stage2_39[20],stage2_38[32],stage2_37[40],stage2_36[51],stage2_35[87]}
   );
   gpc615_5 gpc5336 (
      {stage1_35[148], stage1_35[149], stage1_35[150], stage1_35[151], stage1_35[152]},
      {stage1_36[95]},
      {stage1_37[126], stage1_37[127], stage1_37[128], stage1_37[129], stage1_37[130], stage1_37[131]},
      {stage2_39[21],stage2_38[33],stage2_37[41],stage2_36[52],stage2_35[88]}
   );
   gpc615_5 gpc5337 (
      {stage1_35[153], stage1_35[154], stage1_35[155], stage1_35[156], stage1_35[157]},
      {stage1_36[96]},
      {stage1_37[132], stage1_37[133], stage1_37[134], stage1_37[135], stage1_37[136], stage1_37[137]},
      {stage2_39[22],stage2_38[34],stage2_37[42],stage2_36[53],stage2_35[89]}
   );
   gpc615_5 gpc5338 (
      {stage1_35[158], stage1_35[159], stage1_35[160], stage1_35[161], stage1_35[162]},
      {stage1_36[97]},
      {stage1_37[138], stage1_37[139], stage1_37[140], stage1_37[141], stage1_37[142], stage1_37[143]},
      {stage2_39[23],stage2_38[35],stage2_37[43],stage2_36[54],stage2_35[90]}
   );
   gpc615_5 gpc5339 (
      {stage1_35[163], stage1_35[164], stage1_35[165], stage1_35[166], stage1_35[167]},
      {stage1_36[98]},
      {stage1_37[144], stage1_37[145], stage1_37[146], stage1_37[147], stage1_37[148], stage1_37[149]},
      {stage2_39[24],stage2_38[36],stage2_37[44],stage2_36[55],stage2_35[91]}
   );
   gpc615_5 gpc5340 (
      {stage1_35[168], stage1_35[169], stage1_35[170], stage1_35[171], stage1_35[172]},
      {stage1_36[99]},
      {stage1_37[150], stage1_37[151], stage1_37[152], stage1_37[153], stage1_37[154], stage1_37[155]},
      {stage2_39[25],stage2_38[37],stage2_37[45],stage2_36[56],stage2_35[92]}
   );
   gpc615_5 gpc5341 (
      {stage1_35[173], stage1_35[174], stage1_35[175], stage1_35[176], stage1_35[177]},
      {stage1_36[100]},
      {stage1_37[156], stage1_37[157], stage1_37[158], stage1_37[159], stage1_37[160], stage1_37[161]},
      {stage2_39[26],stage2_38[38],stage2_37[46],stage2_36[57],stage2_35[93]}
   );
   gpc1406_5 gpc5342 (
      {stage1_36[101], stage1_36[102], stage1_36[103], stage1_36[104], stage1_36[105], stage1_36[106]},
      {stage1_38[0], stage1_38[1], stage1_38[2], stage1_38[3]},
      {stage1_39[0]},
      {stage2_40[0],stage2_39[27],stage2_38[39],stage2_37[47],stage2_36[58]}
   );
   gpc606_5 gpc5343 (
      {stage1_36[107], stage1_36[108], stage1_36[109], stage1_36[110], stage1_36[111], stage1_36[112]},
      {stage1_38[4], stage1_38[5], stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9]},
      {stage2_40[1],stage2_39[28],stage2_38[40],stage2_37[48],stage2_36[59]}
   );
   gpc606_5 gpc5344 (
      {stage1_36[113], stage1_36[114], stage1_36[115], stage1_36[116], stage1_36[117], stage1_36[118]},
      {stage1_38[10], stage1_38[11], stage1_38[12], stage1_38[13], stage1_38[14], stage1_38[15]},
      {stage2_40[2],stage2_39[29],stage2_38[41],stage2_37[49],stage2_36[60]}
   );
   gpc606_5 gpc5345 (
      {stage1_36[119], stage1_36[120], stage1_36[121], stage1_36[122], stage1_36[123], stage1_36[124]},
      {stage1_38[16], stage1_38[17], stage1_38[18], stage1_38[19], stage1_38[20], stage1_38[21]},
      {stage2_40[3],stage2_39[30],stage2_38[42],stage2_37[50],stage2_36[61]}
   );
   gpc606_5 gpc5346 (
      {stage1_36[125], stage1_36[126], stage1_36[127], stage1_36[128], stage1_36[129], stage1_36[130]},
      {stage1_38[22], stage1_38[23], stage1_38[24], stage1_38[25], stage1_38[26], stage1_38[27]},
      {stage2_40[4],stage2_39[31],stage2_38[43],stage2_37[51],stage2_36[62]}
   );
   gpc606_5 gpc5347 (
      {stage1_36[131], stage1_36[132], stage1_36[133], stage1_36[134], stage1_36[135], stage1_36[136]},
      {stage1_38[28], stage1_38[29], stage1_38[30], stage1_38[31], stage1_38[32], stage1_38[33]},
      {stage2_40[5],stage2_39[32],stage2_38[44],stage2_37[52],stage2_36[63]}
   );
   gpc606_5 gpc5348 (
      {stage1_36[137], stage1_36[138], stage1_36[139], stage1_36[140], stage1_36[141], stage1_36[142]},
      {stage1_38[34], stage1_38[35], stage1_38[36], stage1_38[37], stage1_38[38], stage1_38[39]},
      {stage2_40[6],stage2_39[33],stage2_38[45],stage2_37[53],stage2_36[64]}
   );
   gpc606_5 gpc5349 (
      {stage1_36[143], stage1_36[144], stage1_36[145], stage1_36[146], stage1_36[147], stage1_36[148]},
      {stage1_38[40], stage1_38[41], stage1_38[42], stage1_38[43], stage1_38[44], stage1_38[45]},
      {stage2_40[7],stage2_39[34],stage2_38[46],stage2_37[54],stage2_36[65]}
   );
   gpc606_5 gpc5350 (
      {stage1_36[149], stage1_36[150], stage1_36[151], stage1_36[152], stage1_36[153], stage1_36[154]},
      {stage1_38[46], stage1_38[47], stage1_38[48], stage1_38[49], stage1_38[50], stage1_38[51]},
      {stage2_40[8],stage2_39[35],stage2_38[47],stage2_37[55],stage2_36[66]}
   );
   gpc606_5 gpc5351 (
      {stage1_36[155], stage1_36[156], stage1_36[157], stage1_36[158], stage1_36[159], stage1_36[160]},
      {stage1_38[52], stage1_38[53], stage1_38[54], stage1_38[55], stage1_38[56], stage1_38[57]},
      {stage2_40[9],stage2_39[36],stage2_38[48],stage2_37[56],stage2_36[67]}
   );
   gpc606_5 gpc5352 (
      {stage1_36[161], stage1_36[162], stage1_36[163], stage1_36[164], stage1_36[165], stage1_36[166]},
      {stage1_38[58], stage1_38[59], stage1_38[60], stage1_38[61], stage1_38[62], stage1_38[63]},
      {stage2_40[10],stage2_39[37],stage2_38[49],stage2_37[57],stage2_36[68]}
   );
   gpc606_5 gpc5353 (
      {stage1_36[167], stage1_36[168], stage1_36[169], stage1_36[170], stage1_36[171], stage1_36[172]},
      {stage1_38[64], stage1_38[65], stage1_38[66], stage1_38[67], stage1_38[68], stage1_38[69]},
      {stage2_40[11],stage2_39[38],stage2_38[50],stage2_37[58],stage2_36[69]}
   );
   gpc606_5 gpc5354 (
      {stage1_36[173], stage1_36[174], stage1_36[175], stage1_36[176], stage1_36[177], stage1_36[178]},
      {stage1_38[70], stage1_38[71], stage1_38[72], stage1_38[73], stage1_38[74], stage1_38[75]},
      {stage2_40[12],stage2_39[39],stage2_38[51],stage2_37[59],stage2_36[70]}
   );
   gpc606_5 gpc5355 (
      {stage1_36[179], stage1_36[180], stage1_36[181], stage1_36[182], stage1_36[183], stage1_36[184]},
      {stage1_38[76], stage1_38[77], stage1_38[78], stage1_38[79], stage1_38[80], stage1_38[81]},
      {stage2_40[13],stage2_39[40],stage2_38[52],stage2_37[60],stage2_36[71]}
   );
   gpc606_5 gpc5356 (
      {stage1_36[185], stage1_36[186], stage1_36[187], stage1_36[188], stage1_36[189], stage1_36[190]},
      {stage1_38[82], stage1_38[83], stage1_38[84], stage1_38[85], stage1_38[86], stage1_38[87]},
      {stage2_40[14],stage2_39[41],stage2_38[53],stage2_37[61],stage2_36[72]}
   );
   gpc606_5 gpc5357 (
      {stage1_36[191], stage1_36[192], stage1_36[193], stage1_36[194], stage1_36[195], stage1_36[196]},
      {stage1_38[88], stage1_38[89], stage1_38[90], stage1_38[91], stage1_38[92], stage1_38[93]},
      {stage2_40[15],stage2_39[42],stage2_38[54],stage2_37[62],stage2_36[73]}
   );
   gpc606_5 gpc5358 (
      {stage1_36[197], stage1_36[198], stage1_36[199], stage1_36[200], stage1_36[201], 1'b0},
      {stage1_38[94], stage1_38[95], stage1_38[96], stage1_38[97], stage1_38[98], stage1_38[99]},
      {stage2_40[16],stage2_39[43],stage2_38[55],stage2_37[63],stage2_36[74]}
   );
   gpc606_5 gpc5359 (
      {stage1_37[162], stage1_37[163], stage1_37[164], stage1_37[165], stage1_37[166], stage1_37[167]},
      {stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5], stage1_39[6]},
      {stage2_41[0],stage2_40[17],stage2_39[44],stage2_38[56],stage2_37[64]}
   );
   gpc606_5 gpc5360 (
      {stage1_37[168], stage1_37[169], stage1_37[170], stage1_37[171], stage1_37[172], stage1_37[173]},
      {stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11], stage1_39[12]},
      {stage2_41[1],stage2_40[18],stage2_39[45],stage2_38[57],stage2_37[65]}
   );
   gpc606_5 gpc5361 (
      {stage1_37[174], stage1_37[175], stage1_37[176], stage1_37[177], stage1_37[178], stage1_37[179]},
      {stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17], stage1_39[18]},
      {stage2_41[2],stage2_40[19],stage2_39[46],stage2_38[58],stage2_37[66]}
   );
   gpc606_5 gpc5362 (
      {stage1_37[180], stage1_37[181], stage1_37[182], stage1_37[183], stage1_37[184], stage1_37[185]},
      {stage1_39[19], stage1_39[20], stage1_39[21], stage1_39[22], stage1_39[23], stage1_39[24]},
      {stage2_41[3],stage2_40[20],stage2_39[47],stage2_38[59],stage2_37[67]}
   );
   gpc606_5 gpc5363 (
      {stage1_37[186], stage1_37[187], stage1_37[188], stage1_37[189], stage1_37[190], stage1_37[191]},
      {stage1_39[25], stage1_39[26], stage1_39[27], stage1_39[28], stage1_39[29], stage1_39[30]},
      {stage2_41[4],stage2_40[21],stage2_39[48],stage2_38[60],stage2_37[68]}
   );
   gpc606_5 gpc5364 (
      {stage1_37[192], stage1_37[193], stage1_37[194], stage1_37[195], stage1_37[196], stage1_37[197]},
      {stage1_39[31], stage1_39[32], stage1_39[33], stage1_39[34], stage1_39[35], stage1_39[36]},
      {stage2_41[5],stage2_40[22],stage2_39[49],stage2_38[61],stage2_37[69]}
   );
   gpc606_5 gpc5365 (
      {stage1_37[198], stage1_37[199], stage1_37[200], stage1_37[201], stage1_37[202], stage1_37[203]},
      {stage1_39[37], stage1_39[38], stage1_39[39], stage1_39[40], stage1_39[41], stage1_39[42]},
      {stage2_41[6],stage2_40[23],stage2_39[50],stage2_38[62],stage2_37[70]}
   );
   gpc606_5 gpc5366 (
      {stage1_37[204], stage1_37[205], stage1_37[206], stage1_37[207], stage1_37[208], stage1_37[209]},
      {stage1_39[43], stage1_39[44], stage1_39[45], stage1_39[46], stage1_39[47], stage1_39[48]},
      {stage2_41[7],stage2_40[24],stage2_39[51],stage2_38[63],stage2_37[71]}
   );
   gpc606_5 gpc5367 (
      {stage1_37[210], stage1_37[211], stage1_37[212], stage1_37[213], stage1_37[214], stage1_37[215]},
      {stage1_39[49], stage1_39[50], stage1_39[51], stage1_39[52], stage1_39[53], stage1_39[54]},
      {stage2_41[8],stage2_40[25],stage2_39[52],stage2_38[64],stage2_37[72]}
   );
   gpc606_5 gpc5368 (
      {stage1_37[216], stage1_37[217], stage1_37[218], stage1_37[219], stage1_37[220], stage1_37[221]},
      {stage1_39[55], stage1_39[56], stage1_39[57], stage1_39[58], stage1_39[59], stage1_39[60]},
      {stage2_41[9],stage2_40[26],stage2_39[53],stage2_38[65],stage2_37[73]}
   );
   gpc606_5 gpc5369 (
      {stage1_37[222], stage1_37[223], stage1_37[224], stage1_37[225], stage1_37[226], stage1_37[227]},
      {stage1_39[61], stage1_39[62], stage1_39[63], stage1_39[64], stage1_39[65], stage1_39[66]},
      {stage2_41[10],stage2_40[27],stage2_39[54],stage2_38[66],stage2_37[74]}
   );
   gpc606_5 gpc5370 (
      {stage1_37[228], stage1_37[229], stage1_37[230], stage1_37[231], stage1_37[232], stage1_37[233]},
      {stage1_39[67], stage1_39[68], stage1_39[69], stage1_39[70], stage1_39[71], stage1_39[72]},
      {stage2_41[11],stage2_40[28],stage2_39[55],stage2_38[67],stage2_37[75]}
   );
   gpc606_5 gpc5371 (
      {stage1_37[234], stage1_37[235], stage1_37[236], stage1_37[237], stage1_37[238], stage1_37[239]},
      {stage1_39[73], stage1_39[74], stage1_39[75], stage1_39[76], stage1_39[77], stage1_39[78]},
      {stage2_41[12],stage2_40[29],stage2_39[56],stage2_38[68],stage2_37[76]}
   );
   gpc606_5 gpc5372 (
      {stage1_37[240], stage1_37[241], stage1_37[242], stage1_37[243], stage1_37[244], stage1_37[245]},
      {stage1_39[79], stage1_39[80], stage1_39[81], stage1_39[82], stage1_39[83], stage1_39[84]},
      {stage2_41[13],stage2_40[30],stage2_39[57],stage2_38[69],stage2_37[77]}
   );
   gpc606_5 gpc5373 (
      {stage1_37[246], stage1_37[247], stage1_37[248], stage1_37[249], stage1_37[250], stage1_37[251]},
      {stage1_39[85], stage1_39[86], stage1_39[87], stage1_39[88], stage1_39[89], stage1_39[90]},
      {stage2_41[14],stage2_40[31],stage2_39[58],stage2_38[70],stage2_37[78]}
   );
   gpc606_5 gpc5374 (
      {stage1_37[252], stage1_37[253], stage1_37[254], stage1_37[255], stage1_37[256], stage1_37[257]},
      {stage1_39[91], stage1_39[92], stage1_39[93], stage1_39[94], stage1_39[95], stage1_39[96]},
      {stage2_41[15],stage2_40[32],stage2_39[59],stage2_38[71],stage2_37[79]}
   );
   gpc606_5 gpc5375 (
      {stage1_37[258], stage1_37[259], stage1_37[260], stage1_37[261], stage1_37[262], stage1_37[263]},
      {stage1_39[97], stage1_39[98], stage1_39[99], stage1_39[100], stage1_39[101], stage1_39[102]},
      {stage2_41[16],stage2_40[33],stage2_39[60],stage2_38[72],stage2_37[80]}
   );
   gpc606_5 gpc5376 (
      {stage1_37[264], stage1_37[265], stage1_37[266], stage1_37[267], stage1_37[268], stage1_37[269]},
      {stage1_39[103], stage1_39[104], stage1_39[105], stage1_39[106], stage1_39[107], stage1_39[108]},
      {stage2_41[17],stage2_40[34],stage2_39[61],stage2_38[73],stage2_37[81]}
   );
   gpc606_5 gpc5377 (
      {stage1_37[270], stage1_37[271], stage1_37[272], stage1_37[273], stage1_37[274], stage1_37[275]},
      {stage1_39[109], stage1_39[110], stage1_39[111], stage1_39[112], stage1_39[113], stage1_39[114]},
      {stage2_41[18],stage2_40[35],stage2_39[62],stage2_38[74],stage2_37[82]}
   );
   gpc606_5 gpc5378 (
      {stage1_37[276], stage1_37[277], stage1_37[278], stage1_37[279], stage1_37[280], stage1_37[281]},
      {stage1_39[115], stage1_39[116], stage1_39[117], stage1_39[118], stage1_39[119], stage1_39[120]},
      {stage2_41[19],stage2_40[36],stage2_39[63],stage2_38[75],stage2_37[83]}
   );
   gpc606_5 gpc5379 (
      {stage1_37[282], stage1_37[283], stage1_37[284], stage1_37[285], stage1_37[286], stage1_37[287]},
      {stage1_39[121], stage1_39[122], stage1_39[123], stage1_39[124], stage1_39[125], stage1_39[126]},
      {stage2_41[20],stage2_40[37],stage2_39[64],stage2_38[76],stage2_37[84]}
   );
   gpc606_5 gpc5380 (
      {stage1_37[288], stage1_37[289], stage1_37[290], stage1_37[291], stage1_37[292], stage1_37[293]},
      {stage1_39[127], stage1_39[128], stage1_39[129], stage1_39[130], stage1_39[131], stage1_39[132]},
      {stage2_41[21],stage2_40[38],stage2_39[65],stage2_38[77],stage2_37[85]}
   );
   gpc606_5 gpc5381 (
      {stage1_37[294], stage1_37[295], stage1_37[296], stage1_37[297], stage1_37[298], stage1_37[299]},
      {stage1_39[133], stage1_39[134], stage1_39[135], stage1_39[136], stage1_39[137], stage1_39[138]},
      {stage2_41[22],stage2_40[39],stage2_39[66],stage2_38[78],stage2_37[86]}
   );
   gpc606_5 gpc5382 (
      {stage1_37[300], stage1_37[301], stage1_37[302], stage1_37[303], stage1_37[304], stage1_37[305]},
      {stage1_39[139], stage1_39[140], stage1_39[141], stage1_39[142], stage1_39[143], stage1_39[144]},
      {stage2_41[23],stage2_40[40],stage2_39[67],stage2_38[79],stage2_37[87]}
   );
   gpc606_5 gpc5383 (
      {stage1_38[100], stage1_38[101], stage1_38[102], stage1_38[103], stage1_38[104], stage1_38[105]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[24],stage2_40[41],stage2_39[68],stage2_38[80]}
   );
   gpc615_5 gpc5384 (
      {stage1_38[106], stage1_38[107], stage1_38[108], stage1_38[109], stage1_38[110]},
      {stage1_39[145]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[25],stage2_40[42],stage2_39[69],stage2_38[81]}
   );
   gpc615_5 gpc5385 (
      {stage1_38[111], stage1_38[112], stage1_38[113], stage1_38[114], stage1_38[115]},
      {stage1_39[146]},
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17]},
      {stage2_42[2],stage2_41[26],stage2_40[43],stage2_39[70],stage2_38[82]}
   );
   gpc615_5 gpc5386 (
      {stage1_38[116], stage1_38[117], stage1_38[118], stage1_38[119], stage1_38[120]},
      {stage1_39[147]},
      {stage1_40[18], stage1_40[19], stage1_40[20], stage1_40[21], stage1_40[22], stage1_40[23]},
      {stage2_42[3],stage2_41[27],stage2_40[44],stage2_39[71],stage2_38[83]}
   );
   gpc615_5 gpc5387 (
      {stage1_38[121], stage1_38[122], stage1_38[123], stage1_38[124], stage1_38[125]},
      {stage1_39[148]},
      {stage1_40[24], stage1_40[25], stage1_40[26], stage1_40[27], stage1_40[28], stage1_40[29]},
      {stage2_42[4],stage2_41[28],stage2_40[45],stage2_39[72],stage2_38[84]}
   );
   gpc615_5 gpc5388 (
      {stage1_38[126], stage1_38[127], stage1_38[128], stage1_38[129], stage1_38[130]},
      {stage1_39[149]},
      {stage1_40[30], stage1_40[31], stage1_40[32], stage1_40[33], stage1_40[34], stage1_40[35]},
      {stage2_42[5],stage2_41[29],stage2_40[46],stage2_39[73],stage2_38[85]}
   );
   gpc615_5 gpc5389 (
      {stage1_38[131], stage1_38[132], stage1_38[133], stage1_38[134], stage1_38[135]},
      {stage1_39[150]},
      {stage1_40[36], stage1_40[37], stage1_40[38], stage1_40[39], stage1_40[40], stage1_40[41]},
      {stage2_42[6],stage2_41[30],stage2_40[47],stage2_39[74],stage2_38[86]}
   );
   gpc615_5 gpc5390 (
      {stage1_38[136], stage1_38[137], stage1_38[138], stage1_38[139], stage1_38[140]},
      {stage1_39[151]},
      {stage1_40[42], stage1_40[43], stage1_40[44], stage1_40[45], stage1_40[46], stage1_40[47]},
      {stage2_42[7],stage2_41[31],stage2_40[48],stage2_39[75],stage2_38[87]}
   );
   gpc615_5 gpc5391 (
      {stage1_38[141], stage1_38[142], stage1_38[143], stage1_38[144], stage1_38[145]},
      {stage1_39[152]},
      {stage1_40[48], stage1_40[49], stage1_40[50], stage1_40[51], stage1_40[52], stage1_40[53]},
      {stage2_42[8],stage2_41[32],stage2_40[49],stage2_39[76],stage2_38[88]}
   );
   gpc615_5 gpc5392 (
      {stage1_38[146], stage1_38[147], stage1_38[148], stage1_38[149], stage1_38[150]},
      {stage1_39[153]},
      {stage1_40[54], stage1_40[55], stage1_40[56], stage1_40[57], stage1_40[58], stage1_40[59]},
      {stage2_42[9],stage2_41[33],stage2_40[50],stage2_39[77],stage2_38[89]}
   );
   gpc615_5 gpc5393 (
      {stage1_38[151], stage1_38[152], stage1_38[153], stage1_38[154], stage1_38[155]},
      {stage1_39[154]},
      {stage1_40[60], stage1_40[61], stage1_40[62], stage1_40[63], stage1_40[64], stage1_40[65]},
      {stage2_42[10],stage2_41[34],stage2_40[51],stage2_39[78],stage2_38[90]}
   );
   gpc615_5 gpc5394 (
      {stage1_38[156], stage1_38[157], stage1_38[158], stage1_38[159], stage1_38[160]},
      {stage1_39[155]},
      {stage1_40[66], stage1_40[67], stage1_40[68], stage1_40[69], stage1_40[70], stage1_40[71]},
      {stage2_42[11],stage2_41[35],stage2_40[52],stage2_39[79],stage2_38[91]}
   );
   gpc615_5 gpc5395 (
      {stage1_38[161], stage1_38[162], stage1_38[163], stage1_38[164], stage1_38[165]},
      {stage1_39[156]},
      {stage1_40[72], stage1_40[73], stage1_40[74], stage1_40[75], stage1_40[76], stage1_40[77]},
      {stage2_42[12],stage2_41[36],stage2_40[53],stage2_39[80],stage2_38[92]}
   );
   gpc615_5 gpc5396 (
      {stage1_38[166], stage1_38[167], stage1_38[168], stage1_38[169], stage1_38[170]},
      {stage1_39[157]},
      {stage1_40[78], stage1_40[79], stage1_40[80], stage1_40[81], stage1_40[82], stage1_40[83]},
      {stage2_42[13],stage2_41[37],stage2_40[54],stage2_39[81],stage2_38[93]}
   );
   gpc615_5 gpc5397 (
      {stage1_38[171], stage1_38[172], stage1_38[173], stage1_38[174], stage1_38[175]},
      {stage1_39[158]},
      {stage1_40[84], stage1_40[85], stage1_40[86], stage1_40[87], stage1_40[88], stage1_40[89]},
      {stage2_42[14],stage2_41[38],stage2_40[55],stage2_39[82],stage2_38[94]}
   );
   gpc615_5 gpc5398 (
      {stage1_38[176], stage1_38[177], stage1_38[178], stage1_38[179], stage1_38[180]},
      {stage1_39[159]},
      {stage1_40[90], stage1_40[91], stage1_40[92], stage1_40[93], stage1_40[94], stage1_40[95]},
      {stage2_42[15],stage2_41[39],stage2_40[56],stage2_39[83],stage2_38[95]}
   );
   gpc615_5 gpc5399 (
      {stage1_38[181], stage1_38[182], stage1_38[183], stage1_38[184], stage1_38[185]},
      {stage1_39[160]},
      {stage1_40[96], stage1_40[97], stage1_40[98], stage1_40[99], stage1_40[100], stage1_40[101]},
      {stage2_42[16],stage2_41[40],stage2_40[57],stage2_39[84],stage2_38[96]}
   );
   gpc615_5 gpc5400 (
      {stage1_38[186], stage1_38[187], stage1_38[188], stage1_38[189], stage1_38[190]},
      {stage1_39[161]},
      {stage1_40[102], stage1_40[103], stage1_40[104], stage1_40[105], stage1_40[106], stage1_40[107]},
      {stage2_42[17],stage2_41[41],stage2_40[58],stage2_39[85],stage2_38[97]}
   );
   gpc615_5 gpc5401 (
      {stage1_38[191], stage1_38[192], stage1_38[193], stage1_38[194], stage1_38[195]},
      {stage1_39[162]},
      {stage1_40[108], stage1_40[109], stage1_40[110], stage1_40[111], stage1_40[112], stage1_40[113]},
      {stage2_42[18],stage2_41[42],stage2_40[59],stage2_39[86],stage2_38[98]}
   );
   gpc615_5 gpc5402 (
      {stage1_38[196], stage1_38[197], stage1_38[198], stage1_38[199], stage1_38[200]},
      {stage1_39[163]},
      {stage1_40[114], stage1_40[115], stage1_40[116], stage1_40[117], stage1_40[118], stage1_40[119]},
      {stage2_42[19],stage2_41[43],stage2_40[60],stage2_39[87],stage2_38[99]}
   );
   gpc615_5 gpc5403 (
      {stage1_38[201], stage1_38[202], stage1_38[203], stage1_38[204], stage1_38[205]},
      {stage1_39[164]},
      {stage1_40[120], stage1_40[121], stage1_40[122], stage1_40[123], stage1_40[124], stage1_40[125]},
      {stage2_42[20],stage2_41[44],stage2_40[61],stage2_39[88],stage2_38[100]}
   );
   gpc615_5 gpc5404 (
      {stage1_38[206], stage1_38[207], stage1_38[208], stage1_38[209], stage1_38[210]},
      {stage1_39[165]},
      {stage1_40[126], stage1_40[127], stage1_40[128], stage1_40[129], stage1_40[130], stage1_40[131]},
      {stage2_42[21],stage2_41[45],stage2_40[62],stage2_39[89],stage2_38[101]}
   );
   gpc615_5 gpc5405 (
      {stage1_38[211], stage1_38[212], stage1_38[213], stage1_38[214], stage1_38[215]},
      {stage1_39[166]},
      {stage1_40[132], stage1_40[133], stage1_40[134], stage1_40[135], stage1_40[136], stage1_40[137]},
      {stage2_42[22],stage2_41[46],stage2_40[63],stage2_39[90],stage2_38[102]}
   );
   gpc615_5 gpc5406 (
      {stage1_38[216], stage1_38[217], stage1_38[218], stage1_38[219], stage1_38[220]},
      {stage1_39[167]},
      {stage1_40[138], stage1_40[139], stage1_40[140], stage1_40[141], stage1_40[142], stage1_40[143]},
      {stage2_42[23],stage2_41[47],stage2_40[64],stage2_39[91],stage2_38[103]}
   );
   gpc615_5 gpc5407 (
      {stage1_38[221], stage1_38[222], stage1_38[223], stage1_38[224], stage1_38[225]},
      {stage1_39[168]},
      {stage1_40[144], stage1_40[145], stage1_40[146], stage1_40[147], stage1_40[148], stage1_40[149]},
      {stage2_42[24],stage2_41[48],stage2_40[65],stage2_39[92],stage2_38[104]}
   );
   gpc615_5 gpc5408 (
      {stage1_38[226], stage1_38[227], stage1_38[228], stage1_38[229], stage1_38[230]},
      {stage1_39[169]},
      {stage1_40[150], stage1_40[151], stage1_40[152], stage1_40[153], stage1_40[154], stage1_40[155]},
      {stage2_42[25],stage2_41[49],stage2_40[66],stage2_39[93],stage2_38[105]}
   );
   gpc606_5 gpc5409 (
      {stage1_40[156], stage1_40[157], stage1_40[158], stage1_40[159], stage1_40[160], stage1_40[161]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[0],stage2_42[26],stage2_41[50],stage2_40[67]}
   );
   gpc606_5 gpc5410 (
      {stage1_40[162], stage1_40[163], stage1_40[164], stage1_40[165], stage1_40[166], stage1_40[167]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[1],stage2_42[27],stage2_41[51],stage2_40[68]}
   );
   gpc606_5 gpc5411 (
      {stage1_40[168], stage1_40[169], stage1_40[170], stage1_40[171], stage1_40[172], stage1_40[173]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[2],stage2_42[28],stage2_41[52],stage2_40[69]}
   );
   gpc606_5 gpc5412 (
      {stage1_40[174], stage1_40[175], stage1_40[176], stage1_40[177], stage1_40[178], stage1_40[179]},
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage2_44[3],stage2_43[3],stage2_42[29],stage2_41[53],stage2_40[70]}
   );
   gpc606_5 gpc5413 (
      {stage1_40[180], stage1_40[181], stage1_40[182], stage1_40[183], stage1_40[184], stage1_40[185]},
      {stage1_42[24], stage1_42[25], stage1_42[26], stage1_42[27], stage1_42[28], stage1_42[29]},
      {stage2_44[4],stage2_43[4],stage2_42[30],stage2_41[54],stage2_40[71]}
   );
   gpc606_5 gpc5414 (
      {stage1_40[186], stage1_40[187], stage1_40[188], stage1_40[189], stage1_40[190], stage1_40[191]},
      {stage1_42[30], stage1_42[31], stage1_42[32], stage1_42[33], stage1_42[34], stage1_42[35]},
      {stage2_44[5],stage2_43[5],stage2_42[31],stage2_41[55],stage2_40[72]}
   );
   gpc606_5 gpc5415 (
      {stage1_40[192], stage1_40[193], stage1_40[194], stage1_40[195], stage1_40[196], stage1_40[197]},
      {stage1_42[36], stage1_42[37], stage1_42[38], stage1_42[39], stage1_42[40], stage1_42[41]},
      {stage2_44[6],stage2_43[6],stage2_42[32],stage2_41[56],stage2_40[73]}
   );
   gpc606_5 gpc5416 (
      {stage1_40[198], stage1_40[199], stage1_40[200], stage1_40[201], stage1_40[202], stage1_40[203]},
      {stage1_42[42], stage1_42[43], stage1_42[44], stage1_42[45], stage1_42[46], stage1_42[47]},
      {stage2_44[7],stage2_43[7],stage2_42[33],stage2_41[57],stage2_40[74]}
   );
   gpc606_5 gpc5417 (
      {stage1_40[204], stage1_40[205], stage1_40[206], stage1_40[207], stage1_40[208], stage1_40[209]},
      {stage1_42[48], stage1_42[49], stage1_42[50], stage1_42[51], stage1_42[52], stage1_42[53]},
      {stage2_44[8],stage2_43[8],stage2_42[34],stage2_41[58],stage2_40[75]}
   );
   gpc606_5 gpc5418 (
      {stage1_40[210], stage1_40[211], stage1_40[212], stage1_40[213], stage1_40[214], stage1_40[215]},
      {stage1_42[54], stage1_42[55], stage1_42[56], stage1_42[57], stage1_42[58], stage1_42[59]},
      {stage2_44[9],stage2_43[9],stage2_42[35],stage2_41[59],stage2_40[76]}
   );
   gpc615_5 gpc5419 (
      {stage1_40[216], stage1_40[217], stage1_40[218], stage1_40[219], stage1_40[220]},
      {stage1_41[0]},
      {stage1_42[60], stage1_42[61], stage1_42[62], stage1_42[63], stage1_42[64], stage1_42[65]},
      {stage2_44[10],stage2_43[10],stage2_42[36],stage2_41[60],stage2_40[77]}
   );
   gpc615_5 gpc5420 (
      {stage1_40[221], stage1_40[222], stage1_40[223], stage1_40[224], stage1_40[225]},
      {stage1_41[1]},
      {stage1_42[66], stage1_42[67], stage1_42[68], stage1_42[69], stage1_42[70], stage1_42[71]},
      {stage2_44[11],stage2_43[11],stage2_42[37],stage2_41[61],stage2_40[78]}
   );
   gpc615_5 gpc5421 (
      {stage1_40[226], stage1_40[227], stage1_40[228], stage1_40[229], stage1_40[230]},
      {stage1_41[2]},
      {stage1_42[72], stage1_42[73], stage1_42[74], stage1_42[75], stage1_42[76], stage1_42[77]},
      {stage2_44[12],stage2_43[12],stage2_42[38],stage2_41[62],stage2_40[79]}
   );
   gpc615_5 gpc5422 (
      {stage1_40[231], stage1_40[232], stage1_40[233], stage1_40[234], stage1_40[235]},
      {stage1_41[3]},
      {stage1_42[78], stage1_42[79], stage1_42[80], stage1_42[81], stage1_42[82], stage1_42[83]},
      {stage2_44[13],stage2_43[13],stage2_42[39],stage2_41[63],stage2_40[80]}
   );
   gpc615_5 gpc5423 (
      {stage1_40[236], stage1_40[237], stage1_40[238], stage1_40[239], stage1_40[240]},
      {stage1_41[4]},
      {stage1_42[84], stage1_42[85], stage1_42[86], stage1_42[87], stage1_42[88], stage1_42[89]},
      {stage2_44[14],stage2_43[14],stage2_42[40],stage2_41[64],stage2_40[81]}
   );
   gpc615_5 gpc5424 (
      {stage1_40[241], stage1_40[242], stage1_40[243], stage1_40[244], stage1_40[245]},
      {stage1_41[5]},
      {stage1_42[90], stage1_42[91], stage1_42[92], stage1_42[93], stage1_42[94], stage1_42[95]},
      {stage2_44[15],stage2_43[15],stage2_42[41],stage2_41[65],stage2_40[82]}
   );
   gpc615_5 gpc5425 (
      {stage1_40[246], stage1_40[247], stage1_40[248], stage1_40[249], stage1_40[250]},
      {stage1_41[6]},
      {stage1_42[96], stage1_42[97], stage1_42[98], stage1_42[99], stage1_42[100], stage1_42[101]},
      {stage2_44[16],stage2_43[16],stage2_42[42],stage2_41[66],stage2_40[83]}
   );
   gpc615_5 gpc5426 (
      {stage1_40[251], stage1_40[252], stage1_40[253], stage1_40[254], stage1_40[255]},
      {stage1_41[7]},
      {stage1_42[102], stage1_42[103], stage1_42[104], stage1_42[105], stage1_42[106], stage1_42[107]},
      {stage2_44[17],stage2_43[17],stage2_42[43],stage2_41[67],stage2_40[84]}
   );
   gpc615_5 gpc5427 (
      {stage1_40[256], stage1_40[257], stage1_40[258], stage1_40[259], stage1_40[260]},
      {stage1_41[8]},
      {stage1_42[108], stage1_42[109], stage1_42[110], stage1_42[111], stage1_42[112], stage1_42[113]},
      {stage2_44[18],stage2_43[18],stage2_42[44],stage2_41[68],stage2_40[85]}
   );
   gpc615_5 gpc5428 (
      {stage1_40[261], stage1_40[262], stage1_40[263], stage1_40[264], stage1_40[265]},
      {stage1_41[9]},
      {stage1_42[114], stage1_42[115], stage1_42[116], stage1_42[117], stage1_42[118], stage1_42[119]},
      {stage2_44[19],stage2_43[19],stage2_42[45],stage2_41[69],stage2_40[86]}
   );
   gpc615_5 gpc5429 (
      {stage1_40[266], stage1_40[267], stage1_40[268], stage1_40[269], stage1_40[270]},
      {stage1_41[10]},
      {stage1_42[120], stage1_42[121], stage1_42[122], stage1_42[123], stage1_42[124], stage1_42[125]},
      {stage2_44[20],stage2_43[20],stage2_42[46],stage2_41[70],stage2_40[87]}
   );
   gpc615_5 gpc5430 (
      {stage1_40[271], stage1_40[272], stage1_40[273], stage1_40[274], stage1_40[275]},
      {stage1_41[11]},
      {stage1_42[126], stage1_42[127], stage1_42[128], stage1_42[129], stage1_42[130], stage1_42[131]},
      {stage2_44[21],stage2_43[21],stage2_42[47],stage2_41[71],stage2_40[88]}
   );
   gpc615_5 gpc5431 (
      {stage1_40[276], stage1_40[277], stage1_40[278], stage1_40[279], stage1_40[280]},
      {stage1_41[12]},
      {stage1_42[132], stage1_42[133], stage1_42[134], stage1_42[135], stage1_42[136], stage1_42[137]},
      {stage2_44[22],stage2_43[22],stage2_42[48],stage2_41[72],stage2_40[89]}
   );
   gpc606_5 gpc5432 (
      {stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17], stage1_41[18]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[23],stage2_43[23],stage2_42[49],stage2_41[73]}
   );
   gpc606_5 gpc5433 (
      {stage1_41[19], stage1_41[20], stage1_41[21], stage1_41[22], stage1_41[23], stage1_41[24]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[24],stage2_43[24],stage2_42[50],stage2_41[74]}
   );
   gpc606_5 gpc5434 (
      {stage1_41[25], stage1_41[26], stage1_41[27], stage1_41[28], stage1_41[29], stage1_41[30]},
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16], stage1_43[17]},
      {stage2_45[2],stage2_44[25],stage2_43[25],stage2_42[51],stage2_41[75]}
   );
   gpc606_5 gpc5435 (
      {stage1_41[31], stage1_41[32], stage1_41[33], stage1_41[34], stage1_41[35], stage1_41[36]},
      {stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21], stage1_43[22], stage1_43[23]},
      {stage2_45[3],stage2_44[26],stage2_43[26],stage2_42[52],stage2_41[76]}
   );
   gpc606_5 gpc5436 (
      {stage1_41[37], stage1_41[38], stage1_41[39], stage1_41[40], stage1_41[41], stage1_41[42]},
      {stage1_43[24], stage1_43[25], stage1_43[26], stage1_43[27], stage1_43[28], stage1_43[29]},
      {stage2_45[4],stage2_44[27],stage2_43[27],stage2_42[53],stage2_41[77]}
   );
   gpc615_5 gpc5437 (
      {stage1_41[43], stage1_41[44], stage1_41[45], stage1_41[46], stage1_41[47]},
      {stage1_42[138]},
      {stage1_43[30], stage1_43[31], stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35]},
      {stage2_45[5],stage2_44[28],stage2_43[28],stage2_42[54],stage2_41[78]}
   );
   gpc615_5 gpc5438 (
      {stage1_41[48], stage1_41[49], stage1_41[50], stage1_41[51], stage1_41[52]},
      {stage1_42[139]},
      {stage1_43[36], stage1_43[37], stage1_43[38], stage1_43[39], stage1_43[40], stage1_43[41]},
      {stage2_45[6],stage2_44[29],stage2_43[29],stage2_42[55],stage2_41[79]}
   );
   gpc615_5 gpc5439 (
      {stage1_41[53], stage1_41[54], stage1_41[55], stage1_41[56], stage1_41[57]},
      {stage1_42[140]},
      {stage1_43[42], stage1_43[43], stage1_43[44], stage1_43[45], stage1_43[46], stage1_43[47]},
      {stage2_45[7],stage2_44[30],stage2_43[30],stage2_42[56],stage2_41[80]}
   );
   gpc615_5 gpc5440 (
      {stage1_41[58], stage1_41[59], stage1_41[60], stage1_41[61], stage1_41[62]},
      {stage1_42[141]},
      {stage1_43[48], stage1_43[49], stage1_43[50], stage1_43[51], stage1_43[52], stage1_43[53]},
      {stage2_45[8],stage2_44[31],stage2_43[31],stage2_42[57],stage2_41[81]}
   );
   gpc615_5 gpc5441 (
      {stage1_41[63], stage1_41[64], stage1_41[65], stage1_41[66], stage1_41[67]},
      {stage1_42[142]},
      {stage1_43[54], stage1_43[55], stage1_43[56], stage1_43[57], stage1_43[58], stage1_43[59]},
      {stage2_45[9],stage2_44[32],stage2_43[32],stage2_42[58],stage2_41[82]}
   );
   gpc615_5 gpc5442 (
      {stage1_41[68], stage1_41[69], stage1_41[70], stage1_41[71], stage1_41[72]},
      {stage1_42[143]},
      {stage1_43[60], stage1_43[61], stage1_43[62], stage1_43[63], stage1_43[64], stage1_43[65]},
      {stage2_45[10],stage2_44[33],stage2_43[33],stage2_42[59],stage2_41[83]}
   );
   gpc615_5 gpc5443 (
      {stage1_41[73], stage1_41[74], stage1_41[75], stage1_41[76], stage1_41[77]},
      {stage1_42[144]},
      {stage1_43[66], stage1_43[67], stage1_43[68], stage1_43[69], stage1_43[70], stage1_43[71]},
      {stage2_45[11],stage2_44[34],stage2_43[34],stage2_42[60],stage2_41[84]}
   );
   gpc615_5 gpc5444 (
      {stage1_41[78], stage1_41[79], stage1_41[80], stage1_41[81], stage1_41[82]},
      {stage1_42[145]},
      {stage1_43[72], stage1_43[73], stage1_43[74], stage1_43[75], stage1_43[76], stage1_43[77]},
      {stage2_45[12],stage2_44[35],stage2_43[35],stage2_42[61],stage2_41[85]}
   );
   gpc615_5 gpc5445 (
      {stage1_41[83], stage1_41[84], stage1_41[85], stage1_41[86], stage1_41[87]},
      {stage1_42[146]},
      {stage1_43[78], stage1_43[79], stage1_43[80], stage1_43[81], stage1_43[82], stage1_43[83]},
      {stage2_45[13],stage2_44[36],stage2_43[36],stage2_42[62],stage2_41[86]}
   );
   gpc615_5 gpc5446 (
      {stage1_41[88], stage1_41[89], stage1_41[90], stage1_41[91], stage1_41[92]},
      {stage1_42[147]},
      {stage1_43[84], stage1_43[85], stage1_43[86], stage1_43[87], stage1_43[88], stage1_43[89]},
      {stage2_45[14],stage2_44[37],stage2_43[37],stage2_42[63],stage2_41[87]}
   );
   gpc615_5 gpc5447 (
      {stage1_41[93], stage1_41[94], stage1_41[95], stage1_41[96], stage1_41[97]},
      {stage1_42[148]},
      {stage1_43[90], stage1_43[91], stage1_43[92], stage1_43[93], stage1_43[94], stage1_43[95]},
      {stage2_45[15],stage2_44[38],stage2_43[38],stage2_42[64],stage2_41[88]}
   );
   gpc615_5 gpc5448 (
      {stage1_41[98], stage1_41[99], stage1_41[100], stage1_41[101], stage1_41[102]},
      {stage1_42[149]},
      {stage1_43[96], stage1_43[97], stage1_43[98], stage1_43[99], stage1_43[100], stage1_43[101]},
      {stage2_45[16],stage2_44[39],stage2_43[39],stage2_42[65],stage2_41[89]}
   );
   gpc615_5 gpc5449 (
      {stage1_41[103], stage1_41[104], stage1_41[105], stage1_41[106], stage1_41[107]},
      {stage1_42[150]},
      {stage1_43[102], stage1_43[103], stage1_43[104], stage1_43[105], stage1_43[106], stage1_43[107]},
      {stage2_45[17],stage2_44[40],stage2_43[40],stage2_42[66],stage2_41[90]}
   );
   gpc615_5 gpc5450 (
      {stage1_41[108], stage1_41[109], stage1_41[110], stage1_41[111], stage1_41[112]},
      {stage1_42[151]},
      {stage1_43[108], stage1_43[109], stage1_43[110], stage1_43[111], stage1_43[112], stage1_43[113]},
      {stage2_45[18],stage2_44[41],stage2_43[41],stage2_42[67],stage2_41[91]}
   );
   gpc615_5 gpc5451 (
      {stage1_41[113], stage1_41[114], stage1_41[115], stage1_41[116], stage1_41[117]},
      {stage1_42[152]},
      {stage1_43[114], stage1_43[115], stage1_43[116], stage1_43[117], stage1_43[118], stage1_43[119]},
      {stage2_45[19],stage2_44[42],stage2_43[42],stage2_42[68],stage2_41[92]}
   );
   gpc615_5 gpc5452 (
      {stage1_41[118], stage1_41[119], stage1_41[120], stage1_41[121], stage1_41[122]},
      {stage1_42[153]},
      {stage1_43[120], stage1_43[121], stage1_43[122], stage1_43[123], stage1_43[124], stage1_43[125]},
      {stage2_45[20],stage2_44[43],stage2_43[43],stage2_42[69],stage2_41[93]}
   );
   gpc615_5 gpc5453 (
      {stage1_41[123], stage1_41[124], stage1_41[125], stage1_41[126], stage1_41[127]},
      {stage1_42[154]},
      {stage1_43[126], stage1_43[127], stage1_43[128], stage1_43[129], stage1_43[130], stage1_43[131]},
      {stage2_45[21],stage2_44[44],stage2_43[44],stage2_42[70],stage2_41[94]}
   );
   gpc615_5 gpc5454 (
      {stage1_41[128], stage1_41[129], stage1_41[130], stage1_41[131], stage1_41[132]},
      {stage1_42[155]},
      {stage1_43[132], stage1_43[133], stage1_43[134], stage1_43[135], stage1_43[136], stage1_43[137]},
      {stage2_45[22],stage2_44[45],stage2_43[45],stage2_42[71],stage2_41[95]}
   );
   gpc615_5 gpc5455 (
      {stage1_41[133], stage1_41[134], stage1_41[135], stage1_41[136], stage1_41[137]},
      {stage1_42[156]},
      {stage1_43[138], stage1_43[139], stage1_43[140], stage1_43[141], stage1_43[142], stage1_43[143]},
      {stage2_45[23],stage2_44[46],stage2_43[46],stage2_42[72],stage2_41[96]}
   );
   gpc615_5 gpc5456 (
      {stage1_41[138], stage1_41[139], stage1_41[140], stage1_41[141], stage1_41[142]},
      {stage1_42[157]},
      {stage1_43[144], stage1_43[145], stage1_43[146], stage1_43[147], stage1_43[148], stage1_43[149]},
      {stage2_45[24],stage2_44[47],stage2_43[47],stage2_42[73],stage2_41[97]}
   );
   gpc615_5 gpc5457 (
      {stage1_41[143], stage1_41[144], stage1_41[145], stage1_41[146], stage1_41[147]},
      {stage1_42[158]},
      {stage1_43[150], stage1_43[151], stage1_43[152], stage1_43[153], stage1_43[154], stage1_43[155]},
      {stage2_45[25],stage2_44[48],stage2_43[48],stage2_42[74],stage2_41[98]}
   );
   gpc615_5 gpc5458 (
      {stage1_41[148], stage1_41[149], stage1_41[150], stage1_41[151], stage1_41[152]},
      {stage1_42[159]},
      {stage1_43[156], stage1_43[157], stage1_43[158], stage1_43[159], stage1_43[160], stage1_43[161]},
      {stage2_45[26],stage2_44[49],stage2_43[49],stage2_42[75],stage2_41[99]}
   );
   gpc615_5 gpc5459 (
      {stage1_41[153], stage1_41[154], stage1_41[155], stage1_41[156], stage1_41[157]},
      {stage1_42[160]},
      {stage1_43[162], stage1_43[163], stage1_43[164], stage1_43[165], stage1_43[166], stage1_43[167]},
      {stage2_45[27],stage2_44[50],stage2_43[50],stage2_42[76],stage2_41[100]}
   );
   gpc615_5 gpc5460 (
      {stage1_41[158], stage1_41[159], stage1_41[160], stage1_41[161], stage1_41[162]},
      {stage1_42[161]},
      {stage1_43[168], stage1_43[169], stage1_43[170], stage1_43[171], stage1_43[172], stage1_43[173]},
      {stage2_45[28],stage2_44[51],stage2_43[51],stage2_42[77],stage2_41[101]}
   );
   gpc615_5 gpc5461 (
      {stage1_41[163], stage1_41[164], stage1_41[165], stage1_41[166], stage1_41[167]},
      {stage1_42[162]},
      {stage1_43[174], stage1_43[175], stage1_43[176], stage1_43[177], stage1_43[178], stage1_43[179]},
      {stage2_45[29],stage2_44[52],stage2_43[52],stage2_42[78],stage2_41[102]}
   );
   gpc615_5 gpc5462 (
      {stage1_42[163], stage1_42[164], stage1_42[165], stage1_42[166], stage1_42[167]},
      {stage1_43[180]},
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage2_46[0],stage2_45[30],stage2_44[53],stage2_43[53],stage2_42[79]}
   );
   gpc615_5 gpc5463 (
      {stage1_43[181], stage1_43[182], stage1_43[183], stage1_43[184], stage1_43[185]},
      {stage1_44[6]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[1],stage2_45[31],stage2_44[54],stage2_43[54]}
   );
   gpc615_5 gpc5464 (
      {stage1_43[186], stage1_43[187], stage1_43[188], stage1_43[189], stage1_43[190]},
      {stage1_44[7]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[2],stage2_45[32],stage2_44[55],stage2_43[55]}
   );
   gpc615_5 gpc5465 (
      {stage1_43[191], stage1_43[192], stage1_43[193], stage1_43[194], stage1_43[195]},
      {stage1_44[8]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[3],stage2_45[33],stage2_44[56],stage2_43[56]}
   );
   gpc615_5 gpc5466 (
      {stage1_43[196], stage1_43[197], stage1_43[198], stage1_43[199], stage1_43[200]},
      {stage1_44[9]},
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage2_47[3],stage2_46[4],stage2_45[34],stage2_44[57],stage2_43[57]}
   );
   gpc615_5 gpc5467 (
      {stage1_43[201], stage1_43[202], stage1_43[203], stage1_43[204], stage1_43[205]},
      {stage1_44[10]},
      {stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27], stage1_45[28], stage1_45[29]},
      {stage2_47[4],stage2_46[5],stage2_45[35],stage2_44[58],stage2_43[58]}
   );
   gpc615_5 gpc5468 (
      {stage1_43[206], stage1_43[207], stage1_43[208], stage1_43[209], stage1_43[210]},
      {stage1_44[11]},
      {stage1_45[30], stage1_45[31], stage1_45[32], stage1_45[33], stage1_45[34], stage1_45[35]},
      {stage2_47[5],stage2_46[6],stage2_45[36],stage2_44[59],stage2_43[59]}
   );
   gpc615_5 gpc5469 (
      {stage1_43[211], stage1_43[212], stage1_43[213], stage1_43[214], stage1_43[215]},
      {stage1_44[12]},
      {stage1_45[36], stage1_45[37], stage1_45[38], stage1_45[39], stage1_45[40], stage1_45[41]},
      {stage2_47[6],stage2_46[7],stage2_45[37],stage2_44[60],stage2_43[60]}
   );
   gpc615_5 gpc5470 (
      {stage1_43[216], stage1_43[217], stage1_43[218], stage1_43[219], stage1_43[220]},
      {stage1_44[13]},
      {stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45], stage1_45[46], stage1_45[47]},
      {stage2_47[7],stage2_46[8],stage2_45[38],stage2_44[61],stage2_43[61]}
   );
   gpc615_5 gpc5471 (
      {stage1_43[221], stage1_43[222], stage1_43[223], stage1_43[224], stage1_43[225]},
      {stage1_44[14]},
      {stage1_45[48], stage1_45[49], stage1_45[50], stage1_45[51], stage1_45[52], stage1_45[53]},
      {stage2_47[8],stage2_46[9],stage2_45[39],stage2_44[62],stage2_43[62]}
   );
   gpc615_5 gpc5472 (
      {stage1_43[226], stage1_43[227], stage1_43[228], stage1_43[229], stage1_43[230]},
      {stage1_44[15]},
      {stage1_45[54], stage1_45[55], stage1_45[56], stage1_45[57], stage1_45[58], stage1_45[59]},
      {stage2_47[9],stage2_46[10],stage2_45[40],stage2_44[63],stage2_43[63]}
   );
   gpc615_5 gpc5473 (
      {stage1_43[231], stage1_43[232], stage1_43[233], stage1_43[234], stage1_43[235]},
      {stage1_44[16]},
      {stage1_45[60], stage1_45[61], stage1_45[62], stage1_45[63], stage1_45[64], stage1_45[65]},
      {stage2_47[10],stage2_46[11],stage2_45[41],stage2_44[64],stage2_43[64]}
   );
   gpc615_5 gpc5474 (
      {stage1_43[236], stage1_43[237], stage1_43[238], stage1_43[239], stage1_43[240]},
      {stage1_44[17]},
      {stage1_45[66], stage1_45[67], stage1_45[68], stage1_45[69], stage1_45[70], stage1_45[71]},
      {stage2_47[11],stage2_46[12],stage2_45[42],stage2_44[65],stage2_43[65]}
   );
   gpc606_5 gpc5475 (
      {stage1_44[18], stage1_44[19], stage1_44[20], stage1_44[21], stage1_44[22], stage1_44[23]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[12],stage2_46[13],stage2_45[43],stage2_44[66]}
   );
   gpc606_5 gpc5476 (
      {stage1_44[24], stage1_44[25], stage1_44[26], stage1_44[27], stage1_44[28], stage1_44[29]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[13],stage2_46[14],stage2_45[44],stage2_44[67]}
   );
   gpc606_5 gpc5477 (
      {stage1_44[30], stage1_44[31], stage1_44[32], stage1_44[33], stage1_44[34], stage1_44[35]},
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16], stage1_46[17]},
      {stage2_48[2],stage2_47[14],stage2_46[15],stage2_45[45],stage2_44[68]}
   );
   gpc606_5 gpc5478 (
      {stage1_44[36], stage1_44[37], stage1_44[38], stage1_44[39], stage1_44[40], stage1_44[41]},
      {stage1_46[18], stage1_46[19], stage1_46[20], stage1_46[21], stage1_46[22], stage1_46[23]},
      {stage2_48[3],stage2_47[15],stage2_46[16],stage2_45[46],stage2_44[69]}
   );
   gpc606_5 gpc5479 (
      {stage1_44[42], stage1_44[43], stage1_44[44], stage1_44[45], stage1_44[46], stage1_44[47]},
      {stage1_46[24], stage1_46[25], stage1_46[26], stage1_46[27], stage1_46[28], stage1_46[29]},
      {stage2_48[4],stage2_47[16],stage2_46[17],stage2_45[47],stage2_44[70]}
   );
   gpc606_5 gpc5480 (
      {stage1_44[48], stage1_44[49], stage1_44[50], stage1_44[51], stage1_44[52], stage1_44[53]},
      {stage1_46[30], stage1_46[31], stage1_46[32], stage1_46[33], stage1_46[34], stage1_46[35]},
      {stage2_48[5],stage2_47[17],stage2_46[18],stage2_45[48],stage2_44[71]}
   );
   gpc606_5 gpc5481 (
      {stage1_44[54], stage1_44[55], stage1_44[56], stage1_44[57], stage1_44[58], stage1_44[59]},
      {stage1_46[36], stage1_46[37], stage1_46[38], stage1_46[39], stage1_46[40], stage1_46[41]},
      {stage2_48[6],stage2_47[18],stage2_46[19],stage2_45[49],stage2_44[72]}
   );
   gpc606_5 gpc5482 (
      {stage1_44[60], stage1_44[61], stage1_44[62], stage1_44[63], stage1_44[64], stage1_44[65]},
      {stage1_46[42], stage1_46[43], stage1_46[44], stage1_46[45], stage1_46[46], stage1_46[47]},
      {stage2_48[7],stage2_47[19],stage2_46[20],stage2_45[50],stage2_44[73]}
   );
   gpc606_5 gpc5483 (
      {stage1_44[66], stage1_44[67], stage1_44[68], stage1_44[69], stage1_44[70], stage1_44[71]},
      {stage1_46[48], stage1_46[49], stage1_46[50], stage1_46[51], stage1_46[52], stage1_46[53]},
      {stage2_48[8],stage2_47[20],stage2_46[21],stage2_45[51],stage2_44[74]}
   );
   gpc606_5 gpc5484 (
      {stage1_44[72], stage1_44[73], stage1_44[74], stage1_44[75], stage1_44[76], stage1_44[77]},
      {stage1_46[54], stage1_46[55], stage1_46[56], stage1_46[57], stage1_46[58], stage1_46[59]},
      {stage2_48[9],stage2_47[21],stage2_46[22],stage2_45[52],stage2_44[75]}
   );
   gpc606_5 gpc5485 (
      {stage1_44[78], stage1_44[79], stage1_44[80], stage1_44[81], stage1_44[82], stage1_44[83]},
      {stage1_46[60], stage1_46[61], stage1_46[62], stage1_46[63], stage1_46[64], stage1_46[65]},
      {stage2_48[10],stage2_47[22],stage2_46[23],stage2_45[53],stage2_44[76]}
   );
   gpc606_5 gpc5486 (
      {stage1_44[84], stage1_44[85], stage1_44[86], stage1_44[87], stage1_44[88], stage1_44[89]},
      {stage1_46[66], stage1_46[67], stage1_46[68], stage1_46[69], stage1_46[70], stage1_46[71]},
      {stage2_48[11],stage2_47[23],stage2_46[24],stage2_45[54],stage2_44[77]}
   );
   gpc606_5 gpc5487 (
      {stage1_44[90], stage1_44[91], stage1_44[92], stage1_44[93], stage1_44[94], stage1_44[95]},
      {stage1_46[72], stage1_46[73], stage1_46[74], stage1_46[75], stage1_46[76], stage1_46[77]},
      {stage2_48[12],stage2_47[24],stage2_46[25],stage2_45[55],stage2_44[78]}
   );
   gpc606_5 gpc5488 (
      {stage1_44[96], stage1_44[97], stage1_44[98], stage1_44[99], stage1_44[100], stage1_44[101]},
      {stage1_46[78], stage1_46[79], stage1_46[80], stage1_46[81], stage1_46[82], stage1_46[83]},
      {stage2_48[13],stage2_47[25],stage2_46[26],stage2_45[56],stage2_44[79]}
   );
   gpc606_5 gpc5489 (
      {stage1_44[102], stage1_44[103], stage1_44[104], stage1_44[105], stage1_44[106], stage1_44[107]},
      {stage1_46[84], stage1_46[85], stage1_46[86], stage1_46[87], stage1_46[88], stage1_46[89]},
      {stage2_48[14],stage2_47[26],stage2_46[27],stage2_45[57],stage2_44[80]}
   );
   gpc606_5 gpc5490 (
      {stage1_44[108], stage1_44[109], stage1_44[110], stage1_44[111], stage1_44[112], stage1_44[113]},
      {stage1_46[90], stage1_46[91], stage1_46[92], stage1_46[93], stage1_46[94], stage1_46[95]},
      {stage2_48[15],stage2_47[27],stage2_46[28],stage2_45[58],stage2_44[81]}
   );
   gpc606_5 gpc5491 (
      {stage1_44[114], stage1_44[115], stage1_44[116], stage1_44[117], stage1_44[118], stage1_44[119]},
      {stage1_46[96], stage1_46[97], stage1_46[98], stage1_46[99], stage1_46[100], stage1_46[101]},
      {stage2_48[16],stage2_47[28],stage2_46[29],stage2_45[59],stage2_44[82]}
   );
   gpc606_5 gpc5492 (
      {stage1_44[120], stage1_44[121], stage1_44[122], stage1_44[123], stage1_44[124], stage1_44[125]},
      {stage1_46[102], stage1_46[103], stage1_46[104], stage1_46[105], stage1_46[106], stage1_46[107]},
      {stage2_48[17],stage2_47[29],stage2_46[30],stage2_45[60],stage2_44[83]}
   );
   gpc606_5 gpc5493 (
      {stage1_44[126], stage1_44[127], stage1_44[128], stage1_44[129], stage1_44[130], stage1_44[131]},
      {stage1_46[108], stage1_46[109], stage1_46[110], stage1_46[111], stage1_46[112], stage1_46[113]},
      {stage2_48[18],stage2_47[30],stage2_46[31],stage2_45[61],stage2_44[84]}
   );
   gpc606_5 gpc5494 (
      {stage1_44[132], stage1_44[133], stage1_44[134], stage1_44[135], stage1_44[136], stage1_44[137]},
      {stage1_46[114], stage1_46[115], stage1_46[116], stage1_46[117], stage1_46[118], stage1_46[119]},
      {stage2_48[19],stage2_47[31],stage2_46[32],stage2_45[62],stage2_44[85]}
   );
   gpc606_5 gpc5495 (
      {stage1_44[138], stage1_44[139], stage1_44[140], stage1_44[141], stage1_44[142], stage1_44[143]},
      {stage1_46[120], stage1_46[121], stage1_46[122], stage1_46[123], stage1_46[124], stage1_46[125]},
      {stage2_48[20],stage2_47[32],stage2_46[33],stage2_45[63],stage2_44[86]}
   );
   gpc606_5 gpc5496 (
      {stage1_44[144], stage1_44[145], stage1_44[146], stage1_44[147], stage1_44[148], stage1_44[149]},
      {stage1_46[126], stage1_46[127], stage1_46[128], stage1_46[129], stage1_46[130], stage1_46[131]},
      {stage2_48[21],stage2_47[33],stage2_46[34],stage2_45[64],stage2_44[87]}
   );
   gpc606_5 gpc5497 (
      {stage1_44[150], stage1_44[151], stage1_44[152], stage1_44[153], stage1_44[154], stage1_44[155]},
      {stage1_46[132], stage1_46[133], stage1_46[134], stage1_46[135], stage1_46[136], stage1_46[137]},
      {stage2_48[22],stage2_47[34],stage2_46[35],stage2_45[65],stage2_44[88]}
   );
   gpc606_5 gpc5498 (
      {stage1_44[156], stage1_44[157], stage1_44[158], stage1_44[159], stage1_44[160], stage1_44[161]},
      {stage1_46[138], stage1_46[139], stage1_46[140], stage1_46[141], stage1_46[142], stage1_46[143]},
      {stage2_48[23],stage2_47[35],stage2_46[36],stage2_45[66],stage2_44[89]}
   );
   gpc606_5 gpc5499 (
      {stage1_44[162], stage1_44[163], stage1_44[164], stage1_44[165], stage1_44[166], stage1_44[167]},
      {stage1_46[144], stage1_46[145], stage1_46[146], stage1_46[147], stage1_46[148], stage1_46[149]},
      {stage2_48[24],stage2_47[36],stage2_46[37],stage2_45[67],stage2_44[90]}
   );
   gpc606_5 gpc5500 (
      {stage1_44[168], stage1_44[169], stage1_44[170], stage1_44[171], stage1_44[172], stage1_44[173]},
      {stage1_46[150], stage1_46[151], stage1_46[152], stage1_46[153], stage1_46[154], stage1_46[155]},
      {stage2_48[25],stage2_47[37],stage2_46[38],stage2_45[68],stage2_44[91]}
   );
   gpc606_5 gpc5501 (
      {stage1_44[174], stage1_44[175], stage1_44[176], stage1_44[177], stage1_44[178], stage1_44[179]},
      {stage1_46[156], stage1_46[157], stage1_46[158], stage1_46[159], stage1_46[160], stage1_46[161]},
      {stage2_48[26],stage2_47[38],stage2_46[39],stage2_45[69],stage2_44[92]}
   );
   gpc606_5 gpc5502 (
      {stage1_44[180], stage1_44[181], stage1_44[182], stage1_44[183], stage1_44[184], stage1_44[185]},
      {stage1_46[162], stage1_46[163], stage1_46[164], stage1_46[165], stage1_46[166], stage1_46[167]},
      {stage2_48[27],stage2_47[39],stage2_46[40],stage2_45[70],stage2_44[93]}
   );
   gpc606_5 gpc5503 (
      {stage1_44[186], stage1_44[187], stage1_44[188], stage1_44[189], stage1_44[190], stage1_44[191]},
      {stage1_46[168], stage1_46[169], stage1_46[170], stage1_46[171], stage1_46[172], stage1_46[173]},
      {stage2_48[28],stage2_47[40],stage2_46[41],stage2_45[71],stage2_44[94]}
   );
   gpc606_5 gpc5504 (
      {stage1_44[192], stage1_44[193], stage1_44[194], stage1_44[195], stage1_44[196], stage1_44[197]},
      {stage1_46[174], stage1_46[175], stage1_46[176], stage1_46[177], stage1_46[178], stage1_46[179]},
      {stage2_48[29],stage2_47[41],stage2_46[42],stage2_45[72],stage2_44[95]}
   );
   gpc606_5 gpc5505 (
      {stage1_44[198], stage1_44[199], stage1_44[200], stage1_44[201], stage1_44[202], stage1_44[203]},
      {stage1_46[180], stage1_46[181], stage1_46[182], stage1_46[183], stage1_46[184], stage1_46[185]},
      {stage2_48[30],stage2_47[42],stage2_46[43],stage2_45[73],stage2_44[96]}
   );
   gpc606_5 gpc5506 (
      {stage1_44[204], stage1_44[205], stage1_44[206], stage1_44[207], stage1_44[208], stage1_44[209]},
      {stage1_46[186], stage1_46[187], stage1_46[188], stage1_46[189], stage1_46[190], stage1_46[191]},
      {stage2_48[31],stage2_47[43],stage2_46[44],stage2_45[74],stage2_44[97]}
   );
   gpc606_5 gpc5507 (
      {stage1_44[210], stage1_44[211], stage1_44[212], stage1_44[213], stage1_44[214], stage1_44[215]},
      {stage1_46[192], stage1_46[193], stage1_46[194], stage1_46[195], stage1_46[196], stage1_46[197]},
      {stage2_48[32],stage2_47[44],stage2_46[45],stage2_45[75],stage2_44[98]}
   );
   gpc606_5 gpc5508 (
      {stage1_44[216], stage1_44[217], stage1_44[218], stage1_44[219], stage1_44[220], stage1_44[221]},
      {stage1_46[198], stage1_46[199], stage1_46[200], stage1_46[201], stage1_46[202], stage1_46[203]},
      {stage2_48[33],stage2_47[45],stage2_46[46],stage2_45[76],stage2_44[99]}
   );
   gpc606_5 gpc5509 (
      {stage1_44[222], stage1_44[223], stage1_44[224], stage1_44[225], stage1_44[226], stage1_44[227]},
      {stage1_46[204], stage1_46[205], stage1_46[206], stage1_46[207], stage1_46[208], stage1_46[209]},
      {stage2_48[34],stage2_47[46],stage2_46[47],stage2_45[77],stage2_44[100]}
   );
   gpc606_5 gpc5510 (
      {stage1_44[228], stage1_44[229], stage1_44[230], stage1_44[231], stage1_44[232], stage1_44[233]},
      {stage1_46[210], stage1_46[211], stage1_46[212], stage1_46[213], stage1_46[214], stage1_46[215]},
      {stage2_48[35],stage2_47[47],stage2_46[48],stage2_45[78],stage2_44[101]}
   );
   gpc606_5 gpc5511 (
      {stage1_44[234], stage1_44[235], stage1_44[236], stage1_44[237], stage1_44[238], stage1_44[239]},
      {stage1_46[216], stage1_46[217], stage1_46[218], stage1_46[219], stage1_46[220], stage1_46[221]},
      {stage2_48[36],stage2_47[48],stage2_46[49],stage2_45[79],stage2_44[102]}
   );
   gpc606_5 gpc5512 (
      {stage1_45[72], stage1_45[73], stage1_45[74], stage1_45[75], stage1_45[76], stage1_45[77]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[37],stage2_47[49],stage2_46[50],stage2_45[80]}
   );
   gpc606_5 gpc5513 (
      {stage1_45[78], stage1_45[79], stage1_45[80], stage1_45[81], stage1_45[82], stage1_45[83]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[38],stage2_47[50],stage2_46[51],stage2_45[81]}
   );
   gpc615_5 gpc5514 (
      {stage1_45[84], stage1_45[85], stage1_45[86], stage1_45[87], stage1_45[88]},
      {stage1_46[222]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[39],stage2_47[51],stage2_46[52],stage2_45[82]}
   );
   gpc615_5 gpc5515 (
      {stage1_45[89], stage1_45[90], stage1_45[91], stage1_45[92], stage1_45[93]},
      {stage1_46[223]},
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage2_49[3],stage2_48[40],stage2_47[52],stage2_46[53],stage2_45[83]}
   );
   gpc615_5 gpc5516 (
      {stage1_45[94], stage1_45[95], stage1_45[96], stage1_45[97], stage1_45[98]},
      {stage1_46[224]},
      {stage1_47[24], stage1_47[25], stage1_47[26], stage1_47[27], stage1_47[28], stage1_47[29]},
      {stage2_49[4],stage2_48[41],stage2_47[53],stage2_46[54],stage2_45[84]}
   );
   gpc615_5 gpc5517 (
      {stage1_45[99], stage1_45[100], stage1_45[101], stage1_45[102], stage1_45[103]},
      {stage1_46[225]},
      {stage1_47[30], stage1_47[31], stage1_47[32], stage1_47[33], stage1_47[34], stage1_47[35]},
      {stage2_49[5],stage2_48[42],stage2_47[54],stage2_46[55],stage2_45[85]}
   );
   gpc615_5 gpc5518 (
      {stage1_45[104], stage1_45[105], stage1_45[106], stage1_45[107], stage1_45[108]},
      {stage1_46[226]},
      {stage1_47[36], stage1_47[37], stage1_47[38], stage1_47[39], stage1_47[40], stage1_47[41]},
      {stage2_49[6],stage2_48[43],stage2_47[55],stage2_46[56],stage2_45[86]}
   );
   gpc615_5 gpc5519 (
      {stage1_45[109], stage1_45[110], stage1_45[111], stage1_45[112], stage1_45[113]},
      {stage1_46[227]},
      {stage1_47[42], stage1_47[43], stage1_47[44], stage1_47[45], stage1_47[46], stage1_47[47]},
      {stage2_49[7],stage2_48[44],stage2_47[56],stage2_46[57],stage2_45[87]}
   );
   gpc615_5 gpc5520 (
      {stage1_45[114], stage1_45[115], stage1_45[116], stage1_45[117], stage1_45[118]},
      {stage1_46[228]},
      {stage1_47[48], stage1_47[49], stage1_47[50], stage1_47[51], stage1_47[52], stage1_47[53]},
      {stage2_49[8],stage2_48[45],stage2_47[57],stage2_46[58],stage2_45[88]}
   );
   gpc615_5 gpc5521 (
      {stage1_45[119], stage1_45[120], stage1_45[121], stage1_45[122], stage1_45[123]},
      {stage1_46[229]},
      {stage1_47[54], stage1_47[55], stage1_47[56], stage1_47[57], stage1_47[58], stage1_47[59]},
      {stage2_49[9],stage2_48[46],stage2_47[58],stage2_46[59],stage2_45[89]}
   );
   gpc615_5 gpc5522 (
      {stage1_45[124], stage1_45[125], stage1_45[126], stage1_45[127], stage1_45[128]},
      {stage1_46[230]},
      {stage1_47[60], stage1_47[61], stage1_47[62], stage1_47[63], stage1_47[64], stage1_47[65]},
      {stage2_49[10],stage2_48[47],stage2_47[59],stage2_46[60],stage2_45[90]}
   );
   gpc615_5 gpc5523 (
      {stage1_45[129], stage1_45[130], stage1_45[131], stage1_45[132], stage1_45[133]},
      {stage1_46[231]},
      {stage1_47[66], stage1_47[67], stage1_47[68], stage1_47[69], stage1_47[70], stage1_47[71]},
      {stage2_49[11],stage2_48[48],stage2_47[60],stage2_46[61],stage2_45[91]}
   );
   gpc615_5 gpc5524 (
      {stage1_45[134], stage1_45[135], stage1_45[136], stage1_45[137], stage1_45[138]},
      {stage1_46[232]},
      {stage1_47[72], stage1_47[73], stage1_47[74], stage1_47[75], stage1_47[76], stage1_47[77]},
      {stage2_49[12],stage2_48[49],stage2_47[61],stage2_46[62],stage2_45[92]}
   );
   gpc615_5 gpc5525 (
      {stage1_45[139], stage1_45[140], stage1_45[141], stage1_45[142], stage1_45[143]},
      {stage1_46[233]},
      {stage1_47[78], stage1_47[79], stage1_47[80], stage1_47[81], stage1_47[82], stage1_47[83]},
      {stage2_49[13],stage2_48[50],stage2_47[62],stage2_46[63],stage2_45[93]}
   );
   gpc615_5 gpc5526 (
      {stage1_45[144], stage1_45[145], stage1_45[146], stage1_45[147], stage1_45[148]},
      {stage1_46[234]},
      {stage1_47[84], stage1_47[85], stage1_47[86], stage1_47[87], stage1_47[88], stage1_47[89]},
      {stage2_49[14],stage2_48[51],stage2_47[63],stage2_46[64],stage2_45[94]}
   );
   gpc615_5 gpc5527 (
      {stage1_45[149], stage1_45[150], stage1_45[151], stage1_45[152], stage1_45[153]},
      {stage1_46[235]},
      {stage1_47[90], stage1_47[91], stage1_47[92], stage1_47[93], stage1_47[94], stage1_47[95]},
      {stage2_49[15],stage2_48[52],stage2_47[64],stage2_46[65],stage2_45[95]}
   );
   gpc615_5 gpc5528 (
      {stage1_45[154], stage1_45[155], stage1_45[156], stage1_45[157], stage1_45[158]},
      {stage1_46[236]},
      {stage1_47[96], stage1_47[97], stage1_47[98], stage1_47[99], stage1_47[100], stage1_47[101]},
      {stage2_49[16],stage2_48[53],stage2_47[65],stage2_46[66],stage2_45[96]}
   );
   gpc615_5 gpc5529 (
      {stage1_45[159], stage1_45[160], stage1_45[161], stage1_45[162], stage1_45[163]},
      {stage1_46[237]},
      {stage1_47[102], stage1_47[103], stage1_47[104], stage1_47[105], stage1_47[106], stage1_47[107]},
      {stage2_49[17],stage2_48[54],stage2_47[66],stage2_46[67],stage2_45[97]}
   );
   gpc615_5 gpc5530 (
      {stage1_45[164], stage1_45[165], stage1_45[166], stage1_45[167], stage1_45[168]},
      {stage1_46[238]},
      {stage1_47[108], stage1_47[109], stage1_47[110], stage1_47[111], stage1_47[112], stage1_47[113]},
      {stage2_49[18],stage2_48[55],stage2_47[67],stage2_46[68],stage2_45[98]}
   );
   gpc615_5 gpc5531 (
      {stage1_45[169], stage1_45[170], stage1_45[171], stage1_45[172], stage1_45[173]},
      {stage1_46[239]},
      {stage1_47[114], stage1_47[115], stage1_47[116], stage1_47[117], stage1_47[118], stage1_47[119]},
      {stage2_49[19],stage2_48[56],stage2_47[68],stage2_46[69],stage2_45[99]}
   );
   gpc615_5 gpc5532 (
      {stage1_45[174], stage1_45[175], stage1_45[176], stage1_45[177], stage1_45[178]},
      {stage1_46[240]},
      {stage1_47[120], stage1_47[121], stage1_47[122], stage1_47[123], stage1_47[124], stage1_47[125]},
      {stage2_49[20],stage2_48[57],stage2_47[69],stage2_46[70],stage2_45[100]}
   );
   gpc615_5 gpc5533 (
      {stage1_45[179], stage1_45[180], stage1_45[181], stage1_45[182], stage1_45[183]},
      {stage1_46[241]},
      {stage1_47[126], stage1_47[127], stage1_47[128], stage1_47[129], stage1_47[130], stage1_47[131]},
      {stage2_49[21],stage2_48[58],stage2_47[70],stage2_46[71],stage2_45[101]}
   );
   gpc615_5 gpc5534 (
      {stage1_45[184], stage1_45[185], stage1_45[186], stage1_45[187], stage1_45[188]},
      {stage1_46[242]},
      {stage1_47[132], stage1_47[133], stage1_47[134], stage1_47[135], stage1_47[136], stage1_47[137]},
      {stage2_49[22],stage2_48[59],stage2_47[71],stage2_46[72],stage2_45[102]}
   );
   gpc615_5 gpc5535 (
      {stage1_45[189], stage1_45[190], stage1_45[191], stage1_45[192], stage1_45[193]},
      {stage1_46[243]},
      {stage1_47[138], stage1_47[139], stage1_47[140], stage1_47[141], stage1_47[142], stage1_47[143]},
      {stage2_49[23],stage2_48[60],stage2_47[72],stage2_46[73],stage2_45[103]}
   );
   gpc615_5 gpc5536 (
      {stage1_45[194], stage1_45[195], stage1_45[196], stage1_45[197], stage1_45[198]},
      {stage1_46[244]},
      {stage1_47[144], stage1_47[145], stage1_47[146], stage1_47[147], stage1_47[148], stage1_47[149]},
      {stage2_49[24],stage2_48[61],stage2_47[73],stage2_46[74],stage2_45[104]}
   );
   gpc615_5 gpc5537 (
      {stage1_46[245], stage1_46[246], stage1_46[247], stage1_46[248], stage1_46[249]},
      {stage1_47[150]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[25],stage2_48[62],stage2_47[74],stage2_46[75]}
   );
   gpc615_5 gpc5538 (
      {stage1_46[250], stage1_46[251], stage1_46[252], stage1_46[253], stage1_46[254]},
      {stage1_47[151]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[26],stage2_48[63],stage2_47[75],stage2_46[76]}
   );
   gpc615_5 gpc5539 (
      {stage1_46[255], stage1_46[256], stage1_46[257], stage1_46[258], stage1_46[259]},
      {stage1_47[152]},
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage2_50[2],stage2_49[27],stage2_48[64],stage2_47[76],stage2_46[77]}
   );
   gpc615_5 gpc5540 (
      {stage1_46[260], stage1_46[261], stage1_46[262], stage1_46[263], stage1_46[264]},
      {stage1_47[153]},
      {stage1_48[18], stage1_48[19], stage1_48[20], stage1_48[21], stage1_48[22], stage1_48[23]},
      {stage2_50[3],stage2_49[28],stage2_48[65],stage2_47[77],stage2_46[78]}
   );
   gpc615_5 gpc5541 (
      {stage1_46[265], stage1_46[266], stage1_46[267], stage1_46[268], stage1_46[269]},
      {stage1_47[154]},
      {stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27], stage1_48[28], stage1_48[29]},
      {stage2_50[4],stage2_49[29],stage2_48[66],stage2_47[78],stage2_46[79]}
   );
   gpc615_5 gpc5542 (
      {stage1_46[270], stage1_46[271], stage1_46[272], stage1_46[273], stage1_46[274]},
      {stage1_47[155]},
      {stage1_48[30], stage1_48[31], stage1_48[32], stage1_48[33], stage1_48[34], stage1_48[35]},
      {stage2_50[5],stage2_49[30],stage2_48[67],stage2_47[79],stage2_46[80]}
   );
   gpc615_5 gpc5543 (
      {stage1_46[275], stage1_46[276], stage1_46[277], stage1_46[278], stage1_46[279]},
      {stage1_47[156]},
      {stage1_48[36], stage1_48[37], stage1_48[38], stage1_48[39], stage1_48[40], stage1_48[41]},
      {stage2_50[6],stage2_49[31],stage2_48[68],stage2_47[80],stage2_46[81]}
   );
   gpc615_5 gpc5544 (
      {stage1_46[280], stage1_46[281], stage1_46[282], stage1_46[283], stage1_46[284]},
      {stage1_47[157]},
      {stage1_48[42], stage1_48[43], stage1_48[44], stage1_48[45], stage1_48[46], stage1_48[47]},
      {stage2_50[7],stage2_49[32],stage2_48[69],stage2_47[81],stage2_46[82]}
   );
   gpc615_5 gpc5545 (
      {stage1_46[285], stage1_46[286], stage1_46[287], stage1_46[288], stage1_46[289]},
      {stage1_47[158]},
      {stage1_48[48], stage1_48[49], stage1_48[50], stage1_48[51], stage1_48[52], stage1_48[53]},
      {stage2_50[8],stage2_49[33],stage2_48[70],stage2_47[82],stage2_46[83]}
   );
   gpc615_5 gpc5546 (
      {stage1_46[290], stage1_46[291], stage1_46[292], stage1_46[293], stage1_46[294]},
      {stage1_47[159]},
      {stage1_48[54], stage1_48[55], stage1_48[56], stage1_48[57], stage1_48[58], stage1_48[59]},
      {stage2_50[9],stage2_49[34],stage2_48[71],stage2_47[83],stage2_46[84]}
   );
   gpc615_5 gpc5547 (
      {stage1_47[160], stage1_47[161], stage1_47[162], stage1_47[163], stage1_47[164]},
      {stage1_48[60]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[10],stage2_49[35],stage2_48[72],stage2_47[84]}
   );
   gpc615_5 gpc5548 (
      {stage1_47[165], stage1_47[166], stage1_47[167], stage1_47[168], stage1_47[169]},
      {stage1_48[61]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[11],stage2_49[36],stage2_48[73],stage2_47[85]}
   );
   gpc615_5 gpc5549 (
      {stage1_47[170], stage1_47[171], stage1_47[172], stage1_47[173], stage1_47[174]},
      {stage1_48[62]},
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage2_51[2],stage2_50[12],stage2_49[37],stage2_48[74],stage2_47[86]}
   );
   gpc615_5 gpc5550 (
      {stage1_47[175], stage1_47[176], stage1_47[177], stage1_47[178], stage1_47[179]},
      {stage1_48[63]},
      {stage1_49[18], stage1_49[19], stage1_49[20], stage1_49[21], stage1_49[22], stage1_49[23]},
      {stage2_51[3],stage2_50[13],stage2_49[38],stage2_48[75],stage2_47[87]}
   );
   gpc615_5 gpc5551 (
      {stage1_47[180], stage1_47[181], stage1_47[182], stage1_47[183], stage1_47[184]},
      {stage1_48[64]},
      {stage1_49[24], stage1_49[25], stage1_49[26], stage1_49[27], stage1_49[28], stage1_49[29]},
      {stage2_51[4],stage2_50[14],stage2_49[39],stage2_48[76],stage2_47[88]}
   );
   gpc615_5 gpc5552 (
      {stage1_47[185], stage1_47[186], stage1_47[187], stage1_47[188], stage1_47[189]},
      {stage1_48[65]},
      {stage1_49[30], stage1_49[31], stage1_49[32], stage1_49[33], stage1_49[34], stage1_49[35]},
      {stage2_51[5],stage2_50[15],stage2_49[40],stage2_48[77],stage2_47[89]}
   );
   gpc615_5 gpc5553 (
      {stage1_47[190], stage1_47[191], stage1_47[192], stage1_47[193], stage1_47[194]},
      {stage1_48[66]},
      {stage1_49[36], stage1_49[37], stage1_49[38], stage1_49[39], stage1_49[40], stage1_49[41]},
      {stage2_51[6],stage2_50[16],stage2_49[41],stage2_48[78],stage2_47[90]}
   );
   gpc615_5 gpc5554 (
      {stage1_47[195], stage1_47[196], stage1_47[197], stage1_47[198], stage1_47[199]},
      {stage1_48[67]},
      {stage1_49[42], stage1_49[43], stage1_49[44], stage1_49[45], stage1_49[46], stage1_49[47]},
      {stage2_51[7],stage2_50[17],stage2_49[42],stage2_48[79],stage2_47[91]}
   );
   gpc615_5 gpc5555 (
      {stage1_47[200], stage1_47[201], stage1_47[202], stage1_47[203], stage1_47[204]},
      {stage1_48[68]},
      {stage1_49[48], stage1_49[49], stage1_49[50], stage1_49[51], stage1_49[52], stage1_49[53]},
      {stage2_51[8],stage2_50[18],stage2_49[43],stage2_48[80],stage2_47[92]}
   );
   gpc615_5 gpc5556 (
      {stage1_47[205], stage1_47[206], stage1_47[207], stage1_47[208], stage1_47[209]},
      {stage1_48[69]},
      {stage1_49[54], stage1_49[55], stage1_49[56], stage1_49[57], stage1_49[58], stage1_49[59]},
      {stage2_51[9],stage2_50[19],stage2_49[44],stage2_48[81],stage2_47[93]}
   );
   gpc615_5 gpc5557 (
      {stage1_47[210], stage1_47[211], stage1_47[212], stage1_47[213], stage1_47[214]},
      {stage1_48[70]},
      {stage1_49[60], stage1_49[61], stage1_49[62], stage1_49[63], stage1_49[64], stage1_49[65]},
      {stage2_51[10],stage2_50[20],stage2_49[45],stage2_48[82],stage2_47[94]}
   );
   gpc615_5 gpc5558 (
      {stage1_47[215], stage1_47[216], stage1_47[217], stage1_47[218], stage1_47[219]},
      {stage1_48[71]},
      {stage1_49[66], stage1_49[67], stage1_49[68], stage1_49[69], stage1_49[70], stage1_49[71]},
      {stage2_51[11],stage2_50[21],stage2_49[46],stage2_48[83],stage2_47[95]}
   );
   gpc615_5 gpc5559 (
      {stage1_47[220], stage1_47[221], stage1_47[222], stage1_47[223], stage1_47[224]},
      {stage1_48[72]},
      {stage1_49[72], stage1_49[73], stage1_49[74], stage1_49[75], stage1_49[76], stage1_49[77]},
      {stage2_51[12],stage2_50[22],stage2_49[47],stage2_48[84],stage2_47[96]}
   );
   gpc615_5 gpc5560 (
      {stage1_47[225], stage1_47[226], stage1_47[227], stage1_47[228], stage1_47[229]},
      {stage1_48[73]},
      {stage1_49[78], stage1_49[79], stage1_49[80], stage1_49[81], stage1_49[82], stage1_49[83]},
      {stage2_51[13],stage2_50[23],stage2_49[48],stage2_48[85],stage2_47[97]}
   );
   gpc606_5 gpc5561 (
      {stage1_48[74], stage1_48[75], stage1_48[76], stage1_48[77], stage1_48[78], stage1_48[79]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[14],stage2_50[24],stage2_49[49],stage2_48[86]}
   );
   gpc606_5 gpc5562 (
      {stage1_48[80], stage1_48[81], stage1_48[82], stage1_48[83], stage1_48[84], stage1_48[85]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[1],stage2_51[15],stage2_50[25],stage2_49[50],stage2_48[87]}
   );
   gpc606_5 gpc5563 (
      {stage1_48[86], stage1_48[87], stage1_48[88], stage1_48[89], stage1_48[90], stage1_48[91]},
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16], stage1_50[17]},
      {stage2_52[2],stage2_51[16],stage2_50[26],stage2_49[51],stage2_48[88]}
   );
   gpc606_5 gpc5564 (
      {stage1_48[92], stage1_48[93], stage1_48[94], stage1_48[95], stage1_48[96], stage1_48[97]},
      {stage1_50[18], stage1_50[19], stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23]},
      {stage2_52[3],stage2_51[17],stage2_50[27],stage2_49[52],stage2_48[89]}
   );
   gpc606_5 gpc5565 (
      {stage1_48[98], stage1_48[99], stage1_48[100], stage1_48[101], stage1_48[102], stage1_48[103]},
      {stage1_50[24], stage1_50[25], stage1_50[26], stage1_50[27], stage1_50[28], stage1_50[29]},
      {stage2_52[4],stage2_51[18],stage2_50[28],stage2_49[53],stage2_48[90]}
   );
   gpc606_5 gpc5566 (
      {stage1_48[104], stage1_48[105], stage1_48[106], stage1_48[107], stage1_48[108], stage1_48[109]},
      {stage1_50[30], stage1_50[31], stage1_50[32], stage1_50[33], stage1_50[34], stage1_50[35]},
      {stage2_52[5],stage2_51[19],stage2_50[29],stage2_49[54],stage2_48[91]}
   );
   gpc606_5 gpc5567 (
      {stage1_48[110], stage1_48[111], stage1_48[112], stage1_48[113], stage1_48[114], stage1_48[115]},
      {stage1_50[36], stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40], stage1_50[41]},
      {stage2_52[6],stage2_51[20],stage2_50[30],stage2_49[55],stage2_48[92]}
   );
   gpc606_5 gpc5568 (
      {stage1_48[116], stage1_48[117], stage1_48[118], stage1_48[119], stage1_48[120], stage1_48[121]},
      {stage1_50[42], stage1_50[43], stage1_50[44], stage1_50[45], stage1_50[46], stage1_50[47]},
      {stage2_52[7],stage2_51[21],stage2_50[31],stage2_49[56],stage2_48[93]}
   );
   gpc615_5 gpc5569 (
      {stage1_48[122], stage1_48[123], stage1_48[124], stage1_48[125], stage1_48[126]},
      {stage1_49[84]},
      {stage1_50[48], stage1_50[49], stage1_50[50], stage1_50[51], stage1_50[52], stage1_50[53]},
      {stage2_52[8],stage2_51[22],stage2_50[32],stage2_49[57],stage2_48[94]}
   );
   gpc615_5 gpc5570 (
      {stage1_48[127], stage1_48[128], stage1_48[129], stage1_48[130], stage1_48[131]},
      {stage1_49[85]},
      {stage1_50[54], stage1_50[55], stage1_50[56], stage1_50[57], stage1_50[58], stage1_50[59]},
      {stage2_52[9],stage2_51[23],stage2_50[33],stage2_49[58],stage2_48[95]}
   );
   gpc615_5 gpc5571 (
      {stage1_48[132], stage1_48[133], stage1_48[134], stage1_48[135], stage1_48[136]},
      {stage1_49[86]},
      {stage1_50[60], stage1_50[61], stage1_50[62], stage1_50[63], stage1_50[64], stage1_50[65]},
      {stage2_52[10],stage2_51[24],stage2_50[34],stage2_49[59],stage2_48[96]}
   );
   gpc615_5 gpc5572 (
      {stage1_48[137], stage1_48[138], stage1_48[139], stage1_48[140], stage1_48[141]},
      {stage1_49[87]},
      {stage1_50[66], stage1_50[67], stage1_50[68], stage1_50[69], stage1_50[70], stage1_50[71]},
      {stage2_52[11],stage2_51[25],stage2_50[35],stage2_49[60],stage2_48[97]}
   );
   gpc615_5 gpc5573 (
      {stage1_48[142], stage1_48[143], stage1_48[144], stage1_48[145], stage1_48[146]},
      {stage1_49[88]},
      {stage1_50[72], stage1_50[73], stage1_50[74], stage1_50[75], stage1_50[76], stage1_50[77]},
      {stage2_52[12],stage2_51[26],stage2_50[36],stage2_49[61],stage2_48[98]}
   );
   gpc615_5 gpc5574 (
      {stage1_48[147], stage1_48[148], stage1_48[149], stage1_48[150], stage1_48[151]},
      {stage1_49[89]},
      {stage1_50[78], stage1_50[79], stage1_50[80], stage1_50[81], stage1_50[82], stage1_50[83]},
      {stage2_52[13],stage2_51[27],stage2_50[37],stage2_49[62],stage2_48[99]}
   );
   gpc615_5 gpc5575 (
      {stage1_48[152], stage1_48[153], stage1_48[154], stage1_48[155], stage1_48[156]},
      {stage1_49[90]},
      {stage1_50[84], stage1_50[85], stage1_50[86], stage1_50[87], stage1_50[88], stage1_50[89]},
      {stage2_52[14],stage2_51[28],stage2_50[38],stage2_49[63],stage2_48[100]}
   );
   gpc615_5 gpc5576 (
      {stage1_48[157], stage1_48[158], stage1_48[159], stage1_48[160], stage1_48[161]},
      {stage1_49[91]},
      {stage1_50[90], stage1_50[91], stage1_50[92], stage1_50[93], stage1_50[94], stage1_50[95]},
      {stage2_52[15],stage2_51[29],stage2_50[39],stage2_49[64],stage2_48[101]}
   );
   gpc615_5 gpc5577 (
      {stage1_48[162], stage1_48[163], stage1_48[164], stage1_48[165], stage1_48[166]},
      {stage1_49[92]},
      {stage1_50[96], stage1_50[97], stage1_50[98], stage1_50[99], stage1_50[100], stage1_50[101]},
      {stage2_52[16],stage2_51[30],stage2_50[40],stage2_49[65],stage2_48[102]}
   );
   gpc615_5 gpc5578 (
      {stage1_48[167], stage1_48[168], stage1_48[169], stage1_48[170], stage1_48[171]},
      {stage1_49[93]},
      {stage1_50[102], stage1_50[103], stage1_50[104], stage1_50[105], stage1_50[106], stage1_50[107]},
      {stage2_52[17],stage2_51[31],stage2_50[41],stage2_49[66],stage2_48[103]}
   );
   gpc606_5 gpc5579 (
      {stage1_49[94], stage1_49[95], stage1_49[96], stage1_49[97], stage1_49[98], stage1_49[99]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[18],stage2_51[32],stage2_50[42],stage2_49[67]}
   );
   gpc606_5 gpc5580 (
      {stage1_49[100], stage1_49[101], stage1_49[102], stage1_49[103], stage1_49[104], stage1_49[105]},
      {stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage2_53[1],stage2_52[19],stage2_51[33],stage2_50[43],stage2_49[68]}
   );
   gpc606_5 gpc5581 (
      {stage1_49[106], stage1_49[107], stage1_49[108], stage1_49[109], stage1_49[110], stage1_49[111]},
      {stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15], stage1_51[16], stage1_51[17]},
      {stage2_53[2],stage2_52[20],stage2_51[34],stage2_50[44],stage2_49[69]}
   );
   gpc606_5 gpc5582 (
      {stage1_49[112], stage1_49[113], stage1_49[114], stage1_49[115], stage1_49[116], stage1_49[117]},
      {stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21], stage1_51[22], stage1_51[23]},
      {stage2_53[3],stage2_52[21],stage2_51[35],stage2_50[45],stage2_49[70]}
   );
   gpc606_5 gpc5583 (
      {stage1_49[118], stage1_49[119], stage1_49[120], stage1_49[121], stage1_49[122], stage1_49[123]},
      {stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27], stage1_51[28], stage1_51[29]},
      {stage2_53[4],stage2_52[22],stage2_51[36],stage2_50[46],stage2_49[71]}
   );
   gpc606_5 gpc5584 (
      {stage1_49[124], stage1_49[125], stage1_49[126], stage1_49[127], stage1_49[128], stage1_49[129]},
      {stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33], stage1_51[34], stage1_51[35]},
      {stage2_53[5],stage2_52[23],stage2_51[37],stage2_50[47],stage2_49[72]}
   );
   gpc606_5 gpc5585 (
      {stage1_49[130], stage1_49[131], stage1_49[132], stage1_49[133], stage1_49[134], stage1_49[135]},
      {stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39], stage1_51[40], stage1_51[41]},
      {stage2_53[6],stage2_52[24],stage2_51[38],stage2_50[48],stage2_49[73]}
   );
   gpc606_5 gpc5586 (
      {stage1_49[136], stage1_49[137], stage1_49[138], stage1_49[139], stage1_49[140], stage1_49[141]},
      {stage1_51[42], stage1_51[43], stage1_51[44], stage1_51[45], stage1_51[46], stage1_51[47]},
      {stage2_53[7],stage2_52[25],stage2_51[39],stage2_50[49],stage2_49[74]}
   );
   gpc606_5 gpc5587 (
      {stage1_49[142], stage1_49[143], stage1_49[144], stage1_49[145], stage1_49[146], stage1_49[147]},
      {stage1_51[48], stage1_51[49], stage1_51[50], stage1_51[51], stage1_51[52], stage1_51[53]},
      {stage2_53[8],stage2_52[26],stage2_51[40],stage2_50[50],stage2_49[75]}
   );
   gpc606_5 gpc5588 (
      {stage1_49[148], stage1_49[149], stage1_49[150], stage1_49[151], stage1_49[152], stage1_49[153]},
      {stage1_51[54], stage1_51[55], stage1_51[56], stage1_51[57], stage1_51[58], stage1_51[59]},
      {stage2_53[9],stage2_52[27],stage2_51[41],stage2_50[51],stage2_49[76]}
   );
   gpc2135_5 gpc5589 (
      {stage1_50[108], stage1_50[109], stage1_50[110], stage1_50[111], stage1_50[112]},
      {stage1_51[60], stage1_51[61], stage1_51[62]},
      {stage1_52[0]},
      {stage1_53[0], stage1_53[1]},
      {stage2_54[0],stage2_53[10],stage2_52[28],stage2_51[42],stage2_50[52]}
   );
   gpc1163_5 gpc5590 (
      {stage1_50[113], stage1_50[114], stage1_50[115]},
      {stage1_51[63], stage1_51[64], stage1_51[65], stage1_51[66], stage1_51[67], stage1_51[68]},
      {stage1_52[1]},
      {stage1_53[2]},
      {stage2_54[1],stage2_53[11],stage2_52[29],stage2_51[43],stage2_50[53]}
   );
   gpc1163_5 gpc5591 (
      {stage1_50[116], stage1_50[117], stage1_50[118]},
      {stage1_51[69], stage1_51[70], stage1_51[71], stage1_51[72], stage1_51[73], stage1_51[74]},
      {stage1_52[2]},
      {stage1_53[3]},
      {stage2_54[2],stage2_53[12],stage2_52[30],stage2_51[44],stage2_50[54]}
   );
   gpc1163_5 gpc5592 (
      {stage1_50[119], stage1_50[120], stage1_50[121]},
      {stage1_51[75], stage1_51[76], stage1_51[77], stage1_51[78], stage1_51[79], stage1_51[80]},
      {stage1_52[3]},
      {stage1_53[4]},
      {stage2_54[3],stage2_53[13],stage2_52[31],stage2_51[45],stage2_50[55]}
   );
   gpc1163_5 gpc5593 (
      {stage1_50[122], stage1_50[123], stage1_50[124]},
      {stage1_51[81], stage1_51[82], stage1_51[83], stage1_51[84], stage1_51[85], stage1_51[86]},
      {stage1_52[4]},
      {stage1_53[5]},
      {stage2_54[4],stage2_53[14],stage2_52[32],stage2_51[46],stage2_50[56]}
   );
   gpc1163_5 gpc5594 (
      {stage1_50[125], stage1_50[126], stage1_50[127]},
      {stage1_51[87], stage1_51[88], stage1_51[89], stage1_51[90], stage1_51[91], stage1_51[92]},
      {stage1_52[5]},
      {stage1_53[6]},
      {stage2_54[5],stage2_53[15],stage2_52[33],stage2_51[47],stage2_50[57]}
   );
   gpc1163_5 gpc5595 (
      {stage1_50[128], stage1_50[129], stage1_50[130]},
      {stage1_51[93], stage1_51[94], stage1_51[95], stage1_51[96], stage1_51[97], stage1_51[98]},
      {stage1_52[6]},
      {stage1_53[7]},
      {stage2_54[6],stage2_53[16],stage2_52[34],stage2_51[48],stage2_50[58]}
   );
   gpc1163_5 gpc5596 (
      {stage1_50[131], stage1_50[132], stage1_50[133]},
      {stage1_51[99], stage1_51[100], stage1_51[101], stage1_51[102], stage1_51[103], stage1_51[104]},
      {stage1_52[7]},
      {stage1_53[8]},
      {stage2_54[7],stage2_53[17],stage2_52[35],stage2_51[49],stage2_50[59]}
   );
   gpc1163_5 gpc5597 (
      {stage1_50[134], stage1_50[135], stage1_50[136]},
      {stage1_51[105], stage1_51[106], stage1_51[107], stage1_51[108], stage1_51[109], stage1_51[110]},
      {stage1_52[8]},
      {stage1_53[9]},
      {stage2_54[8],stage2_53[18],stage2_52[36],stage2_51[50],stage2_50[60]}
   );
   gpc1163_5 gpc5598 (
      {stage1_50[137], stage1_50[138], stage1_50[139]},
      {stage1_51[111], stage1_51[112], stage1_51[113], stage1_51[114], stage1_51[115], stage1_51[116]},
      {stage1_52[9]},
      {stage1_53[10]},
      {stage2_54[9],stage2_53[19],stage2_52[37],stage2_51[51],stage2_50[61]}
   );
   gpc1163_5 gpc5599 (
      {stage1_50[140], stage1_50[141], stage1_50[142]},
      {stage1_51[117], stage1_51[118], stage1_51[119], stage1_51[120], stage1_51[121], stage1_51[122]},
      {stage1_52[10]},
      {stage1_53[11]},
      {stage2_54[10],stage2_53[20],stage2_52[38],stage2_51[52],stage2_50[62]}
   );
   gpc1163_5 gpc5600 (
      {stage1_50[143], stage1_50[144], stage1_50[145]},
      {stage1_51[123], stage1_51[124], stage1_51[125], stage1_51[126], stage1_51[127], stage1_51[128]},
      {stage1_52[11]},
      {stage1_53[12]},
      {stage2_54[11],stage2_53[21],stage2_52[39],stage2_51[53],stage2_50[63]}
   );
   gpc1163_5 gpc5601 (
      {stage1_50[146], stage1_50[147], stage1_50[148]},
      {stage1_51[129], stage1_51[130], stage1_51[131], stage1_51[132], stage1_51[133], stage1_51[134]},
      {stage1_52[12]},
      {stage1_53[13]},
      {stage2_54[12],stage2_53[22],stage2_52[40],stage2_51[54],stage2_50[64]}
   );
   gpc1163_5 gpc5602 (
      {stage1_50[149], stage1_50[150], stage1_50[151]},
      {stage1_51[135], stage1_51[136], stage1_51[137], stage1_51[138], stage1_51[139], stage1_51[140]},
      {stage1_52[13]},
      {stage1_53[14]},
      {stage2_54[13],stage2_53[23],stage2_52[41],stage2_51[55],stage2_50[65]}
   );
   gpc1163_5 gpc5603 (
      {stage1_50[152], stage1_50[153], stage1_50[154]},
      {stage1_51[141], stage1_51[142], stage1_51[143], stage1_51[144], stage1_51[145], stage1_51[146]},
      {stage1_52[14]},
      {stage1_53[15]},
      {stage2_54[14],stage2_53[24],stage2_52[42],stage2_51[56],stage2_50[66]}
   );
   gpc1163_5 gpc5604 (
      {stage1_50[155], stage1_50[156], stage1_50[157]},
      {stage1_51[147], stage1_51[148], stage1_51[149], stage1_51[150], stage1_51[151], stage1_51[152]},
      {stage1_52[15]},
      {stage1_53[16]},
      {stage2_54[15],stage2_53[25],stage2_52[43],stage2_51[57],stage2_50[67]}
   );
   gpc1163_5 gpc5605 (
      {stage1_50[158], stage1_50[159], stage1_50[160]},
      {stage1_51[153], stage1_51[154], stage1_51[155], stage1_51[156], stage1_51[157], stage1_51[158]},
      {stage1_52[16]},
      {stage1_53[17]},
      {stage2_54[16],stage2_53[26],stage2_52[44],stage2_51[58],stage2_50[68]}
   );
   gpc1163_5 gpc5606 (
      {stage1_50[161], stage1_50[162], stage1_50[163]},
      {stage1_51[159], stage1_51[160], stage1_51[161], stage1_51[162], stage1_51[163], stage1_51[164]},
      {stage1_52[17]},
      {stage1_53[18]},
      {stage2_54[17],stage2_53[27],stage2_52[45],stage2_51[59],stage2_50[69]}
   );
   gpc1163_5 gpc5607 (
      {stage1_50[164], stage1_50[165], stage1_50[166]},
      {stage1_51[165], stage1_51[166], stage1_51[167], stage1_51[168], stage1_51[169], stage1_51[170]},
      {stage1_52[18]},
      {stage1_53[19]},
      {stage2_54[18],stage2_53[28],stage2_52[46],stage2_51[60],stage2_50[70]}
   );
   gpc1163_5 gpc5608 (
      {stage1_50[167], stage1_50[168], stage1_50[169]},
      {stage1_51[171], stage1_51[172], stage1_51[173], stage1_51[174], stage1_51[175], stage1_51[176]},
      {stage1_52[19]},
      {stage1_53[20]},
      {stage2_54[19],stage2_53[29],stage2_52[47],stage2_51[61],stage2_50[71]}
   );
   gpc1163_5 gpc5609 (
      {stage1_50[170], stage1_50[171], stage1_50[172]},
      {stage1_51[177], stage1_51[178], stage1_51[179], stage1_51[180], stage1_51[181], stage1_51[182]},
      {stage1_52[20]},
      {stage1_53[21]},
      {stage2_54[20],stage2_53[30],stage2_52[48],stage2_51[62],stage2_50[72]}
   );
   gpc1163_5 gpc5610 (
      {stage1_50[173], stage1_50[174], stage1_50[175]},
      {stage1_51[183], stage1_51[184], stage1_51[185], stage1_51[186], stage1_51[187], stage1_51[188]},
      {stage1_52[21]},
      {stage1_53[22]},
      {stage2_54[21],stage2_53[31],stage2_52[49],stage2_51[63],stage2_50[73]}
   );
   gpc1163_5 gpc5611 (
      {stage1_50[176], stage1_50[177], stage1_50[178]},
      {stage1_51[189], stage1_51[190], stage1_51[191], stage1_51[192], stage1_51[193], stage1_51[194]},
      {stage1_52[22]},
      {stage1_53[23]},
      {stage2_54[22],stage2_53[32],stage2_52[50],stage2_51[64],stage2_50[74]}
   );
   gpc606_5 gpc5612 (
      {stage1_51[195], stage1_51[196], stage1_51[197], stage1_51[198], stage1_51[199], stage1_51[200]},
      {stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27], stage1_53[28], stage1_53[29]},
      {stage2_55[0],stage2_54[23],stage2_53[33],stage2_52[51],stage2_51[65]}
   );
   gpc615_5 gpc5613 (
      {stage1_51[201], stage1_51[202], stage1_51[203], stage1_51[204], stage1_51[205]},
      {stage1_52[23]},
      {stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33], stage1_53[34], stage1_53[35]},
      {stage2_55[1],stage2_54[24],stage2_53[34],stage2_52[52],stage2_51[66]}
   );
   gpc615_5 gpc5614 (
      {stage1_51[206], stage1_51[207], stage1_51[208], stage1_51[209], stage1_51[210]},
      {stage1_52[24]},
      {stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39], stage1_53[40], stage1_53[41]},
      {stage2_55[2],stage2_54[25],stage2_53[35],stage2_52[53],stage2_51[67]}
   );
   gpc615_5 gpc5615 (
      {stage1_51[211], stage1_51[212], stage1_51[213], stage1_51[214], stage1_51[215]},
      {stage1_52[25]},
      {stage1_53[42], stage1_53[43], stage1_53[44], stage1_53[45], stage1_53[46], stage1_53[47]},
      {stage2_55[3],stage2_54[26],stage2_53[36],stage2_52[54],stage2_51[68]}
   );
   gpc615_5 gpc5616 (
      {stage1_51[216], stage1_51[217], stage1_51[218], stage1_51[219], stage1_51[220]},
      {stage1_52[26]},
      {stage1_53[48], stage1_53[49], stage1_53[50], stage1_53[51], stage1_53[52], stage1_53[53]},
      {stage2_55[4],stage2_54[27],stage2_53[37],stage2_52[55],stage2_51[69]}
   );
   gpc615_5 gpc5617 (
      {stage1_51[221], stage1_51[222], stage1_51[223], stage1_51[224], stage1_51[225]},
      {stage1_52[27]},
      {stage1_53[54], stage1_53[55], stage1_53[56], stage1_53[57], stage1_53[58], stage1_53[59]},
      {stage2_55[5],stage2_54[28],stage2_53[38],stage2_52[56],stage2_51[70]}
   );
   gpc615_5 gpc5618 (
      {stage1_51[226], stage1_51[227], stage1_51[228], stage1_51[229], stage1_51[230]},
      {stage1_52[28]},
      {stage1_53[60], stage1_53[61], stage1_53[62], stage1_53[63], stage1_53[64], stage1_53[65]},
      {stage2_55[6],stage2_54[29],stage2_53[39],stage2_52[57],stage2_51[71]}
   );
   gpc615_5 gpc5619 (
      {stage1_51[231], stage1_51[232], stage1_51[233], stage1_51[234], stage1_51[235]},
      {stage1_52[29]},
      {stage1_53[66], stage1_53[67], stage1_53[68], stage1_53[69], stage1_53[70], stage1_53[71]},
      {stage2_55[7],stage2_54[30],stage2_53[40],stage2_52[58],stage2_51[72]}
   );
   gpc615_5 gpc5620 (
      {stage1_51[236], stage1_51[237], stage1_51[238], stage1_51[239], stage1_51[240]},
      {stage1_52[30]},
      {stage1_53[72], stage1_53[73], stage1_53[74], stage1_53[75], stage1_53[76], stage1_53[77]},
      {stage2_55[8],stage2_54[31],stage2_53[41],stage2_52[59],stage2_51[73]}
   );
   gpc615_5 gpc5621 (
      {stage1_51[241], stage1_51[242], stage1_51[243], stage1_51[244], stage1_51[245]},
      {stage1_52[31]},
      {stage1_53[78], stage1_53[79], stage1_53[80], stage1_53[81], stage1_53[82], stage1_53[83]},
      {stage2_55[9],stage2_54[32],stage2_53[42],stage2_52[60],stage2_51[74]}
   );
   gpc615_5 gpc5622 (
      {stage1_51[246], stage1_51[247], stage1_51[248], stage1_51[249], stage1_51[250]},
      {stage1_52[32]},
      {stage1_53[84], stage1_53[85], stage1_53[86], stage1_53[87], stage1_53[88], stage1_53[89]},
      {stage2_55[10],stage2_54[33],stage2_53[43],stage2_52[61],stage2_51[75]}
   );
   gpc615_5 gpc5623 (
      {stage1_51[251], stage1_51[252], stage1_51[253], stage1_51[254], stage1_51[255]},
      {stage1_52[33]},
      {stage1_53[90], stage1_53[91], stage1_53[92], stage1_53[93], stage1_53[94], stage1_53[95]},
      {stage2_55[11],stage2_54[34],stage2_53[44],stage2_52[62],stage2_51[76]}
   );
   gpc615_5 gpc5624 (
      {stage1_51[256], stage1_51[257], stage1_51[258], stage1_51[259], stage1_51[260]},
      {stage1_52[34]},
      {stage1_53[96], stage1_53[97], stage1_53[98], stage1_53[99], stage1_53[100], stage1_53[101]},
      {stage2_55[12],stage2_54[35],stage2_53[45],stage2_52[63],stage2_51[77]}
   );
   gpc615_5 gpc5625 (
      {stage1_51[261], stage1_51[262], stage1_51[263], stage1_51[264], stage1_51[265]},
      {stage1_52[35]},
      {stage1_53[102], stage1_53[103], stage1_53[104], stage1_53[105], stage1_53[106], stage1_53[107]},
      {stage2_55[13],stage2_54[36],stage2_53[46],stage2_52[64],stage2_51[78]}
   );
   gpc606_5 gpc5626 (
      {stage1_52[36], stage1_52[37], stage1_52[38], stage1_52[39], stage1_52[40], stage1_52[41]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[14],stage2_54[37],stage2_53[47],stage2_52[65]}
   );
   gpc606_5 gpc5627 (
      {stage1_52[42], stage1_52[43], stage1_52[44], stage1_52[45], stage1_52[46], stage1_52[47]},
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10], stage1_54[11]},
      {stage2_56[1],stage2_55[15],stage2_54[38],stage2_53[48],stage2_52[66]}
   );
   gpc606_5 gpc5628 (
      {stage1_52[48], stage1_52[49], stage1_52[50], stage1_52[51], stage1_52[52], stage1_52[53]},
      {stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15], stage1_54[16], stage1_54[17]},
      {stage2_56[2],stage2_55[16],stage2_54[39],stage2_53[49],stage2_52[67]}
   );
   gpc606_5 gpc5629 (
      {stage1_52[54], stage1_52[55], stage1_52[56], stage1_52[57], stage1_52[58], stage1_52[59]},
      {stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21], stage1_54[22], stage1_54[23]},
      {stage2_56[3],stage2_55[17],stage2_54[40],stage2_53[50],stage2_52[68]}
   );
   gpc606_5 gpc5630 (
      {stage1_52[60], stage1_52[61], stage1_52[62], stage1_52[63], stage1_52[64], stage1_52[65]},
      {stage1_54[24], stage1_54[25], stage1_54[26], stage1_54[27], stage1_54[28], stage1_54[29]},
      {stage2_56[4],stage2_55[18],stage2_54[41],stage2_53[51],stage2_52[69]}
   );
   gpc606_5 gpc5631 (
      {stage1_52[66], stage1_52[67], stage1_52[68], stage1_52[69], stage1_52[70], stage1_52[71]},
      {stage1_54[30], stage1_54[31], stage1_54[32], stage1_54[33], stage1_54[34], stage1_54[35]},
      {stage2_56[5],stage2_55[19],stage2_54[42],stage2_53[52],stage2_52[70]}
   );
   gpc606_5 gpc5632 (
      {stage1_52[72], stage1_52[73], stage1_52[74], stage1_52[75], stage1_52[76], stage1_52[77]},
      {stage1_54[36], stage1_54[37], stage1_54[38], stage1_54[39], stage1_54[40], stage1_54[41]},
      {stage2_56[6],stage2_55[20],stage2_54[43],stage2_53[53],stage2_52[71]}
   );
   gpc606_5 gpc5633 (
      {stage1_52[78], stage1_52[79], stage1_52[80], stage1_52[81], stage1_52[82], stage1_52[83]},
      {stage1_54[42], stage1_54[43], stage1_54[44], stage1_54[45], stage1_54[46], stage1_54[47]},
      {stage2_56[7],stage2_55[21],stage2_54[44],stage2_53[54],stage2_52[72]}
   );
   gpc606_5 gpc5634 (
      {stage1_52[84], stage1_52[85], stage1_52[86], stage1_52[87], stage1_52[88], stage1_52[89]},
      {stage1_54[48], stage1_54[49], stage1_54[50], stage1_54[51], stage1_54[52], stage1_54[53]},
      {stage2_56[8],stage2_55[22],stage2_54[45],stage2_53[55],stage2_52[73]}
   );
   gpc606_5 gpc5635 (
      {stage1_52[90], stage1_52[91], stage1_52[92], stage1_52[93], stage1_52[94], stage1_52[95]},
      {stage1_54[54], stage1_54[55], stage1_54[56], stage1_54[57], stage1_54[58], stage1_54[59]},
      {stage2_56[9],stage2_55[23],stage2_54[46],stage2_53[56],stage2_52[74]}
   );
   gpc606_5 gpc5636 (
      {stage1_52[96], stage1_52[97], stage1_52[98], stage1_52[99], stage1_52[100], stage1_52[101]},
      {stage1_54[60], stage1_54[61], stage1_54[62], stage1_54[63], stage1_54[64], stage1_54[65]},
      {stage2_56[10],stage2_55[24],stage2_54[47],stage2_53[57],stage2_52[75]}
   );
   gpc615_5 gpc5637 (
      {stage1_52[102], stage1_52[103], stage1_52[104], stage1_52[105], stage1_52[106]},
      {stage1_53[108]},
      {stage1_54[66], stage1_54[67], stage1_54[68], stage1_54[69], stage1_54[70], stage1_54[71]},
      {stage2_56[11],stage2_55[25],stage2_54[48],stage2_53[58],stage2_52[76]}
   );
   gpc615_5 gpc5638 (
      {stage1_52[107], stage1_52[108], stage1_52[109], stage1_52[110], stage1_52[111]},
      {stage1_53[109]},
      {stage1_54[72], stage1_54[73], stage1_54[74], stage1_54[75], stage1_54[76], stage1_54[77]},
      {stage2_56[12],stage2_55[26],stage2_54[49],stage2_53[59],stage2_52[77]}
   );
   gpc615_5 gpc5639 (
      {stage1_52[112], stage1_52[113], stage1_52[114], stage1_52[115], stage1_52[116]},
      {stage1_53[110]},
      {stage1_54[78], stage1_54[79], stage1_54[80], stage1_54[81], stage1_54[82], stage1_54[83]},
      {stage2_56[13],stage2_55[27],stage2_54[50],stage2_53[60],stage2_52[78]}
   );
   gpc615_5 gpc5640 (
      {stage1_52[117], stage1_52[118], stage1_52[119], stage1_52[120], stage1_52[121]},
      {stage1_53[111]},
      {stage1_54[84], stage1_54[85], stage1_54[86], stage1_54[87], stage1_54[88], stage1_54[89]},
      {stage2_56[14],stage2_55[28],stage2_54[51],stage2_53[61],stage2_52[79]}
   );
   gpc615_5 gpc5641 (
      {stage1_52[122], stage1_52[123], stage1_52[124], stage1_52[125], stage1_52[126]},
      {stage1_53[112]},
      {stage1_54[90], stage1_54[91], stage1_54[92], stage1_54[93], stage1_54[94], stage1_54[95]},
      {stage2_56[15],stage2_55[29],stage2_54[52],stage2_53[62],stage2_52[80]}
   );
   gpc615_5 gpc5642 (
      {stage1_52[127], stage1_52[128], stage1_52[129], stage1_52[130], stage1_52[131]},
      {stage1_53[113]},
      {stage1_54[96], stage1_54[97], stage1_54[98], stage1_54[99], stage1_54[100], stage1_54[101]},
      {stage2_56[16],stage2_55[30],stage2_54[53],stage2_53[63],stage2_52[81]}
   );
   gpc615_5 gpc5643 (
      {stage1_52[132], stage1_52[133], stage1_52[134], stage1_52[135], stage1_52[136]},
      {stage1_53[114]},
      {stage1_54[102], stage1_54[103], stage1_54[104], stage1_54[105], stage1_54[106], stage1_54[107]},
      {stage2_56[17],stage2_55[31],stage2_54[54],stage2_53[64],stage2_52[82]}
   );
   gpc615_5 gpc5644 (
      {stage1_52[137], stage1_52[138], stage1_52[139], stage1_52[140], stage1_52[141]},
      {stage1_53[115]},
      {stage1_54[108], stage1_54[109], stage1_54[110], stage1_54[111], stage1_54[112], stage1_54[113]},
      {stage2_56[18],stage2_55[32],stage2_54[55],stage2_53[65],stage2_52[83]}
   );
   gpc615_5 gpc5645 (
      {stage1_52[142], stage1_52[143], stage1_52[144], stage1_52[145], stage1_52[146]},
      {stage1_53[116]},
      {stage1_54[114], stage1_54[115], stage1_54[116], stage1_54[117], stage1_54[118], stage1_54[119]},
      {stage2_56[19],stage2_55[33],stage2_54[56],stage2_53[66],stage2_52[84]}
   );
   gpc615_5 gpc5646 (
      {stage1_52[147], stage1_52[148], stage1_52[149], stage1_52[150], stage1_52[151]},
      {stage1_53[117]},
      {stage1_54[120], stage1_54[121], stage1_54[122], stage1_54[123], stage1_54[124], stage1_54[125]},
      {stage2_56[20],stage2_55[34],stage2_54[57],stage2_53[67],stage2_52[85]}
   );
   gpc615_5 gpc5647 (
      {stage1_52[152], stage1_52[153], stage1_52[154], stage1_52[155], stage1_52[156]},
      {stage1_53[118]},
      {stage1_54[126], stage1_54[127], stage1_54[128], stage1_54[129], stage1_54[130], stage1_54[131]},
      {stage2_56[21],stage2_55[35],stage2_54[58],stage2_53[68],stage2_52[86]}
   );
   gpc615_5 gpc5648 (
      {stage1_52[157], stage1_52[158], stage1_52[159], stage1_52[160], stage1_52[161]},
      {stage1_53[119]},
      {stage1_54[132], stage1_54[133], stage1_54[134], stage1_54[135], stage1_54[136], stage1_54[137]},
      {stage2_56[22],stage2_55[36],stage2_54[59],stage2_53[69],stage2_52[87]}
   );
   gpc615_5 gpc5649 (
      {stage1_52[162], stage1_52[163], stage1_52[164], stage1_52[165], stage1_52[166]},
      {stage1_53[120]},
      {stage1_54[138], stage1_54[139], stage1_54[140], stage1_54[141], stage1_54[142], stage1_54[143]},
      {stage2_56[23],stage2_55[37],stage2_54[60],stage2_53[70],stage2_52[88]}
   );
   gpc615_5 gpc5650 (
      {stage1_52[167], stage1_52[168], stage1_52[169], stage1_52[170], stage1_52[171]},
      {stage1_53[121]},
      {stage1_54[144], stage1_54[145], stage1_54[146], stage1_54[147], stage1_54[148], stage1_54[149]},
      {stage2_56[24],stage2_55[38],stage2_54[61],stage2_53[71],stage2_52[89]}
   );
   gpc615_5 gpc5651 (
      {stage1_52[172], stage1_52[173], stage1_52[174], stage1_52[175], stage1_52[176]},
      {stage1_53[122]},
      {stage1_54[150], stage1_54[151], stage1_54[152], stage1_54[153], stage1_54[154], stage1_54[155]},
      {stage2_56[25],stage2_55[39],stage2_54[62],stage2_53[72],stage2_52[90]}
   );
   gpc615_5 gpc5652 (
      {stage1_52[177], stage1_52[178], stage1_52[179], stage1_52[180], stage1_52[181]},
      {stage1_53[123]},
      {stage1_54[156], stage1_54[157], stage1_54[158], stage1_54[159], stage1_54[160], stage1_54[161]},
      {stage2_56[26],stage2_55[40],stage2_54[63],stage2_53[73],stage2_52[91]}
   );
   gpc615_5 gpc5653 (
      {stage1_52[182], stage1_52[183], stage1_52[184], stage1_52[185], stage1_52[186]},
      {stage1_53[124]},
      {stage1_54[162], stage1_54[163], stage1_54[164], stage1_54[165], stage1_54[166], stage1_54[167]},
      {stage2_56[27],stage2_55[41],stage2_54[64],stage2_53[74],stage2_52[92]}
   );
   gpc615_5 gpc5654 (
      {stage1_53[125], stage1_53[126], stage1_53[127], stage1_53[128], stage1_53[129]},
      {stage1_54[168]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[28],stage2_55[42],stage2_54[65],stage2_53[75]}
   );
   gpc606_5 gpc5655 (
      {stage1_54[169], stage1_54[170], stage1_54[171], stage1_54[172], stage1_54[173], stage1_54[174]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[1],stage2_56[29],stage2_55[43],stage2_54[66]}
   );
   gpc606_5 gpc5656 (
      {stage1_54[175], stage1_54[176], stage1_54[177], stage1_54[178], stage1_54[179], stage1_54[180]},
      {stage1_56[6], stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage2_58[1],stage2_57[2],stage2_56[30],stage2_55[44],stage2_54[67]}
   );
   gpc606_5 gpc5657 (
      {stage1_54[181], stage1_54[182], stage1_54[183], stage1_54[184], stage1_54[185], stage1_54[186]},
      {stage1_56[12], stage1_56[13], stage1_56[14], stage1_56[15], stage1_56[16], stage1_56[17]},
      {stage2_58[2],stage2_57[3],stage2_56[31],stage2_55[45],stage2_54[68]}
   );
   gpc606_5 gpc5658 (
      {stage1_54[187], stage1_54[188], stage1_54[189], stage1_54[190], stage1_54[191], stage1_54[192]},
      {stage1_56[18], stage1_56[19], stage1_56[20], stage1_56[21], stage1_56[22], stage1_56[23]},
      {stage2_58[3],stage2_57[4],stage2_56[32],stage2_55[46],stage2_54[69]}
   );
   gpc615_5 gpc5659 (
      {stage1_54[193], stage1_54[194], stage1_54[195], stage1_54[196], stage1_54[197]},
      {stage1_55[6]},
      {stage1_56[24], stage1_56[25], stage1_56[26], stage1_56[27], stage1_56[28], stage1_56[29]},
      {stage2_58[4],stage2_57[5],stage2_56[33],stage2_55[47],stage2_54[70]}
   );
   gpc615_5 gpc5660 (
      {stage1_54[198], stage1_54[199], stage1_54[200], stage1_54[201], stage1_54[202]},
      {stage1_55[7]},
      {stage1_56[30], stage1_56[31], stage1_56[32], stage1_56[33], stage1_56[34], stage1_56[35]},
      {stage2_58[5],stage2_57[6],stage2_56[34],stage2_55[48],stage2_54[71]}
   );
   gpc2135_5 gpc5661 (
      {stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11], stage1_55[12]},
      {stage1_56[36], stage1_56[37], stage1_56[38]},
      {stage1_57[0]},
      {stage1_58[0], stage1_58[1]},
      {stage2_59[0],stage2_58[6],stage2_57[7],stage2_56[35],stage2_55[49]}
   );
   gpc2135_5 gpc5662 (
      {stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage1_56[39], stage1_56[40], stage1_56[41]},
      {stage1_57[1]},
      {stage1_58[2], stage1_58[3]},
      {stage2_59[1],stage2_58[7],stage2_57[8],stage2_56[36],stage2_55[50]}
   );
   gpc2135_5 gpc5663 (
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22]},
      {stage1_56[42], stage1_56[43], stage1_56[44]},
      {stage1_57[2]},
      {stage1_58[4], stage1_58[5]},
      {stage2_59[2],stage2_58[8],stage2_57[9],stage2_56[37],stage2_55[51]}
   );
   gpc2135_5 gpc5664 (
      {stage1_55[23], stage1_55[24], stage1_55[25], stage1_55[26], stage1_55[27]},
      {stage1_56[45], stage1_56[46], stage1_56[47]},
      {stage1_57[3]},
      {stage1_58[6], stage1_58[7]},
      {stage2_59[3],stage2_58[9],stage2_57[10],stage2_56[38],stage2_55[52]}
   );
   gpc2135_5 gpc5665 (
      {stage1_55[28], stage1_55[29], stage1_55[30], stage1_55[31], stage1_55[32]},
      {stage1_56[48], stage1_56[49], stage1_56[50]},
      {stage1_57[4]},
      {stage1_58[8], stage1_58[9]},
      {stage2_59[4],stage2_58[10],stage2_57[11],stage2_56[39],stage2_55[53]}
   );
   gpc2135_5 gpc5666 (
      {stage1_55[33], stage1_55[34], stage1_55[35], stage1_55[36], stage1_55[37]},
      {stage1_56[51], stage1_56[52], stage1_56[53]},
      {stage1_57[5]},
      {stage1_58[10], stage1_58[11]},
      {stage2_59[5],stage2_58[11],stage2_57[12],stage2_56[40],stage2_55[54]}
   );
   gpc2135_5 gpc5667 (
      {stage1_55[38], stage1_55[39], stage1_55[40], stage1_55[41], stage1_55[42]},
      {stage1_56[54], stage1_56[55], stage1_56[56]},
      {stage1_57[6]},
      {stage1_58[12], stage1_58[13]},
      {stage2_59[6],stage2_58[12],stage2_57[13],stage2_56[41],stage2_55[55]}
   );
   gpc2135_5 gpc5668 (
      {stage1_55[43], stage1_55[44], stage1_55[45], stage1_55[46], stage1_55[47]},
      {stage1_56[57], stage1_56[58], stage1_56[59]},
      {stage1_57[7]},
      {stage1_58[14], stage1_58[15]},
      {stage2_59[7],stage2_58[13],stage2_57[14],stage2_56[42],stage2_55[56]}
   );
   gpc2135_5 gpc5669 (
      {stage1_55[48], stage1_55[49], stage1_55[50], stage1_55[51], stage1_55[52]},
      {stage1_56[60], stage1_56[61], stage1_56[62]},
      {stage1_57[8]},
      {stage1_58[16], stage1_58[17]},
      {stage2_59[8],stage2_58[14],stage2_57[15],stage2_56[43],stage2_55[57]}
   );
   gpc2135_5 gpc5670 (
      {stage1_55[53], stage1_55[54], stage1_55[55], stage1_55[56], stage1_55[57]},
      {stage1_56[63], stage1_56[64], stage1_56[65]},
      {stage1_57[9]},
      {stage1_58[18], stage1_58[19]},
      {stage2_59[9],stage2_58[15],stage2_57[16],stage2_56[44],stage2_55[58]}
   );
   gpc2135_5 gpc5671 (
      {stage1_55[58], stage1_55[59], stage1_55[60], stage1_55[61], stage1_55[62]},
      {stage1_56[66], stage1_56[67], stage1_56[68]},
      {stage1_57[10]},
      {stage1_58[20], stage1_58[21]},
      {stage2_59[10],stage2_58[16],stage2_57[17],stage2_56[45],stage2_55[59]}
   );
   gpc2135_5 gpc5672 (
      {stage1_55[63], stage1_55[64], stage1_55[65], stage1_55[66], stage1_55[67]},
      {stage1_56[69], stage1_56[70], stage1_56[71]},
      {stage1_57[11]},
      {stage1_58[22], stage1_58[23]},
      {stage2_59[11],stage2_58[17],stage2_57[18],stage2_56[46],stage2_55[60]}
   );
   gpc2135_5 gpc5673 (
      {stage1_55[68], stage1_55[69], stage1_55[70], stage1_55[71], stage1_55[72]},
      {stage1_56[72], stage1_56[73], stage1_56[74]},
      {stage1_57[12]},
      {stage1_58[24], stage1_58[25]},
      {stage2_59[12],stage2_58[18],stage2_57[19],stage2_56[47],stage2_55[61]}
   );
   gpc2135_5 gpc5674 (
      {stage1_55[73], stage1_55[74], stage1_55[75], stage1_55[76], stage1_55[77]},
      {stage1_56[75], stage1_56[76], stage1_56[77]},
      {stage1_57[13]},
      {stage1_58[26], stage1_58[27]},
      {stage2_59[13],stage2_58[19],stage2_57[20],stage2_56[48],stage2_55[62]}
   );
   gpc2135_5 gpc5675 (
      {stage1_55[78], stage1_55[79], stage1_55[80], stage1_55[81], stage1_55[82]},
      {stage1_56[78], stage1_56[79], stage1_56[80]},
      {stage1_57[14]},
      {stage1_58[28], stage1_58[29]},
      {stage2_59[14],stage2_58[20],stage2_57[21],stage2_56[49],stage2_55[63]}
   );
   gpc2135_5 gpc5676 (
      {stage1_55[83], stage1_55[84], stage1_55[85], stage1_55[86], stage1_55[87]},
      {stage1_56[81], stage1_56[82], stage1_56[83]},
      {stage1_57[15]},
      {stage1_58[30], stage1_58[31]},
      {stage2_59[15],stage2_58[21],stage2_57[22],stage2_56[50],stage2_55[64]}
   );
   gpc2135_5 gpc5677 (
      {stage1_55[88], stage1_55[89], stage1_55[90], stage1_55[91], stage1_55[92]},
      {stage1_56[84], stage1_56[85], stage1_56[86]},
      {stage1_57[16]},
      {stage1_58[32], stage1_58[33]},
      {stage2_59[16],stage2_58[22],stage2_57[23],stage2_56[51],stage2_55[65]}
   );
   gpc2135_5 gpc5678 (
      {stage1_55[93], stage1_55[94], stage1_55[95], stage1_55[96], stage1_55[97]},
      {stage1_56[87], stage1_56[88], stage1_56[89]},
      {stage1_57[17]},
      {stage1_58[34], stage1_58[35]},
      {stage2_59[17],stage2_58[23],stage2_57[24],stage2_56[52],stage2_55[66]}
   );
   gpc606_5 gpc5679 (
      {stage1_55[98], stage1_55[99], stage1_55[100], stage1_55[101], stage1_55[102], stage1_55[103]},
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22], stage1_57[23]},
      {stage2_59[18],stage2_58[24],stage2_57[25],stage2_56[53],stage2_55[67]}
   );
   gpc606_5 gpc5680 (
      {stage1_55[104], stage1_55[105], stage1_55[106], stage1_55[107], stage1_55[108], stage1_55[109]},
      {stage1_57[24], stage1_57[25], stage1_57[26], stage1_57[27], stage1_57[28], stage1_57[29]},
      {stage2_59[19],stage2_58[25],stage2_57[26],stage2_56[54],stage2_55[68]}
   );
   gpc606_5 gpc5681 (
      {stage1_55[110], stage1_55[111], stage1_55[112], stage1_55[113], stage1_55[114], stage1_55[115]},
      {stage1_57[30], stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35]},
      {stage2_59[20],stage2_58[26],stage2_57[27],stage2_56[55],stage2_55[69]}
   );
   gpc606_5 gpc5682 (
      {stage1_55[116], stage1_55[117], stage1_55[118], stage1_55[119], stage1_55[120], stage1_55[121]},
      {stage1_57[36], stage1_57[37], stage1_57[38], stage1_57[39], stage1_57[40], stage1_57[41]},
      {stage2_59[21],stage2_58[27],stage2_57[28],stage2_56[56],stage2_55[70]}
   );
   gpc606_5 gpc5683 (
      {stage1_55[122], stage1_55[123], stage1_55[124], stage1_55[125], stage1_55[126], stage1_55[127]},
      {stage1_57[42], stage1_57[43], stage1_57[44], stage1_57[45], stage1_57[46], stage1_57[47]},
      {stage2_59[22],stage2_58[28],stage2_57[29],stage2_56[57],stage2_55[71]}
   );
   gpc606_5 gpc5684 (
      {stage1_55[128], stage1_55[129], stage1_55[130], stage1_55[131], stage1_55[132], stage1_55[133]},
      {stage1_57[48], stage1_57[49], stage1_57[50], stage1_57[51], stage1_57[52], stage1_57[53]},
      {stage2_59[23],stage2_58[29],stage2_57[30],stage2_56[58],stage2_55[72]}
   );
   gpc606_5 gpc5685 (
      {stage1_55[134], stage1_55[135], stage1_55[136], stage1_55[137], stage1_55[138], stage1_55[139]},
      {stage1_57[54], stage1_57[55], stage1_57[56], stage1_57[57], stage1_57[58], stage1_57[59]},
      {stage2_59[24],stage2_58[30],stage2_57[31],stage2_56[59],stage2_55[73]}
   );
   gpc606_5 gpc5686 (
      {stage1_55[140], stage1_55[141], stage1_55[142], stage1_55[143], stage1_55[144], stage1_55[145]},
      {stage1_57[60], stage1_57[61], stage1_57[62], stage1_57[63], stage1_57[64], stage1_57[65]},
      {stage2_59[25],stage2_58[31],stage2_57[32],stage2_56[60],stage2_55[74]}
   );
   gpc606_5 gpc5687 (
      {stage1_55[146], stage1_55[147], stage1_55[148], stage1_55[149], stage1_55[150], stage1_55[151]},
      {stage1_57[66], stage1_57[67], stage1_57[68], stage1_57[69], stage1_57[70], stage1_57[71]},
      {stage2_59[26],stage2_58[32],stage2_57[33],stage2_56[61],stage2_55[75]}
   );
   gpc606_5 gpc5688 (
      {stage1_55[152], stage1_55[153], stage1_55[154], stage1_55[155], stage1_55[156], stage1_55[157]},
      {stage1_57[72], stage1_57[73], stage1_57[74], stage1_57[75], stage1_57[76], stage1_57[77]},
      {stage2_59[27],stage2_58[33],stage2_57[34],stage2_56[62],stage2_55[76]}
   );
   gpc606_5 gpc5689 (
      {stage1_55[158], stage1_55[159], stage1_55[160], stage1_55[161], stage1_55[162], stage1_55[163]},
      {stage1_57[78], stage1_57[79], stage1_57[80], stage1_57[81], stage1_57[82], stage1_57[83]},
      {stage2_59[28],stage2_58[34],stage2_57[35],stage2_56[63],stage2_55[77]}
   );
   gpc606_5 gpc5690 (
      {stage1_55[164], stage1_55[165], stage1_55[166], stage1_55[167], stage1_55[168], stage1_55[169]},
      {stage1_57[84], stage1_57[85], stage1_57[86], stage1_57[87], stage1_57[88], stage1_57[89]},
      {stage2_59[29],stage2_58[35],stage2_57[36],stage2_56[64],stage2_55[78]}
   );
   gpc606_5 gpc5691 (
      {stage1_55[170], stage1_55[171], stage1_55[172], stage1_55[173], stage1_55[174], stage1_55[175]},
      {stage1_57[90], stage1_57[91], stage1_57[92], stage1_57[93], stage1_57[94], stage1_57[95]},
      {stage2_59[30],stage2_58[36],stage2_57[37],stage2_56[65],stage2_55[79]}
   );
   gpc606_5 gpc5692 (
      {stage1_55[176], stage1_55[177], stage1_55[178], stage1_55[179], stage1_55[180], stage1_55[181]},
      {stage1_57[96], stage1_57[97], stage1_57[98], stage1_57[99], stage1_57[100], stage1_57[101]},
      {stage2_59[31],stage2_58[37],stage2_57[38],stage2_56[66],stage2_55[80]}
   );
   gpc606_5 gpc5693 (
      {stage1_55[182], stage1_55[183], stage1_55[184], stage1_55[185], stage1_55[186], stage1_55[187]},
      {stage1_57[102], stage1_57[103], stage1_57[104], stage1_57[105], stage1_57[106], stage1_57[107]},
      {stage2_59[32],stage2_58[38],stage2_57[39],stage2_56[67],stage2_55[81]}
   );
   gpc606_5 gpc5694 (
      {stage1_55[188], stage1_55[189], stage1_55[190], stage1_55[191], stage1_55[192], stage1_55[193]},
      {stage1_57[108], stage1_57[109], stage1_57[110], stage1_57[111], stage1_57[112], stage1_57[113]},
      {stage2_59[33],stage2_58[39],stage2_57[40],stage2_56[68],stage2_55[82]}
   );
   gpc606_5 gpc5695 (
      {stage1_55[194], stage1_55[195], stage1_55[196], stage1_55[197], stage1_55[198], stage1_55[199]},
      {stage1_57[114], stage1_57[115], stage1_57[116], stage1_57[117], stage1_57[118], stage1_57[119]},
      {stage2_59[34],stage2_58[40],stage2_57[41],stage2_56[69],stage2_55[83]}
   );
   gpc606_5 gpc5696 (
      {stage1_55[200], stage1_55[201], stage1_55[202], stage1_55[203], stage1_55[204], stage1_55[205]},
      {stage1_57[120], stage1_57[121], stage1_57[122], stage1_57[123], stage1_57[124], stage1_57[125]},
      {stage2_59[35],stage2_58[41],stage2_57[42],stage2_56[70],stage2_55[84]}
   );
   gpc606_5 gpc5697 (
      {stage1_55[206], stage1_55[207], stage1_55[208], stage1_55[209], stage1_55[210], stage1_55[211]},
      {stage1_57[126], stage1_57[127], stage1_57[128], stage1_57[129], stage1_57[130], stage1_57[131]},
      {stage2_59[36],stage2_58[42],stage2_57[43],stage2_56[71],stage2_55[85]}
   );
   gpc606_5 gpc5698 (
      {stage1_55[212], stage1_55[213], stage1_55[214], stage1_55[215], stage1_55[216], stage1_55[217]},
      {stage1_57[132], stage1_57[133], stage1_57[134], stage1_57[135], stage1_57[136], stage1_57[137]},
      {stage2_59[37],stage2_58[43],stage2_57[44],stage2_56[72],stage2_55[86]}
   );
   gpc606_5 gpc5699 (
      {stage1_55[218], stage1_55[219], stage1_55[220], stage1_55[221], stage1_55[222], stage1_55[223]},
      {stage1_57[138], stage1_57[139], stage1_57[140], stage1_57[141], stage1_57[142], stage1_57[143]},
      {stage2_59[38],stage2_58[44],stage2_57[45],stage2_56[73],stage2_55[87]}
   );
   gpc606_5 gpc5700 (
      {stage1_55[224], stage1_55[225], stage1_55[226], stage1_55[227], stage1_55[228], stage1_55[229]},
      {stage1_57[144], stage1_57[145], stage1_57[146], stage1_57[147], stage1_57[148], stage1_57[149]},
      {stage2_59[39],stage2_58[45],stage2_57[46],stage2_56[74],stage2_55[88]}
   );
   gpc606_5 gpc5701 (
      {stage1_55[230], stage1_55[231], stage1_55[232], stage1_55[233], stage1_55[234], stage1_55[235]},
      {stage1_57[150], stage1_57[151], stage1_57[152], stage1_57[153], stage1_57[154], stage1_57[155]},
      {stage2_59[40],stage2_58[46],stage2_57[47],stage2_56[75],stage2_55[89]}
   );
   gpc606_5 gpc5702 (
      {stage1_55[236], stage1_55[237], stage1_55[238], stage1_55[239], stage1_55[240], stage1_55[241]},
      {stage1_57[156], stage1_57[157], stage1_57[158], stage1_57[159], stage1_57[160], stage1_57[161]},
      {stage2_59[41],stage2_58[47],stage2_57[48],stage2_56[76],stage2_55[90]}
   );
   gpc606_5 gpc5703 (
      {stage1_55[242], stage1_55[243], stage1_55[244], stage1_55[245], stage1_55[246], stage1_55[247]},
      {stage1_57[162], stage1_57[163], stage1_57[164], stage1_57[165], stage1_57[166], stage1_57[167]},
      {stage2_59[42],stage2_58[48],stage2_57[49],stage2_56[77],stage2_55[91]}
   );
   gpc606_5 gpc5704 (
      {stage1_55[248], stage1_55[249], stage1_55[250], stage1_55[251], stage1_55[252], stage1_55[253]},
      {stage1_57[168], stage1_57[169], stage1_57[170], stage1_57[171], stage1_57[172], stage1_57[173]},
      {stage2_59[43],stage2_58[49],stage2_57[50],stage2_56[78],stage2_55[92]}
   );
   gpc606_5 gpc5705 (
      {stage1_56[90], stage1_56[91], stage1_56[92], stage1_56[93], stage1_56[94], stage1_56[95]},
      {stage1_58[36], stage1_58[37], stage1_58[38], stage1_58[39], stage1_58[40], stage1_58[41]},
      {stage2_60[0],stage2_59[44],stage2_58[50],stage2_57[51],stage2_56[79]}
   );
   gpc606_5 gpc5706 (
      {stage1_56[96], stage1_56[97], stage1_56[98], stage1_56[99], stage1_56[100], stage1_56[101]},
      {stage1_58[42], stage1_58[43], stage1_58[44], stage1_58[45], stage1_58[46], stage1_58[47]},
      {stage2_60[1],stage2_59[45],stage2_58[51],stage2_57[52],stage2_56[80]}
   );
   gpc606_5 gpc5707 (
      {stage1_56[102], stage1_56[103], stage1_56[104], stage1_56[105], stage1_56[106], stage1_56[107]},
      {stage1_58[48], stage1_58[49], stage1_58[50], stage1_58[51], stage1_58[52], stage1_58[53]},
      {stage2_60[2],stage2_59[46],stage2_58[52],stage2_57[53],stage2_56[81]}
   );
   gpc606_5 gpc5708 (
      {stage1_56[108], stage1_56[109], stage1_56[110], stage1_56[111], stage1_56[112], stage1_56[113]},
      {stage1_58[54], stage1_58[55], stage1_58[56], stage1_58[57], stage1_58[58], stage1_58[59]},
      {stage2_60[3],stage2_59[47],stage2_58[53],stage2_57[54],stage2_56[82]}
   );
   gpc606_5 gpc5709 (
      {stage1_56[114], stage1_56[115], stage1_56[116], stage1_56[117], stage1_56[118], stage1_56[119]},
      {stage1_58[60], stage1_58[61], stage1_58[62], stage1_58[63], stage1_58[64], stage1_58[65]},
      {stage2_60[4],stage2_59[48],stage2_58[54],stage2_57[55],stage2_56[83]}
   );
   gpc606_5 gpc5710 (
      {stage1_56[120], stage1_56[121], stage1_56[122], stage1_56[123], stage1_56[124], stage1_56[125]},
      {stage1_58[66], stage1_58[67], stage1_58[68], stage1_58[69], stage1_58[70], stage1_58[71]},
      {stage2_60[5],stage2_59[49],stage2_58[55],stage2_57[56],stage2_56[84]}
   );
   gpc606_5 gpc5711 (
      {stage1_56[126], stage1_56[127], stage1_56[128], stage1_56[129], stage1_56[130], stage1_56[131]},
      {stage1_58[72], stage1_58[73], stage1_58[74], stage1_58[75], stage1_58[76], stage1_58[77]},
      {stage2_60[6],stage2_59[50],stage2_58[56],stage2_57[57],stage2_56[85]}
   );
   gpc606_5 gpc5712 (
      {stage1_56[132], stage1_56[133], stage1_56[134], stage1_56[135], stage1_56[136], stage1_56[137]},
      {stage1_58[78], stage1_58[79], stage1_58[80], stage1_58[81], stage1_58[82], stage1_58[83]},
      {stage2_60[7],stage2_59[51],stage2_58[57],stage2_57[58],stage2_56[86]}
   );
   gpc606_5 gpc5713 (
      {stage1_56[138], stage1_56[139], stage1_56[140], stage1_56[141], stage1_56[142], stage1_56[143]},
      {stage1_58[84], stage1_58[85], stage1_58[86], stage1_58[87], stage1_58[88], stage1_58[89]},
      {stage2_60[8],stage2_59[52],stage2_58[58],stage2_57[59],stage2_56[87]}
   );
   gpc615_5 gpc5714 (
      {stage1_56[144], stage1_56[145], stage1_56[146], stage1_56[147], stage1_56[148]},
      {stage1_57[174]},
      {stage1_58[90], stage1_58[91], stage1_58[92], stage1_58[93], stage1_58[94], stage1_58[95]},
      {stage2_60[9],stage2_59[53],stage2_58[59],stage2_57[60],stage2_56[88]}
   );
   gpc615_5 gpc5715 (
      {stage1_56[149], stage1_56[150], stage1_56[151], stage1_56[152], stage1_56[153]},
      {stage1_57[175]},
      {stage1_58[96], stage1_58[97], stage1_58[98], stage1_58[99], stage1_58[100], stage1_58[101]},
      {stage2_60[10],stage2_59[54],stage2_58[60],stage2_57[61],stage2_56[89]}
   );
   gpc615_5 gpc5716 (
      {stage1_56[154], stage1_56[155], stage1_56[156], stage1_56[157], stage1_56[158]},
      {stage1_57[176]},
      {stage1_58[102], stage1_58[103], stage1_58[104], stage1_58[105], stage1_58[106], stage1_58[107]},
      {stage2_60[11],stage2_59[55],stage2_58[61],stage2_57[62],stage2_56[90]}
   );
   gpc615_5 gpc5717 (
      {stage1_56[159], stage1_56[160], stage1_56[161], stage1_56[162], stage1_56[163]},
      {stage1_57[177]},
      {stage1_58[108], stage1_58[109], stage1_58[110], stage1_58[111], stage1_58[112], stage1_58[113]},
      {stage2_60[12],stage2_59[56],stage2_58[62],stage2_57[63],stage2_56[91]}
   );
   gpc606_5 gpc5718 (
      {stage1_57[178], stage1_57[179], stage1_57[180], stage1_57[181], stage1_57[182], stage1_57[183]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[13],stage2_59[57],stage2_58[63],stage2_57[64]}
   );
   gpc615_5 gpc5719 (
      {stage1_57[184], stage1_57[185], stage1_57[186], stage1_57[187], stage1_57[188]},
      {stage1_58[114]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[14],stage2_59[58],stage2_58[64],stage2_57[65]}
   );
   gpc615_5 gpc5720 (
      {stage1_58[115], stage1_58[116], stage1_58[117], stage1_58[118], stage1_58[119]},
      {stage1_59[12]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[2],stage2_60[15],stage2_59[59],stage2_58[65]}
   );
   gpc615_5 gpc5721 (
      {stage1_58[120], stage1_58[121], stage1_58[122], stage1_58[123], stage1_58[124]},
      {stage1_59[13]},
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage2_62[1],stage2_61[3],stage2_60[16],stage2_59[60],stage2_58[66]}
   );
   gpc615_5 gpc5722 (
      {stage1_58[125], stage1_58[126], stage1_58[127], stage1_58[128], stage1_58[129]},
      {stage1_59[14]},
      {stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage2_62[2],stage2_61[4],stage2_60[17],stage2_59[61],stage2_58[67]}
   );
   gpc615_5 gpc5723 (
      {stage1_58[130], stage1_58[131], stage1_58[132], stage1_58[133], stage1_58[134]},
      {stage1_59[15]},
      {stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21], stage1_60[22], stage1_60[23]},
      {stage2_62[3],stage2_61[5],stage2_60[18],stage2_59[62],stage2_58[68]}
   );
   gpc615_5 gpc5724 (
      {stage1_58[135], stage1_58[136], stage1_58[137], stage1_58[138], stage1_58[139]},
      {stage1_59[16]},
      {stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27], stage1_60[28], stage1_60[29]},
      {stage2_62[4],stage2_61[6],stage2_60[19],stage2_59[63],stage2_58[69]}
   );
   gpc615_5 gpc5725 (
      {stage1_58[140], stage1_58[141], stage1_58[142], stage1_58[143], stage1_58[144]},
      {stage1_59[17]},
      {stage1_60[30], stage1_60[31], stage1_60[32], stage1_60[33], stage1_60[34], stage1_60[35]},
      {stage2_62[5],stage2_61[7],stage2_60[20],stage2_59[64],stage2_58[70]}
   );
   gpc615_5 gpc5726 (
      {stage1_58[145], stage1_58[146], stage1_58[147], stage1_58[148], stage1_58[149]},
      {stage1_59[18]},
      {stage1_60[36], stage1_60[37], stage1_60[38], stage1_60[39], stage1_60[40], stage1_60[41]},
      {stage2_62[6],stage2_61[8],stage2_60[21],stage2_59[65],stage2_58[71]}
   );
   gpc615_5 gpc5727 (
      {stage1_58[150], stage1_58[151], stage1_58[152], stage1_58[153], stage1_58[154]},
      {stage1_59[19]},
      {stage1_60[42], stage1_60[43], stage1_60[44], stage1_60[45], stage1_60[46], stage1_60[47]},
      {stage2_62[7],stage2_61[9],stage2_60[22],stage2_59[66],stage2_58[72]}
   );
   gpc615_5 gpc5728 (
      {stage1_58[155], stage1_58[156], stage1_58[157], stage1_58[158], stage1_58[159]},
      {stage1_59[20]},
      {stage1_60[48], stage1_60[49], stage1_60[50], stage1_60[51], stage1_60[52], stage1_60[53]},
      {stage2_62[8],stage2_61[10],stage2_60[23],stage2_59[67],stage2_58[73]}
   );
   gpc615_5 gpc5729 (
      {stage1_58[160], stage1_58[161], stage1_58[162], stage1_58[163], stage1_58[164]},
      {stage1_59[21]},
      {stage1_60[54], stage1_60[55], stage1_60[56], stage1_60[57], stage1_60[58], stage1_60[59]},
      {stage2_62[9],stage2_61[11],stage2_60[24],stage2_59[68],stage2_58[74]}
   );
   gpc615_5 gpc5730 (
      {stage1_58[165], stage1_58[166], stage1_58[167], stage1_58[168], stage1_58[169]},
      {stage1_59[22]},
      {stage1_60[60], stage1_60[61], stage1_60[62], stage1_60[63], stage1_60[64], stage1_60[65]},
      {stage2_62[10],stage2_61[12],stage2_60[25],stage2_59[69],stage2_58[75]}
   );
   gpc615_5 gpc5731 (
      {stage1_58[170], stage1_58[171], stage1_58[172], stage1_58[173], stage1_58[174]},
      {stage1_59[23]},
      {stage1_60[66], stage1_60[67], stage1_60[68], stage1_60[69], stage1_60[70], stage1_60[71]},
      {stage2_62[11],stage2_61[13],stage2_60[26],stage2_59[70],stage2_58[76]}
   );
   gpc615_5 gpc5732 (
      {stage1_58[175], stage1_58[176], stage1_58[177], stage1_58[178], stage1_58[179]},
      {stage1_59[24]},
      {stage1_60[72], stage1_60[73], stage1_60[74], stage1_60[75], stage1_60[76], stage1_60[77]},
      {stage2_62[12],stage2_61[14],stage2_60[27],stage2_59[71],stage2_58[77]}
   );
   gpc615_5 gpc5733 (
      {stage1_58[180], stage1_58[181], stage1_58[182], stage1_58[183], stage1_58[184]},
      {stage1_59[25]},
      {stage1_60[78], stage1_60[79], stage1_60[80], stage1_60[81], stage1_60[82], stage1_60[83]},
      {stage2_62[13],stage2_61[15],stage2_60[28],stage2_59[72],stage2_58[78]}
   );
   gpc615_5 gpc5734 (
      {stage1_58[185], stage1_58[186], stage1_58[187], stage1_58[188], stage1_58[189]},
      {stage1_59[26]},
      {stage1_60[84], stage1_60[85], stage1_60[86], stage1_60[87], stage1_60[88], stage1_60[89]},
      {stage2_62[14],stage2_61[16],stage2_60[29],stage2_59[73],stage2_58[79]}
   );
   gpc615_5 gpc5735 (
      {stage1_58[190], stage1_58[191], stage1_58[192], stage1_58[193], stage1_58[194]},
      {stage1_59[27]},
      {stage1_60[90], stage1_60[91], stage1_60[92], stage1_60[93], stage1_60[94], stage1_60[95]},
      {stage2_62[15],stage2_61[17],stage2_60[30],stage2_59[74],stage2_58[80]}
   );
   gpc615_5 gpc5736 (
      {stage1_58[195], stage1_58[196], stage1_58[197], stage1_58[198], stage1_58[199]},
      {stage1_59[28]},
      {stage1_60[96], stage1_60[97], stage1_60[98], stage1_60[99], stage1_60[100], stage1_60[101]},
      {stage2_62[16],stage2_61[18],stage2_60[31],stage2_59[75],stage2_58[81]}
   );
   gpc615_5 gpc5737 (
      {stage1_58[200], stage1_58[201], stage1_58[202], stage1_58[203], stage1_58[204]},
      {stage1_59[29]},
      {stage1_60[102], stage1_60[103], stage1_60[104], stage1_60[105], stage1_60[106], stage1_60[107]},
      {stage2_62[17],stage2_61[19],stage2_60[32],stage2_59[76],stage2_58[82]}
   );
   gpc615_5 gpc5738 (
      {stage1_58[205], stage1_58[206], stage1_58[207], stage1_58[208], stage1_58[209]},
      {stage1_59[30]},
      {stage1_60[108], stage1_60[109], stage1_60[110], stage1_60[111], stage1_60[112], stage1_60[113]},
      {stage2_62[18],stage2_61[20],stage2_60[33],stage2_59[77],stage2_58[83]}
   );
   gpc615_5 gpc5739 (
      {stage1_58[210], stage1_58[211], stage1_58[212], stage1_58[213], stage1_58[214]},
      {stage1_59[31]},
      {stage1_60[114], stage1_60[115], stage1_60[116], stage1_60[117], stage1_60[118], stage1_60[119]},
      {stage2_62[19],stage2_61[21],stage2_60[34],stage2_59[78],stage2_58[84]}
   );
   gpc615_5 gpc5740 (
      {stage1_58[215], stage1_58[216], stage1_58[217], stage1_58[218], stage1_58[219]},
      {stage1_59[32]},
      {stage1_60[120], stage1_60[121], stage1_60[122], stage1_60[123], stage1_60[124], stage1_60[125]},
      {stage2_62[20],stage2_61[22],stage2_60[35],stage2_59[79],stage2_58[85]}
   );
   gpc2135_5 gpc5741 (
      {stage1_59[33], stage1_59[34], stage1_59[35], stage1_59[36], stage1_59[37]},
      {stage1_60[126], stage1_60[127], stage1_60[128]},
      {stage1_61[0]},
      {stage1_62[0], stage1_62[1]},
      {stage2_63[0],stage2_62[21],stage2_61[23],stage2_60[36],stage2_59[80]}
   );
   gpc606_5 gpc5742 (
      {stage1_59[38], stage1_59[39], stage1_59[40], stage1_59[41], stage1_59[42], stage1_59[43]},
      {stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5], stage1_61[6]},
      {stage2_63[1],stage2_62[22],stage2_61[24],stage2_60[37],stage2_59[81]}
   );
   gpc606_5 gpc5743 (
      {stage1_59[44], stage1_59[45], stage1_59[46], stage1_59[47], stage1_59[48], stage1_59[49]},
      {stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11], stage1_61[12]},
      {stage2_63[2],stage2_62[23],stage2_61[25],stage2_60[38],stage2_59[82]}
   );
   gpc606_5 gpc5744 (
      {stage1_59[50], stage1_59[51], stage1_59[52], stage1_59[53], stage1_59[54], stage1_59[55]},
      {stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17], stage1_61[18]},
      {stage2_63[3],stage2_62[24],stage2_61[26],stage2_60[39],stage2_59[83]}
   );
   gpc606_5 gpc5745 (
      {stage1_59[56], stage1_59[57], stage1_59[58], stage1_59[59], stage1_59[60], stage1_59[61]},
      {stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23], stage1_61[24]},
      {stage2_63[4],stage2_62[25],stage2_61[27],stage2_60[40],stage2_59[84]}
   );
   gpc606_5 gpc5746 (
      {stage1_59[62], stage1_59[63], stage1_59[64], stage1_59[65], stage1_59[66], stage1_59[67]},
      {stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29], stage1_61[30]},
      {stage2_63[5],stage2_62[26],stage2_61[28],stage2_60[41],stage2_59[85]}
   );
   gpc606_5 gpc5747 (
      {stage1_59[68], stage1_59[69], stage1_59[70], stage1_59[71], stage1_59[72], stage1_59[73]},
      {stage1_61[31], stage1_61[32], stage1_61[33], stage1_61[34], stage1_61[35], stage1_61[36]},
      {stage2_63[6],stage2_62[27],stage2_61[29],stage2_60[42],stage2_59[86]}
   );
   gpc606_5 gpc5748 (
      {stage1_59[74], stage1_59[75], stage1_59[76], stage1_59[77], stage1_59[78], stage1_59[79]},
      {stage1_61[37], stage1_61[38], stage1_61[39], stage1_61[40], stage1_61[41], stage1_61[42]},
      {stage2_63[7],stage2_62[28],stage2_61[30],stage2_60[43],stage2_59[87]}
   );
   gpc606_5 gpc5749 (
      {stage1_59[80], stage1_59[81], stage1_59[82], stage1_59[83], stage1_59[84], stage1_59[85]},
      {stage1_61[43], stage1_61[44], stage1_61[45], stage1_61[46], stage1_61[47], stage1_61[48]},
      {stage2_63[8],stage2_62[29],stage2_61[31],stage2_60[44],stage2_59[88]}
   );
   gpc606_5 gpc5750 (
      {stage1_59[86], stage1_59[87], stage1_59[88], stage1_59[89], stage1_59[90], stage1_59[91]},
      {stage1_61[49], stage1_61[50], stage1_61[51], stage1_61[52], stage1_61[53], stage1_61[54]},
      {stage2_63[9],stage2_62[30],stage2_61[32],stage2_60[45],stage2_59[89]}
   );
   gpc606_5 gpc5751 (
      {stage1_59[92], stage1_59[93], stage1_59[94], stage1_59[95], stage1_59[96], stage1_59[97]},
      {stage1_61[55], stage1_61[56], stage1_61[57], stage1_61[58], stage1_61[59], stage1_61[60]},
      {stage2_63[10],stage2_62[31],stage2_61[33],stage2_60[46],stage2_59[90]}
   );
   gpc606_5 gpc5752 (
      {stage1_59[98], stage1_59[99], stage1_59[100], stage1_59[101], stage1_59[102], stage1_59[103]},
      {stage1_61[61], stage1_61[62], stage1_61[63], stage1_61[64], stage1_61[65], stage1_61[66]},
      {stage2_63[11],stage2_62[32],stage2_61[34],stage2_60[47],stage2_59[91]}
   );
   gpc606_5 gpc5753 (
      {stage1_59[104], stage1_59[105], stage1_59[106], stage1_59[107], stage1_59[108], stage1_59[109]},
      {stage1_61[67], stage1_61[68], stage1_61[69], stage1_61[70], stage1_61[71], stage1_61[72]},
      {stage2_63[12],stage2_62[33],stage2_61[35],stage2_60[48],stage2_59[92]}
   );
   gpc606_5 gpc5754 (
      {stage1_59[110], stage1_59[111], stage1_59[112], stage1_59[113], stage1_59[114], stage1_59[115]},
      {stage1_61[73], stage1_61[74], stage1_61[75], stage1_61[76], stage1_61[77], stage1_61[78]},
      {stage2_63[13],stage2_62[34],stage2_61[36],stage2_60[49],stage2_59[93]}
   );
   gpc606_5 gpc5755 (
      {stage1_59[116], stage1_59[117], stage1_59[118], stage1_59[119], stage1_59[120], stage1_59[121]},
      {stage1_61[79], stage1_61[80], stage1_61[81], stage1_61[82], stage1_61[83], stage1_61[84]},
      {stage2_63[14],stage2_62[35],stage2_61[37],stage2_60[50],stage2_59[94]}
   );
   gpc606_5 gpc5756 (
      {stage1_59[122], stage1_59[123], stage1_59[124], stage1_59[125], stage1_59[126], stage1_59[127]},
      {stage1_61[85], stage1_61[86], stage1_61[87], stage1_61[88], stage1_61[89], stage1_61[90]},
      {stage2_63[15],stage2_62[36],stage2_61[38],stage2_60[51],stage2_59[95]}
   );
   gpc606_5 gpc5757 (
      {stage1_59[128], stage1_59[129], stage1_59[130], stage1_59[131], stage1_59[132], stage1_59[133]},
      {stage1_61[91], stage1_61[92], stage1_61[93], stage1_61[94], stage1_61[95], stage1_61[96]},
      {stage2_63[16],stage2_62[37],stage2_61[39],stage2_60[52],stage2_59[96]}
   );
   gpc606_5 gpc5758 (
      {stage1_59[134], stage1_59[135], stage1_59[136], stage1_59[137], stage1_59[138], stage1_59[139]},
      {stage1_61[97], stage1_61[98], stage1_61[99], stage1_61[100], stage1_61[101], stage1_61[102]},
      {stage2_63[17],stage2_62[38],stage2_61[40],stage2_60[53],stage2_59[97]}
   );
   gpc606_5 gpc5759 (
      {stage1_59[140], stage1_59[141], stage1_59[142], stage1_59[143], stage1_59[144], stage1_59[145]},
      {stage1_61[103], stage1_61[104], stage1_61[105], stage1_61[106], stage1_61[107], stage1_61[108]},
      {stage2_63[18],stage2_62[39],stage2_61[41],stage2_60[54],stage2_59[98]}
   );
   gpc606_5 gpc5760 (
      {stage1_59[146], stage1_59[147], stage1_59[148], stage1_59[149], stage1_59[150], stage1_59[151]},
      {stage1_61[109], stage1_61[110], stage1_61[111], stage1_61[112], stage1_61[113], stage1_61[114]},
      {stage2_63[19],stage2_62[40],stage2_61[42],stage2_60[55],stage2_59[99]}
   );
   gpc606_5 gpc5761 (
      {stage1_59[152], stage1_59[153], stage1_59[154], stage1_59[155], stage1_59[156], stage1_59[157]},
      {stage1_61[115], stage1_61[116], stage1_61[117], stage1_61[118], stage1_61[119], stage1_61[120]},
      {stage2_63[20],stage2_62[41],stage2_61[43],stage2_60[56],stage2_59[100]}
   );
   gpc606_5 gpc5762 (
      {stage1_59[158], stage1_59[159], stage1_59[160], stage1_59[161], stage1_59[162], stage1_59[163]},
      {stage1_61[121], stage1_61[122], stage1_61[123], stage1_61[124], stage1_61[125], stage1_61[126]},
      {stage2_63[21],stage2_62[42],stage2_61[44],stage2_60[57],stage2_59[101]}
   );
   gpc606_5 gpc5763 (
      {stage1_59[164], stage1_59[165], stage1_59[166], stage1_59[167], stage1_59[168], stage1_59[169]},
      {stage1_61[127], stage1_61[128], stage1_61[129], stage1_61[130], stage1_61[131], stage1_61[132]},
      {stage2_63[22],stage2_62[43],stage2_61[45],stage2_60[58],stage2_59[102]}
   );
   gpc606_5 gpc5764 (
      {stage1_59[170], stage1_59[171], stage1_59[172], stage1_59[173], stage1_59[174], stage1_59[175]},
      {stage1_61[133], stage1_61[134], stage1_61[135], stage1_61[136], stage1_61[137], stage1_61[138]},
      {stage2_63[23],stage2_62[44],stage2_61[46],stage2_60[59],stage2_59[103]}
   );
   gpc606_5 gpc5765 (
      {stage1_59[176], stage1_59[177], stage1_59[178], stage1_59[179], stage1_59[180], stage1_59[181]},
      {stage1_61[139], stage1_61[140], stage1_61[141], stage1_61[142], stage1_61[143], stage1_61[144]},
      {stage2_63[24],stage2_62[45],stage2_61[47],stage2_60[60],stage2_59[104]}
   );
   gpc606_5 gpc5766 (
      {stage1_59[182], stage1_59[183], stage1_59[184], stage1_59[185], stage1_59[186], stage1_59[187]},
      {stage1_61[145], stage1_61[146], stage1_61[147], stage1_61[148], stage1_61[149], stage1_61[150]},
      {stage2_63[25],stage2_62[46],stage2_61[48],stage2_60[61],stage2_59[105]}
   );
   gpc606_5 gpc5767 (
      {stage1_59[188], stage1_59[189], stage1_59[190], stage1_59[191], stage1_59[192], stage1_59[193]},
      {stage1_61[151], stage1_61[152], stage1_61[153], stage1_61[154], stage1_61[155], stage1_61[156]},
      {stage2_63[26],stage2_62[47],stage2_61[49],stage2_60[62],stage2_59[106]}
   );
   gpc606_5 gpc5768 (
      {stage1_59[194], stage1_59[195], stage1_59[196], stage1_59[197], stage1_59[198], stage1_59[199]},
      {stage1_61[157], stage1_61[158], stage1_61[159], stage1_61[160], stage1_61[161], stage1_61[162]},
      {stage2_63[27],stage2_62[48],stage2_61[50],stage2_60[63],stage2_59[107]}
   );
   gpc615_5 gpc5769 (
      {stage1_59[200], stage1_59[201], stage1_59[202], stage1_59[203], stage1_59[204]},
      {stage1_60[129]},
      {stage1_61[163], stage1_61[164], stage1_61[165], stage1_61[166], stage1_61[167], stage1_61[168]},
      {stage2_63[28],stage2_62[49],stage2_61[51],stage2_60[64],stage2_59[108]}
   );
   gpc606_5 gpc5770 (
      {stage1_60[130], stage1_60[131], stage1_60[132], stage1_60[133], stage1_60[134], stage1_60[135]},
      {stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5], stage1_62[6], stage1_62[7]},
      {stage2_64[0],stage2_63[29],stage2_62[50],stage2_61[52],stage2_60[65]}
   );
   gpc606_5 gpc5771 (
      {stage1_60[136], stage1_60[137], stage1_60[138], stage1_60[139], stage1_60[140], stage1_60[141]},
      {stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11], stage1_62[12], stage1_62[13]},
      {stage2_64[1],stage2_63[30],stage2_62[51],stage2_61[53],stage2_60[66]}
   );
   gpc606_5 gpc5772 (
      {stage1_60[142], stage1_60[143], stage1_60[144], stage1_60[145], stage1_60[146], stage1_60[147]},
      {stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17], stage1_62[18], stage1_62[19]},
      {stage2_64[2],stage2_63[31],stage2_62[52],stage2_61[54],stage2_60[67]}
   );
   gpc606_5 gpc5773 (
      {stage1_60[148], stage1_60[149], stage1_60[150], stage1_60[151], stage1_60[152], stage1_60[153]},
      {stage1_62[20], stage1_62[21], stage1_62[22], stage1_62[23], stage1_62[24], stage1_62[25]},
      {stage2_64[3],stage2_63[32],stage2_62[53],stage2_61[55],stage2_60[68]}
   );
   gpc606_5 gpc5774 (
      {stage1_60[154], stage1_60[155], stage1_60[156], stage1_60[157], stage1_60[158], stage1_60[159]},
      {stage1_62[26], stage1_62[27], stage1_62[28], stage1_62[29], stage1_62[30], stage1_62[31]},
      {stage2_64[4],stage2_63[33],stage2_62[54],stage2_61[56],stage2_60[69]}
   );
   gpc606_5 gpc5775 (
      {stage1_60[160], stage1_60[161], stage1_60[162], stage1_60[163], stage1_60[164], stage1_60[165]},
      {stage1_62[32], stage1_62[33], stage1_62[34], stage1_62[35], stage1_62[36], stage1_62[37]},
      {stage2_64[5],stage2_63[34],stage2_62[55],stage2_61[57],stage2_60[70]}
   );
   gpc606_5 gpc5776 (
      {stage1_60[166], stage1_60[167], stage1_60[168], stage1_60[169], stage1_60[170], stage1_60[171]},
      {stage1_62[38], stage1_62[39], stage1_62[40], stage1_62[41], stage1_62[42], stage1_62[43]},
      {stage2_64[6],stage2_63[35],stage2_62[56],stage2_61[58],stage2_60[71]}
   );
   gpc606_5 gpc5777 (
      {stage1_60[172], stage1_60[173], stage1_60[174], stage1_60[175], stage1_60[176], stage1_60[177]},
      {stage1_62[44], stage1_62[45], stage1_62[46], stage1_62[47], stage1_62[48], stage1_62[49]},
      {stage2_64[7],stage2_63[36],stage2_62[57],stage2_61[59],stage2_60[72]}
   );
   gpc606_5 gpc5778 (
      {stage1_60[178], stage1_60[179], stage1_60[180], stage1_60[181], stage1_60[182], stage1_60[183]},
      {stage1_62[50], stage1_62[51], stage1_62[52], stage1_62[53], stage1_62[54], stage1_62[55]},
      {stage2_64[8],stage2_63[37],stage2_62[58],stage2_61[60],stage2_60[73]}
   );
   gpc615_5 gpc5779 (
      {stage1_60[184], stage1_60[185], stage1_60[186], stage1_60[187], stage1_60[188]},
      {stage1_61[169]},
      {stage1_62[56], stage1_62[57], stage1_62[58], stage1_62[59], stage1_62[60], stage1_62[61]},
      {stage2_64[9],stage2_63[38],stage2_62[59],stage2_61[61],stage2_60[74]}
   );
   gpc615_5 gpc5780 (
      {stage1_60[189], stage1_60[190], stage1_60[191], stage1_60[192], stage1_60[193]},
      {stage1_61[170]},
      {stage1_62[62], stage1_62[63], stage1_62[64], stage1_62[65], stage1_62[66], stage1_62[67]},
      {stage2_64[10],stage2_63[39],stage2_62[60],stage2_61[62],stage2_60[75]}
   );
   gpc615_5 gpc5781 (
      {stage1_60[194], stage1_60[195], stage1_60[196], stage1_60[197], stage1_60[198]},
      {stage1_61[171]},
      {stage1_62[68], stage1_62[69], stage1_62[70], stage1_62[71], stage1_62[72], stage1_62[73]},
      {stage2_64[11],stage2_63[40],stage2_62[61],stage2_61[63],stage2_60[76]}
   );
   gpc615_5 gpc5782 (
      {stage1_60[199], stage1_60[200], stage1_60[201], stage1_60[202], stage1_60[203]},
      {stage1_61[172]},
      {stage1_62[74], stage1_62[75], stage1_62[76], stage1_62[77], stage1_62[78], stage1_62[79]},
      {stage2_64[12],stage2_63[41],stage2_62[62],stage2_61[64],stage2_60[77]}
   );
   gpc615_5 gpc5783 (
      {stage1_60[204], stage1_60[205], stage1_60[206], stage1_60[207], stage1_60[208]},
      {stage1_61[173]},
      {stage1_62[80], stage1_62[81], stage1_62[82], stage1_62[83], stage1_62[84], stage1_62[85]},
      {stage2_64[13],stage2_63[42],stage2_62[63],stage2_61[65],stage2_60[78]}
   );
   gpc615_5 gpc5784 (
      {stage1_61[174], stage1_61[175], stage1_61[176], stage1_61[177], stage1_61[178]},
      {stage1_62[86]},
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5]},
      {stage2_65[0],stage2_64[14],stage2_63[43],stage2_62[64],stage2_61[66]}
   );
   gpc615_5 gpc5785 (
      {stage1_61[179], stage1_61[180], stage1_61[181], stage1_61[182], stage1_61[183]},
      {stage1_62[87]},
      {stage1_63[6], stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11]},
      {stage2_65[1],stage2_64[15],stage2_63[44],stage2_62[65],stage2_61[67]}
   );
   gpc615_5 gpc5786 (
      {stage1_61[184], stage1_61[185], stage1_61[186], stage1_61[187], stage1_61[188]},
      {stage1_62[88]},
      {stage1_63[12], stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17]},
      {stage2_65[2],stage2_64[16],stage2_63[45],stage2_62[66],stage2_61[68]}
   );
   gpc615_5 gpc5787 (
      {stage1_61[189], stage1_61[190], stage1_61[191], stage1_61[192], stage1_61[193]},
      {stage1_62[89]},
      {stage1_63[18], stage1_63[19], stage1_63[20], stage1_63[21], stage1_63[22], stage1_63[23]},
      {stage2_65[3],stage2_64[17],stage2_63[46],stage2_62[67],stage2_61[69]}
   );
   gpc615_5 gpc5788 (
      {stage1_61[194], stage1_61[195], stage1_61[196], stage1_61[197], stage1_61[198]},
      {stage1_62[90]},
      {stage1_63[24], stage1_63[25], stage1_63[26], stage1_63[27], stage1_63[28], stage1_63[29]},
      {stage2_65[4],stage2_64[18],stage2_63[47],stage2_62[68],stage2_61[70]}
   );
   gpc615_5 gpc5789 (
      {stage1_61[199], stage1_61[200], stage1_61[201], stage1_61[202], stage1_61[203]},
      {stage1_62[91]},
      {stage1_63[30], stage1_63[31], stage1_63[32], stage1_63[33], stage1_63[34], stage1_63[35]},
      {stage2_65[5],stage2_64[19],stage2_63[48],stage2_62[69],stage2_61[71]}
   );
   gpc615_5 gpc5790 (
      {stage1_61[204], stage1_61[205], stage1_61[206], stage1_61[207], stage1_61[208]},
      {stage1_62[92]},
      {stage1_63[36], stage1_63[37], stage1_63[38], stage1_63[39], stage1_63[40], stage1_63[41]},
      {stage2_65[6],stage2_64[20],stage2_63[49],stage2_62[70],stage2_61[72]}
   );
   gpc615_5 gpc5791 (
      {stage1_61[209], stage1_61[210], stage1_61[211], stage1_61[212], stage1_61[213]},
      {stage1_62[93]},
      {stage1_63[42], stage1_63[43], stage1_63[44], stage1_63[45], stage1_63[46], stage1_63[47]},
      {stage2_65[7],stage2_64[21],stage2_63[50],stage2_62[71],stage2_61[73]}
   );
   gpc615_5 gpc5792 (
      {stage1_61[214], stage1_61[215], stage1_61[216], stage1_61[217], stage1_61[218]},
      {stage1_62[94]},
      {stage1_63[48], stage1_63[49], stage1_63[50], stage1_63[51], stage1_63[52], stage1_63[53]},
      {stage2_65[8],stage2_64[22],stage2_63[51],stage2_62[72],stage2_61[74]}
   );
   gpc1163_5 gpc5793 (
      {stage1_62[95], stage1_62[96], stage1_62[97]},
      {stage1_63[54], stage1_63[55], stage1_63[56], stage1_63[57], stage1_63[58], stage1_63[59]},
      {stage1_64[0]},
      {stage1_65[0]},
      {stage2_66[0],stage2_65[9],stage2_64[23],stage2_63[52],stage2_62[73]}
   );
   gpc1163_5 gpc5794 (
      {stage1_62[98], stage1_62[99], stage1_62[100]},
      {stage1_63[60], stage1_63[61], stage1_63[62], stage1_63[63], stage1_63[64], stage1_63[65]},
      {stage1_64[1]},
      {stage1_65[1]},
      {stage2_66[1],stage2_65[10],stage2_64[24],stage2_63[53],stage2_62[74]}
   );
   gpc1163_5 gpc5795 (
      {stage1_62[101], stage1_62[102], stage1_62[103]},
      {stage1_63[66], stage1_63[67], stage1_63[68], stage1_63[69], stage1_63[70], stage1_63[71]},
      {stage1_64[2]},
      {stage1_65[2]},
      {stage2_66[2],stage2_65[11],stage2_64[25],stage2_63[54],stage2_62[75]}
   );
   gpc1163_5 gpc5796 (
      {stage1_62[104], stage1_62[105], stage1_62[106]},
      {stage1_63[72], stage1_63[73], stage1_63[74], stage1_63[75], stage1_63[76], stage1_63[77]},
      {stage1_64[3]},
      {stage1_65[3]},
      {stage2_66[3],stage2_65[12],stage2_64[26],stage2_63[55],stage2_62[76]}
   );
   gpc1163_5 gpc5797 (
      {stage1_62[107], stage1_62[108], stage1_62[109]},
      {stage1_63[78], stage1_63[79], stage1_63[80], stage1_63[81], stage1_63[82], stage1_63[83]},
      {stage1_64[4]},
      {stage1_65[4]},
      {stage2_66[4],stage2_65[13],stage2_64[27],stage2_63[56],stage2_62[77]}
   );
   gpc1163_5 gpc5798 (
      {stage1_62[110], stage1_62[111], stage1_62[112]},
      {stage1_63[84], stage1_63[85], stage1_63[86], stage1_63[87], stage1_63[88], stage1_63[89]},
      {stage1_64[5]},
      {stage1_65[5]},
      {stage2_66[5],stage2_65[14],stage2_64[28],stage2_63[57],stage2_62[78]}
   );
   gpc1163_5 gpc5799 (
      {stage1_62[113], stage1_62[114], stage1_62[115]},
      {stage1_63[90], stage1_63[91], stage1_63[92], stage1_63[93], stage1_63[94], stage1_63[95]},
      {stage1_64[6]},
      {stage1_65[6]},
      {stage2_66[6],stage2_65[15],stage2_64[29],stage2_63[58],stage2_62[79]}
   );
   gpc1163_5 gpc5800 (
      {stage1_62[116], stage1_62[117], stage1_62[118]},
      {stage1_63[96], stage1_63[97], stage1_63[98], stage1_63[99], stage1_63[100], stage1_63[101]},
      {stage1_64[7]},
      {stage1_65[7]},
      {stage2_66[7],stage2_65[16],stage2_64[30],stage2_63[59],stage2_62[80]}
   );
   gpc1163_5 gpc5801 (
      {stage1_62[119], stage1_62[120], stage1_62[121]},
      {stage1_63[102], stage1_63[103], stage1_63[104], stage1_63[105], stage1_63[106], stage1_63[107]},
      {stage1_64[8]},
      {stage1_65[8]},
      {stage2_66[8],stage2_65[17],stage2_64[31],stage2_63[60],stage2_62[81]}
   );
   gpc1163_5 gpc5802 (
      {stage1_62[122], stage1_62[123], stage1_62[124]},
      {stage1_63[108], stage1_63[109], stage1_63[110], stage1_63[111], stage1_63[112], stage1_63[113]},
      {stage1_64[9]},
      {stage1_65[9]},
      {stage2_66[9],stage2_65[18],stage2_64[32],stage2_63[61],stage2_62[82]}
   );
   gpc1163_5 gpc5803 (
      {stage1_62[125], stage1_62[126], stage1_62[127]},
      {stage1_63[114], stage1_63[115], stage1_63[116], stage1_63[117], stage1_63[118], stage1_63[119]},
      {stage1_64[10]},
      {stage1_65[10]},
      {stage2_66[10],stage2_65[19],stage2_64[33],stage2_63[62],stage2_62[83]}
   );
   gpc1163_5 gpc5804 (
      {stage1_62[128], stage1_62[129], stage1_62[130]},
      {stage1_63[120], stage1_63[121], stage1_63[122], stage1_63[123], stage1_63[124], stage1_63[125]},
      {stage1_64[11]},
      {stage1_65[11]},
      {stage2_66[11],stage2_65[20],stage2_64[34],stage2_63[63],stage2_62[84]}
   );
   gpc1163_5 gpc5805 (
      {stage1_62[131], stage1_62[132], stage1_62[133]},
      {stage1_63[126], stage1_63[127], stage1_63[128], stage1_63[129], stage1_63[130], stage1_63[131]},
      {stage1_64[12]},
      {stage1_65[12]},
      {stage2_66[12],stage2_65[21],stage2_64[35],stage2_63[64],stage2_62[85]}
   );
   gpc1163_5 gpc5806 (
      {stage1_62[134], stage1_62[135], stage1_62[136]},
      {stage1_63[132], stage1_63[133], stage1_63[134], stage1_63[135], stage1_63[136], stage1_63[137]},
      {stage1_64[13]},
      {stage1_65[13]},
      {stage2_66[13],stage2_65[22],stage2_64[36],stage2_63[65],stage2_62[86]}
   );
   gpc1163_5 gpc5807 (
      {stage1_62[137], stage1_62[138], stage1_62[139]},
      {stage1_63[138], stage1_63[139], stage1_63[140], stage1_63[141], stage1_63[142], stage1_63[143]},
      {stage1_64[14]},
      {stage1_65[14]},
      {stage2_66[14],stage2_65[23],stage2_64[37],stage2_63[66],stage2_62[87]}
   );
   gpc1163_5 gpc5808 (
      {stage1_62[140], stage1_62[141], stage1_62[142]},
      {stage1_63[144], stage1_63[145], stage1_63[146], stage1_63[147], stage1_63[148], stage1_63[149]},
      {stage1_64[15]},
      {stage1_65[15]},
      {stage2_66[15],stage2_65[24],stage2_64[38],stage2_63[67],stage2_62[88]}
   );
   gpc1163_5 gpc5809 (
      {stage1_62[143], stage1_62[144], stage1_62[145]},
      {stage1_63[150], stage1_63[151], stage1_63[152], stage1_63[153], stage1_63[154], stage1_63[155]},
      {stage1_64[16]},
      {stage1_65[16]},
      {stage2_66[16],stage2_65[25],stage2_64[39],stage2_63[68],stage2_62[89]}
   );
   gpc1163_5 gpc5810 (
      {stage1_62[146], stage1_62[147], stage1_62[148]},
      {stage1_63[156], stage1_63[157], stage1_63[158], stage1_63[159], stage1_63[160], stage1_63[161]},
      {stage1_64[17]},
      {stage1_65[17]},
      {stage2_66[17],stage2_65[26],stage2_64[40],stage2_63[69],stage2_62[90]}
   );
   gpc1163_5 gpc5811 (
      {stage1_62[149], stage1_62[150], stage1_62[151]},
      {stage1_63[162], stage1_63[163], stage1_63[164], stage1_63[165], stage1_63[166], stage1_63[167]},
      {stage1_64[18]},
      {stage1_65[18]},
      {stage2_66[18],stage2_65[27],stage2_64[41],stage2_63[70],stage2_62[91]}
   );
   gpc1163_5 gpc5812 (
      {stage1_62[152], stage1_62[153], stage1_62[154]},
      {stage1_63[168], stage1_63[169], stage1_63[170], stage1_63[171], stage1_63[172], stage1_63[173]},
      {stage1_64[19]},
      {stage1_65[19]},
      {stage2_66[19],stage2_65[28],stage2_64[42],stage2_63[71],stage2_62[92]}
   );
   gpc1163_5 gpc5813 (
      {stage1_62[155], stage1_62[156], stage1_62[157]},
      {stage1_63[174], stage1_63[175], stage1_63[176], stage1_63[177], stage1_63[178], stage1_63[179]},
      {stage1_64[20]},
      {stage1_65[20]},
      {stage2_66[20],stage2_65[29],stage2_64[43],stage2_63[72],stage2_62[93]}
   );
   gpc1163_5 gpc5814 (
      {stage1_62[158], stage1_62[159], stage1_62[160]},
      {stage1_63[180], stage1_63[181], stage1_63[182], stage1_63[183], stage1_63[184], stage1_63[185]},
      {stage1_64[21]},
      {stage1_65[21]},
      {stage2_66[21],stage2_65[30],stage2_64[44],stage2_63[73],stage2_62[94]}
   );
   gpc1163_5 gpc5815 (
      {stage1_62[161], stage1_62[162], stage1_62[163]},
      {stage1_63[186], stage1_63[187], stage1_63[188], stage1_63[189], stage1_63[190], stage1_63[191]},
      {stage1_64[22]},
      {stage1_65[22]},
      {stage2_66[22],stage2_65[31],stage2_64[45],stage2_63[74],stage2_62[95]}
   );
   gpc1163_5 gpc5816 (
      {stage1_62[164], stage1_62[165], stage1_62[166]},
      {stage1_63[192], stage1_63[193], stage1_63[194], stage1_63[195], stage1_63[196], stage1_63[197]},
      {stage1_64[23]},
      {stage1_65[23]},
      {stage2_66[23],stage2_65[32],stage2_64[46],stage2_63[75],stage2_62[96]}
   );
   gpc1163_5 gpc5817 (
      {stage1_62[167], stage1_62[168], stage1_62[169]},
      {stage1_63[198], stage1_63[199], stage1_63[200], stage1_63[201], stage1_63[202], stage1_63[203]},
      {stage1_64[24]},
      {stage1_65[24]},
      {stage2_66[24],stage2_65[33],stage2_64[47],stage2_63[76],stage2_62[97]}
   );
   gpc1163_5 gpc5818 (
      {stage1_62[170], stage1_62[171], stage1_62[172]},
      {stage1_63[204], stage1_63[205], stage1_63[206], stage1_63[207], stage1_63[208], stage1_63[209]},
      {stage1_64[25]},
      {stage1_65[25]},
      {stage2_66[25],stage2_65[34],stage2_64[48],stage2_63[77],stage2_62[98]}
   );
   gpc1163_5 gpc5819 (
      {stage1_62[173], stage1_62[174], stage1_62[175]},
      {stage1_63[210], stage1_63[211], stage1_63[212], stage1_63[213], stage1_63[214], stage1_63[215]},
      {stage1_64[26]},
      {stage1_65[26]},
      {stage2_66[26],stage2_65[35],stage2_64[49],stage2_63[78],stage2_62[99]}
   );
   gpc1163_5 gpc5820 (
      {stage1_62[176], stage1_62[177], stage1_62[178]},
      {stage1_63[216], stage1_63[217], stage1_63[218], stage1_63[219], stage1_63[220], stage1_63[221]},
      {stage1_64[27]},
      {stage1_65[27]},
      {stage2_66[27],stage2_65[36],stage2_64[50],stage2_63[79],stage2_62[100]}
   );
   gpc1163_5 gpc5821 (
      {stage1_62[179], stage1_62[180], stage1_62[181]},
      {stage1_63[222], stage1_63[223], stage1_63[224], stage1_63[225], stage1_63[226], stage1_63[227]},
      {stage1_64[28]},
      {stage1_65[28]},
      {stage2_66[28],stage2_65[37],stage2_64[51],stage2_63[80],stage2_62[101]}
   );
   gpc615_5 gpc5822 (
      {stage1_62[182], stage1_62[183], stage1_62[184], stage1_62[185], stage1_62[186]},
      {stage1_63[228]},
      {stage1_64[29], stage1_64[30], stage1_64[31], stage1_64[32], stage1_64[33], stage1_64[34]},
      {stage2_66[29],stage2_65[38],stage2_64[52],stage2_63[81],stage2_62[102]}
   );
   gpc615_5 gpc5823 (
      {stage1_62[187], stage1_62[188], stage1_62[189], stage1_62[190], stage1_62[191]},
      {stage1_63[229]},
      {stage1_64[35], stage1_64[36], stage1_64[37], stage1_64[38], stage1_64[39], stage1_64[40]},
      {stage2_66[30],stage2_65[39],stage2_64[53],stage2_63[82],stage2_62[103]}
   );
   gpc135_4 gpc5824 (
      {stage1_63[230], stage1_63[231], stage1_63[232], stage1_63[233], stage1_63[234]},
      {stage1_64[41], stage1_64[42], stage1_64[43]},
      {stage1_65[29]},
      {stage2_66[31],stage2_65[40],stage2_64[54],stage2_63[83]}
   );
   gpc135_4 gpc5825 (
      {stage1_63[235], stage1_63[236], stage1_63[237], stage1_63[238], stage1_63[239]},
      {stage1_64[44], stage1_64[45], stage1_64[46]},
      {stage1_65[30]},
      {stage2_66[32],stage2_65[41],stage2_64[55],stage2_63[84]}
   );
   gpc207_4 gpc5826 (
      {stage1_63[240], stage1_63[241], stage1_63[242], stage1_63[243], stage1_63[244], stage1_63[245], stage1_63[246]},
      {stage1_65[31], stage1_65[32]},
      {stage2_66[33],stage2_65[42],stage2_64[56],stage2_63[85]}
   );
   gpc207_4 gpc5827 (
      {stage1_63[247], stage1_63[248], stage1_63[249], stage1_63[250], stage1_63[251], stage1_63[252], stage1_63[253]},
      {stage1_65[33], stage1_65[34]},
      {stage2_66[34],stage2_65[43],stage2_64[57],stage2_63[86]}
   );
   gpc207_4 gpc5828 (
      {stage1_63[254], stage1_63[255], stage1_63[256], stage1_63[257], stage1_63[258], stage1_63[259], stage1_63[260]},
      {stage1_65[35], stage1_65[36]},
      {stage2_66[35],stage2_65[44],stage2_64[58],stage2_63[87]}
   );
   gpc207_4 gpc5829 (
      {stage1_63[261], stage1_63[262], stage1_63[263], stage1_63[264], stage1_63[265], stage1_63[266], stage1_63[267]},
      {stage1_65[37], stage1_65[38]},
      {stage2_66[36],stage2_65[45],stage2_64[59],stage2_63[88]}
   );
   gpc207_4 gpc5830 (
      {stage1_63[268], stage1_63[269], stage1_63[270], stage1_63[271], stage1_63[272], stage1_63[273], stage1_63[274]},
      {stage1_65[39], stage1_65[40]},
      {stage2_66[37],stage2_65[46],stage2_64[60],stage2_63[89]}
   );
   gpc207_4 gpc5831 (
      {stage1_63[275], stage1_63[276], stage1_63[277], stage1_63[278], stage1_63[279], stage1_63[280], stage1_63[281]},
      {stage1_65[41], stage1_65[42]},
      {stage2_66[38],stage2_65[47],stage2_64[61],stage2_63[90]}
   );
   gpc207_4 gpc5832 (
      {stage1_63[282], stage1_63[283], stage1_63[284], stage1_63[285], stage1_63[286], stage1_63[287], stage1_63[288]},
      {stage1_65[43], stage1_65[44]},
      {stage2_66[39],stage2_65[48],stage2_64[62],stage2_63[91]}
   );
   gpc207_4 gpc5833 (
      {stage1_63[289], stage1_63[290], stage1_63[291], stage1_63[292], stage1_63[293], stage1_63[294], stage1_63[295]},
      {stage1_65[45], stage1_65[46]},
      {stage2_66[40],stage2_65[49],stage2_64[63],stage2_63[92]}
   );
   gpc207_4 gpc5834 (
      {stage1_63[296], stage1_63[297], stage1_63[298], stage1_63[299], stage1_63[300], stage1_63[301], stage1_63[302]},
      {stage1_65[47], stage1_65[48]},
      {stage2_66[41],stage2_65[50],stage2_64[64],stage2_63[93]}
   );
   gpc1_1 gpc5835 (
      {stage1_0[108]},
      {stage2_0[21]}
   );
   gpc1_1 gpc5836 (
      {stage1_0[109]},
      {stage2_0[22]}
   );
   gpc1_1 gpc5837 (
      {stage1_0[110]},
      {stage2_0[23]}
   );
   gpc1_1 gpc5838 (
      {stage1_0[111]},
      {stage2_0[24]}
   );
   gpc1_1 gpc5839 (
      {stage1_0[112]},
      {stage2_0[25]}
   );
   gpc1_1 gpc5840 (
      {stage1_0[113]},
      {stage2_0[26]}
   );
   gpc1_1 gpc5841 (
      {stage1_0[114]},
      {stage2_0[27]}
   );
   gpc1_1 gpc5842 (
      {stage1_0[115]},
      {stage2_0[28]}
   );
   gpc1_1 gpc5843 (
      {stage1_0[116]},
      {stage2_0[29]}
   );
   gpc1_1 gpc5844 (
      {stage1_0[117]},
      {stage2_0[30]}
   );
   gpc1_1 gpc5845 (
      {stage1_0[118]},
      {stage2_0[31]}
   );
   gpc1_1 gpc5846 (
      {stage1_0[119]},
      {stage2_0[32]}
   );
   gpc1_1 gpc5847 (
      {stage1_0[120]},
      {stage2_0[33]}
   );
   gpc1_1 gpc5848 (
      {stage1_0[121]},
      {stage2_0[34]}
   );
   gpc1_1 gpc5849 (
      {stage1_0[122]},
      {stage2_0[35]}
   );
   gpc1_1 gpc5850 (
      {stage1_0[123]},
      {stage2_0[36]}
   );
   gpc1_1 gpc5851 (
      {stage1_0[124]},
      {stage2_0[37]}
   );
   gpc1_1 gpc5852 (
      {stage1_1[168]},
      {stage2_1[46]}
   );
   gpc1_1 gpc5853 (
      {stage1_1[169]},
      {stage2_1[47]}
   );
   gpc1_1 gpc5854 (
      {stage1_1[170]},
      {stage2_1[48]}
   );
   gpc1_1 gpc5855 (
      {stage1_1[171]},
      {stage2_1[49]}
   );
   gpc1_1 gpc5856 (
      {stage1_1[172]},
      {stage2_1[50]}
   );
   gpc1_1 gpc5857 (
      {stage1_1[173]},
      {stage2_1[51]}
   );
   gpc1_1 gpc5858 (
      {stage1_1[174]},
      {stage2_1[52]}
   );
   gpc1_1 gpc5859 (
      {stage1_1[175]},
      {stage2_1[53]}
   );
   gpc1_1 gpc5860 (
      {stage1_2[144]},
      {stage2_2[49]}
   );
   gpc1_1 gpc5861 (
      {stage1_2[145]},
      {stage2_2[50]}
   );
   gpc1_1 gpc5862 (
      {stage1_2[146]},
      {stage2_2[51]}
   );
   gpc1_1 gpc5863 (
      {stage1_2[147]},
      {stage2_2[52]}
   );
   gpc1_1 gpc5864 (
      {stage1_2[148]},
      {stage2_2[53]}
   );
   gpc1_1 gpc5865 (
      {stage1_2[149]},
      {stage2_2[54]}
   );
   gpc1_1 gpc5866 (
      {stage1_2[150]},
      {stage2_2[55]}
   );
   gpc1_1 gpc5867 (
      {stage1_2[151]},
      {stage2_2[56]}
   );
   gpc1_1 gpc5868 (
      {stage1_2[152]},
      {stage2_2[57]}
   );
   gpc1_1 gpc5869 (
      {stage1_2[153]},
      {stage2_2[58]}
   );
   gpc1_1 gpc5870 (
      {stage1_2[154]},
      {stage2_2[59]}
   );
   gpc1_1 gpc5871 (
      {stage1_2[155]},
      {stage2_2[60]}
   );
   gpc1_1 gpc5872 (
      {stage1_2[156]},
      {stage2_2[61]}
   );
   gpc1_1 gpc5873 (
      {stage1_2[157]},
      {stage2_2[62]}
   );
   gpc1_1 gpc5874 (
      {stage1_3[150]},
      {stage2_3[49]}
   );
   gpc1_1 gpc5875 (
      {stage1_3[151]},
      {stage2_3[50]}
   );
   gpc1_1 gpc5876 (
      {stage1_3[152]},
      {stage2_3[51]}
   );
   gpc1_1 gpc5877 (
      {stage1_3[153]},
      {stage2_3[52]}
   );
   gpc1_1 gpc5878 (
      {stage1_3[154]},
      {stage2_3[53]}
   );
   gpc1_1 gpc5879 (
      {stage1_3[155]},
      {stage2_3[54]}
   );
   gpc1_1 gpc5880 (
      {stage1_3[156]},
      {stage2_3[55]}
   );
   gpc1_1 gpc5881 (
      {stage1_3[157]},
      {stage2_3[56]}
   );
   gpc1_1 gpc5882 (
      {stage1_3[158]},
      {stage2_3[57]}
   );
   gpc1_1 gpc5883 (
      {stage1_3[159]},
      {stage2_3[58]}
   );
   gpc1_1 gpc5884 (
      {stage1_3[160]},
      {stage2_3[59]}
   );
   gpc1_1 gpc5885 (
      {stage1_3[161]},
      {stage2_3[60]}
   );
   gpc1_1 gpc5886 (
      {stage1_3[162]},
      {stage2_3[61]}
   );
   gpc1_1 gpc5887 (
      {stage1_3[163]},
      {stage2_3[62]}
   );
   gpc1_1 gpc5888 (
      {stage1_3[164]},
      {stage2_3[63]}
   );
   gpc1_1 gpc5889 (
      {stage1_3[165]},
      {stage2_3[64]}
   );
   gpc1_1 gpc5890 (
      {stage1_3[166]},
      {stage2_3[65]}
   );
   gpc1_1 gpc5891 (
      {stage1_3[167]},
      {stage2_3[66]}
   );
   gpc1_1 gpc5892 (
      {stage1_3[168]},
      {stage2_3[67]}
   );
   gpc1_1 gpc5893 (
      {stage1_3[169]},
      {stage2_3[68]}
   );
   gpc1_1 gpc5894 (
      {stage1_3[170]},
      {stage2_3[69]}
   );
   gpc1_1 gpc5895 (
      {stage1_3[171]},
      {stage2_3[70]}
   );
   gpc1_1 gpc5896 (
      {stage1_3[172]},
      {stage2_3[71]}
   );
   gpc1_1 gpc5897 (
      {stage1_3[173]},
      {stage2_3[72]}
   );
   gpc1_1 gpc5898 (
      {stage1_3[174]},
      {stage2_3[73]}
   );
   gpc1_1 gpc5899 (
      {stage1_3[175]},
      {stage2_3[74]}
   );
   gpc1_1 gpc5900 (
      {stage1_3[176]},
      {stage2_3[75]}
   );
   gpc1_1 gpc5901 (
      {stage1_3[177]},
      {stage2_3[76]}
   );
   gpc1_1 gpc5902 (
      {stage1_3[178]},
      {stage2_3[77]}
   );
   gpc1_1 gpc5903 (
      {stage1_3[179]},
      {stage2_3[78]}
   );
   gpc1_1 gpc5904 (
      {stage1_3[180]},
      {stage2_3[79]}
   );
   gpc1_1 gpc5905 (
      {stage1_3[181]},
      {stage2_3[80]}
   );
   gpc1_1 gpc5906 (
      {stage1_3[182]},
      {stage2_3[81]}
   );
   gpc1_1 gpc5907 (
      {stage1_3[183]},
      {stage2_3[82]}
   );
   gpc1_1 gpc5908 (
      {stage1_3[184]},
      {stage2_3[83]}
   );
   gpc1_1 gpc5909 (
      {stage1_3[185]},
      {stage2_3[84]}
   );
   gpc1_1 gpc5910 (
      {stage1_3[186]},
      {stage2_3[85]}
   );
   gpc1_1 gpc5911 (
      {stage1_3[187]},
      {stage2_3[86]}
   );
   gpc1_1 gpc5912 (
      {stage1_3[188]},
      {stage2_3[87]}
   );
   gpc1_1 gpc5913 (
      {stage1_3[189]},
      {stage2_3[88]}
   );
   gpc1_1 gpc5914 (
      {stage1_3[190]},
      {stage2_3[89]}
   );
   gpc1_1 gpc5915 (
      {stage1_3[191]},
      {stage2_3[90]}
   );
   gpc1_1 gpc5916 (
      {stage1_3[192]},
      {stage2_3[91]}
   );
   gpc1_1 gpc5917 (
      {stage1_3[193]},
      {stage2_3[92]}
   );
   gpc1_1 gpc5918 (
      {stage1_3[194]},
      {stage2_3[93]}
   );
   gpc1_1 gpc5919 (
      {stage1_3[195]},
      {stage2_3[94]}
   );
   gpc1_1 gpc5920 (
      {stage1_3[196]},
      {stage2_3[95]}
   );
   gpc1_1 gpc5921 (
      {stage1_3[197]},
      {stage2_3[96]}
   );
   gpc1_1 gpc5922 (
      {stage1_3[198]},
      {stage2_3[97]}
   );
   gpc1_1 gpc5923 (
      {stage1_3[199]},
      {stage2_3[98]}
   );
   gpc1_1 gpc5924 (
      {stage1_3[200]},
      {stage2_3[99]}
   );
   gpc1_1 gpc5925 (
      {stage1_3[201]},
      {stage2_3[100]}
   );
   gpc1_1 gpc5926 (
      {stage1_3[202]},
      {stage2_3[101]}
   );
   gpc1_1 gpc5927 (
      {stage1_3[203]},
      {stage2_3[102]}
   );
   gpc1_1 gpc5928 (
      {stage1_3[204]},
      {stage2_3[103]}
   );
   gpc1_1 gpc5929 (
      {stage1_3[205]},
      {stage2_3[104]}
   );
   gpc1_1 gpc5930 (
      {stage1_3[206]},
      {stage2_3[105]}
   );
   gpc1_1 gpc5931 (
      {stage1_3[207]},
      {stage2_3[106]}
   );
   gpc1_1 gpc5932 (
      {stage1_3[208]},
      {stage2_3[107]}
   );
   gpc1_1 gpc5933 (
      {stage1_3[209]},
      {stage2_3[108]}
   );
   gpc1_1 gpc5934 (
      {stage1_3[210]},
      {stage2_3[109]}
   );
   gpc1_1 gpc5935 (
      {stage1_3[211]},
      {stage2_3[110]}
   );
   gpc1_1 gpc5936 (
      {stage1_3[212]},
      {stage2_3[111]}
   );
   gpc1_1 gpc5937 (
      {stage1_3[213]},
      {stage2_3[112]}
   );
   gpc1_1 gpc5938 (
      {stage1_3[214]},
      {stage2_3[113]}
   );
   gpc1_1 gpc5939 (
      {stage1_4[195]},
      {stage2_4[79]}
   );
   gpc1_1 gpc5940 (
      {stage1_4[196]},
      {stage2_4[80]}
   );
   gpc1_1 gpc5941 (
      {stage1_4[197]},
      {stage2_4[81]}
   );
   gpc1_1 gpc5942 (
      {stage1_4[198]},
      {stage2_4[82]}
   );
   gpc1_1 gpc5943 (
      {stage1_4[199]},
      {stage2_4[83]}
   );
   gpc1_1 gpc5944 (
      {stage1_4[200]},
      {stage2_4[84]}
   );
   gpc1_1 gpc5945 (
      {stage1_4[201]},
      {stage2_4[85]}
   );
   gpc1_1 gpc5946 (
      {stage1_4[202]},
      {stage2_4[86]}
   );
   gpc1_1 gpc5947 (
      {stage1_4[203]},
      {stage2_4[87]}
   );
   gpc1_1 gpc5948 (
      {stage1_4[204]},
      {stage2_4[88]}
   );
   gpc1_1 gpc5949 (
      {stage1_4[205]},
      {stage2_4[89]}
   );
   gpc1_1 gpc5950 (
      {stage1_4[206]},
      {stage2_4[90]}
   );
   gpc1_1 gpc5951 (
      {stage1_4[207]},
      {stage2_4[91]}
   );
   gpc1_1 gpc5952 (
      {stage1_4[208]},
      {stage2_4[92]}
   );
   gpc1_1 gpc5953 (
      {stage1_4[209]},
      {stage2_4[93]}
   );
   gpc1_1 gpc5954 (
      {stage1_4[210]},
      {stage2_4[94]}
   );
   gpc1_1 gpc5955 (
      {stage1_4[211]},
      {stage2_4[95]}
   );
   gpc1_1 gpc5956 (
      {stage1_4[212]},
      {stage2_4[96]}
   );
   gpc1_1 gpc5957 (
      {stage1_4[213]},
      {stage2_4[97]}
   );
   gpc1_1 gpc5958 (
      {stage1_4[214]},
      {stage2_4[98]}
   );
   gpc1_1 gpc5959 (
      {stage1_4[215]},
      {stage2_4[99]}
   );
   gpc1_1 gpc5960 (
      {stage1_4[216]},
      {stage2_4[100]}
   );
   gpc1_1 gpc5961 (
      {stage1_4[217]},
      {stage2_4[101]}
   );
   gpc1_1 gpc5962 (
      {stage1_4[218]},
      {stage2_4[102]}
   );
   gpc1_1 gpc5963 (
      {stage1_4[219]},
      {stage2_4[103]}
   );
   gpc1_1 gpc5964 (
      {stage1_4[220]},
      {stage2_4[104]}
   );
   gpc1_1 gpc5965 (
      {stage1_4[221]},
      {stage2_4[105]}
   );
   gpc1_1 gpc5966 (
      {stage1_4[222]},
      {stage2_4[106]}
   );
   gpc1_1 gpc5967 (
      {stage1_4[223]},
      {stage2_4[107]}
   );
   gpc1_1 gpc5968 (
      {stage1_4[224]},
      {stage2_4[108]}
   );
   gpc1_1 gpc5969 (
      {stage1_4[225]},
      {stage2_4[109]}
   );
   gpc1_1 gpc5970 (
      {stage1_4[226]},
      {stage2_4[110]}
   );
   gpc1_1 gpc5971 (
      {stage1_4[227]},
      {stage2_4[111]}
   );
   gpc1_1 gpc5972 (
      {stage1_5[124]},
      {stage2_5[78]}
   );
   gpc1_1 gpc5973 (
      {stage1_5[125]},
      {stage2_5[79]}
   );
   gpc1_1 gpc5974 (
      {stage1_5[126]},
      {stage2_5[80]}
   );
   gpc1_1 gpc5975 (
      {stage1_5[127]},
      {stage2_5[81]}
   );
   gpc1_1 gpc5976 (
      {stage1_5[128]},
      {stage2_5[82]}
   );
   gpc1_1 gpc5977 (
      {stage1_5[129]},
      {stage2_5[83]}
   );
   gpc1_1 gpc5978 (
      {stage1_5[130]},
      {stage2_5[84]}
   );
   gpc1_1 gpc5979 (
      {stage1_5[131]},
      {stage2_5[85]}
   );
   gpc1_1 gpc5980 (
      {stage1_5[132]},
      {stage2_5[86]}
   );
   gpc1_1 gpc5981 (
      {stage1_5[133]},
      {stage2_5[87]}
   );
   gpc1_1 gpc5982 (
      {stage1_5[134]},
      {stage2_5[88]}
   );
   gpc1_1 gpc5983 (
      {stage1_5[135]},
      {stage2_5[89]}
   );
   gpc1_1 gpc5984 (
      {stage1_5[136]},
      {stage2_5[90]}
   );
   gpc1_1 gpc5985 (
      {stage1_5[137]},
      {stage2_5[91]}
   );
   gpc1_1 gpc5986 (
      {stage1_5[138]},
      {stage2_5[92]}
   );
   gpc1_1 gpc5987 (
      {stage1_5[139]},
      {stage2_5[93]}
   );
   gpc1_1 gpc5988 (
      {stage1_5[140]},
      {stage2_5[94]}
   );
   gpc1_1 gpc5989 (
      {stage1_5[141]},
      {stage2_5[95]}
   );
   gpc1_1 gpc5990 (
      {stage1_5[142]},
      {stage2_5[96]}
   );
   gpc1_1 gpc5991 (
      {stage1_5[143]},
      {stage2_5[97]}
   );
   gpc1_1 gpc5992 (
      {stage1_5[144]},
      {stage2_5[98]}
   );
   gpc1_1 gpc5993 (
      {stage1_5[145]},
      {stage2_5[99]}
   );
   gpc1_1 gpc5994 (
      {stage1_5[146]},
      {stage2_5[100]}
   );
   gpc1_1 gpc5995 (
      {stage1_5[147]},
      {stage2_5[101]}
   );
   gpc1_1 gpc5996 (
      {stage1_5[148]},
      {stage2_5[102]}
   );
   gpc1_1 gpc5997 (
      {stage1_5[149]},
      {stage2_5[103]}
   );
   gpc1_1 gpc5998 (
      {stage1_5[150]},
      {stage2_5[104]}
   );
   gpc1_1 gpc5999 (
      {stage1_5[151]},
      {stage2_5[105]}
   );
   gpc1_1 gpc6000 (
      {stage1_5[152]},
      {stage2_5[106]}
   );
   gpc1_1 gpc6001 (
      {stage1_5[153]},
      {stage2_5[107]}
   );
   gpc1_1 gpc6002 (
      {stage1_5[154]},
      {stage2_5[108]}
   );
   gpc1_1 gpc6003 (
      {stage1_5[155]},
      {stage2_5[109]}
   );
   gpc1_1 gpc6004 (
      {stage1_5[156]},
      {stage2_5[110]}
   );
   gpc1_1 gpc6005 (
      {stage1_5[157]},
      {stage2_5[111]}
   );
   gpc1_1 gpc6006 (
      {stage1_5[158]},
      {stage2_5[112]}
   );
   gpc1_1 gpc6007 (
      {stage1_5[159]},
      {stage2_5[113]}
   );
   gpc1_1 gpc6008 (
      {stage1_5[160]},
      {stage2_5[114]}
   );
   gpc1_1 gpc6009 (
      {stage1_5[161]},
      {stage2_5[115]}
   );
   gpc1_1 gpc6010 (
      {stage1_5[162]},
      {stage2_5[116]}
   );
   gpc1_1 gpc6011 (
      {stage1_5[163]},
      {stage2_5[117]}
   );
   gpc1_1 gpc6012 (
      {stage1_5[164]},
      {stage2_5[118]}
   );
   gpc1_1 gpc6013 (
      {stage1_5[165]},
      {stage2_5[119]}
   );
   gpc1_1 gpc6014 (
      {stage1_5[166]},
      {stage2_5[120]}
   );
   gpc1_1 gpc6015 (
      {stage1_5[167]},
      {stage2_5[121]}
   );
   gpc1_1 gpc6016 (
      {stage1_5[168]},
      {stage2_5[122]}
   );
   gpc1_1 gpc6017 (
      {stage1_5[169]},
      {stage2_5[123]}
   );
   gpc1_1 gpc6018 (
      {stage1_5[170]},
      {stage2_5[124]}
   );
   gpc1_1 gpc6019 (
      {stage1_5[171]},
      {stage2_5[125]}
   );
   gpc1_1 gpc6020 (
      {stage1_5[172]},
      {stage2_5[126]}
   );
   gpc1_1 gpc6021 (
      {stage1_5[173]},
      {stage2_5[127]}
   );
   gpc1_1 gpc6022 (
      {stage1_5[174]},
      {stage2_5[128]}
   );
   gpc1_1 gpc6023 (
      {stage1_5[175]},
      {stage2_5[129]}
   );
   gpc1_1 gpc6024 (
      {stage1_5[176]},
      {stage2_5[130]}
   );
   gpc1_1 gpc6025 (
      {stage1_5[177]},
      {stage2_5[131]}
   );
   gpc1_1 gpc6026 (
      {stage1_5[178]},
      {stage2_5[132]}
   );
   gpc1_1 gpc6027 (
      {stage1_5[179]},
      {stage2_5[133]}
   );
   gpc1_1 gpc6028 (
      {stage1_5[180]},
      {stage2_5[134]}
   );
   gpc1_1 gpc6029 (
      {stage1_5[181]},
      {stage2_5[135]}
   );
   gpc1_1 gpc6030 (
      {stage1_5[182]},
      {stage2_5[136]}
   );
   gpc1_1 gpc6031 (
      {stage1_5[183]},
      {stage2_5[137]}
   );
   gpc1_1 gpc6032 (
      {stage1_5[184]},
      {stage2_5[138]}
   );
   gpc1_1 gpc6033 (
      {stage1_5[185]},
      {stage2_5[139]}
   );
   gpc1_1 gpc6034 (
      {stage1_5[186]},
      {stage2_5[140]}
   );
   gpc1_1 gpc6035 (
      {stage1_5[187]},
      {stage2_5[141]}
   );
   gpc1_1 gpc6036 (
      {stage1_5[188]},
      {stage2_5[142]}
   );
   gpc1_1 gpc6037 (
      {stage1_5[189]},
      {stage2_5[143]}
   );
   gpc1_1 gpc6038 (
      {stage1_5[190]},
      {stage2_5[144]}
   );
   gpc1_1 gpc6039 (
      {stage1_5[191]},
      {stage2_5[145]}
   );
   gpc1_1 gpc6040 (
      {stage1_5[192]},
      {stage2_5[146]}
   );
   gpc1_1 gpc6041 (
      {stage1_5[193]},
      {stage2_5[147]}
   );
   gpc1_1 gpc6042 (
      {stage1_5[194]},
      {stage2_5[148]}
   );
   gpc1_1 gpc6043 (
      {stage1_5[195]},
      {stage2_5[149]}
   );
   gpc1_1 gpc6044 (
      {stage1_5[196]},
      {stage2_5[150]}
   );
   gpc1_1 gpc6045 (
      {stage1_5[197]},
      {stage2_5[151]}
   );
   gpc1_1 gpc6046 (
      {stage1_6[175]},
      {stage2_6[53]}
   );
   gpc1_1 gpc6047 (
      {stage1_6[176]},
      {stage2_6[54]}
   );
   gpc1_1 gpc6048 (
      {stage1_6[177]},
      {stage2_6[55]}
   );
   gpc1_1 gpc6049 (
      {stage1_6[178]},
      {stage2_6[56]}
   );
   gpc1_1 gpc6050 (
      {stage1_6[179]},
      {stage2_6[57]}
   );
   gpc1_1 gpc6051 (
      {stage1_6[180]},
      {stage2_6[58]}
   );
   gpc1_1 gpc6052 (
      {stage1_6[181]},
      {stage2_6[59]}
   );
   gpc1_1 gpc6053 (
      {stage1_6[182]},
      {stage2_6[60]}
   );
   gpc1_1 gpc6054 (
      {stage1_6[183]},
      {stage2_6[61]}
   );
   gpc1_1 gpc6055 (
      {stage1_6[184]},
      {stage2_6[62]}
   );
   gpc1_1 gpc6056 (
      {stage1_6[185]},
      {stage2_6[63]}
   );
   gpc1_1 gpc6057 (
      {stage1_6[186]},
      {stage2_6[64]}
   );
   gpc1_1 gpc6058 (
      {stage1_6[187]},
      {stage2_6[65]}
   );
   gpc1_1 gpc6059 (
      {stage1_6[188]},
      {stage2_6[66]}
   );
   gpc1_1 gpc6060 (
      {stage1_6[189]},
      {stage2_6[67]}
   );
   gpc1_1 gpc6061 (
      {stage1_6[190]},
      {stage2_6[68]}
   );
   gpc1_1 gpc6062 (
      {stage1_6[191]},
      {stage2_6[69]}
   );
   gpc1_1 gpc6063 (
      {stage1_6[192]},
      {stage2_6[70]}
   );
   gpc1_1 gpc6064 (
      {stage1_6[193]},
      {stage2_6[71]}
   );
   gpc1_1 gpc6065 (
      {stage1_6[194]},
      {stage2_6[72]}
   );
   gpc1_1 gpc6066 (
      {stage1_6[195]},
      {stage2_6[73]}
   );
   gpc1_1 gpc6067 (
      {stage1_6[196]},
      {stage2_6[74]}
   );
   gpc1_1 gpc6068 (
      {stage1_6[197]},
      {stage2_6[75]}
   );
   gpc1_1 gpc6069 (
      {stage1_6[198]},
      {stage2_6[76]}
   );
   gpc1_1 gpc6070 (
      {stage1_6[199]},
      {stage2_6[77]}
   );
   gpc1_1 gpc6071 (
      {stage1_6[200]},
      {stage2_6[78]}
   );
   gpc1_1 gpc6072 (
      {stage1_6[201]},
      {stage2_6[79]}
   );
   gpc1_1 gpc6073 (
      {stage1_6[202]},
      {stage2_6[80]}
   );
   gpc1_1 gpc6074 (
      {stage1_6[203]},
      {stage2_6[81]}
   );
   gpc1_1 gpc6075 (
      {stage1_6[204]},
      {stage2_6[82]}
   );
   gpc1_1 gpc6076 (
      {stage1_6[205]},
      {stage2_6[83]}
   );
   gpc1_1 gpc6077 (
      {stage1_6[206]},
      {stage2_6[84]}
   );
   gpc1_1 gpc6078 (
      {stage1_6[207]},
      {stage2_6[85]}
   );
   gpc1_1 gpc6079 (
      {stage1_6[208]},
      {stage2_6[86]}
   );
   gpc1_1 gpc6080 (
      {stage1_6[209]},
      {stage2_6[87]}
   );
   gpc1_1 gpc6081 (
      {stage1_6[210]},
      {stage2_6[88]}
   );
   gpc1_1 gpc6082 (
      {stage1_6[211]},
      {stage2_6[89]}
   );
   gpc1_1 gpc6083 (
      {stage1_6[212]},
      {stage2_6[90]}
   );
   gpc1_1 gpc6084 (
      {stage1_6[213]},
      {stage2_6[91]}
   );
   gpc1_1 gpc6085 (
      {stage1_7[217]},
      {stage2_7[69]}
   );
   gpc1_1 gpc6086 (
      {stage1_7[218]},
      {stage2_7[70]}
   );
   gpc1_1 gpc6087 (
      {stage1_7[219]},
      {stage2_7[71]}
   );
   gpc1_1 gpc6088 (
      {stage1_7[220]},
      {stage2_7[72]}
   );
   gpc1_1 gpc6089 (
      {stage1_8[134]},
      {stage2_8[88]}
   );
   gpc1_1 gpc6090 (
      {stage1_8[135]},
      {stage2_8[89]}
   );
   gpc1_1 gpc6091 (
      {stage1_8[136]},
      {stage2_8[90]}
   );
   gpc1_1 gpc6092 (
      {stage1_8[137]},
      {stage2_8[91]}
   );
   gpc1_1 gpc6093 (
      {stage1_8[138]},
      {stage2_8[92]}
   );
   gpc1_1 gpc6094 (
      {stage1_8[139]},
      {stage2_8[93]}
   );
   gpc1_1 gpc6095 (
      {stage1_8[140]},
      {stage2_8[94]}
   );
   gpc1_1 gpc6096 (
      {stage1_8[141]},
      {stage2_8[95]}
   );
   gpc1_1 gpc6097 (
      {stage1_8[142]},
      {stage2_8[96]}
   );
   gpc1_1 gpc6098 (
      {stage1_8[143]},
      {stage2_8[97]}
   );
   gpc1_1 gpc6099 (
      {stage1_8[144]},
      {stage2_8[98]}
   );
   gpc1_1 gpc6100 (
      {stage1_8[145]},
      {stage2_8[99]}
   );
   gpc1_1 gpc6101 (
      {stage1_8[146]},
      {stage2_8[100]}
   );
   gpc1_1 gpc6102 (
      {stage1_8[147]},
      {stage2_8[101]}
   );
   gpc1_1 gpc6103 (
      {stage1_8[148]},
      {stage2_8[102]}
   );
   gpc1_1 gpc6104 (
      {stage1_8[149]},
      {stage2_8[103]}
   );
   gpc1_1 gpc6105 (
      {stage1_8[150]},
      {stage2_8[104]}
   );
   gpc1_1 gpc6106 (
      {stage1_8[151]},
      {stage2_8[105]}
   );
   gpc1_1 gpc6107 (
      {stage1_8[152]},
      {stage2_8[106]}
   );
   gpc1_1 gpc6108 (
      {stage1_8[153]},
      {stage2_8[107]}
   );
   gpc1_1 gpc6109 (
      {stage1_8[154]},
      {stage2_8[108]}
   );
   gpc1_1 gpc6110 (
      {stage1_8[155]},
      {stage2_8[109]}
   );
   gpc1_1 gpc6111 (
      {stage1_8[156]},
      {stage2_8[110]}
   );
   gpc1_1 gpc6112 (
      {stage1_8[157]},
      {stage2_8[111]}
   );
   gpc1_1 gpc6113 (
      {stage1_8[158]},
      {stage2_8[112]}
   );
   gpc1_1 gpc6114 (
      {stage1_8[159]},
      {stage2_8[113]}
   );
   gpc1_1 gpc6115 (
      {stage1_8[160]},
      {stage2_8[114]}
   );
   gpc1_1 gpc6116 (
      {stage1_8[161]},
      {stage2_8[115]}
   );
   gpc1_1 gpc6117 (
      {stage1_8[162]},
      {stage2_8[116]}
   );
   gpc1_1 gpc6118 (
      {stage1_8[163]},
      {stage2_8[117]}
   );
   gpc1_1 gpc6119 (
      {stage1_8[164]},
      {stage2_8[118]}
   );
   gpc1_1 gpc6120 (
      {stage1_8[165]},
      {stage2_8[119]}
   );
   gpc1_1 gpc6121 (
      {stage1_8[166]},
      {stage2_8[120]}
   );
   gpc1_1 gpc6122 (
      {stage1_8[167]},
      {stage2_8[121]}
   );
   gpc1_1 gpc6123 (
      {stage1_8[168]},
      {stage2_8[122]}
   );
   gpc1_1 gpc6124 (
      {stage1_8[169]},
      {stage2_8[123]}
   );
   gpc1_1 gpc6125 (
      {stage1_8[170]},
      {stage2_8[124]}
   );
   gpc1_1 gpc6126 (
      {stage1_8[171]},
      {stage2_8[125]}
   );
   gpc1_1 gpc6127 (
      {stage1_8[172]},
      {stage2_8[126]}
   );
   gpc1_1 gpc6128 (
      {stage1_8[173]},
      {stage2_8[127]}
   );
   gpc1_1 gpc6129 (
      {stage1_8[174]},
      {stage2_8[128]}
   );
   gpc1_1 gpc6130 (
      {stage1_8[175]},
      {stage2_8[129]}
   );
   gpc1_1 gpc6131 (
      {stage1_8[176]},
      {stage2_8[130]}
   );
   gpc1_1 gpc6132 (
      {stage1_8[177]},
      {stage2_8[131]}
   );
   gpc1_1 gpc6133 (
      {stage1_8[178]},
      {stage2_8[132]}
   );
   gpc1_1 gpc6134 (
      {stage1_8[179]},
      {stage2_8[133]}
   );
   gpc1_1 gpc6135 (
      {stage1_8[180]},
      {stage2_8[134]}
   );
   gpc1_1 gpc6136 (
      {stage1_8[181]},
      {stage2_8[135]}
   );
   gpc1_1 gpc6137 (
      {stage1_8[182]},
      {stage2_8[136]}
   );
   gpc1_1 gpc6138 (
      {stage1_8[183]},
      {stage2_8[137]}
   );
   gpc1_1 gpc6139 (
      {stage1_8[184]},
      {stage2_8[138]}
   );
   gpc1_1 gpc6140 (
      {stage1_8[185]},
      {stage2_8[139]}
   );
   gpc1_1 gpc6141 (
      {stage1_8[186]},
      {stage2_8[140]}
   );
   gpc1_1 gpc6142 (
      {stage1_8[187]},
      {stage2_8[141]}
   );
   gpc1_1 gpc6143 (
      {stage1_8[188]},
      {stage2_8[142]}
   );
   gpc1_1 gpc6144 (
      {stage1_8[189]},
      {stage2_8[143]}
   );
   gpc1_1 gpc6145 (
      {stage1_8[190]},
      {stage2_8[144]}
   );
   gpc1_1 gpc6146 (
      {stage1_8[191]},
      {stage2_8[145]}
   );
   gpc1_1 gpc6147 (
      {stage1_8[192]},
      {stage2_8[146]}
   );
   gpc1_1 gpc6148 (
      {stage1_8[193]},
      {stage2_8[147]}
   );
   gpc1_1 gpc6149 (
      {stage1_8[194]},
      {stage2_8[148]}
   );
   gpc1_1 gpc6150 (
      {stage1_8[195]},
      {stage2_8[149]}
   );
   gpc1_1 gpc6151 (
      {stage1_8[196]},
      {stage2_8[150]}
   );
   gpc1_1 gpc6152 (
      {stage1_8[197]},
      {stage2_8[151]}
   );
   gpc1_1 gpc6153 (
      {stage1_8[198]},
      {stage2_8[152]}
   );
   gpc1_1 gpc6154 (
      {stage1_8[199]},
      {stage2_8[153]}
   );
   gpc1_1 gpc6155 (
      {stage1_8[200]},
      {stage2_8[154]}
   );
   gpc1_1 gpc6156 (
      {stage1_8[201]},
      {stage2_8[155]}
   );
   gpc1_1 gpc6157 (
      {stage1_8[202]},
      {stage2_8[156]}
   );
   gpc1_1 gpc6158 (
      {stage1_8[203]},
      {stage2_8[157]}
   );
   gpc1_1 gpc6159 (
      {stage1_8[204]},
      {stage2_8[158]}
   );
   gpc1_1 gpc6160 (
      {stage1_8[205]},
      {stage2_8[159]}
   );
   gpc1_1 gpc6161 (
      {stage1_9[132]},
      {stage2_9[61]}
   );
   gpc1_1 gpc6162 (
      {stage1_9[133]},
      {stage2_9[62]}
   );
   gpc1_1 gpc6163 (
      {stage1_9[134]},
      {stage2_9[63]}
   );
   gpc1_1 gpc6164 (
      {stage1_9[135]},
      {stage2_9[64]}
   );
   gpc1_1 gpc6165 (
      {stage1_9[136]},
      {stage2_9[65]}
   );
   gpc1_1 gpc6166 (
      {stage1_9[137]},
      {stage2_9[66]}
   );
   gpc1_1 gpc6167 (
      {stage1_9[138]},
      {stage2_9[67]}
   );
   gpc1_1 gpc6168 (
      {stage1_9[139]},
      {stage2_9[68]}
   );
   gpc1_1 gpc6169 (
      {stage1_9[140]},
      {stage2_9[69]}
   );
   gpc1_1 gpc6170 (
      {stage1_9[141]},
      {stage2_9[70]}
   );
   gpc1_1 gpc6171 (
      {stage1_9[142]},
      {stage2_9[71]}
   );
   gpc1_1 gpc6172 (
      {stage1_9[143]},
      {stage2_9[72]}
   );
   gpc1_1 gpc6173 (
      {stage1_9[144]},
      {stage2_9[73]}
   );
   gpc1_1 gpc6174 (
      {stage1_9[145]},
      {stage2_9[74]}
   );
   gpc1_1 gpc6175 (
      {stage1_9[146]},
      {stage2_9[75]}
   );
   gpc1_1 gpc6176 (
      {stage1_9[147]},
      {stage2_9[76]}
   );
   gpc1_1 gpc6177 (
      {stage1_9[148]},
      {stage2_9[77]}
   );
   gpc1_1 gpc6178 (
      {stage1_9[149]},
      {stage2_9[78]}
   );
   gpc1_1 gpc6179 (
      {stage1_9[150]},
      {stage2_9[79]}
   );
   gpc1_1 gpc6180 (
      {stage1_9[151]},
      {stage2_9[80]}
   );
   gpc1_1 gpc6181 (
      {stage1_9[152]},
      {stage2_9[81]}
   );
   gpc1_1 gpc6182 (
      {stage1_9[153]},
      {stage2_9[82]}
   );
   gpc1_1 gpc6183 (
      {stage1_9[154]},
      {stage2_9[83]}
   );
   gpc1_1 gpc6184 (
      {stage1_9[155]},
      {stage2_9[84]}
   );
   gpc1_1 gpc6185 (
      {stage1_9[156]},
      {stage2_9[85]}
   );
   gpc1_1 gpc6186 (
      {stage1_9[157]},
      {stage2_9[86]}
   );
   gpc1_1 gpc6187 (
      {stage1_9[158]},
      {stage2_9[87]}
   );
   gpc1_1 gpc6188 (
      {stage1_9[159]},
      {stage2_9[88]}
   );
   gpc1_1 gpc6189 (
      {stage1_9[160]},
      {stage2_9[89]}
   );
   gpc1_1 gpc6190 (
      {stage1_9[161]},
      {stage2_9[90]}
   );
   gpc1_1 gpc6191 (
      {stage1_9[162]},
      {stage2_9[91]}
   );
   gpc1_1 gpc6192 (
      {stage1_9[163]},
      {stage2_9[92]}
   );
   gpc1_1 gpc6193 (
      {stage1_9[164]},
      {stage2_9[93]}
   );
   gpc1_1 gpc6194 (
      {stage1_9[165]},
      {stage2_9[94]}
   );
   gpc1_1 gpc6195 (
      {stage1_9[166]},
      {stage2_9[95]}
   );
   gpc1_1 gpc6196 (
      {stage1_9[167]},
      {stage2_9[96]}
   );
   gpc1_1 gpc6197 (
      {stage1_9[168]},
      {stage2_9[97]}
   );
   gpc1_1 gpc6198 (
      {stage1_9[169]},
      {stage2_9[98]}
   );
   gpc1_1 gpc6199 (
      {stage1_9[170]},
      {stage2_9[99]}
   );
   gpc1_1 gpc6200 (
      {stage1_9[171]},
      {stage2_9[100]}
   );
   gpc1_1 gpc6201 (
      {stage1_9[172]},
      {stage2_9[101]}
   );
   gpc1_1 gpc6202 (
      {stage1_9[173]},
      {stage2_9[102]}
   );
   gpc1_1 gpc6203 (
      {stage1_9[174]},
      {stage2_9[103]}
   );
   gpc1_1 gpc6204 (
      {stage1_9[175]},
      {stage2_9[104]}
   );
   gpc1_1 gpc6205 (
      {stage1_9[176]},
      {stage2_9[105]}
   );
   gpc1_1 gpc6206 (
      {stage1_9[177]},
      {stage2_9[106]}
   );
   gpc1_1 gpc6207 (
      {stage1_9[178]},
      {stage2_9[107]}
   );
   gpc1_1 gpc6208 (
      {stage1_9[179]},
      {stage2_9[108]}
   );
   gpc1_1 gpc6209 (
      {stage1_9[180]},
      {stage2_9[109]}
   );
   gpc1_1 gpc6210 (
      {stage1_9[181]},
      {stage2_9[110]}
   );
   gpc1_1 gpc6211 (
      {stage1_9[182]},
      {stage2_9[111]}
   );
   gpc1_1 gpc6212 (
      {stage1_9[183]},
      {stage2_9[112]}
   );
   gpc1_1 gpc6213 (
      {stage1_9[184]},
      {stage2_9[113]}
   );
   gpc1_1 gpc6214 (
      {stage1_9[185]},
      {stage2_9[114]}
   );
   gpc1_1 gpc6215 (
      {stage1_9[186]},
      {stage2_9[115]}
   );
   gpc1_1 gpc6216 (
      {stage1_9[187]},
      {stage2_9[116]}
   );
   gpc1_1 gpc6217 (
      {stage1_9[188]},
      {stage2_9[117]}
   );
   gpc1_1 gpc6218 (
      {stage1_9[189]},
      {stage2_9[118]}
   );
   gpc1_1 gpc6219 (
      {stage1_9[190]},
      {stage2_9[119]}
   );
   gpc1_1 gpc6220 (
      {stage1_9[191]},
      {stage2_9[120]}
   );
   gpc1_1 gpc6221 (
      {stage1_9[192]},
      {stage2_9[121]}
   );
   gpc1_1 gpc6222 (
      {stage1_9[193]},
      {stage2_9[122]}
   );
   gpc1_1 gpc6223 (
      {stage1_9[194]},
      {stage2_9[123]}
   );
   gpc1_1 gpc6224 (
      {stage1_9[195]},
      {stage2_9[124]}
   );
   gpc1_1 gpc6225 (
      {stage1_9[196]},
      {stage2_9[125]}
   );
   gpc1_1 gpc6226 (
      {stage1_9[197]},
      {stage2_9[126]}
   );
   gpc1_1 gpc6227 (
      {stage1_9[198]},
      {stage2_9[127]}
   );
   gpc1_1 gpc6228 (
      {stage1_9[199]},
      {stage2_9[128]}
   );
   gpc1_1 gpc6229 (
      {stage1_9[200]},
      {stage2_9[129]}
   );
   gpc1_1 gpc6230 (
      {stage1_9[201]},
      {stage2_9[130]}
   );
   gpc1_1 gpc6231 (
      {stage1_9[202]},
      {stage2_9[131]}
   );
   gpc1_1 gpc6232 (
      {stage1_9[203]},
      {stage2_9[132]}
   );
   gpc1_1 gpc6233 (
      {stage1_9[204]},
      {stage2_9[133]}
   );
   gpc1_1 gpc6234 (
      {stage1_9[205]},
      {stage2_9[134]}
   );
   gpc1_1 gpc6235 (
      {stage1_9[206]},
      {stage2_9[135]}
   );
   gpc1_1 gpc6236 (
      {stage1_9[207]},
      {stage2_9[136]}
   );
   gpc1_1 gpc6237 (
      {stage1_9[208]},
      {stage2_9[137]}
   );
   gpc1_1 gpc6238 (
      {stage1_9[209]},
      {stage2_9[138]}
   );
   gpc1_1 gpc6239 (
      {stage1_9[210]},
      {stage2_9[139]}
   );
   gpc1_1 gpc6240 (
      {stage1_9[211]},
      {stage2_9[140]}
   );
   gpc1_1 gpc6241 (
      {stage1_9[212]},
      {stage2_9[141]}
   );
   gpc1_1 gpc6242 (
      {stage1_9[213]},
      {stage2_9[142]}
   );
   gpc1_1 gpc6243 (
      {stage1_10[175]},
      {stage2_10[54]}
   );
   gpc1_1 gpc6244 (
      {stage1_10[176]},
      {stage2_10[55]}
   );
   gpc1_1 gpc6245 (
      {stage1_10[177]},
      {stage2_10[56]}
   );
   gpc1_1 gpc6246 (
      {stage1_10[178]},
      {stage2_10[57]}
   );
   gpc1_1 gpc6247 (
      {stage1_10[179]},
      {stage2_10[58]}
   );
   gpc1_1 gpc6248 (
      {stage1_10[180]},
      {stage2_10[59]}
   );
   gpc1_1 gpc6249 (
      {stage1_10[181]},
      {stage2_10[60]}
   );
   gpc1_1 gpc6250 (
      {stage1_10[182]},
      {stage2_10[61]}
   );
   gpc1_1 gpc6251 (
      {stage1_10[183]},
      {stage2_10[62]}
   );
   gpc1_1 gpc6252 (
      {stage1_10[184]},
      {stage2_10[63]}
   );
   gpc1_1 gpc6253 (
      {stage1_10[185]},
      {stage2_10[64]}
   );
   gpc1_1 gpc6254 (
      {stage1_10[186]},
      {stage2_10[65]}
   );
   gpc1_1 gpc6255 (
      {stage1_10[187]},
      {stage2_10[66]}
   );
   gpc1_1 gpc6256 (
      {stage1_10[188]},
      {stage2_10[67]}
   );
   gpc1_1 gpc6257 (
      {stage1_10[189]},
      {stage2_10[68]}
   );
   gpc1_1 gpc6258 (
      {stage1_10[190]},
      {stage2_10[69]}
   );
   gpc1_1 gpc6259 (
      {stage1_10[191]},
      {stage2_10[70]}
   );
   gpc1_1 gpc6260 (
      {stage1_10[192]},
      {stage2_10[71]}
   );
   gpc1_1 gpc6261 (
      {stage1_10[193]},
      {stage2_10[72]}
   );
   gpc1_1 gpc6262 (
      {stage1_10[194]},
      {stage2_10[73]}
   );
   gpc1_1 gpc6263 (
      {stage1_10[195]},
      {stage2_10[74]}
   );
   gpc1_1 gpc6264 (
      {stage1_10[196]},
      {stage2_10[75]}
   );
   gpc1_1 gpc6265 (
      {stage1_10[197]},
      {stage2_10[76]}
   );
   gpc1_1 gpc6266 (
      {stage1_10[198]},
      {stage2_10[77]}
   );
   gpc1_1 gpc6267 (
      {stage1_10[199]},
      {stage2_10[78]}
   );
   gpc1_1 gpc6268 (
      {stage1_10[200]},
      {stage2_10[79]}
   );
   gpc1_1 gpc6269 (
      {stage1_10[201]},
      {stage2_10[80]}
   );
   gpc1_1 gpc6270 (
      {stage1_10[202]},
      {stage2_10[81]}
   );
   gpc1_1 gpc6271 (
      {stage1_10[203]},
      {stage2_10[82]}
   );
   gpc1_1 gpc6272 (
      {stage1_10[204]},
      {stage2_10[83]}
   );
   gpc1_1 gpc6273 (
      {stage1_10[205]},
      {stage2_10[84]}
   );
   gpc1_1 gpc6274 (
      {stage1_10[206]},
      {stage2_10[85]}
   );
   gpc1_1 gpc6275 (
      {stage1_10[207]},
      {stage2_10[86]}
   );
   gpc1_1 gpc6276 (
      {stage1_10[208]},
      {stage2_10[87]}
   );
   gpc1_1 gpc6277 (
      {stage1_10[209]},
      {stage2_10[88]}
   );
   gpc1_1 gpc6278 (
      {stage1_10[210]},
      {stage2_10[89]}
   );
   gpc1_1 gpc6279 (
      {stage1_10[211]},
      {stage2_10[90]}
   );
   gpc1_1 gpc6280 (
      {stage1_10[212]},
      {stage2_10[91]}
   );
   gpc1_1 gpc6281 (
      {stage1_10[213]},
      {stage2_10[92]}
   );
   gpc1_1 gpc6282 (
      {stage1_10[214]},
      {stage2_10[93]}
   );
   gpc1_1 gpc6283 (
      {stage1_10[215]},
      {stage2_10[94]}
   );
   gpc1_1 gpc6284 (
      {stage1_10[216]},
      {stage2_10[95]}
   );
   gpc1_1 gpc6285 (
      {stage1_10[217]},
      {stage2_10[96]}
   );
   gpc1_1 gpc6286 (
      {stage1_10[218]},
      {stage2_10[97]}
   );
   gpc1_1 gpc6287 (
      {stage1_10[219]},
      {stage2_10[98]}
   );
   gpc1_1 gpc6288 (
      {stage1_10[220]},
      {stage2_10[99]}
   );
   gpc1_1 gpc6289 (
      {stage1_10[221]},
      {stage2_10[100]}
   );
   gpc1_1 gpc6290 (
      {stage1_10[222]},
      {stage2_10[101]}
   );
   gpc1_1 gpc6291 (
      {stage1_10[223]},
      {stage2_10[102]}
   );
   gpc1_1 gpc6292 (
      {stage1_10[224]},
      {stage2_10[103]}
   );
   gpc1_1 gpc6293 (
      {stage1_10[225]},
      {stage2_10[104]}
   );
   gpc1_1 gpc6294 (
      {stage1_10[226]},
      {stage2_10[105]}
   );
   gpc1_1 gpc6295 (
      {stage1_10[227]},
      {stage2_10[106]}
   );
   gpc1_1 gpc6296 (
      {stage1_10[228]},
      {stage2_10[107]}
   );
   gpc1_1 gpc6297 (
      {stage1_10[229]},
      {stage2_10[108]}
   );
   gpc1_1 gpc6298 (
      {stage1_10[230]},
      {stage2_10[109]}
   );
   gpc1_1 gpc6299 (
      {stage1_10[231]},
      {stage2_10[110]}
   );
   gpc1_1 gpc6300 (
      {stage1_10[232]},
      {stage2_10[111]}
   );
   gpc1_1 gpc6301 (
      {stage1_10[233]},
      {stage2_10[112]}
   );
   gpc1_1 gpc6302 (
      {stage1_10[234]},
      {stage2_10[113]}
   );
   gpc1_1 gpc6303 (
      {stage1_10[235]},
      {stage2_10[114]}
   );
   gpc1_1 gpc6304 (
      {stage1_10[236]},
      {stage2_10[115]}
   );
   gpc1_1 gpc6305 (
      {stage1_10[237]},
      {stage2_10[116]}
   );
   gpc1_1 gpc6306 (
      {stage1_10[238]},
      {stage2_10[117]}
   );
   gpc1_1 gpc6307 (
      {stage1_10[239]},
      {stage2_10[118]}
   );
   gpc1_1 gpc6308 (
      {stage1_10[240]},
      {stage2_10[119]}
   );
   gpc1_1 gpc6309 (
      {stage1_10[241]},
      {stage2_10[120]}
   );
   gpc1_1 gpc6310 (
      {stage1_10[242]},
      {stage2_10[121]}
   );
   gpc1_1 gpc6311 (
      {stage1_10[243]},
      {stage2_10[122]}
   );
   gpc1_1 gpc6312 (
      {stage1_10[244]},
      {stage2_10[123]}
   );
   gpc1_1 gpc6313 (
      {stage1_10[245]},
      {stage2_10[124]}
   );
   gpc1_1 gpc6314 (
      {stage1_10[246]},
      {stage2_10[125]}
   );
   gpc1_1 gpc6315 (
      {stage1_10[247]},
      {stage2_10[126]}
   );
   gpc1_1 gpc6316 (
      {stage1_10[248]},
      {stage2_10[127]}
   );
   gpc1_1 gpc6317 (
      {stage1_10[249]},
      {stage2_10[128]}
   );
   gpc1_1 gpc6318 (
      {stage1_10[250]},
      {stage2_10[129]}
   );
   gpc1_1 gpc6319 (
      {stage1_10[251]},
      {stage2_10[130]}
   );
   gpc1_1 gpc6320 (
      {stage1_10[252]},
      {stage2_10[131]}
   );
   gpc1_1 gpc6321 (
      {stage1_10[253]},
      {stage2_10[132]}
   );
   gpc1_1 gpc6322 (
      {stage1_10[254]},
      {stage2_10[133]}
   );
   gpc1_1 gpc6323 (
      {stage1_10[255]},
      {stage2_10[134]}
   );
   gpc1_1 gpc6324 (
      {stage1_10[256]},
      {stage2_10[135]}
   );
   gpc1_1 gpc6325 (
      {stage1_10[257]},
      {stage2_10[136]}
   );
   gpc1_1 gpc6326 (
      {stage1_10[258]},
      {stage2_10[137]}
   );
   gpc1_1 gpc6327 (
      {stage1_10[259]},
      {stage2_10[138]}
   );
   gpc1_1 gpc6328 (
      {stage1_10[260]},
      {stage2_10[139]}
   );
   gpc1_1 gpc6329 (
      {stage1_10[261]},
      {stage2_10[140]}
   );
   gpc1_1 gpc6330 (
      {stage1_10[262]},
      {stage2_10[141]}
   );
   gpc1_1 gpc6331 (
      {stage1_10[263]},
      {stage2_10[142]}
   );
   gpc1_1 gpc6332 (
      {stage1_10[264]},
      {stage2_10[143]}
   );
   gpc1_1 gpc6333 (
      {stage1_10[265]},
      {stage2_10[144]}
   );
   gpc1_1 gpc6334 (
      {stage1_10[266]},
      {stage2_10[145]}
   );
   gpc1_1 gpc6335 (
      {stage1_10[267]},
      {stage2_10[146]}
   );
   gpc1_1 gpc6336 (
      {stage1_10[268]},
      {stage2_10[147]}
   );
   gpc1_1 gpc6337 (
      {stage1_10[269]},
      {stage2_10[148]}
   );
   gpc1_1 gpc6338 (
      {stage1_10[270]},
      {stage2_10[149]}
   );
   gpc1_1 gpc6339 (
      {stage1_10[271]},
      {stage2_10[150]}
   );
   gpc1_1 gpc6340 (
      {stage1_10[272]},
      {stage2_10[151]}
   );
   gpc1_1 gpc6341 (
      {stage1_10[273]},
      {stage2_10[152]}
   );
   gpc1_1 gpc6342 (
      {stage1_10[274]},
      {stage2_10[153]}
   );
   gpc1_1 gpc6343 (
      {stage1_10[275]},
      {stage2_10[154]}
   );
   gpc1_1 gpc6344 (
      {stage1_10[276]},
      {stage2_10[155]}
   );
   gpc1_1 gpc6345 (
      {stage1_10[277]},
      {stage2_10[156]}
   );
   gpc1_1 gpc6346 (
      {stage1_10[278]},
      {stage2_10[157]}
   );
   gpc1_1 gpc6347 (
      {stage1_10[279]},
      {stage2_10[158]}
   );
   gpc1_1 gpc6348 (
      {stage1_10[280]},
      {stage2_10[159]}
   );
   gpc1_1 gpc6349 (
      {stage1_10[281]},
      {stage2_10[160]}
   );
   gpc1_1 gpc6350 (
      {stage1_10[282]},
      {stage2_10[161]}
   );
   gpc1_1 gpc6351 (
      {stage1_10[283]},
      {stage2_10[162]}
   );
   gpc1_1 gpc6352 (
      {stage1_10[284]},
      {stage2_10[163]}
   );
   gpc1_1 gpc6353 (
      {stage1_11[228]},
      {stage2_11[90]}
   );
   gpc1_1 gpc6354 (
      {stage1_11[229]},
      {stage2_11[91]}
   );
   gpc1_1 gpc6355 (
      {stage1_11[230]},
      {stage2_11[92]}
   );
   gpc1_1 gpc6356 (
      {stage1_11[231]},
      {stage2_11[93]}
   );
   gpc1_1 gpc6357 (
      {stage1_11[232]},
      {stage2_11[94]}
   );
   gpc1_1 gpc6358 (
      {stage1_11[233]},
      {stage2_11[95]}
   );
   gpc1_1 gpc6359 (
      {stage1_11[234]},
      {stage2_11[96]}
   );
   gpc1_1 gpc6360 (
      {stage1_11[235]},
      {stage2_11[97]}
   );
   gpc1_1 gpc6361 (
      {stage1_11[236]},
      {stage2_11[98]}
   );
   gpc1_1 gpc6362 (
      {stage1_11[237]},
      {stage2_11[99]}
   );
   gpc1_1 gpc6363 (
      {stage1_11[238]},
      {stage2_11[100]}
   );
   gpc1_1 gpc6364 (
      {stage1_11[239]},
      {stage2_11[101]}
   );
   gpc1_1 gpc6365 (
      {stage1_11[240]},
      {stage2_11[102]}
   );
   gpc1_1 gpc6366 (
      {stage1_11[241]},
      {stage2_11[103]}
   );
   gpc1_1 gpc6367 (
      {stage1_11[242]},
      {stage2_11[104]}
   );
   gpc1_1 gpc6368 (
      {stage1_11[243]},
      {stage2_11[105]}
   );
   gpc1_1 gpc6369 (
      {stage1_11[244]},
      {stage2_11[106]}
   );
   gpc1_1 gpc6370 (
      {stage1_11[245]},
      {stage2_11[107]}
   );
   gpc1_1 gpc6371 (
      {stage1_11[246]},
      {stage2_11[108]}
   );
   gpc1_1 gpc6372 (
      {stage1_11[247]},
      {stage2_11[109]}
   );
   gpc1_1 gpc6373 (
      {stage1_11[248]},
      {stage2_11[110]}
   );
   gpc1_1 gpc6374 (
      {stage1_11[249]},
      {stage2_11[111]}
   );
   gpc1_1 gpc6375 (
      {stage1_11[250]},
      {stage2_11[112]}
   );
   gpc1_1 gpc6376 (
      {stage1_11[251]},
      {stage2_11[113]}
   );
   gpc1_1 gpc6377 (
      {stage1_11[252]},
      {stage2_11[114]}
   );
   gpc1_1 gpc6378 (
      {stage1_11[253]},
      {stage2_11[115]}
   );
   gpc1_1 gpc6379 (
      {stage1_11[254]},
      {stage2_11[116]}
   );
   gpc1_1 gpc6380 (
      {stage1_11[255]},
      {stage2_11[117]}
   );
   gpc1_1 gpc6381 (
      {stage1_11[256]},
      {stage2_11[118]}
   );
   gpc1_1 gpc6382 (
      {stage1_11[257]},
      {stage2_11[119]}
   );
   gpc1_1 gpc6383 (
      {stage1_11[258]},
      {stage2_11[120]}
   );
   gpc1_1 gpc6384 (
      {stage1_11[259]},
      {stage2_11[121]}
   );
   gpc1_1 gpc6385 (
      {stage1_11[260]},
      {stage2_11[122]}
   );
   gpc1_1 gpc6386 (
      {stage1_11[261]},
      {stage2_11[123]}
   );
   gpc1_1 gpc6387 (
      {stage1_11[262]},
      {stage2_11[124]}
   );
   gpc1_1 gpc6388 (
      {stage1_11[263]},
      {stage2_11[125]}
   );
   gpc1_1 gpc6389 (
      {stage1_11[264]},
      {stage2_11[126]}
   );
   gpc1_1 gpc6390 (
      {stage1_11[265]},
      {stage2_11[127]}
   );
   gpc1_1 gpc6391 (
      {stage1_11[266]},
      {stage2_11[128]}
   );
   gpc1_1 gpc6392 (
      {stage1_11[267]},
      {stage2_11[129]}
   );
   gpc1_1 gpc6393 (
      {stage1_11[268]},
      {stage2_11[130]}
   );
   gpc1_1 gpc6394 (
      {stage1_11[269]},
      {stage2_11[131]}
   );
   gpc1_1 gpc6395 (
      {stage1_11[270]},
      {stage2_11[132]}
   );
   gpc1_1 gpc6396 (
      {stage1_11[271]},
      {stage2_11[133]}
   );
   gpc1_1 gpc6397 (
      {stage1_11[272]},
      {stage2_11[134]}
   );
   gpc1_1 gpc6398 (
      {stage1_11[273]},
      {stage2_11[135]}
   );
   gpc1_1 gpc6399 (
      {stage1_11[274]},
      {stage2_11[136]}
   );
   gpc1_1 gpc6400 (
      {stage1_11[275]},
      {stage2_11[137]}
   );
   gpc1_1 gpc6401 (
      {stage1_11[276]},
      {stage2_11[138]}
   );
   gpc1_1 gpc6402 (
      {stage1_12[163]},
      {stage2_12[81]}
   );
   gpc1_1 gpc6403 (
      {stage1_12[164]},
      {stage2_12[82]}
   );
   gpc1_1 gpc6404 (
      {stage1_12[165]},
      {stage2_12[83]}
   );
   gpc1_1 gpc6405 (
      {stage1_12[166]},
      {stage2_12[84]}
   );
   gpc1_1 gpc6406 (
      {stage1_12[167]},
      {stage2_12[85]}
   );
   gpc1_1 gpc6407 (
      {stage1_12[168]},
      {stage2_12[86]}
   );
   gpc1_1 gpc6408 (
      {stage1_12[169]},
      {stage2_12[87]}
   );
   gpc1_1 gpc6409 (
      {stage1_12[170]},
      {stage2_12[88]}
   );
   gpc1_1 gpc6410 (
      {stage1_12[171]},
      {stage2_12[89]}
   );
   gpc1_1 gpc6411 (
      {stage1_12[172]},
      {stage2_12[90]}
   );
   gpc1_1 gpc6412 (
      {stage1_12[173]},
      {stage2_12[91]}
   );
   gpc1_1 gpc6413 (
      {stage1_12[174]},
      {stage2_12[92]}
   );
   gpc1_1 gpc6414 (
      {stage1_12[175]},
      {stage2_12[93]}
   );
   gpc1_1 gpc6415 (
      {stage1_12[176]},
      {stage2_12[94]}
   );
   gpc1_1 gpc6416 (
      {stage1_12[177]},
      {stage2_12[95]}
   );
   gpc1_1 gpc6417 (
      {stage1_12[178]},
      {stage2_12[96]}
   );
   gpc1_1 gpc6418 (
      {stage1_12[179]},
      {stage2_12[97]}
   );
   gpc1_1 gpc6419 (
      {stage1_12[180]},
      {stage2_12[98]}
   );
   gpc1_1 gpc6420 (
      {stage1_12[181]},
      {stage2_12[99]}
   );
   gpc1_1 gpc6421 (
      {stage1_12[182]},
      {stage2_12[100]}
   );
   gpc1_1 gpc6422 (
      {stage1_12[183]},
      {stage2_12[101]}
   );
   gpc1_1 gpc6423 (
      {stage1_12[184]},
      {stage2_12[102]}
   );
   gpc1_1 gpc6424 (
      {stage1_12[185]},
      {stage2_12[103]}
   );
   gpc1_1 gpc6425 (
      {stage1_12[186]},
      {stage2_12[104]}
   );
   gpc1_1 gpc6426 (
      {stage1_12[187]},
      {stage2_12[105]}
   );
   gpc1_1 gpc6427 (
      {stage1_12[188]},
      {stage2_12[106]}
   );
   gpc1_1 gpc6428 (
      {stage1_14[217]},
      {stage2_14[106]}
   );
   gpc1_1 gpc6429 (
      {stage1_14[218]},
      {stage2_14[107]}
   );
   gpc1_1 gpc6430 (
      {stage1_15[123]},
      {stage2_15[93]}
   );
   gpc1_1 gpc6431 (
      {stage1_15[124]},
      {stage2_15[94]}
   );
   gpc1_1 gpc6432 (
      {stage1_15[125]},
      {stage2_15[95]}
   );
   gpc1_1 gpc6433 (
      {stage1_15[126]},
      {stage2_15[96]}
   );
   gpc1_1 gpc6434 (
      {stage1_15[127]},
      {stage2_15[97]}
   );
   gpc1_1 gpc6435 (
      {stage1_15[128]},
      {stage2_15[98]}
   );
   gpc1_1 gpc6436 (
      {stage1_15[129]},
      {stage2_15[99]}
   );
   gpc1_1 gpc6437 (
      {stage1_15[130]},
      {stage2_15[100]}
   );
   gpc1_1 gpc6438 (
      {stage1_15[131]},
      {stage2_15[101]}
   );
   gpc1_1 gpc6439 (
      {stage1_15[132]},
      {stage2_15[102]}
   );
   gpc1_1 gpc6440 (
      {stage1_15[133]},
      {stage2_15[103]}
   );
   gpc1_1 gpc6441 (
      {stage1_15[134]},
      {stage2_15[104]}
   );
   gpc1_1 gpc6442 (
      {stage1_15[135]},
      {stage2_15[105]}
   );
   gpc1_1 gpc6443 (
      {stage1_15[136]},
      {stage2_15[106]}
   );
   gpc1_1 gpc6444 (
      {stage1_15[137]},
      {stage2_15[107]}
   );
   gpc1_1 gpc6445 (
      {stage1_15[138]},
      {stage2_15[108]}
   );
   gpc1_1 gpc6446 (
      {stage1_15[139]},
      {stage2_15[109]}
   );
   gpc1_1 gpc6447 (
      {stage1_15[140]},
      {stage2_15[110]}
   );
   gpc1_1 gpc6448 (
      {stage1_15[141]},
      {stage2_15[111]}
   );
   gpc1_1 gpc6449 (
      {stage1_15[142]},
      {stage2_15[112]}
   );
   gpc1_1 gpc6450 (
      {stage1_15[143]},
      {stage2_15[113]}
   );
   gpc1_1 gpc6451 (
      {stage1_15[144]},
      {stage2_15[114]}
   );
   gpc1_1 gpc6452 (
      {stage1_15[145]},
      {stage2_15[115]}
   );
   gpc1_1 gpc6453 (
      {stage1_15[146]},
      {stage2_15[116]}
   );
   gpc1_1 gpc6454 (
      {stage1_15[147]},
      {stage2_15[117]}
   );
   gpc1_1 gpc6455 (
      {stage1_15[148]},
      {stage2_15[118]}
   );
   gpc1_1 gpc6456 (
      {stage1_15[149]},
      {stage2_15[119]}
   );
   gpc1_1 gpc6457 (
      {stage1_15[150]},
      {stage2_15[120]}
   );
   gpc1_1 gpc6458 (
      {stage1_15[151]},
      {stage2_15[121]}
   );
   gpc1_1 gpc6459 (
      {stage1_15[152]},
      {stage2_15[122]}
   );
   gpc1_1 gpc6460 (
      {stage1_15[153]},
      {stage2_15[123]}
   );
   gpc1_1 gpc6461 (
      {stage1_15[154]},
      {stage2_15[124]}
   );
   gpc1_1 gpc6462 (
      {stage1_15[155]},
      {stage2_15[125]}
   );
   gpc1_1 gpc6463 (
      {stage1_15[156]},
      {stage2_15[126]}
   );
   gpc1_1 gpc6464 (
      {stage1_15[157]},
      {stage2_15[127]}
   );
   gpc1_1 gpc6465 (
      {stage1_15[158]},
      {stage2_15[128]}
   );
   gpc1_1 gpc6466 (
      {stage1_15[159]},
      {stage2_15[129]}
   );
   gpc1_1 gpc6467 (
      {stage1_15[160]},
      {stage2_15[130]}
   );
   gpc1_1 gpc6468 (
      {stage1_15[161]},
      {stage2_15[131]}
   );
   gpc1_1 gpc6469 (
      {stage1_15[162]},
      {stage2_15[132]}
   );
   gpc1_1 gpc6470 (
      {stage1_15[163]},
      {stage2_15[133]}
   );
   gpc1_1 gpc6471 (
      {stage1_15[164]},
      {stage2_15[134]}
   );
   gpc1_1 gpc6472 (
      {stage1_15[165]},
      {stage2_15[135]}
   );
   gpc1_1 gpc6473 (
      {stage1_15[166]},
      {stage2_15[136]}
   );
   gpc1_1 gpc6474 (
      {stage1_15[167]},
      {stage2_15[137]}
   );
   gpc1_1 gpc6475 (
      {stage1_15[168]},
      {stage2_15[138]}
   );
   gpc1_1 gpc6476 (
      {stage1_15[169]},
      {stage2_15[139]}
   );
   gpc1_1 gpc6477 (
      {stage1_15[170]},
      {stage2_15[140]}
   );
   gpc1_1 gpc6478 (
      {stage1_16[198]},
      {stage2_16[59]}
   );
   gpc1_1 gpc6479 (
      {stage1_16[199]},
      {stage2_16[60]}
   );
   gpc1_1 gpc6480 (
      {stage1_16[200]},
      {stage2_16[61]}
   );
   gpc1_1 gpc6481 (
      {stage1_16[201]},
      {stage2_16[62]}
   );
   gpc1_1 gpc6482 (
      {stage1_16[202]},
      {stage2_16[63]}
   );
   gpc1_1 gpc6483 (
      {stage1_16[203]},
      {stage2_16[64]}
   );
   gpc1_1 gpc6484 (
      {stage1_16[204]},
      {stage2_16[65]}
   );
   gpc1_1 gpc6485 (
      {stage1_16[205]},
      {stage2_16[66]}
   );
   gpc1_1 gpc6486 (
      {stage1_16[206]},
      {stage2_16[67]}
   );
   gpc1_1 gpc6487 (
      {stage1_16[207]},
      {stage2_16[68]}
   );
   gpc1_1 gpc6488 (
      {stage1_16[208]},
      {stage2_16[69]}
   );
   gpc1_1 gpc6489 (
      {stage1_16[209]},
      {stage2_16[70]}
   );
   gpc1_1 gpc6490 (
      {stage1_16[210]},
      {stage2_16[71]}
   );
   gpc1_1 gpc6491 (
      {stage1_16[211]},
      {stage2_16[72]}
   );
   gpc1_1 gpc6492 (
      {stage1_16[212]},
      {stage2_16[73]}
   );
   gpc1_1 gpc6493 (
      {stage1_16[213]},
      {stage2_16[74]}
   );
   gpc1_1 gpc6494 (
      {stage1_16[214]},
      {stage2_16[75]}
   );
   gpc1_1 gpc6495 (
      {stage1_16[215]},
      {stage2_16[76]}
   );
   gpc1_1 gpc6496 (
      {stage1_16[216]},
      {stage2_16[77]}
   );
   gpc1_1 gpc6497 (
      {stage1_16[217]},
      {stage2_16[78]}
   );
   gpc1_1 gpc6498 (
      {stage1_16[218]},
      {stage2_16[79]}
   );
   gpc1_1 gpc6499 (
      {stage1_16[219]},
      {stage2_16[80]}
   );
   gpc1_1 gpc6500 (
      {stage1_16[220]},
      {stage2_16[81]}
   );
   gpc1_1 gpc6501 (
      {stage1_16[221]},
      {stage2_16[82]}
   );
   gpc1_1 gpc6502 (
      {stage1_17[228]},
      {stage2_17[86]}
   );
   gpc1_1 gpc6503 (
      {stage1_18[191]},
      {stage2_18[101]}
   );
   gpc1_1 gpc6504 (
      {stage1_18[192]},
      {stage2_18[102]}
   );
   gpc1_1 gpc6505 (
      {stage1_18[193]},
      {stage2_18[103]}
   );
   gpc1_1 gpc6506 (
      {stage1_18[194]},
      {stage2_18[104]}
   );
   gpc1_1 gpc6507 (
      {stage1_18[195]},
      {stage2_18[105]}
   );
   gpc1_1 gpc6508 (
      {stage1_18[196]},
      {stage2_18[106]}
   );
   gpc1_1 gpc6509 (
      {stage1_18[197]},
      {stage2_18[107]}
   );
   gpc1_1 gpc6510 (
      {stage1_18[198]},
      {stage2_18[108]}
   );
   gpc1_1 gpc6511 (
      {stage1_18[199]},
      {stage2_18[109]}
   );
   gpc1_1 gpc6512 (
      {stage1_18[200]},
      {stage2_18[110]}
   );
   gpc1_1 gpc6513 (
      {stage1_18[201]},
      {stage2_18[111]}
   );
   gpc1_1 gpc6514 (
      {stage1_18[202]},
      {stage2_18[112]}
   );
   gpc1_1 gpc6515 (
      {stage1_18[203]},
      {stage2_18[113]}
   );
   gpc1_1 gpc6516 (
      {stage1_18[204]},
      {stage2_18[114]}
   );
   gpc1_1 gpc6517 (
      {stage1_18[205]},
      {stage2_18[115]}
   );
   gpc1_1 gpc6518 (
      {stage1_18[206]},
      {stage2_18[116]}
   );
   gpc1_1 gpc6519 (
      {stage1_18[207]},
      {stage2_18[117]}
   );
   gpc1_1 gpc6520 (
      {stage1_18[208]},
      {stage2_18[118]}
   );
   gpc1_1 gpc6521 (
      {stage1_19[234]},
      {stage2_19[71]}
   );
   gpc1_1 gpc6522 (
      {stage1_19[235]},
      {stage2_19[72]}
   );
   gpc1_1 gpc6523 (
      {stage1_19[236]},
      {stage2_19[73]}
   );
   gpc1_1 gpc6524 (
      {stage1_19[237]},
      {stage2_19[74]}
   );
   gpc1_1 gpc6525 (
      {stage1_19[238]},
      {stage2_19[75]}
   );
   gpc1_1 gpc6526 (
      {stage1_19[239]},
      {stage2_19[76]}
   );
   gpc1_1 gpc6527 (
      {stage1_19[240]},
      {stage2_19[77]}
   );
   gpc1_1 gpc6528 (
      {stage1_19[241]},
      {stage2_19[78]}
   );
   gpc1_1 gpc6529 (
      {stage1_19[242]},
      {stage2_19[79]}
   );
   gpc1_1 gpc6530 (
      {stage1_19[243]},
      {stage2_19[80]}
   );
   gpc1_1 gpc6531 (
      {stage1_19[244]},
      {stage2_19[81]}
   );
   gpc1_1 gpc6532 (
      {stage1_19[245]},
      {stage2_19[82]}
   );
   gpc1_1 gpc6533 (
      {stage1_19[246]},
      {stage2_19[83]}
   );
   gpc1_1 gpc6534 (
      {stage1_19[247]},
      {stage2_19[84]}
   );
   gpc1_1 gpc6535 (
      {stage1_19[248]},
      {stage2_19[85]}
   );
   gpc1_1 gpc6536 (
      {stage1_19[249]},
      {stage2_19[86]}
   );
   gpc1_1 gpc6537 (
      {stage1_19[250]},
      {stage2_19[87]}
   );
   gpc1_1 gpc6538 (
      {stage1_19[251]},
      {stage2_19[88]}
   );
   gpc1_1 gpc6539 (
      {stage1_19[252]},
      {stage2_19[89]}
   );
   gpc1_1 gpc6540 (
      {stage1_19[253]},
      {stage2_19[90]}
   );
   gpc1_1 gpc6541 (
      {stage1_19[254]},
      {stage2_19[91]}
   );
   gpc1_1 gpc6542 (
      {stage1_19[255]},
      {stage2_19[92]}
   );
   gpc1_1 gpc6543 (
      {stage1_19[256]},
      {stage2_19[93]}
   );
   gpc1_1 gpc6544 (
      {stage1_19[257]},
      {stage2_19[94]}
   );
   gpc1_1 gpc6545 (
      {stage1_19[258]},
      {stage2_19[95]}
   );
   gpc1_1 gpc6546 (
      {stage1_19[259]},
      {stage2_19[96]}
   );
   gpc1_1 gpc6547 (
      {stage1_19[260]},
      {stage2_19[97]}
   );
   gpc1_1 gpc6548 (
      {stage1_19[261]},
      {stage2_19[98]}
   );
   gpc1_1 gpc6549 (
      {stage1_19[262]},
      {stage2_19[99]}
   );
   gpc1_1 gpc6550 (
      {stage1_19[263]},
      {stage2_19[100]}
   );
   gpc1_1 gpc6551 (
      {stage1_19[264]},
      {stage2_19[101]}
   );
   gpc1_1 gpc6552 (
      {stage1_19[265]},
      {stage2_19[102]}
   );
   gpc1_1 gpc6553 (
      {stage1_19[266]},
      {stage2_19[103]}
   );
   gpc1_1 gpc6554 (
      {stage1_19[267]},
      {stage2_19[104]}
   );
   gpc1_1 gpc6555 (
      {stage1_19[268]},
      {stage2_19[105]}
   );
   gpc1_1 gpc6556 (
      {stage1_19[269]},
      {stage2_19[106]}
   );
   gpc1_1 gpc6557 (
      {stage1_19[270]},
      {stage2_19[107]}
   );
   gpc1_1 gpc6558 (
      {stage1_19[271]},
      {stage2_19[108]}
   );
   gpc1_1 gpc6559 (
      {stage1_19[272]},
      {stage2_19[109]}
   );
   gpc1_1 gpc6560 (
      {stage1_19[273]},
      {stage2_19[110]}
   );
   gpc1_1 gpc6561 (
      {stage1_19[274]},
      {stage2_19[111]}
   );
   gpc1_1 gpc6562 (
      {stage1_19[275]},
      {stage2_19[112]}
   );
   gpc1_1 gpc6563 (
      {stage1_20[262]},
      {stage2_20[87]}
   );
   gpc1_1 gpc6564 (
      {stage1_20[263]},
      {stage2_20[88]}
   );
   gpc1_1 gpc6565 (
      {stage1_20[264]},
      {stage2_20[89]}
   );
   gpc1_1 gpc6566 (
      {stage1_20[265]},
      {stage2_20[90]}
   );
   gpc1_1 gpc6567 (
      {stage1_20[266]},
      {stage2_20[91]}
   );
   gpc1_1 gpc6568 (
      {stage1_20[267]},
      {stage2_20[92]}
   );
   gpc1_1 gpc6569 (
      {stage1_21[174]},
      {stage2_21[112]}
   );
   gpc1_1 gpc6570 (
      {stage1_21[175]},
      {stage2_21[113]}
   );
   gpc1_1 gpc6571 (
      {stage1_21[176]},
      {stage2_21[114]}
   );
   gpc1_1 gpc6572 (
      {stage1_21[177]},
      {stage2_21[115]}
   );
   gpc1_1 gpc6573 (
      {stage1_21[178]},
      {stage2_21[116]}
   );
   gpc1_1 gpc6574 (
      {stage1_21[179]},
      {stage2_21[117]}
   );
   gpc1_1 gpc6575 (
      {stage1_21[180]},
      {stage2_21[118]}
   );
   gpc1_1 gpc6576 (
      {stage1_21[181]},
      {stage2_21[119]}
   );
   gpc1_1 gpc6577 (
      {stage1_21[182]},
      {stage2_21[120]}
   );
   gpc1_1 gpc6578 (
      {stage1_21[183]},
      {stage2_21[121]}
   );
   gpc1_1 gpc6579 (
      {stage1_21[184]},
      {stage2_21[122]}
   );
   gpc1_1 gpc6580 (
      {stage1_21[185]},
      {stage2_21[123]}
   );
   gpc1_1 gpc6581 (
      {stage1_21[186]},
      {stage2_21[124]}
   );
   gpc1_1 gpc6582 (
      {stage1_21[187]},
      {stage2_21[125]}
   );
   gpc1_1 gpc6583 (
      {stage1_21[188]},
      {stage2_21[126]}
   );
   gpc1_1 gpc6584 (
      {stage1_21[189]},
      {stage2_21[127]}
   );
   gpc1_1 gpc6585 (
      {stage1_22[145]},
      {stage2_22[82]}
   );
   gpc1_1 gpc6586 (
      {stage1_22[146]},
      {stage2_22[83]}
   );
   gpc1_1 gpc6587 (
      {stage1_22[147]},
      {stage2_22[84]}
   );
   gpc1_1 gpc6588 (
      {stage1_22[148]},
      {stage2_22[85]}
   );
   gpc1_1 gpc6589 (
      {stage1_22[149]},
      {stage2_22[86]}
   );
   gpc1_1 gpc6590 (
      {stage1_22[150]},
      {stage2_22[87]}
   );
   gpc1_1 gpc6591 (
      {stage1_22[151]},
      {stage2_22[88]}
   );
   gpc1_1 gpc6592 (
      {stage1_22[152]},
      {stage2_22[89]}
   );
   gpc1_1 gpc6593 (
      {stage1_22[153]},
      {stage2_22[90]}
   );
   gpc1_1 gpc6594 (
      {stage1_22[154]},
      {stage2_22[91]}
   );
   gpc1_1 gpc6595 (
      {stage1_22[155]},
      {stage2_22[92]}
   );
   gpc1_1 gpc6596 (
      {stage1_22[156]},
      {stage2_22[93]}
   );
   gpc1_1 gpc6597 (
      {stage1_22[157]},
      {stage2_22[94]}
   );
   gpc1_1 gpc6598 (
      {stage1_22[158]},
      {stage2_22[95]}
   );
   gpc1_1 gpc6599 (
      {stage1_22[159]},
      {stage2_22[96]}
   );
   gpc1_1 gpc6600 (
      {stage1_22[160]},
      {stage2_22[97]}
   );
   gpc1_1 gpc6601 (
      {stage1_22[161]},
      {stage2_22[98]}
   );
   gpc1_1 gpc6602 (
      {stage1_22[162]},
      {stage2_22[99]}
   );
   gpc1_1 gpc6603 (
      {stage1_22[163]},
      {stage2_22[100]}
   );
   gpc1_1 gpc6604 (
      {stage1_22[164]},
      {stage2_22[101]}
   );
   gpc1_1 gpc6605 (
      {stage1_22[165]},
      {stage2_22[102]}
   );
   gpc1_1 gpc6606 (
      {stage1_22[166]},
      {stage2_22[103]}
   );
   gpc1_1 gpc6607 (
      {stage1_22[167]},
      {stage2_22[104]}
   );
   gpc1_1 gpc6608 (
      {stage1_22[168]},
      {stage2_22[105]}
   );
   gpc1_1 gpc6609 (
      {stage1_22[169]},
      {stage2_22[106]}
   );
   gpc1_1 gpc6610 (
      {stage1_22[170]},
      {stage2_22[107]}
   );
   gpc1_1 gpc6611 (
      {stage1_24[210]},
      {stage2_24[98]}
   );
   gpc1_1 gpc6612 (
      {stage1_24[211]},
      {stage2_24[99]}
   );
   gpc1_1 gpc6613 (
      {stage1_24[212]},
      {stage2_24[100]}
   );
   gpc1_1 gpc6614 (
      {stage1_24[213]},
      {stage2_24[101]}
   );
   gpc1_1 gpc6615 (
      {stage1_25[175]},
      {stage2_25[87]}
   );
   gpc1_1 gpc6616 (
      {stage1_25[176]},
      {stage2_25[88]}
   );
   gpc1_1 gpc6617 (
      {stage1_25[177]},
      {stage2_25[89]}
   );
   gpc1_1 gpc6618 (
      {stage1_25[178]},
      {stage2_25[90]}
   );
   gpc1_1 gpc6619 (
      {stage1_25[179]},
      {stage2_25[91]}
   );
   gpc1_1 gpc6620 (
      {stage1_25[180]},
      {stage2_25[92]}
   );
   gpc1_1 gpc6621 (
      {stage1_25[181]},
      {stage2_25[93]}
   );
   gpc1_1 gpc6622 (
      {stage1_25[182]},
      {stage2_25[94]}
   );
   gpc1_1 gpc6623 (
      {stage1_25[183]},
      {stage2_25[95]}
   );
   gpc1_1 gpc6624 (
      {stage1_26[248]},
      {stage2_26[82]}
   );
   gpc1_1 gpc6625 (
      {stage1_26[249]},
      {stage2_26[83]}
   );
   gpc1_1 gpc6626 (
      {stage1_26[250]},
      {stage2_26[84]}
   );
   gpc1_1 gpc6627 (
      {stage1_29[216]},
      {stage2_29[74]}
   );
   gpc1_1 gpc6628 (
      {stage1_29[217]},
      {stage2_29[75]}
   );
   gpc1_1 gpc6629 (
      {stage1_29[218]},
      {stage2_29[76]}
   );
   gpc1_1 gpc6630 (
      {stage1_29[219]},
      {stage2_29[77]}
   );
   gpc1_1 gpc6631 (
      {stage1_29[220]},
      {stage2_29[78]}
   );
   gpc1_1 gpc6632 (
      {stage1_29[221]},
      {stage2_29[79]}
   );
   gpc1_1 gpc6633 (
      {stage1_29[222]},
      {stage2_29[80]}
   );
   gpc1_1 gpc6634 (
      {stage1_29[223]},
      {stage2_29[81]}
   );
   gpc1_1 gpc6635 (
      {stage1_29[224]},
      {stage2_29[82]}
   );
   gpc1_1 gpc6636 (
      {stage1_29[225]},
      {stage2_29[83]}
   );
   gpc1_1 gpc6637 (
      {stage1_29[226]},
      {stage2_29[84]}
   );
   gpc1_1 gpc6638 (
      {stage1_29[227]},
      {stage2_29[85]}
   );
   gpc1_1 gpc6639 (
      {stage1_29[228]},
      {stage2_29[86]}
   );
   gpc1_1 gpc6640 (
      {stage1_30[160]},
      {stage2_30[85]}
   );
   gpc1_1 gpc6641 (
      {stage1_30[161]},
      {stage2_30[86]}
   );
   gpc1_1 gpc6642 (
      {stage1_30[162]},
      {stage2_30[87]}
   );
   gpc1_1 gpc6643 (
      {stage1_30[163]},
      {stage2_30[88]}
   );
   gpc1_1 gpc6644 (
      {stage1_30[164]},
      {stage2_30[89]}
   );
   gpc1_1 gpc6645 (
      {stage1_30[165]},
      {stage2_30[90]}
   );
   gpc1_1 gpc6646 (
      {stage1_30[166]},
      {stage2_30[91]}
   );
   gpc1_1 gpc6647 (
      {stage1_30[167]},
      {stage2_30[92]}
   );
   gpc1_1 gpc6648 (
      {stage1_30[168]},
      {stage2_30[93]}
   );
   gpc1_1 gpc6649 (
      {stage1_30[169]},
      {stage2_30[94]}
   );
   gpc1_1 gpc6650 (
      {stage1_30[170]},
      {stage2_30[95]}
   );
   gpc1_1 gpc6651 (
      {stage1_30[171]},
      {stage2_30[96]}
   );
   gpc1_1 gpc6652 (
      {stage1_30[172]},
      {stage2_30[97]}
   );
   gpc1_1 gpc6653 (
      {stage1_30[173]},
      {stage2_30[98]}
   );
   gpc1_1 gpc6654 (
      {stage1_30[174]},
      {stage2_30[99]}
   );
   gpc1_1 gpc6655 (
      {stage1_30[175]},
      {stage2_30[100]}
   );
   gpc1_1 gpc6656 (
      {stage1_30[176]},
      {stage2_30[101]}
   );
   gpc1_1 gpc6657 (
      {stage1_30[177]},
      {stage2_30[102]}
   );
   gpc1_1 gpc6658 (
      {stage1_30[178]},
      {stage2_30[103]}
   );
   gpc1_1 gpc6659 (
      {stage1_30[179]},
      {stage2_30[104]}
   );
   gpc1_1 gpc6660 (
      {stage1_30[180]},
      {stage2_30[105]}
   );
   gpc1_1 gpc6661 (
      {stage1_30[181]},
      {stage2_30[106]}
   );
   gpc1_1 gpc6662 (
      {stage1_30[182]},
      {stage2_30[107]}
   );
   gpc1_1 gpc6663 (
      {stage1_30[183]},
      {stage2_30[108]}
   );
   gpc1_1 gpc6664 (
      {stage1_30[184]},
      {stage2_30[109]}
   );
   gpc1_1 gpc6665 (
      {stage1_30[185]},
      {stage2_30[110]}
   );
   gpc1_1 gpc6666 (
      {stage1_30[186]},
      {stage2_30[111]}
   );
   gpc1_1 gpc6667 (
      {stage1_30[187]},
      {stage2_30[112]}
   );
   gpc1_1 gpc6668 (
      {stage1_30[188]},
      {stage2_30[113]}
   );
   gpc1_1 gpc6669 (
      {stage1_30[189]},
      {stage2_30[114]}
   );
   gpc1_1 gpc6670 (
      {stage1_30[190]},
      {stage2_30[115]}
   );
   gpc1_1 gpc6671 (
      {stage1_30[191]},
      {stage2_30[116]}
   );
   gpc1_1 gpc6672 (
      {stage1_32[189]},
      {stage2_32[78]}
   );
   gpc1_1 gpc6673 (
      {stage1_32[190]},
      {stage2_32[79]}
   );
   gpc1_1 gpc6674 (
      {stage1_32[191]},
      {stage2_32[80]}
   );
   gpc1_1 gpc6675 (
      {stage1_32[192]},
      {stage2_32[81]}
   );
   gpc1_1 gpc6676 (
      {stage1_32[193]},
      {stage2_32[82]}
   );
   gpc1_1 gpc6677 (
      {stage1_32[194]},
      {stage2_32[83]}
   );
   gpc1_1 gpc6678 (
      {stage1_32[195]},
      {stage2_32[84]}
   );
   gpc1_1 gpc6679 (
      {stage1_32[196]},
      {stage2_32[85]}
   );
   gpc1_1 gpc6680 (
      {stage1_32[197]},
      {stage2_32[86]}
   );
   gpc1_1 gpc6681 (
      {stage1_32[198]},
      {stage2_32[87]}
   );
   gpc1_1 gpc6682 (
      {stage1_32[199]},
      {stage2_32[88]}
   );
   gpc1_1 gpc6683 (
      {stage1_32[200]},
      {stage2_32[89]}
   );
   gpc1_1 gpc6684 (
      {stage1_32[201]},
      {stage2_32[90]}
   );
   gpc1_1 gpc6685 (
      {stage1_32[202]},
      {stage2_32[91]}
   );
   gpc1_1 gpc6686 (
      {stage1_32[203]},
      {stage2_32[92]}
   );
   gpc1_1 gpc6687 (
      {stage1_32[204]},
      {stage2_32[93]}
   );
   gpc1_1 gpc6688 (
      {stage1_32[205]},
      {stage2_32[94]}
   );
   gpc1_1 gpc6689 (
      {stage1_32[206]},
      {stage2_32[95]}
   );
   gpc1_1 gpc6690 (
      {stage1_32[207]},
      {stage2_32[96]}
   );
   gpc1_1 gpc6691 (
      {stage1_32[208]},
      {stage2_32[97]}
   );
   gpc1_1 gpc6692 (
      {stage1_32[209]},
      {stage2_32[98]}
   );
   gpc1_1 gpc6693 (
      {stage1_32[210]},
      {stage2_32[99]}
   );
   gpc1_1 gpc6694 (
      {stage1_32[211]},
      {stage2_32[100]}
   );
   gpc1_1 gpc6695 (
      {stage1_32[212]},
      {stage2_32[101]}
   );
   gpc1_1 gpc6696 (
      {stage1_32[213]},
      {stage2_32[102]}
   );
   gpc1_1 gpc6697 (
      {stage1_32[214]},
      {stage2_32[103]}
   );
   gpc1_1 gpc6698 (
      {stage1_32[215]},
      {stage2_32[104]}
   );
   gpc1_1 gpc6699 (
      {stage1_32[216]},
      {stage2_32[105]}
   );
   gpc1_1 gpc6700 (
      {stage1_34[140]},
      {stage2_34[82]}
   );
   gpc1_1 gpc6701 (
      {stage1_34[141]},
      {stage2_34[83]}
   );
   gpc1_1 gpc6702 (
      {stage1_34[142]},
      {stage2_34[84]}
   );
   gpc1_1 gpc6703 (
      {stage1_34[143]},
      {stage2_34[85]}
   );
   gpc1_1 gpc6704 (
      {stage1_34[144]},
      {stage2_34[86]}
   );
   gpc1_1 gpc6705 (
      {stage1_34[145]},
      {stage2_34[87]}
   );
   gpc1_1 gpc6706 (
      {stage1_34[146]},
      {stage2_34[88]}
   );
   gpc1_1 gpc6707 (
      {stage1_34[147]},
      {stage2_34[89]}
   );
   gpc1_1 gpc6708 (
      {stage1_34[148]},
      {stage2_34[90]}
   );
   gpc1_1 gpc6709 (
      {stage1_34[149]},
      {stage2_34[91]}
   );
   gpc1_1 gpc6710 (
      {stage1_34[150]},
      {stage2_34[92]}
   );
   gpc1_1 gpc6711 (
      {stage1_34[151]},
      {stage2_34[93]}
   );
   gpc1_1 gpc6712 (
      {stage1_34[152]},
      {stage2_34[94]}
   );
   gpc1_1 gpc6713 (
      {stage1_34[153]},
      {stage2_34[95]}
   );
   gpc1_1 gpc6714 (
      {stage1_34[154]},
      {stage2_34[96]}
   );
   gpc1_1 gpc6715 (
      {stage1_34[155]},
      {stage2_34[97]}
   );
   gpc1_1 gpc6716 (
      {stage1_34[156]},
      {stage2_34[98]}
   );
   gpc1_1 gpc6717 (
      {stage1_34[157]},
      {stage2_34[99]}
   );
   gpc1_1 gpc6718 (
      {stage1_34[158]},
      {stage2_34[100]}
   );
   gpc1_1 gpc6719 (
      {stage1_34[159]},
      {stage2_34[101]}
   );
   gpc1_1 gpc6720 (
      {stage1_34[160]},
      {stage2_34[102]}
   );
   gpc1_1 gpc6721 (
      {stage1_34[161]},
      {stage2_34[103]}
   );
   gpc1_1 gpc6722 (
      {stage1_34[162]},
      {stage2_34[104]}
   );
   gpc1_1 gpc6723 (
      {stage1_34[163]},
      {stage2_34[105]}
   );
   gpc1_1 gpc6724 (
      {stage1_34[164]},
      {stage2_34[106]}
   );
   gpc1_1 gpc6725 (
      {stage1_34[165]},
      {stage2_34[107]}
   );
   gpc1_1 gpc6726 (
      {stage1_34[166]},
      {stage2_34[108]}
   );
   gpc1_1 gpc6727 (
      {stage1_34[167]},
      {stage2_34[109]}
   );
   gpc1_1 gpc6728 (
      {stage1_34[168]},
      {stage2_34[110]}
   );
   gpc1_1 gpc6729 (
      {stage1_34[169]},
      {stage2_34[111]}
   );
   gpc1_1 gpc6730 (
      {stage1_34[170]},
      {stage2_34[112]}
   );
   gpc1_1 gpc6731 (
      {stage1_34[171]},
      {stage2_34[113]}
   );
   gpc1_1 gpc6732 (
      {stage1_34[172]},
      {stage2_34[114]}
   );
   gpc1_1 gpc6733 (
      {stage1_34[173]},
      {stage2_34[115]}
   );
   gpc1_1 gpc6734 (
      {stage1_34[174]},
      {stage2_34[116]}
   );
   gpc1_1 gpc6735 (
      {stage1_34[175]},
      {stage2_34[117]}
   );
   gpc1_1 gpc6736 (
      {stage1_34[176]},
      {stage2_34[118]}
   );
   gpc1_1 gpc6737 (
      {stage1_34[177]},
      {stage2_34[119]}
   );
   gpc1_1 gpc6738 (
      {stage1_34[178]},
      {stage2_34[120]}
   );
   gpc1_1 gpc6739 (
      {stage1_34[179]},
      {stage2_34[121]}
   );
   gpc1_1 gpc6740 (
      {stage1_34[180]},
      {stage2_34[122]}
   );
   gpc1_1 gpc6741 (
      {stage1_34[181]},
      {stage2_34[123]}
   );
   gpc1_1 gpc6742 (
      {stage1_34[182]},
      {stage2_34[124]}
   );
   gpc1_1 gpc6743 (
      {stage1_34[183]},
      {stage2_34[125]}
   );
   gpc1_1 gpc6744 (
      {stage1_34[184]},
      {stage2_34[126]}
   );
   gpc1_1 gpc6745 (
      {stage1_34[185]},
      {stage2_34[127]}
   );
   gpc1_1 gpc6746 (
      {stage1_34[186]},
      {stage2_34[128]}
   );
   gpc1_1 gpc6747 (
      {stage1_34[187]},
      {stage2_34[129]}
   );
   gpc1_1 gpc6748 (
      {stage1_34[188]},
      {stage2_34[130]}
   );
   gpc1_1 gpc6749 (
      {stage1_34[189]},
      {stage2_34[131]}
   );
   gpc1_1 gpc6750 (
      {stage1_35[178]},
      {stage2_35[94]}
   );
   gpc1_1 gpc6751 (
      {stage1_35[179]},
      {stage2_35[95]}
   );
   gpc1_1 gpc6752 (
      {stage1_35[180]},
      {stage2_35[96]}
   );
   gpc1_1 gpc6753 (
      {stage1_35[181]},
      {stage2_35[97]}
   );
   gpc1_1 gpc6754 (
      {stage1_35[182]},
      {stage2_35[98]}
   );
   gpc1_1 gpc6755 (
      {stage1_35[183]},
      {stage2_35[99]}
   );
   gpc1_1 gpc6756 (
      {stage1_35[184]},
      {stage2_35[100]}
   );
   gpc1_1 gpc6757 (
      {stage1_35[185]},
      {stage2_35[101]}
   );
   gpc1_1 gpc6758 (
      {stage1_35[186]},
      {stage2_35[102]}
   );
   gpc1_1 gpc6759 (
      {stage1_35[187]},
      {stage2_35[103]}
   );
   gpc1_1 gpc6760 (
      {stage1_35[188]},
      {stage2_35[104]}
   );
   gpc1_1 gpc6761 (
      {stage1_35[189]},
      {stage2_35[105]}
   );
   gpc1_1 gpc6762 (
      {stage1_35[190]},
      {stage2_35[106]}
   );
   gpc1_1 gpc6763 (
      {stage1_35[191]},
      {stage2_35[107]}
   );
   gpc1_1 gpc6764 (
      {stage1_35[192]},
      {stage2_35[108]}
   );
   gpc1_1 gpc6765 (
      {stage1_35[193]},
      {stage2_35[109]}
   );
   gpc1_1 gpc6766 (
      {stage1_35[194]},
      {stage2_35[110]}
   );
   gpc1_1 gpc6767 (
      {stage1_35[195]},
      {stage2_35[111]}
   );
   gpc1_1 gpc6768 (
      {stage1_35[196]},
      {stage2_35[112]}
   );
   gpc1_1 gpc6769 (
      {stage1_35[197]},
      {stage2_35[113]}
   );
   gpc1_1 gpc6770 (
      {stage1_35[198]},
      {stage2_35[114]}
   );
   gpc1_1 gpc6771 (
      {stage1_35[199]},
      {stage2_35[115]}
   );
   gpc1_1 gpc6772 (
      {stage1_35[200]},
      {stage2_35[116]}
   );
   gpc1_1 gpc6773 (
      {stage1_35[201]},
      {stage2_35[117]}
   );
   gpc1_1 gpc6774 (
      {stage1_35[202]},
      {stage2_35[118]}
   );
   gpc1_1 gpc6775 (
      {stage1_35[203]},
      {stage2_35[119]}
   );
   gpc1_1 gpc6776 (
      {stage1_35[204]},
      {stage2_35[120]}
   );
   gpc1_1 gpc6777 (
      {stage1_35[205]},
      {stage2_35[121]}
   );
   gpc1_1 gpc6778 (
      {stage1_35[206]},
      {stage2_35[122]}
   );
   gpc1_1 gpc6779 (
      {stage1_35[207]},
      {stage2_35[123]}
   );
   gpc1_1 gpc6780 (
      {stage1_35[208]},
      {stage2_35[124]}
   );
   gpc1_1 gpc6781 (
      {stage1_35[209]},
      {stage2_35[125]}
   );
   gpc1_1 gpc6782 (
      {stage1_35[210]},
      {stage2_35[126]}
   );
   gpc1_1 gpc6783 (
      {stage1_35[211]},
      {stage2_35[127]}
   );
   gpc1_1 gpc6784 (
      {stage1_35[212]},
      {stage2_35[128]}
   );
   gpc1_1 gpc6785 (
      {stage1_35[213]},
      {stage2_35[129]}
   );
   gpc1_1 gpc6786 (
      {stage1_35[214]},
      {stage2_35[130]}
   );
   gpc1_1 gpc6787 (
      {stage1_35[215]},
      {stage2_35[131]}
   );
   gpc1_1 gpc6788 (
      {stage1_35[216]},
      {stage2_35[132]}
   );
   gpc1_1 gpc6789 (
      {stage1_37[306]},
      {stage2_37[88]}
   );
   gpc1_1 gpc6790 (
      {stage1_37[307]},
      {stage2_37[89]}
   );
   gpc1_1 gpc6791 (
      {stage1_38[231]},
      {stage2_38[106]}
   );
   gpc1_1 gpc6792 (
      {stage1_38[232]},
      {stage2_38[107]}
   );
   gpc1_1 gpc6793 (
      {stage1_38[233]},
      {stage2_38[108]}
   );
   gpc1_1 gpc6794 (
      {stage1_38[234]},
      {stage2_38[109]}
   );
   gpc1_1 gpc6795 (
      {stage1_38[235]},
      {stage2_38[110]}
   );
   gpc1_1 gpc6796 (
      {stage1_38[236]},
      {stage2_38[111]}
   );
   gpc1_1 gpc6797 (
      {stage1_38[237]},
      {stage2_38[112]}
   );
   gpc1_1 gpc6798 (
      {stage1_38[238]},
      {stage2_38[113]}
   );
   gpc1_1 gpc6799 (
      {stage1_38[239]},
      {stage2_38[114]}
   );
   gpc1_1 gpc6800 (
      {stage1_38[240]},
      {stage2_38[115]}
   );
   gpc1_1 gpc6801 (
      {stage1_38[241]},
      {stage2_38[116]}
   );
   gpc1_1 gpc6802 (
      {stage1_38[242]},
      {stage2_38[117]}
   );
   gpc1_1 gpc6803 (
      {stage1_38[243]},
      {stage2_38[118]}
   );
   gpc1_1 gpc6804 (
      {stage1_38[244]},
      {stage2_38[119]}
   );
   gpc1_1 gpc6805 (
      {stage1_38[245]},
      {stage2_38[120]}
   );
   gpc1_1 gpc6806 (
      {stage1_38[246]},
      {stage2_38[121]}
   );
   gpc1_1 gpc6807 (
      {stage1_38[247]},
      {stage2_38[122]}
   );
   gpc1_1 gpc6808 (
      {stage1_38[248]},
      {stage2_38[123]}
   );
   gpc1_1 gpc6809 (
      {stage1_38[249]},
      {stage2_38[124]}
   );
   gpc1_1 gpc6810 (
      {stage1_38[250]},
      {stage2_38[125]}
   );
   gpc1_1 gpc6811 (
      {stage1_38[251]},
      {stage2_38[126]}
   );
   gpc1_1 gpc6812 (
      {stage1_38[252]},
      {stage2_38[127]}
   );
   gpc1_1 gpc6813 (
      {stage1_38[253]},
      {stage2_38[128]}
   );
   gpc1_1 gpc6814 (
      {stage1_38[254]},
      {stage2_38[129]}
   );
   gpc1_1 gpc6815 (
      {stage1_38[255]},
      {stage2_38[130]}
   );
   gpc1_1 gpc6816 (
      {stage1_38[256]},
      {stage2_38[131]}
   );
   gpc1_1 gpc6817 (
      {stage1_38[257]},
      {stage2_38[132]}
   );
   gpc1_1 gpc6818 (
      {stage1_38[258]},
      {stage2_38[133]}
   );
   gpc1_1 gpc6819 (
      {stage1_38[259]},
      {stage2_38[134]}
   );
   gpc1_1 gpc6820 (
      {stage1_38[260]},
      {stage2_38[135]}
   );
   gpc1_1 gpc6821 (
      {stage1_38[261]},
      {stage2_38[136]}
   );
   gpc1_1 gpc6822 (
      {stage1_38[262]},
      {stage2_38[137]}
   );
   gpc1_1 gpc6823 (
      {stage1_38[263]},
      {stage2_38[138]}
   );
   gpc1_1 gpc6824 (
      {stage1_38[264]},
      {stage2_38[139]}
   );
   gpc1_1 gpc6825 (
      {stage1_39[170]},
      {stage2_39[94]}
   );
   gpc1_1 gpc6826 (
      {stage1_39[171]},
      {stage2_39[95]}
   );
   gpc1_1 gpc6827 (
      {stage1_39[172]},
      {stage2_39[96]}
   );
   gpc1_1 gpc6828 (
      {stage1_39[173]},
      {stage2_39[97]}
   );
   gpc1_1 gpc6829 (
      {stage1_39[174]},
      {stage2_39[98]}
   );
   gpc1_1 gpc6830 (
      {stage1_39[175]},
      {stage2_39[99]}
   );
   gpc1_1 gpc6831 (
      {stage1_39[176]},
      {stage2_39[100]}
   );
   gpc1_1 gpc6832 (
      {stage1_39[177]},
      {stage2_39[101]}
   );
   gpc1_1 gpc6833 (
      {stage1_39[178]},
      {stage2_39[102]}
   );
   gpc1_1 gpc6834 (
      {stage1_39[179]},
      {stage2_39[103]}
   );
   gpc1_1 gpc6835 (
      {stage1_39[180]},
      {stage2_39[104]}
   );
   gpc1_1 gpc6836 (
      {stage1_39[181]},
      {stage2_39[105]}
   );
   gpc1_1 gpc6837 (
      {stage1_39[182]},
      {stage2_39[106]}
   );
   gpc1_1 gpc6838 (
      {stage1_39[183]},
      {stage2_39[107]}
   );
   gpc1_1 gpc6839 (
      {stage1_39[184]},
      {stage2_39[108]}
   );
   gpc1_1 gpc6840 (
      {stage1_39[185]},
      {stage2_39[109]}
   );
   gpc1_1 gpc6841 (
      {stage1_39[186]},
      {stage2_39[110]}
   );
   gpc1_1 gpc6842 (
      {stage1_39[187]},
      {stage2_39[111]}
   );
   gpc1_1 gpc6843 (
      {stage1_39[188]},
      {stage2_39[112]}
   );
   gpc1_1 gpc6844 (
      {stage1_39[189]},
      {stage2_39[113]}
   );
   gpc1_1 gpc6845 (
      {stage1_39[190]},
      {stage2_39[114]}
   );
   gpc1_1 gpc6846 (
      {stage1_39[191]},
      {stage2_39[115]}
   );
   gpc1_1 gpc6847 (
      {stage1_39[192]},
      {stage2_39[116]}
   );
   gpc1_1 gpc6848 (
      {stage1_39[193]},
      {stage2_39[117]}
   );
   gpc1_1 gpc6849 (
      {stage1_39[194]},
      {stage2_39[118]}
   );
   gpc1_1 gpc6850 (
      {stage1_39[195]},
      {stage2_39[119]}
   );
   gpc1_1 gpc6851 (
      {stage1_39[196]},
      {stage2_39[120]}
   );
   gpc1_1 gpc6852 (
      {stage1_39[197]},
      {stage2_39[121]}
   );
   gpc1_1 gpc6853 (
      {stage1_39[198]},
      {stage2_39[122]}
   );
   gpc1_1 gpc6854 (
      {stage1_39[199]},
      {stage2_39[123]}
   );
   gpc1_1 gpc6855 (
      {stage1_39[200]},
      {stage2_39[124]}
   );
   gpc1_1 gpc6856 (
      {stage1_39[201]},
      {stage2_39[125]}
   );
   gpc1_1 gpc6857 (
      {stage1_39[202]},
      {stage2_39[126]}
   );
   gpc1_1 gpc6858 (
      {stage1_39[203]},
      {stage2_39[127]}
   );
   gpc1_1 gpc6859 (
      {stage1_39[204]},
      {stage2_39[128]}
   );
   gpc1_1 gpc6860 (
      {stage1_39[205]},
      {stage2_39[129]}
   );
   gpc1_1 gpc6861 (
      {stage1_39[206]},
      {stage2_39[130]}
   );
   gpc1_1 gpc6862 (
      {stage1_39[207]},
      {stage2_39[131]}
   );
   gpc1_1 gpc6863 (
      {stage1_39[208]},
      {stage2_39[132]}
   );
   gpc1_1 gpc6864 (
      {stage1_39[209]},
      {stage2_39[133]}
   );
   gpc1_1 gpc6865 (
      {stage1_39[210]},
      {stage2_39[134]}
   );
   gpc1_1 gpc6866 (
      {stage1_39[211]},
      {stage2_39[135]}
   );
   gpc1_1 gpc6867 (
      {stage1_39[212]},
      {stage2_39[136]}
   );
   gpc1_1 gpc6868 (
      {stage1_40[281]},
      {stage2_40[90]}
   );
   gpc1_1 gpc6869 (
      {stage1_40[282]},
      {stage2_40[91]}
   );
   gpc1_1 gpc6870 (
      {stage1_40[283]},
      {stage2_40[92]}
   );
   gpc1_1 gpc6871 (
      {stage1_40[284]},
      {stage2_40[93]}
   );
   gpc1_1 gpc6872 (
      {stage1_40[285]},
      {stage2_40[94]}
   );
   gpc1_1 gpc6873 (
      {stage1_40[286]},
      {stage2_40[95]}
   );
   gpc1_1 gpc6874 (
      {stage1_40[287]},
      {stage2_40[96]}
   );
   gpc1_1 gpc6875 (
      {stage1_40[288]},
      {stage2_40[97]}
   );
   gpc1_1 gpc6876 (
      {stage1_40[289]},
      {stage2_40[98]}
   );
   gpc1_1 gpc6877 (
      {stage1_40[290]},
      {stage2_40[99]}
   );
   gpc1_1 gpc6878 (
      {stage1_40[291]},
      {stage2_40[100]}
   );
   gpc1_1 gpc6879 (
      {stage1_40[292]},
      {stage2_40[101]}
   );
   gpc1_1 gpc6880 (
      {stage1_40[293]},
      {stage2_40[102]}
   );
   gpc1_1 gpc6881 (
      {stage1_40[294]},
      {stage2_40[103]}
   );
   gpc1_1 gpc6882 (
      {stage1_40[295]},
      {stage2_40[104]}
   );
   gpc1_1 gpc6883 (
      {stage1_40[296]},
      {stage2_40[105]}
   );
   gpc1_1 gpc6884 (
      {stage1_40[297]},
      {stage2_40[106]}
   );
   gpc1_1 gpc6885 (
      {stage1_40[298]},
      {stage2_40[107]}
   );
   gpc1_1 gpc6886 (
      {stage1_40[299]},
      {stage2_40[108]}
   );
   gpc1_1 gpc6887 (
      {stage1_40[300]},
      {stage2_40[109]}
   );
   gpc1_1 gpc6888 (
      {stage1_40[301]},
      {stage2_40[110]}
   );
   gpc1_1 gpc6889 (
      {stage1_40[302]},
      {stage2_40[111]}
   );
   gpc1_1 gpc6890 (
      {stage1_40[303]},
      {stage2_40[112]}
   );
   gpc1_1 gpc6891 (
      {stage1_41[168]},
      {stage2_41[103]}
   );
   gpc1_1 gpc6892 (
      {stage1_41[169]},
      {stage2_41[104]}
   );
   gpc1_1 gpc6893 (
      {stage1_41[170]},
      {stage2_41[105]}
   );
   gpc1_1 gpc6894 (
      {stage1_42[168]},
      {stage2_42[80]}
   );
   gpc1_1 gpc6895 (
      {stage1_42[169]},
      {stage2_42[81]}
   );
   gpc1_1 gpc6896 (
      {stage1_42[170]},
      {stage2_42[82]}
   );
   gpc1_1 gpc6897 (
      {stage1_42[171]},
      {stage2_42[83]}
   );
   gpc1_1 gpc6898 (
      {stage1_42[172]},
      {stage2_42[84]}
   );
   gpc1_1 gpc6899 (
      {stage1_42[173]},
      {stage2_42[85]}
   );
   gpc1_1 gpc6900 (
      {stage1_43[241]},
      {stage2_43[66]}
   );
   gpc1_1 gpc6901 (
      {stage1_43[242]},
      {stage2_43[67]}
   );
   gpc1_1 gpc6902 (
      {stage1_43[243]},
      {stage2_43[68]}
   );
   gpc1_1 gpc6903 (
      {stage1_43[244]},
      {stage2_43[69]}
   );
   gpc1_1 gpc6904 (
      {stage1_43[245]},
      {stage2_43[70]}
   );
   gpc1_1 gpc6905 (
      {stage1_43[246]},
      {stage2_43[71]}
   );
   gpc1_1 gpc6906 (
      {stage1_43[247]},
      {stage2_43[72]}
   );
   gpc1_1 gpc6907 (
      {stage1_43[248]},
      {stage2_43[73]}
   );
   gpc1_1 gpc6908 (
      {stage1_43[249]},
      {stage2_43[74]}
   );
   gpc1_1 gpc6909 (
      {stage1_43[250]},
      {stage2_43[75]}
   );
   gpc1_1 gpc6910 (
      {stage1_43[251]},
      {stage2_43[76]}
   );
   gpc1_1 gpc6911 (
      {stage1_43[252]},
      {stage2_43[77]}
   );
   gpc1_1 gpc6912 (
      {stage1_43[253]},
      {stage2_43[78]}
   );
   gpc1_1 gpc6913 (
      {stage1_44[240]},
      {stage2_44[103]}
   );
   gpc1_1 gpc6914 (
      {stage1_44[241]},
      {stage2_44[104]}
   );
   gpc1_1 gpc6915 (
      {stage1_44[242]},
      {stage2_44[105]}
   );
   gpc1_1 gpc6916 (
      {stage1_44[243]},
      {stage2_44[106]}
   );
   gpc1_1 gpc6917 (
      {stage1_44[244]},
      {stage2_44[107]}
   );
   gpc1_1 gpc6918 (
      {stage1_44[245]},
      {stage2_44[108]}
   );
   gpc1_1 gpc6919 (
      {stage1_44[246]},
      {stage2_44[109]}
   );
   gpc1_1 gpc6920 (
      {stage1_44[247]},
      {stage2_44[110]}
   );
   gpc1_1 gpc6921 (
      {stage1_44[248]},
      {stage2_44[111]}
   );
   gpc1_1 gpc6922 (
      {stage1_44[249]},
      {stage2_44[112]}
   );
   gpc1_1 gpc6923 (
      {stage1_44[250]},
      {stage2_44[113]}
   );
   gpc1_1 gpc6924 (
      {stage1_44[251]},
      {stage2_44[114]}
   );
   gpc1_1 gpc6925 (
      {stage1_44[252]},
      {stage2_44[115]}
   );
   gpc1_1 gpc6926 (
      {stage1_44[253]},
      {stage2_44[116]}
   );
   gpc1_1 gpc6927 (
      {stage1_44[254]},
      {stage2_44[117]}
   );
   gpc1_1 gpc6928 (
      {stage1_44[255]},
      {stage2_44[118]}
   );
   gpc1_1 gpc6929 (
      {stage1_45[199]},
      {stage2_45[105]}
   );
   gpc1_1 gpc6930 (
      {stage1_45[200]},
      {stage2_45[106]}
   );
   gpc1_1 gpc6931 (
      {stage1_45[201]},
      {stage2_45[107]}
   );
   gpc1_1 gpc6932 (
      {stage1_45[202]},
      {stage2_45[108]}
   );
   gpc1_1 gpc6933 (
      {stage1_45[203]},
      {stage2_45[109]}
   );
   gpc1_1 gpc6934 (
      {stage1_45[204]},
      {stage2_45[110]}
   );
   gpc1_1 gpc6935 (
      {stage1_45[205]},
      {stage2_45[111]}
   );
   gpc1_1 gpc6936 (
      {stage1_45[206]},
      {stage2_45[112]}
   );
   gpc1_1 gpc6937 (
      {stage1_45[207]},
      {stage2_45[113]}
   );
   gpc1_1 gpc6938 (
      {stage1_45[208]},
      {stage2_45[114]}
   );
   gpc1_1 gpc6939 (
      {stage1_45[209]},
      {stage2_45[115]}
   );
   gpc1_1 gpc6940 (
      {stage1_45[210]},
      {stage2_45[116]}
   );
   gpc1_1 gpc6941 (
      {stage1_45[211]},
      {stage2_45[117]}
   );
   gpc1_1 gpc6942 (
      {stage1_46[295]},
      {stage2_46[85]}
   );
   gpc1_1 gpc6943 (
      {stage1_46[296]},
      {stage2_46[86]}
   );
   gpc1_1 gpc6944 (
      {stage1_46[297]},
      {stage2_46[87]}
   );
   gpc1_1 gpc6945 (
      {stage1_47[230]},
      {stage2_47[98]}
   );
   gpc1_1 gpc6946 (
      {stage1_47[231]},
      {stage2_47[99]}
   );
   gpc1_1 gpc6947 (
      {stage1_47[232]},
      {stage2_47[100]}
   );
   gpc1_1 gpc6948 (
      {stage1_47[233]},
      {stage2_47[101]}
   );
   gpc1_1 gpc6949 (
      {stage1_47[234]},
      {stage2_47[102]}
   );
   gpc1_1 gpc6950 (
      {stage1_47[235]},
      {stage2_47[103]}
   );
   gpc1_1 gpc6951 (
      {stage1_48[172]},
      {stage2_48[104]}
   );
   gpc1_1 gpc6952 (
      {stage1_48[173]},
      {stage2_48[105]}
   );
   gpc1_1 gpc6953 (
      {stage1_48[174]},
      {stage2_48[106]}
   );
   gpc1_1 gpc6954 (
      {stage1_48[175]},
      {stage2_48[107]}
   );
   gpc1_1 gpc6955 (
      {stage1_48[176]},
      {stage2_48[108]}
   );
   gpc1_1 gpc6956 (
      {stage1_48[177]},
      {stage2_48[109]}
   );
   gpc1_1 gpc6957 (
      {stage1_48[178]},
      {stage2_48[110]}
   );
   gpc1_1 gpc6958 (
      {stage1_48[179]},
      {stage2_48[111]}
   );
   gpc1_1 gpc6959 (
      {stage1_48[180]},
      {stage2_48[112]}
   );
   gpc1_1 gpc6960 (
      {stage1_48[181]},
      {stage2_48[113]}
   );
   gpc1_1 gpc6961 (
      {stage1_48[182]},
      {stage2_48[114]}
   );
   gpc1_1 gpc6962 (
      {stage1_48[183]},
      {stage2_48[115]}
   );
   gpc1_1 gpc6963 (
      {stage1_48[184]},
      {stage2_48[116]}
   );
   gpc1_1 gpc6964 (
      {stage1_48[185]},
      {stage2_48[117]}
   );
   gpc1_1 gpc6965 (
      {stage1_48[186]},
      {stage2_48[118]}
   );
   gpc1_1 gpc6966 (
      {stage1_48[187]},
      {stage2_48[119]}
   );
   gpc1_1 gpc6967 (
      {stage1_48[188]},
      {stage2_48[120]}
   );
   gpc1_1 gpc6968 (
      {stage1_48[189]},
      {stage2_48[121]}
   );
   gpc1_1 gpc6969 (
      {stage1_48[190]},
      {stage2_48[122]}
   );
   gpc1_1 gpc6970 (
      {stage1_48[191]},
      {stage2_48[123]}
   );
   gpc1_1 gpc6971 (
      {stage1_48[192]},
      {stage2_48[124]}
   );
   gpc1_1 gpc6972 (
      {stage1_48[193]},
      {stage2_48[125]}
   );
   gpc1_1 gpc6973 (
      {stage1_48[194]},
      {stage2_48[126]}
   );
   gpc1_1 gpc6974 (
      {stage1_48[195]},
      {stage2_48[127]}
   );
   gpc1_1 gpc6975 (
      {stage1_48[196]},
      {stage2_48[128]}
   );
   gpc1_1 gpc6976 (
      {stage1_48[197]},
      {stage2_48[129]}
   );
   gpc1_1 gpc6977 (
      {stage1_49[154]},
      {stage2_49[77]}
   );
   gpc1_1 gpc6978 (
      {stage1_49[155]},
      {stage2_49[78]}
   );
   gpc1_1 gpc6979 (
      {stage1_49[156]},
      {stage2_49[79]}
   );
   gpc1_1 gpc6980 (
      {stage1_49[157]},
      {stage2_49[80]}
   );
   gpc1_1 gpc6981 (
      {stage1_49[158]},
      {stage2_49[81]}
   );
   gpc1_1 gpc6982 (
      {stage1_49[159]},
      {stage2_49[82]}
   );
   gpc1_1 gpc6983 (
      {stage1_49[160]},
      {stage2_49[83]}
   );
   gpc1_1 gpc6984 (
      {stage1_49[161]},
      {stage2_49[84]}
   );
   gpc1_1 gpc6985 (
      {stage1_49[162]},
      {stage2_49[85]}
   );
   gpc1_1 gpc6986 (
      {stage1_49[163]},
      {stage2_49[86]}
   );
   gpc1_1 gpc6987 (
      {stage1_49[164]},
      {stage2_49[87]}
   );
   gpc1_1 gpc6988 (
      {stage1_49[165]},
      {stage2_49[88]}
   );
   gpc1_1 gpc6989 (
      {stage1_49[166]},
      {stage2_49[89]}
   );
   gpc1_1 gpc6990 (
      {stage1_49[167]},
      {stage2_49[90]}
   );
   gpc1_1 gpc6991 (
      {stage1_49[168]},
      {stage2_49[91]}
   );
   gpc1_1 gpc6992 (
      {stage1_49[169]},
      {stage2_49[92]}
   );
   gpc1_1 gpc6993 (
      {stage1_49[170]},
      {stage2_49[93]}
   );
   gpc1_1 gpc6994 (
      {stage1_49[171]},
      {stage2_49[94]}
   );
   gpc1_1 gpc6995 (
      {stage1_49[172]},
      {stage2_49[95]}
   );
   gpc1_1 gpc6996 (
      {stage1_50[179]},
      {stage2_50[75]}
   );
   gpc1_1 gpc6997 (
      {stage1_50[180]},
      {stage2_50[76]}
   );
   gpc1_1 gpc6998 (
      {stage1_50[181]},
      {stage2_50[77]}
   );
   gpc1_1 gpc6999 (
      {stage1_50[182]},
      {stage2_50[78]}
   );
   gpc1_1 gpc7000 (
      {stage1_50[183]},
      {stage2_50[79]}
   );
   gpc1_1 gpc7001 (
      {stage1_50[184]},
      {stage2_50[80]}
   );
   gpc1_1 gpc7002 (
      {stage1_50[185]},
      {stage2_50[81]}
   );
   gpc1_1 gpc7003 (
      {stage1_50[186]},
      {stage2_50[82]}
   );
   gpc1_1 gpc7004 (
      {stage1_50[187]},
      {stage2_50[83]}
   );
   gpc1_1 gpc7005 (
      {stage1_50[188]},
      {stage2_50[84]}
   );
   gpc1_1 gpc7006 (
      {stage1_50[189]},
      {stage2_50[85]}
   );
   gpc1_1 gpc7007 (
      {stage1_51[266]},
      {stage2_51[79]}
   );
   gpc1_1 gpc7008 (
      {stage1_51[267]},
      {stage2_51[80]}
   );
   gpc1_1 gpc7009 (
      {stage1_51[268]},
      {stage2_51[81]}
   );
   gpc1_1 gpc7010 (
      {stage1_51[269]},
      {stage2_51[82]}
   );
   gpc1_1 gpc7011 (
      {stage1_51[270]},
      {stage2_51[83]}
   );
   gpc1_1 gpc7012 (
      {stage1_51[271]},
      {stage2_51[84]}
   );
   gpc1_1 gpc7013 (
      {stage1_51[272]},
      {stage2_51[85]}
   );
   gpc1_1 gpc7014 (
      {stage1_51[273]},
      {stage2_51[86]}
   );
   gpc1_1 gpc7015 (
      {stage1_51[274]},
      {stage2_51[87]}
   );
   gpc1_1 gpc7016 (
      {stage1_52[187]},
      {stage2_52[93]}
   );
   gpc1_1 gpc7017 (
      {stage1_52[188]},
      {stage2_52[94]}
   );
   gpc1_1 gpc7018 (
      {stage1_52[189]},
      {stage2_52[95]}
   );
   gpc1_1 gpc7019 (
      {stage1_52[190]},
      {stage2_52[96]}
   );
   gpc1_1 gpc7020 (
      {stage1_52[191]},
      {stage2_52[97]}
   );
   gpc1_1 gpc7021 (
      {stage1_52[192]},
      {stage2_52[98]}
   );
   gpc1_1 gpc7022 (
      {stage1_52[193]},
      {stage2_52[99]}
   );
   gpc1_1 gpc7023 (
      {stage1_52[194]},
      {stage2_52[100]}
   );
   gpc1_1 gpc7024 (
      {stage1_52[195]},
      {stage2_52[101]}
   );
   gpc1_1 gpc7025 (
      {stage1_52[196]},
      {stage2_52[102]}
   );
   gpc1_1 gpc7026 (
      {stage1_52[197]},
      {stage2_52[103]}
   );
   gpc1_1 gpc7027 (
      {stage1_52[198]},
      {stage2_52[104]}
   );
   gpc1_1 gpc7028 (
      {stage1_53[130]},
      {stage2_53[76]}
   );
   gpc1_1 gpc7029 (
      {stage1_53[131]},
      {stage2_53[77]}
   );
   gpc1_1 gpc7030 (
      {stage1_53[132]},
      {stage2_53[78]}
   );
   gpc1_1 gpc7031 (
      {stage1_53[133]},
      {stage2_53[79]}
   );
   gpc1_1 gpc7032 (
      {stage1_53[134]},
      {stage2_53[80]}
   );
   gpc1_1 gpc7033 (
      {stage1_53[135]},
      {stage2_53[81]}
   );
   gpc1_1 gpc7034 (
      {stage1_53[136]},
      {stage2_53[82]}
   );
   gpc1_1 gpc7035 (
      {stage1_53[137]},
      {stage2_53[83]}
   );
   gpc1_1 gpc7036 (
      {stage1_53[138]},
      {stage2_53[84]}
   );
   gpc1_1 gpc7037 (
      {stage1_53[139]},
      {stage2_53[85]}
   );
   gpc1_1 gpc7038 (
      {stage1_53[140]},
      {stage2_53[86]}
   );
   gpc1_1 gpc7039 (
      {stage1_53[141]},
      {stage2_53[87]}
   );
   gpc1_1 gpc7040 (
      {stage1_53[142]},
      {stage2_53[88]}
   );
   gpc1_1 gpc7041 (
      {stage1_53[143]},
      {stage2_53[89]}
   );
   gpc1_1 gpc7042 (
      {stage1_53[144]},
      {stage2_53[90]}
   );
   gpc1_1 gpc7043 (
      {stage1_53[145]},
      {stage2_53[91]}
   );
   gpc1_1 gpc7044 (
      {stage1_53[146]},
      {stage2_53[92]}
   );
   gpc1_1 gpc7045 (
      {stage1_53[147]},
      {stage2_53[93]}
   );
   gpc1_1 gpc7046 (
      {stage1_53[148]},
      {stage2_53[94]}
   );
   gpc1_1 gpc7047 (
      {stage1_53[149]},
      {stage2_53[95]}
   );
   gpc1_1 gpc7048 (
      {stage1_53[150]},
      {stage2_53[96]}
   );
   gpc1_1 gpc7049 (
      {stage1_53[151]},
      {stage2_53[97]}
   );
   gpc1_1 gpc7050 (
      {stage1_53[152]},
      {stage2_53[98]}
   );
   gpc1_1 gpc7051 (
      {stage1_53[153]},
      {stage2_53[99]}
   );
   gpc1_1 gpc7052 (
      {stage1_53[154]},
      {stage2_53[100]}
   );
   gpc1_1 gpc7053 (
      {stage1_53[155]},
      {stage2_53[101]}
   );
   gpc1_1 gpc7054 (
      {stage1_53[156]},
      {stage2_53[102]}
   );
   gpc1_1 gpc7055 (
      {stage1_53[157]},
      {stage2_53[103]}
   );
   gpc1_1 gpc7056 (
      {stage1_53[158]},
      {stage2_53[104]}
   );
   gpc1_1 gpc7057 (
      {stage1_53[159]},
      {stage2_53[105]}
   );
   gpc1_1 gpc7058 (
      {stage1_53[160]},
      {stage2_53[106]}
   );
   gpc1_1 gpc7059 (
      {stage1_53[161]},
      {stage2_53[107]}
   );
   gpc1_1 gpc7060 (
      {stage1_53[162]},
      {stage2_53[108]}
   );
   gpc1_1 gpc7061 (
      {stage1_53[163]},
      {stage2_53[109]}
   );
   gpc1_1 gpc7062 (
      {stage1_53[164]},
      {stage2_53[110]}
   );
   gpc1_1 gpc7063 (
      {stage1_53[165]},
      {stage2_53[111]}
   );
   gpc1_1 gpc7064 (
      {stage1_53[166]},
      {stage2_53[112]}
   );
   gpc1_1 gpc7065 (
      {stage1_53[167]},
      {stage2_53[113]}
   );
   gpc1_1 gpc7066 (
      {stage1_53[168]},
      {stage2_53[114]}
   );
   gpc1_1 gpc7067 (
      {stage1_54[203]},
      {stage2_54[72]}
   );
   gpc1_1 gpc7068 (
      {stage1_54[204]},
      {stage2_54[73]}
   );
   gpc1_1 gpc7069 (
      {stage1_54[205]},
      {stage2_54[74]}
   );
   gpc1_1 gpc7070 (
      {stage1_54[206]},
      {stage2_54[75]}
   );
   gpc1_1 gpc7071 (
      {stage1_54[207]},
      {stage2_54[76]}
   );
   gpc1_1 gpc7072 (
      {stage1_54[208]},
      {stage2_54[77]}
   );
   gpc1_1 gpc7073 (
      {stage1_54[209]},
      {stage2_54[78]}
   );
   gpc1_1 gpc7074 (
      {stage1_54[210]},
      {stage2_54[79]}
   );
   gpc1_1 gpc7075 (
      {stage1_54[211]},
      {stage2_54[80]}
   );
   gpc1_1 gpc7076 (
      {stage1_54[212]},
      {stage2_54[81]}
   );
   gpc1_1 gpc7077 (
      {stage1_54[213]},
      {stage2_54[82]}
   );
   gpc1_1 gpc7078 (
      {stage1_54[214]},
      {stage2_54[83]}
   );
   gpc1_1 gpc7079 (
      {stage1_54[215]},
      {stage2_54[84]}
   );
   gpc1_1 gpc7080 (
      {stage1_54[216]},
      {stage2_54[85]}
   );
   gpc1_1 gpc7081 (
      {stage1_54[217]},
      {stage2_54[86]}
   );
   gpc1_1 gpc7082 (
      {stage1_54[218]},
      {stage2_54[87]}
   );
   gpc1_1 gpc7083 (
      {stage1_54[219]},
      {stage2_54[88]}
   );
   gpc1_1 gpc7084 (
      {stage1_54[220]},
      {stage2_54[89]}
   );
   gpc1_1 gpc7085 (
      {stage1_54[221]},
      {stage2_54[90]}
   );
   gpc1_1 gpc7086 (
      {stage1_54[222]},
      {stage2_54[91]}
   );
   gpc1_1 gpc7087 (
      {stage1_54[223]},
      {stage2_54[92]}
   );
   gpc1_1 gpc7088 (
      {stage1_54[224]},
      {stage2_54[93]}
   );
   gpc1_1 gpc7089 (
      {stage1_54[225]},
      {stage2_54[94]}
   );
   gpc1_1 gpc7090 (
      {stage1_54[226]},
      {stage2_54[95]}
   );
   gpc1_1 gpc7091 (
      {stage1_54[227]},
      {stage2_54[96]}
   );
   gpc1_1 gpc7092 (
      {stage1_54[228]},
      {stage2_54[97]}
   );
   gpc1_1 gpc7093 (
      {stage1_54[229]},
      {stage2_54[98]}
   );
   gpc1_1 gpc7094 (
      {stage1_54[230]},
      {stage2_54[99]}
   );
   gpc1_1 gpc7095 (
      {stage1_55[254]},
      {stage2_55[93]}
   );
   gpc1_1 gpc7096 (
      {stage1_55[255]},
      {stage2_55[94]}
   );
   gpc1_1 gpc7097 (
      {stage1_55[256]},
      {stage2_55[95]}
   );
   gpc1_1 gpc7098 (
      {stage1_55[257]},
      {stage2_55[96]}
   );
   gpc1_1 gpc7099 (
      {stage1_55[258]},
      {stage2_55[97]}
   );
   gpc1_1 gpc7100 (
      {stage1_55[259]},
      {stage2_55[98]}
   );
   gpc1_1 gpc7101 (
      {stage1_55[260]},
      {stage2_55[99]}
   );
   gpc1_1 gpc7102 (
      {stage1_55[261]},
      {stage2_55[100]}
   );
   gpc1_1 gpc7103 (
      {stage1_55[262]},
      {stage2_55[101]}
   );
   gpc1_1 gpc7104 (
      {stage1_55[263]},
      {stage2_55[102]}
   );
   gpc1_1 gpc7105 (
      {stage1_55[264]},
      {stage2_55[103]}
   );
   gpc1_1 gpc7106 (
      {stage1_55[265]},
      {stage2_55[104]}
   );
   gpc1_1 gpc7107 (
      {stage1_55[266]},
      {stage2_55[105]}
   );
   gpc1_1 gpc7108 (
      {stage1_56[164]},
      {stage2_56[92]}
   );
   gpc1_1 gpc7109 (
      {stage1_56[165]},
      {stage2_56[93]}
   );
   gpc1_1 gpc7110 (
      {stage1_56[166]},
      {stage2_56[94]}
   );
   gpc1_1 gpc7111 (
      {stage1_56[167]},
      {stage2_56[95]}
   );
   gpc1_1 gpc7112 (
      {stage1_56[168]},
      {stage2_56[96]}
   );
   gpc1_1 gpc7113 (
      {stage1_56[169]},
      {stage2_56[97]}
   );
   gpc1_1 gpc7114 (
      {stage1_56[170]},
      {stage2_56[98]}
   );
   gpc1_1 gpc7115 (
      {stage1_56[171]},
      {stage2_56[99]}
   );
   gpc1_1 gpc7116 (
      {stage1_56[172]},
      {stage2_56[100]}
   );
   gpc1_1 gpc7117 (
      {stage1_56[173]},
      {stage2_56[101]}
   );
   gpc1_1 gpc7118 (
      {stage1_56[174]},
      {stage2_56[102]}
   );
   gpc1_1 gpc7119 (
      {stage1_56[175]},
      {stage2_56[103]}
   );
   gpc1_1 gpc7120 (
      {stage1_56[176]},
      {stage2_56[104]}
   );
   gpc1_1 gpc7121 (
      {stage1_56[177]},
      {stage2_56[105]}
   );
   gpc1_1 gpc7122 (
      {stage1_56[178]},
      {stage2_56[106]}
   );
   gpc1_1 gpc7123 (
      {stage1_56[179]},
      {stage2_56[107]}
   );
   gpc1_1 gpc7124 (
      {stage1_56[180]},
      {stage2_56[108]}
   );
   gpc1_1 gpc7125 (
      {stage1_56[181]},
      {stage2_56[109]}
   );
   gpc1_1 gpc7126 (
      {stage1_56[182]},
      {stage2_56[110]}
   );
   gpc1_1 gpc7127 (
      {stage1_56[183]},
      {stage2_56[111]}
   );
   gpc1_1 gpc7128 (
      {stage1_56[184]},
      {stage2_56[112]}
   );
   gpc1_1 gpc7129 (
      {stage1_56[185]},
      {stage2_56[113]}
   );
   gpc1_1 gpc7130 (
      {stage1_56[186]},
      {stage2_56[114]}
   );
   gpc1_1 gpc7131 (
      {stage1_59[205]},
      {stage2_59[109]}
   );
   gpc1_1 gpc7132 (
      {stage1_60[209]},
      {stage2_60[79]}
   );
   gpc1_1 gpc7133 (
      {stage1_60[210]},
      {stage2_60[80]}
   );
   gpc1_1 gpc7134 (
      {stage1_60[211]},
      {stage2_60[81]}
   );
   gpc1_1 gpc7135 (
      {stage1_60[212]},
      {stage2_60[82]}
   );
   gpc1_1 gpc7136 (
      {stage1_60[213]},
      {stage2_60[83]}
   );
   gpc1_1 gpc7137 (
      {stage1_60[214]},
      {stage2_60[84]}
   );
   gpc1_1 gpc7138 (
      {stage1_62[192]},
      {stage2_62[104]}
   );
   gpc1_1 gpc7139 (
      {stage1_63[303]},
      {stage2_63[94]}
   );
   gpc1_1 gpc7140 (
      {stage1_63[304]},
      {stage2_63[95]}
   );
   gpc1_1 gpc7141 (
      {stage1_63[305]},
      {stage2_63[96]}
   );
   gpc1_1 gpc7142 (
      {stage1_63[306]},
      {stage2_63[97]}
   );
   gpc1_1 gpc7143 (
      {stage1_63[307]},
      {stage2_63[98]}
   );
   gpc1_1 gpc7144 (
      {stage1_64[47]},
      {stage2_64[65]}
   );
   gpc1_1 gpc7145 (
      {stage1_64[48]},
      {stage2_64[66]}
   );
   gpc1_1 gpc7146 (
      {stage1_64[49]},
      {stage2_64[67]}
   );
   gpc1_1 gpc7147 (
      {stage1_64[50]},
      {stage2_64[68]}
   );
   gpc1_1 gpc7148 (
      {stage1_64[51]},
      {stage2_64[69]}
   );
   gpc1_1 gpc7149 (
      {stage1_64[52]},
      {stage2_64[70]}
   );
   gpc1_1 gpc7150 (
      {stage1_64[53]},
      {stage2_64[71]}
   );
   gpc1_1 gpc7151 (
      {stage1_64[54]},
      {stage2_64[72]}
   );
   gpc1_1 gpc7152 (
      {stage1_64[55]},
      {stage2_64[73]}
   );
   gpc1_1 gpc7153 (
      {stage1_64[56]},
      {stage2_64[74]}
   );
   gpc1_1 gpc7154 (
      {stage1_64[57]},
      {stage2_64[75]}
   );
   gpc1_1 gpc7155 (
      {stage1_64[58]},
      {stage2_64[76]}
   );
   gpc1_1 gpc7156 (
      {stage1_64[59]},
      {stage2_64[77]}
   );
   gpc1_1 gpc7157 (
      {stage1_64[60]},
      {stage2_64[78]}
   );
   gpc1_1 gpc7158 (
      {stage1_64[61]},
      {stage2_64[79]}
   );
   gpc1_1 gpc7159 (
      {stage1_64[62]},
      {stage2_64[80]}
   );
   gpc1_1 gpc7160 (
      {stage1_64[63]},
      {stage2_64[81]}
   );
   gpc1_1 gpc7161 (
      {stage1_64[64]},
      {stage2_64[82]}
   );
   gpc1_1 gpc7162 (
      {stage1_64[65]},
      {stage2_64[83]}
   );
   gpc1_1 gpc7163 (
      {stage1_64[66]},
      {stage2_64[84]}
   );
   gpc1_1 gpc7164 (
      {stage1_64[67]},
      {stage2_64[85]}
   );
   gpc1_1 gpc7165 (
      {stage1_64[68]},
      {stage2_64[86]}
   );
   gpc1_1 gpc7166 (
      {stage1_64[69]},
      {stage2_64[87]}
   );
   gpc1_1 gpc7167 (
      {stage1_64[70]},
      {stage2_64[88]}
   );
   gpc1_1 gpc7168 (
      {stage1_64[71]},
      {stage2_64[89]}
   );
   gpc1_1 gpc7169 (
      {stage1_64[72]},
      {stage2_64[90]}
   );
   gpc1_1 gpc7170 (
      {stage1_64[73]},
      {stage2_64[91]}
   );
   gpc1_1 gpc7171 (
      {stage1_64[74]},
      {stage2_64[92]}
   );
   gpc1_1 gpc7172 (
      {stage1_64[75]},
      {stage2_64[93]}
   );
   gpc1_1 gpc7173 (
      {stage1_64[76]},
      {stage2_64[94]}
   );
   gpc1_1 gpc7174 (
      {stage1_64[77]},
      {stage2_64[95]}
   );
   gpc1_1 gpc7175 (
      {stage1_64[78]},
      {stage2_64[96]}
   );
   gpc1_1 gpc7176 (
      {stage1_64[79]},
      {stage2_64[97]}
   );
   gpc1_1 gpc7177 (
      {stage1_64[80]},
      {stage2_64[98]}
   );
   gpc1_1 gpc7178 (
      {stage1_64[81]},
      {stage2_64[99]}
   );
   gpc1_1 gpc7179 (
      {stage1_64[82]},
      {stage2_64[100]}
   );
   gpc1_1 gpc7180 (
      {stage1_64[83]},
      {stage2_64[101]}
   );
   gpc1_1 gpc7181 (
      {stage1_64[84]},
      {stage2_64[102]}
   );
   gpc1_1 gpc7182 (
      {stage1_64[85]},
      {stage2_64[103]}
   );
   gpc1_1 gpc7183 (
      {stage1_64[86]},
      {stage2_64[104]}
   );
   gpc1_1 gpc7184 (
      {stage1_64[87]},
      {stage2_64[105]}
   );
   gpc1_1 gpc7185 (
      {stage1_64[88]},
      {stage2_64[106]}
   );
   gpc1_1 gpc7186 (
      {stage1_64[89]},
      {stage2_64[107]}
   );
   gpc1_1 gpc7187 (
      {stage1_64[90]},
      {stage2_64[108]}
   );
   gpc1_1 gpc7188 (
      {stage1_64[91]},
      {stage2_64[109]}
   );
   gpc1_1 gpc7189 (
      {stage1_64[92]},
      {stage2_64[110]}
   );
   gpc1_1 gpc7190 (
      {stage1_64[93]},
      {stage2_64[111]}
   );
   gpc1_1 gpc7191 (
      {stage1_64[94]},
      {stage2_64[112]}
   );
   gpc1_1 gpc7192 (
      {stage1_64[95]},
      {stage2_64[113]}
   );
   gpc1_1 gpc7193 (
      {stage1_64[96]},
      {stage2_64[114]}
   );
   gpc1_1 gpc7194 (
      {stage1_64[97]},
      {stage2_64[115]}
   );
   gpc1_1 gpc7195 (
      {stage1_64[98]},
      {stage2_64[116]}
   );
   gpc1_1 gpc7196 (
      {stage1_64[99]},
      {stage2_64[117]}
   );
   gpc1_1 gpc7197 (
      {stage1_64[100]},
      {stage2_64[118]}
   );
   gpc1_1 gpc7198 (
      {stage1_64[101]},
      {stage2_64[119]}
   );
   gpc1_1 gpc7199 (
      {stage1_64[102]},
      {stage2_64[120]}
   );
   gpc1_1 gpc7200 (
      {stage1_64[103]},
      {stage2_64[121]}
   );
   gpc1_1 gpc7201 (
      {stage1_64[104]},
      {stage2_64[122]}
   );
   gpc1_1 gpc7202 (
      {stage1_64[105]},
      {stage2_64[123]}
   );
   gpc1_1 gpc7203 (
      {stage1_64[106]},
      {stage2_64[124]}
   );
   gpc1_1 gpc7204 (
      {stage1_64[107]},
      {stage2_64[125]}
   );
   gpc1_1 gpc7205 (
      {stage1_64[108]},
      {stage2_64[126]}
   );
   gpc1_1 gpc7206 (
      {stage1_64[109]},
      {stage2_64[127]}
   );
   gpc1_1 gpc7207 (
      {stage1_64[110]},
      {stage2_64[128]}
   );
   gpc1_1 gpc7208 (
      {stage1_64[111]},
      {stage2_64[129]}
   );
   gpc1_1 gpc7209 (
      {stage1_64[112]},
      {stage2_64[130]}
   );
   gpc1_1 gpc7210 (
      {stage1_64[113]},
      {stage2_64[131]}
   );
   gpc1_1 gpc7211 (
      {stage1_64[114]},
      {stage2_64[132]}
   );
   gpc1_1 gpc7212 (
      {stage1_64[115]},
      {stage2_64[133]}
   );
   gpc1_1 gpc7213 (
      {stage1_64[116]},
      {stage2_64[134]}
   );
   gpc1_1 gpc7214 (
      {stage1_64[117]},
      {stage2_64[135]}
   );
   gpc1_1 gpc7215 (
      {stage1_64[118]},
      {stage2_64[136]}
   );
   gpc1_1 gpc7216 (
      {stage1_64[119]},
      {stage2_64[137]}
   );
   gpc1_1 gpc7217 (
      {stage1_64[120]},
      {stage2_64[138]}
   );
   gpc1_1 gpc7218 (
      {stage1_64[121]},
      {stage2_64[139]}
   );
   gpc1_1 gpc7219 (
      {stage1_64[122]},
      {stage2_64[140]}
   );
   gpc1_1 gpc7220 (
      {stage1_64[123]},
      {stage2_64[141]}
   );
   gpc1_1 gpc7221 (
      {stage1_65[49]},
      {stage2_65[51]}
   );
   gpc1_1 gpc7222 (
      {stage1_65[50]},
      {stage2_65[52]}
   );
   gpc1_1 gpc7223 (
      {stage1_65[51]},
      {stage2_65[53]}
   );
   gpc1_1 gpc7224 (
      {stage1_65[52]},
      {stage2_65[54]}
   );
   gpc1_1 gpc7225 (
      {stage1_65[53]},
      {stage2_65[55]}
   );
   gpc1343_5 gpc7226 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3]},
      {stage2_2[0], stage2_2[1], stage2_2[2]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1343_5 gpc7227 (
      {stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7]},
      {stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1343_5 gpc7228 (
      {stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[6], stage2_2[7], stage2_2[8]},
      {stage2_3[2]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc1343_5 gpc7229 (
      {stage2_0[9], stage2_0[10], stage2_0[11]},
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15]},
      {stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage2_3[3]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc2135_5 gpc7230 (
      {stage2_0[12], stage2_0[13], stage2_0[14], stage2_0[15], stage2_0[16]},
      {stage2_1[16], stage2_1[17], stage2_1[18]},
      {stage2_2[12]},
      {stage2_3[4], stage2_3[5]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc606_5 gpc7231 (
      {stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20], stage2_0[21], stage2_0[22]},
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc606_5 gpc7232 (
      {stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23], stage2_1[24]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[0],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc7233 (
      {stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29], stage2_1[30]},
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17]},
      {stage3_5[1],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc7234 (
      {stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35], stage2_1[36]},
      {stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23]},
      {stage3_5[2],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc615_5 gpc7235 (
      {stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_2[19]},
      {stage2_3[24], stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29]},
      {stage3_5[3],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc606_5 gpc7236 (
      {stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24], stage2_2[25]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[4],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc606_5 gpc7237 (
      {stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29], stage2_2[30], stage2_2[31]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[5],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc615_5 gpc7238 (
      {stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34]},
      {stage2_4[12]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[2],stage3_5[6],stage3_4[12],stage3_3[12]}
   );
   gpc615_5 gpc7239 (
      {stage2_3[35], stage2_3[36], stage2_3[37], stage2_3[38], stage2_3[39]},
      {stage2_4[13]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[3],stage3_5[7],stage3_4[13],stage3_3[13]}
   );
   gpc615_5 gpc7240 (
      {stage2_3[40], stage2_3[41], stage2_3[42], stage2_3[43], stage2_3[44]},
      {stage2_4[14]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[4],stage3_5[8],stage3_4[14],stage3_3[14]}
   );
   gpc615_5 gpc7241 (
      {stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48], stage2_3[49]},
      {stage2_4[15]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[5],stage3_5[9],stage3_4[15],stage3_3[15]}
   );
   gpc615_5 gpc7242 (
      {stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53], stage2_3[54]},
      {stage2_4[16]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[6],stage3_5[10],stage3_4[16],stage3_3[16]}
   );
   gpc615_5 gpc7243 (
      {stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58], stage2_3[59]},
      {stage2_4[17]},
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage3_7[5],stage3_6[7],stage3_5[11],stage3_4[17],stage3_3[17]}
   );
   gpc615_5 gpc7244 (
      {stage2_3[60], stage2_3[61], stage2_3[62], stage2_3[63], stage2_3[64]},
      {stage2_4[18]},
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage3_7[6],stage3_6[8],stage3_5[12],stage3_4[18],stage3_3[18]}
   );
   gpc615_5 gpc7245 (
      {stage2_3[65], stage2_3[66], stage2_3[67], stage2_3[68], stage2_3[69]},
      {stage2_4[19]},
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage3_7[7],stage3_6[9],stage3_5[13],stage3_4[19],stage3_3[19]}
   );
   gpc615_5 gpc7246 (
      {stage2_3[70], stage2_3[71], stage2_3[72], stage2_3[73], stage2_3[74]},
      {stage2_4[20]},
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage3_7[8],stage3_6[10],stage3_5[14],stage3_4[20],stage3_3[20]}
   );
   gpc615_5 gpc7247 (
      {stage2_3[75], stage2_3[76], stage2_3[77], stage2_3[78], stage2_3[79]},
      {stage2_4[21]},
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage3_7[9],stage3_6[11],stage3_5[15],stage3_4[21],stage3_3[21]}
   );
   gpc615_5 gpc7248 (
      {stage2_3[80], stage2_3[81], stage2_3[82], stage2_3[83], stage2_3[84]},
      {stage2_4[22]},
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64], stage2_5[65]},
      {stage3_7[10],stage3_6[12],stage3_5[16],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc7249 (
      {stage2_3[85], stage2_3[86], stage2_3[87], stage2_3[88], stage2_3[89]},
      {stage2_4[23]},
      {stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70], stage2_5[71]},
      {stage3_7[11],stage3_6[13],stage3_5[17],stage3_4[23],stage3_3[23]}
   );
   gpc615_5 gpc7250 (
      {stage2_3[90], stage2_3[91], stage2_3[92], stage2_3[93], stage2_3[94]},
      {stage2_4[24]},
      {stage2_5[72], stage2_5[73], stage2_5[74], stage2_5[75], stage2_5[76], stage2_5[77]},
      {stage3_7[12],stage3_6[14],stage3_5[18],stage3_4[24],stage3_3[24]}
   );
   gpc615_5 gpc7251 (
      {stage2_3[95], stage2_3[96], stage2_3[97], stage2_3[98], stage2_3[99]},
      {stage2_4[25]},
      {stage2_5[78], stage2_5[79], stage2_5[80], stage2_5[81], stage2_5[82], stage2_5[83]},
      {stage3_7[13],stage3_6[15],stage3_5[19],stage3_4[25],stage3_3[25]}
   );
   gpc615_5 gpc7252 (
      {stage2_3[100], stage2_3[101], stage2_3[102], stage2_3[103], stage2_3[104]},
      {stage2_4[26]},
      {stage2_5[84], stage2_5[85], stage2_5[86], stage2_5[87], stage2_5[88], stage2_5[89]},
      {stage3_7[14],stage3_6[16],stage3_5[20],stage3_4[26],stage3_3[26]}
   );
   gpc615_5 gpc7253 (
      {stage2_3[105], stage2_3[106], stage2_3[107], stage2_3[108], stage2_3[109]},
      {stage2_4[27]},
      {stage2_5[90], stage2_5[91], stage2_5[92], stage2_5[93], stage2_5[94], stage2_5[95]},
      {stage3_7[15],stage3_6[17],stage3_5[21],stage3_4[27],stage3_3[27]}
   );
   gpc615_5 gpc7254 (
      {stage2_3[110], stage2_3[111], stage2_3[112], stage2_3[113], 1'b0},
      {stage2_4[28]},
      {stage2_5[96], stage2_5[97], stage2_5[98], stage2_5[99], stage2_5[100], stage2_5[101]},
      {stage3_7[16],stage3_6[18],stage3_5[22],stage3_4[28],stage3_3[28]}
   );
   gpc606_5 gpc7255 (
      {stage2_5[102], stage2_5[103], stage2_5[104], stage2_5[105], stage2_5[106], stage2_5[107]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[0],stage3_7[17],stage3_6[19],stage3_5[23]}
   );
   gpc606_5 gpc7256 (
      {stage2_5[108], stage2_5[109], stage2_5[110], stage2_5[111], stage2_5[112], stage2_5[113]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[1],stage3_7[18],stage3_6[20],stage3_5[24]}
   );
   gpc606_5 gpc7257 (
      {stage2_5[114], stage2_5[115], stage2_5[116], stage2_5[117], stage2_5[118], stage2_5[119]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[2],stage3_7[19],stage3_6[21],stage3_5[25]}
   );
   gpc606_5 gpc7258 (
      {stage2_5[120], stage2_5[121], stage2_5[122], stage2_5[123], stage2_5[124], stage2_5[125]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[3],stage3_7[20],stage3_6[22],stage3_5[26]}
   );
   gpc606_5 gpc7259 (
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[4],stage3_8[4],stage3_7[21],stage3_6[23]}
   );
   gpc615_5 gpc7260 (
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10]},
      {stage2_7[24]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[5],stage3_8[5],stage3_7[22],stage3_6[24]}
   );
   gpc615_5 gpc7261 (
      {stage2_6[11], stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15]},
      {stage2_7[25]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[6],stage3_8[6],stage3_7[23],stage3_6[25]}
   );
   gpc615_5 gpc7262 (
      {stage2_6[16], stage2_6[17], stage2_6[18], stage2_6[19], stage2_6[20]},
      {stage2_7[26]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[7],stage3_8[7],stage3_7[24],stage3_6[26]}
   );
   gpc615_5 gpc7263 (
      {stage2_6[21], stage2_6[22], stage2_6[23], stage2_6[24], stage2_6[25]},
      {stage2_7[27]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[8],stage3_8[8],stage3_7[25],stage3_6[27]}
   );
   gpc615_5 gpc7264 (
      {stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29], stage2_6[30]},
      {stage2_7[28]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[9],stage3_8[9],stage3_7[26],stage3_6[28]}
   );
   gpc615_5 gpc7265 (
      {stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage2_7[29]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[10],stage3_8[10],stage3_7[27],stage3_6[29]}
   );
   gpc615_5 gpc7266 (
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40]},
      {stage2_7[30]},
      {stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage3_10[7],stage3_9[11],stage3_8[11],stage3_7[28],stage3_6[30]}
   );
   gpc615_5 gpc7267 (
      {stage2_6[41], stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45]},
      {stage2_7[31]},
      {stage2_8[48], stage2_8[49], stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53]},
      {stage3_10[8],stage3_9[12],stage3_8[12],stage3_7[29],stage3_6[31]}
   );
   gpc615_5 gpc7268 (
      {stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_8[54]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[9],stage3_9[13],stage3_8[13],stage3_7[30]}
   );
   gpc615_5 gpc7269 (
      {stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage2_8[55]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[10],stage3_9[14],stage3_8[14],stage3_7[31]}
   );
   gpc615_5 gpc7270 (
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46]},
      {stage2_8[56]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[11],stage3_9[15],stage3_8[15],stage3_7[32]}
   );
   gpc615_5 gpc7271 (
      {stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51]},
      {stage2_8[57]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[12],stage3_9[16],stage3_8[16],stage3_7[33]}
   );
   gpc615_5 gpc7272 (
      {stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56]},
      {stage2_8[58]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[13],stage3_9[17],stage3_8[17],stage3_7[34]}
   );
   gpc606_5 gpc7273 (
      {stage2_8[59], stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63], stage2_8[64]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[5],stage3_10[14],stage3_9[18],stage3_8[18]}
   );
   gpc606_5 gpc7274 (
      {stage2_8[65], stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[6],stage3_10[15],stage3_9[19],stage3_8[19]}
   );
   gpc606_5 gpc7275 (
      {stage2_8[71], stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75], stage2_8[76]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[7],stage3_10[16],stage3_9[20],stage3_8[20]}
   );
   gpc606_5 gpc7276 (
      {stage2_8[77], stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81], stage2_8[82]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[8],stage3_10[17],stage3_9[21],stage3_8[21]}
   );
   gpc606_5 gpc7277 (
      {stage2_8[83], stage2_8[84], stage2_8[85], stage2_8[86], stage2_8[87], stage2_8[88]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[9],stage3_10[18],stage3_9[22],stage3_8[22]}
   );
   gpc606_5 gpc7278 (
      {stage2_8[89], stage2_8[90], stage2_8[91], stage2_8[92], stage2_8[93], stage2_8[94]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[10],stage3_10[19],stage3_9[23],stage3_8[23]}
   );
   gpc606_5 gpc7279 (
      {stage2_8[95], stage2_8[96], stage2_8[97], stage2_8[98], stage2_8[99], stage2_8[100]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[6],stage3_11[11],stage3_10[20],stage3_9[24],stage3_8[24]}
   );
   gpc606_5 gpc7280 (
      {stage2_8[101], stage2_8[102], stage2_8[103], stage2_8[104], stage2_8[105], stage2_8[106]},
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage3_12[7],stage3_11[12],stage3_10[21],stage3_9[25],stage3_8[25]}
   );
   gpc606_5 gpc7281 (
      {stage2_8[107], stage2_8[108], stage2_8[109], stage2_8[110], stage2_8[111], stage2_8[112]},
      {stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53]},
      {stage3_12[8],stage3_11[13],stage3_10[22],stage3_9[26],stage3_8[26]}
   );
   gpc606_5 gpc7282 (
      {stage2_8[113], stage2_8[114], stage2_8[115], stage2_8[116], stage2_8[117], stage2_8[118]},
      {stage2_10[54], stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59]},
      {stage3_12[9],stage3_11[14],stage3_10[23],stage3_9[27],stage3_8[27]}
   );
   gpc606_5 gpc7283 (
      {stage2_8[119], stage2_8[120], stage2_8[121], stage2_8[122], stage2_8[123], stage2_8[124]},
      {stage2_10[60], stage2_10[61], stage2_10[62], stage2_10[63], stage2_10[64], stage2_10[65]},
      {stage3_12[10],stage3_11[15],stage3_10[24],stage3_9[28],stage3_8[28]}
   );
   gpc606_5 gpc7284 (
      {stage2_8[125], stage2_8[126], stage2_8[127], stage2_8[128], stage2_8[129], stage2_8[130]},
      {stage2_10[66], stage2_10[67], stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71]},
      {stage3_12[11],stage3_11[16],stage3_10[25],stage3_9[29],stage3_8[29]}
   );
   gpc606_5 gpc7285 (
      {stage2_8[131], stage2_8[132], stage2_8[133], stage2_8[134], stage2_8[135], stage2_8[136]},
      {stage2_10[72], stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76], stage2_10[77]},
      {stage3_12[12],stage3_11[17],stage3_10[26],stage3_9[30],stage3_8[30]}
   );
   gpc606_5 gpc7286 (
      {stage2_8[137], stage2_8[138], stage2_8[139], stage2_8[140], stage2_8[141], stage2_8[142]},
      {stage2_10[78], stage2_10[79], stage2_10[80], stage2_10[81], stage2_10[82], stage2_10[83]},
      {stage3_12[13],stage3_11[18],stage3_10[27],stage3_9[31],stage3_8[31]}
   );
   gpc606_5 gpc7287 (
      {stage2_8[143], stage2_8[144], stage2_8[145], stage2_8[146], stage2_8[147], stage2_8[148]},
      {stage2_10[84], stage2_10[85], stage2_10[86], stage2_10[87], stage2_10[88], stage2_10[89]},
      {stage3_12[14],stage3_11[19],stage3_10[28],stage3_9[32],stage3_8[32]}
   );
   gpc606_5 gpc7288 (
      {stage2_8[149], stage2_8[150], stage2_8[151], stage2_8[152], stage2_8[153], stage2_8[154]},
      {stage2_10[90], stage2_10[91], stage2_10[92], stage2_10[93], stage2_10[94], stage2_10[95]},
      {stage3_12[15],stage3_11[20],stage3_10[29],stage3_9[33],stage3_8[33]}
   );
   gpc606_5 gpc7289 (
      {stage2_8[155], stage2_8[156], stage2_8[157], stage2_8[158], stage2_8[159], 1'b0},
      {stage2_10[96], stage2_10[97], stage2_10[98], stage2_10[99], stage2_10[100], stage2_10[101]},
      {stage3_12[16],stage3_11[21],stage3_10[30],stage3_9[34],stage3_8[34]}
   );
   gpc606_5 gpc7290 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[17],stage3_11[22],stage3_10[31],stage3_9[35]}
   );
   gpc606_5 gpc7291 (
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[18],stage3_11[23],stage3_10[32],stage3_9[36]}
   );
   gpc606_5 gpc7292 (
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[19],stage3_11[24],stage3_10[33],stage3_9[37]}
   );
   gpc606_5 gpc7293 (
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[20],stage3_11[25],stage3_10[34],stage3_9[38]}
   );
   gpc606_5 gpc7294 (
      {stage2_9[54], stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage3_13[4],stage3_12[21],stage3_11[26],stage3_10[35],stage3_9[39]}
   );
   gpc606_5 gpc7295 (
      {stage2_9[60], stage2_9[61], stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35]},
      {stage3_13[5],stage3_12[22],stage3_11[27],stage3_10[36],stage3_9[40]}
   );
   gpc606_5 gpc7296 (
      {stage2_9[66], stage2_9[67], stage2_9[68], stage2_9[69], stage2_9[70], stage2_9[71]},
      {stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41]},
      {stage3_13[6],stage3_12[23],stage3_11[28],stage3_10[37],stage3_9[41]}
   );
   gpc606_5 gpc7297 (
      {stage2_9[72], stage2_9[73], stage2_9[74], stage2_9[75], stage2_9[76], stage2_9[77]},
      {stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47]},
      {stage3_13[7],stage3_12[24],stage3_11[29],stage3_10[38],stage3_9[42]}
   );
   gpc606_5 gpc7298 (
      {stage2_9[78], stage2_9[79], stage2_9[80], stage2_9[81], stage2_9[82], stage2_9[83]},
      {stage2_11[48], stage2_11[49], stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53]},
      {stage3_13[8],stage3_12[25],stage3_11[30],stage3_10[39],stage3_9[43]}
   );
   gpc606_5 gpc7299 (
      {stage2_9[84], stage2_9[85], stage2_9[86], stage2_9[87], stage2_9[88], stage2_9[89]},
      {stage2_11[54], stage2_11[55], stage2_11[56], stage2_11[57], stage2_11[58], stage2_11[59]},
      {stage3_13[9],stage3_12[26],stage3_11[31],stage3_10[40],stage3_9[44]}
   );
   gpc606_5 gpc7300 (
      {stage2_9[90], stage2_9[91], stage2_9[92], stage2_9[93], stage2_9[94], stage2_9[95]},
      {stage2_11[60], stage2_11[61], stage2_11[62], stage2_11[63], stage2_11[64], stage2_11[65]},
      {stage3_13[10],stage3_12[27],stage3_11[32],stage3_10[41],stage3_9[45]}
   );
   gpc606_5 gpc7301 (
      {stage2_9[96], stage2_9[97], stage2_9[98], stage2_9[99], stage2_9[100], stage2_9[101]},
      {stage2_11[66], stage2_11[67], stage2_11[68], stage2_11[69], stage2_11[70], stage2_11[71]},
      {stage3_13[11],stage3_12[28],stage3_11[33],stage3_10[42],stage3_9[46]}
   );
   gpc606_5 gpc7302 (
      {stage2_9[102], stage2_9[103], stage2_9[104], stage2_9[105], stage2_9[106], stage2_9[107]},
      {stage2_11[72], stage2_11[73], stage2_11[74], stage2_11[75], stage2_11[76], stage2_11[77]},
      {stage3_13[12],stage3_12[29],stage3_11[34],stage3_10[43],stage3_9[47]}
   );
   gpc606_5 gpc7303 (
      {stage2_9[108], stage2_9[109], stage2_9[110], stage2_9[111], stage2_9[112], stage2_9[113]},
      {stage2_11[78], stage2_11[79], stage2_11[80], stage2_11[81], stage2_11[82], stage2_11[83]},
      {stage3_13[13],stage3_12[30],stage3_11[35],stage3_10[44],stage3_9[48]}
   );
   gpc606_5 gpc7304 (
      {stage2_9[114], stage2_9[115], stage2_9[116], stage2_9[117], stage2_9[118], stage2_9[119]},
      {stage2_11[84], stage2_11[85], stage2_11[86], stage2_11[87], stage2_11[88], stage2_11[89]},
      {stage3_13[14],stage3_12[31],stage3_11[36],stage3_10[45],stage3_9[49]}
   );
   gpc606_5 gpc7305 (
      {stage2_9[120], stage2_9[121], stage2_9[122], stage2_9[123], stage2_9[124], stage2_9[125]},
      {stage2_11[90], stage2_11[91], stage2_11[92], stage2_11[93], stage2_11[94], stage2_11[95]},
      {stage3_13[15],stage3_12[32],stage3_11[37],stage3_10[46],stage3_9[50]}
   );
   gpc606_5 gpc7306 (
      {stage2_9[126], stage2_9[127], stage2_9[128], stage2_9[129], stage2_9[130], stage2_9[131]},
      {stage2_11[96], stage2_11[97], stage2_11[98], stage2_11[99], stage2_11[100], stage2_11[101]},
      {stage3_13[16],stage3_12[33],stage3_11[38],stage3_10[47],stage3_9[51]}
   );
   gpc606_5 gpc7307 (
      {stage2_9[132], stage2_9[133], stage2_9[134], stage2_9[135], stage2_9[136], stage2_9[137]},
      {stage2_11[102], stage2_11[103], stage2_11[104], stage2_11[105], stage2_11[106], stage2_11[107]},
      {stage3_13[17],stage3_12[34],stage3_11[39],stage3_10[48],stage3_9[52]}
   );
   gpc606_5 gpc7308 (
      {stage2_9[138], stage2_9[139], stage2_9[140], stage2_9[141], stage2_9[142], 1'b0},
      {stage2_11[108], stage2_11[109], stage2_11[110], stage2_11[111], stage2_11[112], stage2_11[113]},
      {stage3_13[18],stage3_12[35],stage3_11[40],stage3_10[49],stage3_9[53]}
   );
   gpc615_5 gpc7309 (
      {stage2_10[102], stage2_10[103], stage2_10[104], stage2_10[105], stage2_10[106]},
      {stage2_11[114]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[19],stage3_12[36],stage3_11[41],stage3_10[50]}
   );
   gpc615_5 gpc7310 (
      {stage2_10[107], stage2_10[108], stage2_10[109], stage2_10[110], stage2_10[111]},
      {stage2_11[115]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[20],stage3_12[37],stage3_11[42],stage3_10[51]}
   );
   gpc615_5 gpc7311 (
      {stage2_10[112], stage2_10[113], stage2_10[114], stage2_10[115], stage2_10[116]},
      {stage2_11[116]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[21],stage3_12[38],stage3_11[43],stage3_10[52]}
   );
   gpc615_5 gpc7312 (
      {stage2_11[117], stage2_11[118], stage2_11[119], stage2_11[120], stage2_11[121]},
      {stage2_12[18]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[3],stage3_13[22],stage3_12[39],stage3_11[44]}
   );
   gpc615_5 gpc7313 (
      {stage2_11[122], stage2_11[123], stage2_11[124], stage2_11[125], stage2_11[126]},
      {stage2_12[19]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[4],stage3_13[23],stage3_12[40],stage3_11[45]}
   );
   gpc606_5 gpc7314 (
      {stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[2],stage3_14[5],stage3_13[24],stage3_12[41]}
   );
   gpc606_5 gpc7315 (
      {stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29], stage2_12[30], stage2_12[31]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[3],stage3_14[6],stage3_13[25],stage3_12[42]}
   );
   gpc606_5 gpc7316 (
      {stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35], stage2_12[36], stage2_12[37]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[4],stage3_14[7],stage3_13[26],stage3_12[43]}
   );
   gpc606_5 gpc7317 (
      {stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41], stage2_12[42], stage2_12[43]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[5],stage3_14[8],stage3_13[27],stage3_12[44]}
   );
   gpc606_5 gpc7318 (
      {stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47], stage2_12[48], stage2_12[49]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[6],stage3_14[9],stage3_13[28],stage3_12[45]}
   );
   gpc606_5 gpc7319 (
      {stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53], stage2_12[54], stage2_12[55]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[7],stage3_14[10],stage3_13[29],stage3_12[46]}
   );
   gpc606_5 gpc7320 (
      {stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59], stage2_12[60], stage2_12[61]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[8],stage3_14[11],stage3_13[30],stage3_12[47]}
   );
   gpc606_5 gpc7321 (
      {stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65], stage2_12[66], stage2_12[67]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[9],stage3_14[12],stage3_13[31],stage3_12[48]}
   );
   gpc606_5 gpc7322 (
      {stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71], stage2_12[72], stage2_12[73]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[10],stage3_14[13],stage3_13[32],stage3_12[49]}
   );
   gpc606_5 gpc7323 (
      {stage2_12[74], stage2_12[75], stage2_12[76], stage2_12[77], stage2_12[78], stage2_12[79]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[11],stage3_14[14],stage3_13[33],stage3_12[50]}
   );
   gpc606_5 gpc7324 (
      {stage2_12[80], stage2_12[81], stage2_12[82], stage2_12[83], stage2_12[84], stage2_12[85]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[12],stage3_14[15],stage3_13[34],stage3_12[51]}
   );
   gpc606_5 gpc7325 (
      {stage2_12[86], stage2_12[87], stage2_12[88], stage2_12[89], stage2_12[90], stage2_12[91]},
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage3_16[11],stage3_15[13],stage3_14[16],stage3_13[35],stage3_12[52]}
   );
   gpc606_5 gpc7326 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[12],stage3_15[14],stage3_14[17],stage3_13[36]}
   );
   gpc606_5 gpc7327 (
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[13],stage3_15[15],stage3_14[18],stage3_13[37]}
   );
   gpc606_5 gpc7328 (
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[14],stage3_15[16],stage3_14[19],stage3_13[38]}
   );
   gpc606_5 gpc7329 (
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[15],stage3_15[17],stage3_14[20],stage3_13[39]}
   );
   gpc606_5 gpc7330 (
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[16],stage3_15[18],stage3_14[21],stage3_13[40]}
   );
   gpc606_5 gpc7331 (
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34], stage2_15[35]},
      {stage3_17[5],stage3_16[17],stage3_15[19],stage3_14[22],stage3_13[41]}
   );
   gpc606_5 gpc7332 (
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage2_15[36], stage2_15[37], stage2_15[38], stage2_15[39], stage2_15[40], stage2_15[41]},
      {stage3_17[6],stage3_16[18],stage3_15[20],stage3_14[23],stage3_13[42]}
   );
   gpc606_5 gpc7333 (
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage2_15[42], stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46], stage2_15[47]},
      {stage3_17[7],stage3_16[19],stage3_15[21],stage3_14[24],stage3_13[43]}
   );
   gpc606_5 gpc7334 (
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage2_15[48], stage2_15[49], stage2_15[50], stage2_15[51], stage2_15[52], stage2_15[53]},
      {stage3_17[8],stage3_16[20],stage3_15[22],stage3_14[25],stage3_13[44]}
   );
   gpc606_5 gpc7335 (
      {stage2_14[72], stage2_14[73], stage2_14[74], stage2_14[75], stage2_14[76], stage2_14[77]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[9],stage3_16[21],stage3_15[23],stage3_14[26]}
   );
   gpc606_5 gpc7336 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82], stage2_14[83]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[10],stage3_16[22],stage3_15[24],stage3_14[27]}
   );
   gpc606_5 gpc7337 (
      {stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87], stage2_14[88], stage2_14[89]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[11],stage3_16[23],stage3_15[25],stage3_14[28]}
   );
   gpc606_5 gpc7338 (
      {stage2_14[90], stage2_14[91], stage2_14[92], stage2_14[93], stage2_14[94], stage2_14[95]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[12],stage3_16[24],stage3_15[26],stage3_14[29]}
   );
   gpc606_5 gpc7339 (
      {stage2_14[96], stage2_14[97], stage2_14[98], stage2_14[99], stage2_14[100], stage2_14[101]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[13],stage3_16[25],stage3_15[27],stage3_14[30]}
   );
   gpc606_5 gpc7340 (
      {stage2_14[102], stage2_14[103], stage2_14[104], stage2_14[105], stage2_14[106], stage2_14[107]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[14],stage3_16[26],stage3_15[28],stage3_14[31]}
   );
   gpc207_4 gpc7341 (
      {stage2_15[54], stage2_15[55], stage2_15[56], stage2_15[57], stage2_15[58], stage2_15[59], stage2_15[60]},
      {stage2_17[0], stage2_17[1]},
      {stage3_18[6],stage3_17[15],stage3_16[27],stage3_15[29]}
   );
   gpc207_4 gpc7342 (
      {stage2_15[61], stage2_15[62], stage2_15[63], stage2_15[64], stage2_15[65], stage2_15[66], stage2_15[67]},
      {stage2_17[2], stage2_17[3]},
      {stage3_18[7],stage3_17[16],stage3_16[28],stage3_15[30]}
   );
   gpc615_5 gpc7343 (
      {stage2_15[68], stage2_15[69], stage2_15[70], stage2_15[71], stage2_15[72]},
      {stage2_16[36]},
      {stage2_17[4], stage2_17[5], stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9]},
      {stage3_19[0],stage3_18[8],stage3_17[17],stage3_16[29],stage3_15[31]}
   );
   gpc615_5 gpc7344 (
      {stage2_15[73], stage2_15[74], stage2_15[75], stage2_15[76], stage2_15[77]},
      {stage2_16[37]},
      {stage2_17[10], stage2_17[11], stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15]},
      {stage3_19[1],stage3_18[9],stage3_17[18],stage3_16[30],stage3_15[32]}
   );
   gpc615_5 gpc7345 (
      {stage2_15[78], stage2_15[79], stage2_15[80], stage2_15[81], stage2_15[82]},
      {stage2_16[38]},
      {stage2_17[16], stage2_17[17], stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21]},
      {stage3_19[2],stage3_18[10],stage3_17[19],stage3_16[31],stage3_15[33]}
   );
   gpc615_5 gpc7346 (
      {stage2_15[83], stage2_15[84], stage2_15[85], stage2_15[86], stage2_15[87]},
      {stage2_16[39]},
      {stage2_17[22], stage2_17[23], stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27]},
      {stage3_19[3],stage3_18[11],stage3_17[20],stage3_16[32],stage3_15[34]}
   );
   gpc615_5 gpc7347 (
      {stage2_15[88], stage2_15[89], stage2_15[90], stage2_15[91], stage2_15[92]},
      {stage2_16[40]},
      {stage2_17[28], stage2_17[29], stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33]},
      {stage3_19[4],stage3_18[12],stage3_17[21],stage3_16[33],stage3_15[35]}
   );
   gpc615_5 gpc7348 (
      {stage2_15[93], stage2_15[94], stage2_15[95], stage2_15[96], stage2_15[97]},
      {stage2_16[41]},
      {stage2_17[34], stage2_17[35], stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39]},
      {stage3_19[5],stage3_18[13],stage3_17[22],stage3_16[34],stage3_15[36]}
   );
   gpc615_5 gpc7349 (
      {stage2_15[98], stage2_15[99], stage2_15[100], stage2_15[101], stage2_15[102]},
      {stage2_16[42]},
      {stage2_17[40], stage2_17[41], stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45]},
      {stage3_19[6],stage3_18[14],stage3_17[23],stage3_16[35],stage3_15[37]}
   );
   gpc615_5 gpc7350 (
      {stage2_15[103], stage2_15[104], stage2_15[105], stage2_15[106], stage2_15[107]},
      {stage2_16[43]},
      {stage2_17[46], stage2_17[47], stage2_17[48], stage2_17[49], stage2_17[50], stage2_17[51]},
      {stage3_19[7],stage3_18[15],stage3_17[24],stage3_16[36],stage3_15[38]}
   );
   gpc615_5 gpc7351 (
      {stage2_15[108], stage2_15[109], stage2_15[110], stage2_15[111], stage2_15[112]},
      {stage2_16[44]},
      {stage2_17[52], stage2_17[53], stage2_17[54], stage2_17[55], stage2_17[56], stage2_17[57]},
      {stage3_19[8],stage3_18[16],stage3_17[25],stage3_16[37],stage3_15[39]}
   );
   gpc615_5 gpc7352 (
      {stage2_15[113], stage2_15[114], stage2_15[115], stage2_15[116], stage2_15[117]},
      {stage2_16[45]},
      {stage2_17[58], stage2_17[59], stage2_17[60], stage2_17[61], stage2_17[62], stage2_17[63]},
      {stage3_19[9],stage3_18[17],stage3_17[26],stage3_16[38],stage3_15[40]}
   );
   gpc615_5 gpc7353 (
      {stage2_15[118], stage2_15[119], stage2_15[120], stage2_15[121], stage2_15[122]},
      {stage2_16[46]},
      {stage2_17[64], stage2_17[65], stage2_17[66], stage2_17[67], stage2_17[68], stage2_17[69]},
      {stage3_19[10],stage3_18[18],stage3_17[27],stage3_16[39],stage3_15[41]}
   );
   gpc615_5 gpc7354 (
      {stage2_15[123], stage2_15[124], stage2_15[125], stage2_15[126], stage2_15[127]},
      {stage2_16[47]},
      {stage2_17[70], stage2_17[71], stage2_17[72], stage2_17[73], stage2_17[74], stage2_17[75]},
      {stage3_19[11],stage3_18[19],stage3_17[28],stage3_16[40],stage3_15[42]}
   );
   gpc615_5 gpc7355 (
      {stage2_15[128], stage2_15[129], stage2_15[130], stage2_15[131], stage2_15[132]},
      {stage2_16[48]},
      {stage2_17[76], stage2_17[77], stage2_17[78], stage2_17[79], stage2_17[80], stage2_17[81]},
      {stage3_19[12],stage3_18[20],stage3_17[29],stage3_16[41],stage3_15[43]}
   );
   gpc615_5 gpc7356 (
      {stage2_15[133], stage2_15[134], stage2_15[135], stage2_15[136], stage2_15[137]},
      {stage2_16[49]},
      {stage2_17[82], stage2_17[83], stage2_17[84], stage2_17[85], stage2_17[86], 1'b0},
      {stage3_19[13],stage3_18[21],stage3_17[30],stage3_16[42],stage3_15[44]}
   );
   gpc606_5 gpc7357 (
      {stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53], stage2_16[54], stage2_16[55]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[14],stage3_18[22],stage3_17[31],stage3_16[43]}
   );
   gpc606_5 gpc7358 (
      {stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59], stage2_16[60], stage2_16[61]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[15],stage3_18[23],stage3_17[32],stage3_16[44]}
   );
   gpc606_5 gpc7359 (
      {stage2_16[62], stage2_16[63], stage2_16[64], stage2_16[65], stage2_16[66], stage2_16[67]},
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage3_20[2],stage3_19[16],stage3_18[24],stage3_17[33],stage3_16[45]}
   );
   gpc606_5 gpc7360 (
      {stage2_16[68], stage2_16[69], stage2_16[70], stage2_16[71], stage2_16[72], stage2_16[73]},
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage3_20[3],stage3_19[17],stage3_18[25],stage3_17[34],stage3_16[46]}
   );
   gpc606_5 gpc7361 (
      {stage2_16[74], stage2_16[75], stage2_16[76], stage2_16[77], stage2_16[78], stage2_16[79]},
      {stage2_18[24], stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29]},
      {stage3_20[4],stage3_19[18],stage3_18[26],stage3_17[35],stage3_16[47]}
   );
   gpc2135_5 gpc7362 (
      {stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34]},
      {stage2_19[0], stage2_19[1], stage2_19[2]},
      {stage2_20[0]},
      {stage2_21[0], stage2_21[1]},
      {stage3_22[0],stage3_21[0],stage3_20[5],stage3_19[19],stage3_18[27]}
   );
   gpc2135_5 gpc7363 (
      {stage2_18[35], stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39]},
      {stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage2_20[1]},
      {stage2_21[2], stage2_21[3]},
      {stage3_22[1],stage3_21[1],stage3_20[6],stage3_19[20],stage3_18[28]}
   );
   gpc2135_5 gpc7364 (
      {stage2_18[40], stage2_18[41], stage2_18[42], stage2_18[43], stage2_18[44]},
      {stage2_19[6], stage2_19[7], stage2_19[8]},
      {stage2_20[2]},
      {stage2_21[4], stage2_21[5]},
      {stage3_22[2],stage3_21[2],stage3_20[7],stage3_19[21],stage3_18[29]}
   );
   gpc2135_5 gpc7365 (
      {stage2_18[45], stage2_18[46], stage2_18[47], stage2_18[48], stage2_18[49]},
      {stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage2_20[3]},
      {stage2_21[6], stage2_21[7]},
      {stage3_22[3],stage3_21[3],stage3_20[8],stage3_19[22],stage3_18[30]}
   );
   gpc2135_5 gpc7366 (
      {stage2_18[50], stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54]},
      {stage2_19[12], stage2_19[13], stage2_19[14]},
      {stage2_20[4]},
      {stage2_21[8], stage2_21[9]},
      {stage3_22[4],stage3_21[4],stage3_20[9],stage3_19[23],stage3_18[31]}
   );
   gpc2135_5 gpc7367 (
      {stage2_18[55], stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59]},
      {stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage2_20[5]},
      {stage2_21[10], stage2_21[11]},
      {stage3_22[5],stage3_21[5],stage3_20[10],stage3_19[24],stage3_18[32]}
   );
   gpc2135_5 gpc7368 (
      {stage2_18[60], stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64]},
      {stage2_19[18], stage2_19[19], stage2_19[20]},
      {stage2_20[6]},
      {stage2_21[12], stage2_21[13]},
      {stage3_22[6],stage3_21[6],stage3_20[11],stage3_19[25],stage3_18[33]}
   );
   gpc2135_5 gpc7369 (
      {stage2_18[65], stage2_18[66], stage2_18[67], stage2_18[68], stage2_18[69]},
      {stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage2_20[7]},
      {stage2_21[14], stage2_21[15]},
      {stage3_22[7],stage3_21[7],stage3_20[12],stage3_19[26],stage3_18[34]}
   );
   gpc2135_5 gpc7370 (
      {stage2_18[70], stage2_18[71], stage2_18[72], stage2_18[73], stage2_18[74]},
      {stage2_19[24], stage2_19[25], stage2_19[26]},
      {stage2_20[8]},
      {stage2_21[16], stage2_21[17]},
      {stage3_22[8],stage3_21[8],stage3_20[13],stage3_19[27],stage3_18[35]}
   );
   gpc2135_5 gpc7371 (
      {stage2_18[75], stage2_18[76], stage2_18[77], stage2_18[78], stage2_18[79]},
      {stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage2_20[9]},
      {stage2_21[18], stage2_21[19]},
      {stage3_22[9],stage3_21[9],stage3_20[14],stage3_19[28],stage3_18[36]}
   );
   gpc2135_5 gpc7372 (
      {stage2_18[80], stage2_18[81], stage2_18[82], stage2_18[83], stage2_18[84]},
      {stage2_19[30], stage2_19[31], stage2_19[32]},
      {stage2_20[10]},
      {stage2_21[20], stage2_21[21]},
      {stage3_22[10],stage3_21[10],stage3_20[15],stage3_19[29],stage3_18[37]}
   );
   gpc2135_5 gpc7373 (
      {stage2_18[85], stage2_18[86], stage2_18[87], stage2_18[88], stage2_18[89]},
      {stage2_19[33], stage2_19[34], stage2_19[35]},
      {stage2_20[11]},
      {stage2_21[22], stage2_21[23]},
      {stage3_22[11],stage3_21[11],stage3_20[16],stage3_19[30],stage3_18[38]}
   );
   gpc615_5 gpc7374 (
      {stage2_18[90], stage2_18[91], stage2_18[92], stage2_18[93], stage2_18[94]},
      {stage2_19[36]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[12],stage3_21[12],stage3_20[17],stage3_19[31],stage3_18[39]}
   );
   gpc615_5 gpc7375 (
      {stage2_18[95], stage2_18[96], stage2_18[97], stage2_18[98], stage2_18[99]},
      {stage2_19[37]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[13],stage3_21[13],stage3_20[18],stage3_19[32],stage3_18[40]}
   );
   gpc615_5 gpc7376 (
      {stage2_19[38], stage2_19[39], stage2_19[40], stage2_19[41], stage2_19[42]},
      {stage2_20[24]},
      {stage2_21[24], stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28], stage2_21[29]},
      {stage3_23[0],stage3_22[14],stage3_21[14],stage3_20[19],stage3_19[33]}
   );
   gpc615_5 gpc7377 (
      {stage2_19[43], stage2_19[44], stage2_19[45], stage2_19[46], stage2_19[47]},
      {stage2_20[25]},
      {stage2_21[30], stage2_21[31], stage2_21[32], stage2_21[33], stage2_21[34], stage2_21[35]},
      {stage3_23[1],stage3_22[15],stage3_21[15],stage3_20[20],stage3_19[34]}
   );
   gpc615_5 gpc7378 (
      {stage2_19[48], stage2_19[49], stage2_19[50], stage2_19[51], stage2_19[52]},
      {stage2_20[26]},
      {stage2_21[36], stage2_21[37], stage2_21[38], stage2_21[39], stage2_21[40], stage2_21[41]},
      {stage3_23[2],stage3_22[16],stage3_21[16],stage3_20[21],stage3_19[35]}
   );
   gpc615_5 gpc7379 (
      {stage2_19[53], stage2_19[54], stage2_19[55], stage2_19[56], stage2_19[57]},
      {stage2_20[27]},
      {stage2_21[42], stage2_21[43], stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47]},
      {stage3_23[3],stage3_22[17],stage3_21[17],stage3_20[22],stage3_19[36]}
   );
   gpc615_5 gpc7380 (
      {stage2_19[58], stage2_19[59], stage2_19[60], stage2_19[61], stage2_19[62]},
      {stage2_20[28]},
      {stage2_21[48], stage2_21[49], stage2_21[50], stage2_21[51], stage2_21[52], stage2_21[53]},
      {stage3_23[4],stage3_22[18],stage3_21[18],stage3_20[23],stage3_19[37]}
   );
   gpc615_5 gpc7381 (
      {stage2_19[63], stage2_19[64], stage2_19[65], stage2_19[66], stage2_19[67]},
      {stage2_20[29]},
      {stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57], stage2_21[58], stage2_21[59]},
      {stage3_23[5],stage3_22[19],stage3_21[19],stage3_20[24],stage3_19[38]}
   );
   gpc615_5 gpc7382 (
      {stage2_19[68], stage2_19[69], stage2_19[70], stage2_19[71], stage2_19[72]},
      {stage2_20[30]},
      {stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63], stage2_21[64], stage2_21[65]},
      {stage3_23[6],stage3_22[20],stage3_21[20],stage3_20[25],stage3_19[39]}
   );
   gpc615_5 gpc7383 (
      {stage2_19[73], stage2_19[74], stage2_19[75], stage2_19[76], stage2_19[77]},
      {stage2_20[31]},
      {stage2_21[66], stage2_21[67], stage2_21[68], stage2_21[69], stage2_21[70], stage2_21[71]},
      {stage3_23[7],stage3_22[21],stage3_21[21],stage3_20[26],stage3_19[40]}
   );
   gpc615_5 gpc7384 (
      {stage2_19[78], stage2_19[79], stage2_19[80], stage2_19[81], stage2_19[82]},
      {stage2_20[32]},
      {stage2_21[72], stage2_21[73], stage2_21[74], stage2_21[75], stage2_21[76], stage2_21[77]},
      {stage3_23[8],stage3_22[22],stage3_21[22],stage3_20[27],stage3_19[41]}
   );
   gpc615_5 gpc7385 (
      {stage2_19[83], stage2_19[84], stage2_19[85], stage2_19[86], stage2_19[87]},
      {stage2_20[33]},
      {stage2_21[78], stage2_21[79], stage2_21[80], stage2_21[81], stage2_21[82], stage2_21[83]},
      {stage3_23[9],stage3_22[23],stage3_21[23],stage3_20[28],stage3_19[42]}
   );
   gpc615_5 gpc7386 (
      {stage2_19[88], stage2_19[89], stage2_19[90], stage2_19[91], stage2_19[92]},
      {stage2_20[34]},
      {stage2_21[84], stage2_21[85], stage2_21[86], stage2_21[87], stage2_21[88], stage2_21[89]},
      {stage3_23[10],stage3_22[24],stage3_21[24],stage3_20[29],stage3_19[43]}
   );
   gpc615_5 gpc7387 (
      {stage2_19[93], stage2_19[94], stage2_19[95], stage2_19[96], stage2_19[97]},
      {stage2_20[35]},
      {stage2_21[90], stage2_21[91], stage2_21[92], stage2_21[93], stage2_21[94], stage2_21[95]},
      {stage3_23[11],stage3_22[25],stage3_21[25],stage3_20[30],stage3_19[44]}
   );
   gpc615_5 gpc7388 (
      {stage2_19[98], stage2_19[99], stage2_19[100], stage2_19[101], stage2_19[102]},
      {stage2_20[36]},
      {stage2_21[96], stage2_21[97], stage2_21[98], stage2_21[99], stage2_21[100], stage2_21[101]},
      {stage3_23[12],stage3_22[26],stage3_21[26],stage3_20[31],stage3_19[45]}
   );
   gpc615_5 gpc7389 (
      {stage2_19[103], stage2_19[104], stage2_19[105], stage2_19[106], stage2_19[107]},
      {stage2_20[37]},
      {stage2_21[102], stage2_21[103], stage2_21[104], stage2_21[105], stage2_21[106], stage2_21[107]},
      {stage3_23[13],stage3_22[27],stage3_21[27],stage3_20[32],stage3_19[46]}
   );
   gpc615_5 gpc7390 (
      {stage2_19[108], stage2_19[109], stage2_19[110], stage2_19[111], stage2_19[112]},
      {stage2_20[38]},
      {stage2_21[108], stage2_21[109], stage2_21[110], stage2_21[111], stage2_21[112], stage2_21[113]},
      {stage3_23[14],stage3_22[28],stage3_21[28],stage3_20[33],stage3_19[47]}
   );
   gpc606_5 gpc7391 (
      {stage2_20[39], stage2_20[40], stage2_20[41], stage2_20[42], stage2_20[43], stage2_20[44]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[15],stage3_22[29],stage3_21[29],stage3_20[34]}
   );
   gpc606_5 gpc7392 (
      {stage2_21[114], stage2_21[115], stage2_21[116], stage2_21[117], stage2_21[118], stage2_21[119]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[1],stage3_23[16],stage3_22[30],stage3_21[30]}
   );
   gpc606_5 gpc7393 (
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[1],stage3_24[2],stage3_23[17],stage3_22[31]}
   );
   gpc606_5 gpc7394 (
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[2],stage3_24[3],stage3_23[18],stage3_22[32]}
   );
   gpc606_5 gpc7395 (
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[3],stage3_24[4],stage3_23[19],stage3_22[33]}
   );
   gpc606_5 gpc7396 (
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23]},
      {stage3_26[3],stage3_25[4],stage3_24[5],stage3_23[20],stage3_22[34]}
   );
   gpc615_5 gpc7397 (
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34]},
      {stage2_23[6]},
      {stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29]},
      {stage3_26[4],stage3_25[5],stage3_24[6],stage3_23[21],stage3_22[35]}
   );
   gpc615_5 gpc7398 (
      {stage2_22[35], stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39]},
      {stage2_23[7]},
      {stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34], stage2_24[35]},
      {stage3_26[5],stage3_25[6],stage3_24[7],stage3_23[22],stage3_22[36]}
   );
   gpc615_5 gpc7399 (
      {stage2_22[40], stage2_22[41], stage2_22[42], stage2_22[43], stage2_22[44]},
      {stage2_23[8]},
      {stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40], stage2_24[41]},
      {stage3_26[6],stage3_25[7],stage3_24[8],stage3_23[23],stage3_22[37]}
   );
   gpc615_5 gpc7400 (
      {stage2_22[45], stage2_22[46], stage2_22[47], stage2_22[48], stage2_22[49]},
      {stage2_23[9]},
      {stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46], stage2_24[47]},
      {stage3_26[7],stage3_25[8],stage3_24[9],stage3_23[24],stage3_22[38]}
   );
   gpc615_5 gpc7401 (
      {stage2_22[50], stage2_22[51], stage2_22[52], stage2_22[53], stage2_22[54]},
      {stage2_23[10]},
      {stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52], stage2_24[53]},
      {stage3_26[8],stage3_25[9],stage3_24[10],stage3_23[25],stage3_22[39]}
   );
   gpc615_5 gpc7402 (
      {stage2_22[55], stage2_22[56], stage2_22[57], stage2_22[58], stage2_22[59]},
      {stage2_23[11]},
      {stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58], stage2_24[59]},
      {stage3_26[9],stage3_25[10],stage3_24[11],stage3_23[26],stage3_22[40]}
   );
   gpc615_5 gpc7403 (
      {stage2_22[60], stage2_22[61], stage2_22[62], stage2_22[63], stage2_22[64]},
      {stage2_23[12]},
      {stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64], stage2_24[65]},
      {stage3_26[10],stage3_25[11],stage3_24[12],stage3_23[27],stage3_22[41]}
   );
   gpc615_5 gpc7404 (
      {stage2_22[65], stage2_22[66], stage2_22[67], stage2_22[68], stage2_22[69]},
      {stage2_23[13]},
      {stage2_24[66], stage2_24[67], stage2_24[68], stage2_24[69], stage2_24[70], stage2_24[71]},
      {stage3_26[11],stage3_25[12],stage3_24[13],stage3_23[28],stage3_22[42]}
   );
   gpc615_5 gpc7405 (
      {stage2_22[70], stage2_22[71], stage2_22[72], stage2_22[73], stage2_22[74]},
      {stage2_23[14]},
      {stage2_24[72], stage2_24[73], stage2_24[74], stage2_24[75], stage2_24[76], stage2_24[77]},
      {stage3_26[12],stage3_25[13],stage3_24[14],stage3_23[29],stage3_22[43]}
   );
   gpc615_5 gpc7406 (
      {stage2_22[75], stage2_22[76], stage2_22[77], stage2_22[78], stage2_22[79]},
      {stage2_23[15]},
      {stage2_24[78], stage2_24[79], stage2_24[80], stage2_24[81], stage2_24[82], stage2_24[83]},
      {stage3_26[13],stage3_25[14],stage3_24[15],stage3_23[30],stage3_22[44]}
   );
   gpc2116_5 gpc7407 (
      {stage2_23[16], stage2_23[17], stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21]},
      {stage2_24[84]},
      {stage2_25[0]},
      {stage2_26[0], stage2_26[1]},
      {stage3_27[0],stage3_26[14],stage3_25[15],stage3_24[16],stage3_23[31]}
   );
   gpc615_5 gpc7408 (
      {stage2_23[22], stage2_23[23], stage2_23[24], stage2_23[25], stage2_23[26]},
      {stage2_24[85]},
      {stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5], stage2_25[6]},
      {stage3_27[1],stage3_26[15],stage3_25[16],stage3_24[17],stage3_23[32]}
   );
   gpc615_5 gpc7409 (
      {stage2_23[27], stage2_23[28], stage2_23[29], stage2_23[30], stage2_23[31]},
      {stage2_24[86]},
      {stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11], stage2_25[12]},
      {stage3_27[2],stage3_26[16],stage3_25[17],stage3_24[18],stage3_23[33]}
   );
   gpc615_5 gpc7410 (
      {stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35], stage2_23[36]},
      {stage2_24[87]},
      {stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17], stage2_25[18]},
      {stage3_27[3],stage3_26[17],stage3_25[18],stage3_24[19],stage3_23[34]}
   );
   gpc615_5 gpc7411 (
      {stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40], stage2_23[41]},
      {stage2_24[88]},
      {stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23], stage2_25[24]},
      {stage3_27[4],stage3_26[18],stage3_25[19],stage3_24[20],stage3_23[35]}
   );
   gpc615_5 gpc7412 (
      {stage2_23[42], stage2_23[43], stage2_23[44], stage2_23[45], stage2_23[46]},
      {stage2_24[89]},
      {stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29], stage2_25[30]},
      {stage3_27[5],stage3_26[19],stage3_25[20],stage3_24[21],stage3_23[36]}
   );
   gpc615_5 gpc7413 (
      {stage2_23[47], stage2_23[48], stage2_23[49], stage2_23[50], stage2_23[51]},
      {stage2_24[90]},
      {stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35], stage2_25[36]},
      {stage3_27[6],stage3_26[20],stage3_25[21],stage3_24[22],stage3_23[37]}
   );
   gpc615_5 gpc7414 (
      {stage2_23[52], stage2_23[53], stage2_23[54], stage2_23[55], stage2_23[56]},
      {stage2_24[91]},
      {stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41], stage2_25[42]},
      {stage3_27[7],stage3_26[21],stage3_25[22],stage3_24[23],stage3_23[38]}
   );
   gpc615_5 gpc7415 (
      {stage2_23[57], stage2_23[58], stage2_23[59], stage2_23[60], stage2_23[61]},
      {stage2_24[92]},
      {stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47], stage2_25[48]},
      {stage3_27[8],stage3_26[22],stage3_25[23],stage3_24[24],stage3_23[39]}
   );
   gpc615_5 gpc7416 (
      {stage2_23[62], stage2_23[63], stage2_23[64], stage2_23[65], stage2_23[66]},
      {stage2_24[93]},
      {stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53], stage2_25[54]},
      {stage3_27[9],stage3_26[23],stage3_25[24],stage3_24[25],stage3_23[40]}
   );
   gpc615_5 gpc7417 (
      {stage2_23[67], stage2_23[68], stage2_23[69], stage2_23[70], stage2_23[71]},
      {stage2_24[94]},
      {stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59], stage2_25[60]},
      {stage3_27[10],stage3_26[24],stage3_25[25],stage3_24[26],stage3_23[41]}
   );
   gpc615_5 gpc7418 (
      {stage2_23[72], stage2_23[73], stage2_23[74], stage2_23[75], 1'b0},
      {stage2_24[95]},
      {stage2_25[61], stage2_25[62], stage2_25[63], stage2_25[64], stage2_25[65], stage2_25[66]},
      {stage3_27[11],stage3_26[25],stage3_25[26],stage3_24[27],stage3_23[42]}
   );
   gpc606_5 gpc7419 (
      {stage2_24[96], stage2_24[97], stage2_24[98], stage2_24[99], stage2_24[100], stage2_24[101]},
      {stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5], stage2_26[6], stage2_26[7]},
      {stage3_28[0],stage3_27[12],stage3_26[26],stage3_25[27],stage3_24[28]}
   );
   gpc606_5 gpc7420 (
      {stage2_25[67], stage2_25[68], stage2_25[69], stage2_25[70], stage2_25[71], stage2_25[72]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[1],stage3_27[13],stage3_26[27],stage3_25[28]}
   );
   gpc606_5 gpc7421 (
      {stage2_25[73], stage2_25[74], stage2_25[75], stage2_25[76], stage2_25[77], stage2_25[78]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[2],stage3_27[14],stage3_26[28],stage3_25[29]}
   );
   gpc606_5 gpc7422 (
      {stage2_25[79], stage2_25[80], stage2_25[81], stage2_25[82], stage2_25[83], stage2_25[84]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[3],stage3_27[15],stage3_26[29],stage3_25[30]}
   );
   gpc606_5 gpc7423 (
      {stage2_25[85], stage2_25[86], stage2_25[87], stage2_25[88], stage2_25[89], stage2_25[90]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[4],stage3_27[16],stage3_26[30],stage3_25[31]}
   );
   gpc606_5 gpc7424 (
      {stage2_25[91], stage2_25[92], stage2_25[93], stage2_25[94], stage2_25[95], 1'b0},
      {stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27], stage2_27[28], stage2_27[29]},
      {stage3_29[4],stage3_28[5],stage3_27[17],stage3_26[31],stage3_25[32]}
   );
   gpc135_4 gpc7425 (
      {stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11], stage2_26[12]},
      {stage2_27[30], stage2_27[31], stage2_27[32]},
      {stage2_28[0]},
      {stage3_29[5],stage3_28[6],stage3_27[18],stage3_26[32]}
   );
   gpc135_4 gpc7426 (
      {stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage2_27[33], stage2_27[34], stage2_27[35]},
      {stage2_28[1]},
      {stage3_29[6],stage3_28[7],stage3_27[19],stage3_26[33]}
   );
   gpc135_4 gpc7427 (
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22]},
      {stage2_27[36], stage2_27[37], stage2_27[38]},
      {stage2_28[2]},
      {stage3_29[7],stage3_28[8],stage3_27[20],stage3_26[34]}
   );
   gpc135_4 gpc7428 (
      {stage2_26[23], stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27]},
      {stage2_27[39], stage2_27[40], stage2_27[41]},
      {stage2_28[3]},
      {stage3_29[8],stage3_28[9],stage3_27[21],stage3_26[35]}
   );
   gpc135_4 gpc7429 (
      {stage2_26[28], stage2_26[29], stage2_26[30], stage2_26[31], stage2_26[32]},
      {stage2_27[42], stage2_27[43], stage2_27[44]},
      {stage2_28[4]},
      {stage3_29[9],stage3_28[10],stage3_27[22],stage3_26[36]}
   );
   gpc135_4 gpc7430 (
      {stage2_26[33], stage2_26[34], stage2_26[35], stage2_26[36], stage2_26[37]},
      {stage2_27[45], stage2_27[46], stage2_27[47]},
      {stage2_28[5]},
      {stage3_29[10],stage3_28[11],stage3_27[23],stage3_26[37]}
   );
   gpc135_4 gpc7431 (
      {stage2_26[38], stage2_26[39], stage2_26[40], stage2_26[41], stage2_26[42]},
      {stage2_27[48], stage2_27[49], stage2_27[50]},
      {stage2_28[6]},
      {stage3_29[11],stage3_28[12],stage3_27[24],stage3_26[38]}
   );
   gpc135_4 gpc7432 (
      {stage2_26[43], stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47]},
      {stage2_27[51], stage2_27[52], stage2_27[53]},
      {stage2_28[7]},
      {stage3_29[12],stage3_28[13],stage3_27[25],stage3_26[39]}
   );
   gpc135_4 gpc7433 (
      {stage2_26[48], stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52]},
      {stage2_27[54], stage2_27[55], stage2_27[56]},
      {stage2_28[8]},
      {stage3_29[13],stage3_28[14],stage3_27[26],stage3_26[40]}
   );
   gpc135_4 gpc7434 (
      {stage2_26[53], stage2_26[54], stage2_26[55], stage2_26[56], stage2_26[57]},
      {stage2_27[57], stage2_27[58], stage2_27[59]},
      {stage2_28[9]},
      {stage3_29[14],stage3_28[15],stage3_27[27],stage3_26[41]}
   );
   gpc135_4 gpc7435 (
      {stage2_26[58], stage2_26[59], stage2_26[60], stage2_26[61], stage2_26[62]},
      {stage2_27[60], stage2_27[61], stage2_27[62]},
      {stage2_28[10]},
      {stage3_29[15],stage3_28[16],stage3_27[28],stage3_26[42]}
   );
   gpc135_4 gpc7436 (
      {stage2_26[63], stage2_26[64], stage2_26[65], stage2_26[66], stage2_26[67]},
      {stage2_27[63], stage2_27[64], stage2_27[65]},
      {stage2_28[11]},
      {stage3_29[16],stage3_28[17],stage3_27[29],stage3_26[43]}
   );
   gpc135_4 gpc7437 (
      {stage2_26[68], stage2_26[69], stage2_26[70], stage2_26[71], stage2_26[72]},
      {stage2_27[66], stage2_27[67], stage2_27[68]},
      {stage2_28[12]},
      {stage3_29[17],stage3_28[18],stage3_27[30],stage3_26[44]}
   );
   gpc1343_5 gpc7438 (
      {stage2_26[73], stage2_26[74], stage2_26[75]},
      {stage2_27[69], stage2_27[70], stage2_27[71], stage2_27[72]},
      {stage2_28[13], stage2_28[14], stage2_28[15]},
      {stage2_29[0]},
      {stage3_30[0],stage3_29[18],stage3_28[19],stage3_27[31],stage3_26[45]}
   );
   gpc117_4 gpc7439 (
      {stage2_26[76], stage2_26[77], stage2_26[78], stage2_26[79], stage2_26[80], stage2_26[81], stage2_26[82]},
      {stage2_27[73]},
      {stage2_28[16]},
      {stage3_29[19],stage3_28[20],stage3_27[32],stage3_26[46]}
   );
   gpc7_3 gpc7440 (
      {stage2_27[74], stage2_27[75], stage2_27[76], stage2_27[77], stage2_27[78], stage2_27[79], stage2_27[80]},
      {stage3_29[20],stage3_28[21],stage3_27[33]}
   );
   gpc7_3 gpc7441 (
      {stage2_27[81], stage2_27[82], stage2_27[83], stage2_27[84], stage2_27[85], stage2_27[86], stage2_27[87]},
      {stage3_29[21],stage3_28[22],stage3_27[34]}
   );
   gpc615_5 gpc7442 (
      {stage2_27[88], stage2_27[89], stage2_27[90], stage2_27[91], stage2_27[92]},
      {stage2_28[17]},
      {stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5], stage2_29[6]},
      {stage3_31[0],stage3_30[1],stage3_29[22],stage3_28[23],stage3_27[35]}
   );
   gpc606_5 gpc7443 (
      {stage2_28[18], stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[1],stage3_30[2],stage3_29[23],stage3_28[24]}
   );
   gpc615_5 gpc7444 (
      {stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28]},
      {stage2_29[7]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[2],stage3_30[3],stage3_29[24],stage3_28[25]}
   );
   gpc615_5 gpc7445 (
      {stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33]},
      {stage2_29[8]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[3],stage3_30[4],stage3_29[25],stage3_28[26]}
   );
   gpc615_5 gpc7446 (
      {stage2_28[34], stage2_28[35], stage2_28[36], stage2_28[37], stage2_28[38]},
      {stage2_29[9]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[4],stage3_30[5],stage3_29[26],stage3_28[27]}
   );
   gpc615_5 gpc7447 (
      {stage2_28[39], stage2_28[40], stage2_28[41], stage2_28[42], stage2_28[43]},
      {stage2_29[10]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[5],stage3_30[6],stage3_29[27],stage3_28[28]}
   );
   gpc615_5 gpc7448 (
      {stage2_28[44], stage2_28[45], stage2_28[46], stage2_28[47], stage2_28[48]},
      {stage2_29[11]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage3_32[5],stage3_31[6],stage3_30[7],stage3_29[28],stage3_28[29]}
   );
   gpc615_5 gpc7449 (
      {stage2_28[49], stage2_28[50], stage2_28[51], stage2_28[52], stage2_28[53]},
      {stage2_29[12]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage3_32[6],stage3_31[7],stage3_30[8],stage3_29[29],stage3_28[30]}
   );
   gpc615_5 gpc7450 (
      {stage2_28[54], stage2_28[55], stage2_28[56], stage2_28[57], stage2_28[58]},
      {stage2_29[13]},
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage3_32[7],stage3_31[8],stage3_30[9],stage3_29[30],stage3_28[31]}
   );
   gpc615_5 gpc7451 (
      {stage2_28[59], stage2_28[60], stage2_28[61], stage2_28[62], stage2_28[63]},
      {stage2_29[14]},
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], stage2_30[52], stage2_30[53]},
      {stage3_32[8],stage3_31[9],stage3_30[10],stage3_29[31],stage3_28[32]}
   );
   gpc615_5 gpc7452 (
      {stage2_28[64], stage2_28[65], stage2_28[66], stage2_28[67], stage2_28[68]},
      {stage2_29[15]},
      {stage2_30[54], stage2_30[55], stage2_30[56], stage2_30[57], stage2_30[58], stage2_30[59]},
      {stage3_32[9],stage3_31[10],stage3_30[11],stage3_29[32],stage3_28[33]}
   );
   gpc1163_5 gpc7453 (
      {stage2_29[16], stage2_29[17], stage2_29[18]},
      {stage2_30[60], stage2_30[61], stage2_30[62], stage2_30[63], stage2_30[64], stage2_30[65]},
      {stage2_31[0]},
      {stage2_32[0]},
      {stage3_33[0],stage3_32[10],stage3_31[11],stage3_30[12],stage3_29[33]}
   );
   gpc1163_5 gpc7454 (
      {stage2_29[19], stage2_29[20], stage2_29[21]},
      {stage2_30[66], stage2_30[67], stage2_30[68], stage2_30[69], stage2_30[70], stage2_30[71]},
      {stage2_31[1]},
      {stage2_32[1]},
      {stage3_33[1],stage3_32[11],stage3_31[12],stage3_30[13],stage3_29[34]}
   );
   gpc1163_5 gpc7455 (
      {stage2_29[22], stage2_29[23], stage2_29[24]},
      {stage2_30[72], stage2_30[73], stage2_30[74], stage2_30[75], stage2_30[76], stage2_30[77]},
      {stage2_31[2]},
      {stage2_32[2]},
      {stage3_33[2],stage3_32[12],stage3_31[13],stage3_30[14],stage3_29[35]}
   );
   gpc1163_5 gpc7456 (
      {stage2_29[25], stage2_29[26], stage2_29[27]},
      {stage2_30[78], stage2_30[79], stage2_30[80], stage2_30[81], stage2_30[82], stage2_30[83]},
      {stage2_31[3]},
      {stage2_32[3]},
      {stage3_33[3],stage3_32[13],stage3_31[14],stage3_30[15],stage3_29[36]}
   );
   gpc1163_5 gpc7457 (
      {stage2_29[28], stage2_29[29], stage2_29[30]},
      {stage2_30[84], stage2_30[85], stage2_30[86], stage2_30[87], stage2_30[88], stage2_30[89]},
      {stage2_31[4]},
      {stage2_32[4]},
      {stage3_33[4],stage3_32[14],stage3_31[15],stage3_30[16],stage3_29[37]}
   );
   gpc1163_5 gpc7458 (
      {stage2_29[31], stage2_29[32], stage2_29[33]},
      {stage2_30[90], stage2_30[91], stage2_30[92], stage2_30[93], stage2_30[94], stage2_30[95]},
      {stage2_31[5]},
      {stage2_32[5]},
      {stage3_33[5],stage3_32[15],stage3_31[16],stage3_30[17],stage3_29[38]}
   );
   gpc606_5 gpc7459 (
      {stage2_29[34], stage2_29[35], stage2_29[36], stage2_29[37], stage2_29[38], stage2_29[39]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[6],stage3_32[16],stage3_31[17],stage3_30[18],stage3_29[39]}
   );
   gpc606_5 gpc7460 (
      {stage2_29[40], stage2_29[41], stage2_29[42], stage2_29[43], stage2_29[44], stage2_29[45]},
      {stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17]},
      {stage3_33[7],stage3_32[17],stage3_31[18],stage3_30[19],stage3_29[40]}
   );
   gpc606_5 gpc7461 (
      {stage2_29[46], stage2_29[47], stage2_29[48], stage2_29[49], stage2_29[50], stage2_29[51]},
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage3_33[8],stage3_32[18],stage3_31[19],stage3_30[20],stage3_29[41]}
   );
   gpc606_5 gpc7462 (
      {stage2_29[52], stage2_29[53], stage2_29[54], stage2_29[55], stage2_29[56], stage2_29[57]},
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage3_33[9],stage3_32[19],stage3_31[20],stage3_30[21],stage3_29[42]}
   );
   gpc606_5 gpc7463 (
      {stage2_29[58], stage2_29[59], stage2_29[60], stage2_29[61], stage2_29[62], stage2_29[63]},
      {stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34], stage2_31[35]},
      {stage3_33[10],stage3_32[20],stage3_31[21],stage3_30[22],stage3_29[43]}
   );
   gpc606_5 gpc7464 (
      {stage2_29[64], stage2_29[65], stage2_29[66], stage2_29[67], stage2_29[68], stage2_29[69]},
      {stage2_31[36], stage2_31[37], stage2_31[38], stage2_31[39], stage2_31[40], stage2_31[41]},
      {stage3_33[11],stage3_32[21],stage3_31[22],stage3_30[23],stage3_29[44]}
   );
   gpc606_5 gpc7465 (
      {stage2_29[70], stage2_29[71], stage2_29[72], stage2_29[73], stage2_29[74], stage2_29[75]},
      {stage2_31[42], stage2_31[43], stage2_31[44], stage2_31[45], stage2_31[46], stage2_31[47]},
      {stage3_33[12],stage3_32[22],stage3_31[23],stage3_30[24],stage3_29[45]}
   );
   gpc606_5 gpc7466 (
      {stage2_29[76], stage2_29[77], stage2_29[78], stage2_29[79], stage2_29[80], stage2_29[81]},
      {stage2_31[48], stage2_31[49], stage2_31[50], stage2_31[51], stage2_31[52], stage2_31[53]},
      {stage3_33[13],stage3_32[23],stage3_31[24],stage3_30[25],stage3_29[46]}
   );
   gpc606_5 gpc7467 (
      {stage2_29[82], stage2_29[83], stage2_29[84], stage2_29[85], stage2_29[86], 1'b0},
      {stage2_31[54], stage2_31[55], stage2_31[56], stage2_31[57], stage2_31[58], stage2_31[59]},
      {stage3_33[14],stage3_32[24],stage3_31[25],stage3_30[26],stage3_29[47]}
   );
   gpc207_4 gpc7468 (
      {stage2_30[96], stage2_30[97], stage2_30[98], stage2_30[99], stage2_30[100], stage2_30[101], stage2_30[102]},
      {stage2_32[6], stage2_32[7]},
      {stage3_33[15],stage3_32[25],stage3_31[26],stage3_30[27]}
   );
   gpc615_5 gpc7469 (
      {stage2_31[60], stage2_31[61], stage2_31[62], stage2_31[63], stage2_31[64]},
      {stage2_32[8]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[0],stage3_33[16],stage3_32[26],stage3_31[27]}
   );
   gpc615_5 gpc7470 (
      {stage2_31[65], stage2_31[66], stage2_31[67], stage2_31[68], stage2_31[69]},
      {stage2_32[9]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[1],stage3_33[17],stage3_32[27],stage3_31[28]}
   );
   gpc615_5 gpc7471 (
      {stage2_31[70], stage2_31[71], stage2_31[72], stage2_31[73], stage2_31[74]},
      {stage2_32[10]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[2],stage3_33[18],stage3_32[28],stage3_31[29]}
   );
   gpc615_5 gpc7472 (
      {stage2_31[75], stage2_31[76], stage2_31[77], stage2_31[78], stage2_31[79]},
      {stage2_32[11]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[3],stage3_33[19],stage3_32[29],stage3_31[30]}
   );
   gpc615_5 gpc7473 (
      {stage2_31[80], stage2_31[81], stage2_31[82], stage2_31[83], stage2_31[84]},
      {stage2_32[12]},
      {stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29]},
      {stage3_35[4],stage3_34[4],stage3_33[20],stage3_32[30],stage3_31[31]}
   );
   gpc615_5 gpc7474 (
      {stage2_31[85], stage2_31[86], stage2_31[87], stage2_31[88], stage2_31[89]},
      {stage2_32[13]},
      {stage2_33[30], stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35]},
      {stage3_35[5],stage3_34[5],stage3_33[21],stage3_32[31],stage3_31[32]}
   );
   gpc615_5 gpc7475 (
      {stage2_31[90], stage2_31[91], stage2_31[92], stage2_31[93], stage2_31[94]},
      {stage2_32[14]},
      {stage2_33[36], stage2_33[37], stage2_33[38], stage2_33[39], stage2_33[40], stage2_33[41]},
      {stage3_35[6],stage3_34[6],stage3_33[22],stage3_32[32],stage3_31[33]}
   );
   gpc606_5 gpc7476 (
      {stage2_32[15], stage2_32[16], stage2_32[17], stage2_32[18], stage2_32[19], stage2_32[20]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[7],stage3_34[7],stage3_33[23],stage3_32[33]}
   );
   gpc606_5 gpc7477 (
      {stage2_32[21], stage2_32[22], stage2_32[23], stage2_32[24], stage2_32[25], stage2_32[26]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[8],stage3_34[8],stage3_33[24],stage3_32[34]}
   );
   gpc606_5 gpc7478 (
      {stage2_32[27], stage2_32[28], stage2_32[29], stage2_32[30], stage2_32[31], stage2_32[32]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17]},
      {stage3_36[2],stage3_35[9],stage3_34[9],stage3_33[25],stage3_32[35]}
   );
   gpc606_5 gpc7479 (
      {stage2_32[33], stage2_32[34], stage2_32[35], stage2_32[36], stage2_32[37], stage2_32[38]},
      {stage2_34[18], stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23]},
      {stage3_36[3],stage3_35[10],stage3_34[10],stage3_33[26],stage3_32[36]}
   );
   gpc606_5 gpc7480 (
      {stage2_32[39], stage2_32[40], stage2_32[41], stage2_32[42], stage2_32[43], stage2_32[44]},
      {stage2_34[24], stage2_34[25], stage2_34[26], stage2_34[27], stage2_34[28], stage2_34[29]},
      {stage3_36[4],stage3_35[11],stage3_34[11],stage3_33[27],stage3_32[37]}
   );
   gpc606_5 gpc7481 (
      {stage2_32[45], stage2_32[46], stage2_32[47], stage2_32[48], stage2_32[49], stage2_32[50]},
      {stage2_34[30], stage2_34[31], stage2_34[32], stage2_34[33], stage2_34[34], stage2_34[35]},
      {stage3_36[5],stage3_35[12],stage3_34[12],stage3_33[28],stage3_32[38]}
   );
   gpc606_5 gpc7482 (
      {stage2_32[51], stage2_32[52], stage2_32[53], stage2_32[54], stage2_32[55], stage2_32[56]},
      {stage2_34[36], stage2_34[37], stage2_34[38], stage2_34[39], stage2_34[40], stage2_34[41]},
      {stage3_36[6],stage3_35[13],stage3_34[13],stage3_33[29],stage3_32[39]}
   );
   gpc606_5 gpc7483 (
      {stage2_32[57], stage2_32[58], stage2_32[59], stage2_32[60], stage2_32[61], stage2_32[62]},
      {stage2_34[42], stage2_34[43], stage2_34[44], stage2_34[45], stage2_34[46], stage2_34[47]},
      {stage3_36[7],stage3_35[14],stage3_34[14],stage3_33[30],stage3_32[40]}
   );
   gpc606_5 gpc7484 (
      {stage2_32[63], stage2_32[64], stage2_32[65], stage2_32[66], stage2_32[67], stage2_32[68]},
      {stage2_34[48], stage2_34[49], stage2_34[50], stage2_34[51], stage2_34[52], stage2_34[53]},
      {stage3_36[8],stage3_35[15],stage3_34[15],stage3_33[31],stage3_32[41]}
   );
   gpc606_5 gpc7485 (
      {stage2_32[69], stage2_32[70], stage2_32[71], stage2_32[72], stage2_32[73], stage2_32[74]},
      {stage2_34[54], stage2_34[55], stage2_34[56], stage2_34[57], stage2_34[58], stage2_34[59]},
      {stage3_36[9],stage3_35[16],stage3_34[16],stage3_33[32],stage3_32[42]}
   );
   gpc606_5 gpc7486 (
      {stage2_32[75], stage2_32[76], stage2_32[77], stage2_32[78], stage2_32[79], stage2_32[80]},
      {stage2_34[60], stage2_34[61], stage2_34[62], stage2_34[63], stage2_34[64], stage2_34[65]},
      {stage3_36[10],stage3_35[17],stage3_34[17],stage3_33[33],stage3_32[43]}
   );
   gpc606_5 gpc7487 (
      {stage2_32[81], stage2_32[82], stage2_32[83], stage2_32[84], stage2_32[85], stage2_32[86]},
      {stage2_34[66], stage2_34[67], stage2_34[68], stage2_34[69], stage2_34[70], stage2_34[71]},
      {stage3_36[11],stage3_35[18],stage3_34[18],stage3_33[34],stage3_32[44]}
   );
   gpc606_5 gpc7488 (
      {stage2_32[87], stage2_32[88], stage2_32[89], stage2_32[90], stage2_32[91], stage2_32[92]},
      {stage2_34[72], stage2_34[73], stage2_34[74], stage2_34[75], stage2_34[76], stage2_34[77]},
      {stage3_36[12],stage3_35[19],stage3_34[19],stage3_33[35],stage3_32[45]}
   );
   gpc606_5 gpc7489 (
      {stage2_32[93], stage2_32[94], stage2_32[95], stage2_32[96], stage2_32[97], stage2_32[98]},
      {stage2_34[78], stage2_34[79], stage2_34[80], stage2_34[81], stage2_34[82], stage2_34[83]},
      {stage3_36[13],stage3_35[20],stage3_34[20],stage3_33[36],stage3_32[46]}
   );
   gpc606_5 gpc7490 (
      {stage2_33[42], stage2_33[43], stage2_33[44], stage2_33[45], stage2_33[46], stage2_33[47]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[14],stage3_35[21],stage3_34[21],stage3_33[37]}
   );
   gpc606_5 gpc7491 (
      {stage2_33[48], stage2_33[49], stage2_33[50], stage2_33[51], stage2_33[52], stage2_33[53]},
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11]},
      {stage3_37[1],stage3_36[15],stage3_35[22],stage3_34[22],stage3_33[38]}
   );
   gpc606_5 gpc7492 (
      {stage2_33[54], stage2_33[55], stage2_33[56], stage2_33[57], stage2_33[58], stage2_33[59]},
      {stage2_35[12], stage2_35[13], stage2_35[14], stage2_35[15], stage2_35[16], stage2_35[17]},
      {stage3_37[2],stage3_36[16],stage3_35[23],stage3_34[23],stage3_33[39]}
   );
   gpc606_5 gpc7493 (
      {stage2_33[60], stage2_33[61], stage2_33[62], stage2_33[63], stage2_33[64], stage2_33[65]},
      {stage2_35[18], stage2_35[19], stage2_35[20], stage2_35[21], stage2_35[22], stage2_35[23]},
      {stage3_37[3],stage3_36[17],stage3_35[24],stage3_34[24],stage3_33[40]}
   );
   gpc606_5 gpc7494 (
      {stage2_33[66], stage2_33[67], stage2_33[68], stage2_33[69], stage2_33[70], stage2_33[71]},
      {stage2_35[24], stage2_35[25], stage2_35[26], stage2_35[27], stage2_35[28], stage2_35[29]},
      {stage3_37[4],stage3_36[18],stage3_35[25],stage3_34[25],stage3_33[41]}
   );
   gpc1163_5 gpc7495 (
      {stage2_34[84], stage2_34[85], stage2_34[86]},
      {stage2_35[30], stage2_35[31], stage2_35[32], stage2_35[33], stage2_35[34], stage2_35[35]},
      {stage2_36[0]},
      {stage2_37[0]},
      {stage3_38[0],stage3_37[5],stage3_36[19],stage3_35[26],stage3_34[26]}
   );
   gpc1163_5 gpc7496 (
      {stage2_34[87], stage2_34[88], stage2_34[89]},
      {stage2_35[36], stage2_35[37], stage2_35[38], stage2_35[39], stage2_35[40], stage2_35[41]},
      {stage2_36[1]},
      {stage2_37[1]},
      {stage3_38[1],stage3_37[6],stage3_36[20],stage3_35[27],stage3_34[27]}
   );
   gpc1163_5 gpc7497 (
      {stage2_34[90], stage2_34[91], stage2_34[92]},
      {stage2_35[42], stage2_35[43], stage2_35[44], stage2_35[45], stage2_35[46], stage2_35[47]},
      {stage2_36[2]},
      {stage2_37[2]},
      {stage3_38[2],stage3_37[7],stage3_36[21],stage3_35[28],stage3_34[28]}
   );
   gpc1163_5 gpc7498 (
      {stage2_34[93], stage2_34[94], stage2_34[95]},
      {stage2_35[48], stage2_35[49], stage2_35[50], stage2_35[51], stage2_35[52], stage2_35[53]},
      {stage2_36[3]},
      {stage2_37[3]},
      {stage3_38[3],stage3_37[8],stage3_36[22],stage3_35[29],stage3_34[29]}
   );
   gpc1163_5 gpc7499 (
      {stage2_34[96], stage2_34[97], stage2_34[98]},
      {stage2_35[54], stage2_35[55], stage2_35[56], stage2_35[57], stage2_35[58], stage2_35[59]},
      {stage2_36[4]},
      {stage2_37[4]},
      {stage3_38[4],stage3_37[9],stage3_36[23],stage3_35[30],stage3_34[30]}
   );
   gpc1163_5 gpc7500 (
      {stage2_34[99], stage2_34[100], stage2_34[101]},
      {stage2_35[60], stage2_35[61], stage2_35[62], stage2_35[63], stage2_35[64], stage2_35[65]},
      {stage2_36[5]},
      {stage2_37[5]},
      {stage3_38[5],stage3_37[10],stage3_36[24],stage3_35[31],stage3_34[31]}
   );
   gpc1163_5 gpc7501 (
      {stage2_34[102], stage2_34[103], stage2_34[104]},
      {stage2_35[66], stage2_35[67], stage2_35[68], stage2_35[69], stage2_35[70], stage2_35[71]},
      {stage2_36[6]},
      {stage2_37[6]},
      {stage3_38[6],stage3_37[11],stage3_36[25],stage3_35[32],stage3_34[32]}
   );
   gpc1163_5 gpc7502 (
      {stage2_34[105], stage2_34[106], stage2_34[107]},
      {stage2_35[72], stage2_35[73], stage2_35[74], stage2_35[75], stage2_35[76], stage2_35[77]},
      {stage2_36[7]},
      {stage2_37[7]},
      {stage3_38[7],stage3_37[12],stage3_36[26],stage3_35[33],stage3_34[33]}
   );
   gpc1163_5 gpc7503 (
      {stage2_34[108], stage2_34[109], stage2_34[110]},
      {stage2_35[78], stage2_35[79], stage2_35[80], stage2_35[81], stage2_35[82], stage2_35[83]},
      {stage2_36[8]},
      {stage2_37[8]},
      {stage3_38[8],stage3_37[13],stage3_36[27],stage3_35[34],stage3_34[34]}
   );
   gpc1163_5 gpc7504 (
      {stage2_34[111], stage2_34[112], stage2_34[113]},
      {stage2_35[84], stage2_35[85], stage2_35[86], stage2_35[87], stage2_35[88], stage2_35[89]},
      {stage2_36[9]},
      {stage2_37[9]},
      {stage3_38[9],stage3_37[14],stage3_36[28],stage3_35[35],stage3_34[35]}
   );
   gpc615_5 gpc7505 (
      {stage2_34[114], stage2_34[115], stage2_34[116], stage2_34[117], stage2_34[118]},
      {stage2_35[90]},
      {stage2_36[10], stage2_36[11], stage2_36[12], stage2_36[13], stage2_36[14], stage2_36[15]},
      {stage3_38[10],stage3_37[15],stage3_36[29],stage3_35[36],stage3_34[36]}
   );
   gpc615_5 gpc7506 (
      {stage2_34[119], stage2_34[120], stage2_34[121], stage2_34[122], stage2_34[123]},
      {stage2_35[91]},
      {stage2_36[16], stage2_36[17], stage2_36[18], stage2_36[19], stage2_36[20], stage2_36[21]},
      {stage3_38[11],stage3_37[16],stage3_36[30],stage3_35[37],stage3_34[37]}
   );
   gpc615_5 gpc7507 (
      {stage2_34[124], stage2_34[125], stage2_34[126], stage2_34[127], stage2_34[128]},
      {stage2_35[92]},
      {stage2_36[22], stage2_36[23], stage2_36[24], stage2_36[25], stage2_36[26], stage2_36[27]},
      {stage3_38[12],stage3_37[17],stage3_36[31],stage3_35[38],stage3_34[38]}
   );
   gpc1406_5 gpc7508 (
      {stage2_35[93], stage2_35[94], stage2_35[95], stage2_35[96], stage2_35[97], stage2_35[98]},
      {stage2_37[10], stage2_37[11], stage2_37[12], stage2_37[13]},
      {stage2_38[0]},
      {stage3_39[0],stage3_38[13],stage3_37[18],stage3_36[32],stage3_35[39]}
   );
   gpc1406_5 gpc7509 (
      {stage2_35[99], stage2_35[100], stage2_35[101], stage2_35[102], stage2_35[103], stage2_35[104]},
      {stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage2_38[1]},
      {stage3_39[1],stage3_38[14],stage3_37[19],stage3_36[33],stage3_35[40]}
   );
   gpc615_5 gpc7510 (
      {stage2_35[105], stage2_35[106], stage2_35[107], stage2_35[108], stage2_35[109]},
      {stage2_36[28]},
      {stage2_37[18], stage2_37[19], stage2_37[20], stage2_37[21], stage2_37[22], stage2_37[23]},
      {stage3_39[2],stage3_38[15],stage3_37[20],stage3_36[34],stage3_35[41]}
   );
   gpc615_5 gpc7511 (
      {stage2_35[110], stage2_35[111], stage2_35[112], stage2_35[113], stage2_35[114]},
      {stage2_36[29]},
      {stage2_37[24], stage2_37[25], stage2_37[26], stage2_37[27], stage2_37[28], stage2_37[29]},
      {stage3_39[3],stage3_38[16],stage3_37[21],stage3_36[35],stage3_35[42]}
   );
   gpc615_5 gpc7512 (
      {stage2_35[115], stage2_35[116], stage2_35[117], stage2_35[118], stage2_35[119]},
      {stage2_36[30]},
      {stage2_37[30], stage2_37[31], stage2_37[32], stage2_37[33], stage2_37[34], stage2_37[35]},
      {stage3_39[4],stage3_38[17],stage3_37[22],stage3_36[36],stage3_35[43]}
   );
   gpc606_5 gpc7513 (
      {stage2_36[31], stage2_36[32], stage2_36[33], stage2_36[34], stage2_36[35], stage2_36[36]},
      {stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5], stage2_38[6], stage2_38[7]},
      {stage3_40[0],stage3_39[5],stage3_38[18],stage3_37[23],stage3_36[37]}
   );
   gpc606_5 gpc7514 (
      {stage2_36[37], stage2_36[38], stage2_36[39], stage2_36[40], stage2_36[41], stage2_36[42]},
      {stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11], stage2_38[12], stage2_38[13]},
      {stage3_40[1],stage3_39[6],stage3_38[19],stage3_37[24],stage3_36[38]}
   );
   gpc606_5 gpc7515 (
      {stage2_36[43], stage2_36[44], stage2_36[45], stage2_36[46], stage2_36[47], stage2_36[48]},
      {stage2_38[14], stage2_38[15], stage2_38[16], stage2_38[17], stage2_38[18], stage2_38[19]},
      {stage3_40[2],stage3_39[7],stage3_38[20],stage3_37[25],stage3_36[39]}
   );
   gpc606_5 gpc7516 (
      {stage2_36[49], stage2_36[50], stage2_36[51], stage2_36[52], stage2_36[53], stage2_36[54]},
      {stage2_38[20], stage2_38[21], stage2_38[22], stage2_38[23], stage2_38[24], stage2_38[25]},
      {stage3_40[3],stage3_39[8],stage3_38[21],stage3_37[26],stage3_36[40]}
   );
   gpc606_5 gpc7517 (
      {stage2_36[55], stage2_36[56], stage2_36[57], stage2_36[58], stage2_36[59], stage2_36[60]},
      {stage2_38[26], stage2_38[27], stage2_38[28], stage2_38[29], stage2_38[30], stage2_38[31]},
      {stage3_40[4],stage3_39[9],stage3_38[22],stage3_37[27],stage3_36[41]}
   );
   gpc606_5 gpc7518 (
      {stage2_36[61], stage2_36[62], stage2_36[63], stage2_36[64], stage2_36[65], stage2_36[66]},
      {stage2_38[32], stage2_38[33], stage2_38[34], stage2_38[35], stage2_38[36], stage2_38[37]},
      {stage3_40[5],stage3_39[10],stage3_38[23],stage3_37[28],stage3_36[42]}
   );
   gpc606_5 gpc7519 (
      {stage2_36[67], stage2_36[68], stage2_36[69], stage2_36[70], stage2_36[71], stage2_36[72]},
      {stage2_38[38], stage2_38[39], stage2_38[40], stage2_38[41], stage2_38[42], stage2_38[43]},
      {stage3_40[6],stage3_39[11],stage3_38[24],stage3_37[29],stage3_36[43]}
   );
   gpc606_5 gpc7520 (
      {stage2_37[36], stage2_37[37], stage2_37[38], stage2_37[39], stage2_37[40], stage2_37[41]},
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5]},
      {stage3_41[0],stage3_40[7],stage3_39[12],stage3_38[25],stage3_37[30]}
   );
   gpc606_5 gpc7521 (
      {stage2_37[42], stage2_37[43], stage2_37[44], stage2_37[45], stage2_37[46], stage2_37[47]},
      {stage2_39[6], stage2_39[7], stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11]},
      {stage3_41[1],stage3_40[8],stage3_39[13],stage3_38[26],stage3_37[31]}
   );
   gpc606_5 gpc7522 (
      {stage2_37[48], stage2_37[49], stage2_37[50], stage2_37[51], stage2_37[52], stage2_37[53]},
      {stage2_39[12], stage2_39[13], stage2_39[14], stage2_39[15], stage2_39[16], stage2_39[17]},
      {stage3_41[2],stage3_40[9],stage3_39[14],stage3_38[27],stage3_37[32]}
   );
   gpc615_5 gpc7523 (
      {stage2_37[54], stage2_37[55], stage2_37[56], stage2_37[57], stage2_37[58]},
      {stage2_38[44]},
      {stage2_39[18], stage2_39[19], stage2_39[20], stage2_39[21], stage2_39[22], stage2_39[23]},
      {stage3_41[3],stage3_40[10],stage3_39[15],stage3_38[28],stage3_37[33]}
   );
   gpc615_5 gpc7524 (
      {stage2_37[59], stage2_37[60], stage2_37[61], stage2_37[62], stage2_37[63]},
      {stage2_38[45]},
      {stage2_39[24], stage2_39[25], stage2_39[26], stage2_39[27], stage2_39[28], stage2_39[29]},
      {stage3_41[4],stage3_40[11],stage3_39[16],stage3_38[29],stage3_37[34]}
   );
   gpc615_5 gpc7525 (
      {stage2_37[64], stage2_37[65], stage2_37[66], stage2_37[67], stage2_37[68]},
      {stage2_38[46]},
      {stage2_39[30], stage2_39[31], stage2_39[32], stage2_39[33], stage2_39[34], stage2_39[35]},
      {stage3_41[5],stage3_40[12],stage3_39[17],stage3_38[30],stage3_37[35]}
   );
   gpc615_5 gpc7526 (
      {stage2_37[69], stage2_37[70], stage2_37[71], stage2_37[72], stage2_37[73]},
      {stage2_38[47]},
      {stage2_39[36], stage2_39[37], stage2_39[38], stage2_39[39], stage2_39[40], stage2_39[41]},
      {stage3_41[6],stage3_40[13],stage3_39[18],stage3_38[31],stage3_37[36]}
   );
   gpc606_5 gpc7527 (
      {stage2_38[48], stage2_38[49], stage2_38[50], stage2_38[51], stage2_38[52], stage2_38[53]},
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage3_42[0],stage3_41[7],stage3_40[14],stage3_39[19],stage3_38[32]}
   );
   gpc606_5 gpc7528 (
      {stage2_38[54], stage2_38[55], stage2_38[56], stage2_38[57], stage2_38[58], stage2_38[59]},
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage3_42[1],stage3_41[8],stage3_40[15],stage3_39[20],stage3_38[33]}
   );
   gpc606_5 gpc7529 (
      {stage2_38[60], stage2_38[61], stage2_38[62], stage2_38[63], stage2_38[64], stage2_38[65]},
      {stage2_40[12], stage2_40[13], stage2_40[14], stage2_40[15], stage2_40[16], stage2_40[17]},
      {stage3_42[2],stage3_41[9],stage3_40[16],stage3_39[21],stage3_38[34]}
   );
   gpc606_5 gpc7530 (
      {stage2_38[66], stage2_38[67], stage2_38[68], stage2_38[69], stage2_38[70], stage2_38[71]},
      {stage2_40[18], stage2_40[19], stage2_40[20], stage2_40[21], stage2_40[22], stage2_40[23]},
      {stage3_42[3],stage3_41[10],stage3_40[17],stage3_39[22],stage3_38[35]}
   );
   gpc606_5 gpc7531 (
      {stage2_38[72], stage2_38[73], stage2_38[74], stage2_38[75], stage2_38[76], stage2_38[77]},
      {stage2_40[24], stage2_40[25], stage2_40[26], stage2_40[27], stage2_40[28], stage2_40[29]},
      {stage3_42[4],stage3_41[11],stage3_40[18],stage3_39[23],stage3_38[36]}
   );
   gpc606_5 gpc7532 (
      {stage2_38[78], stage2_38[79], stage2_38[80], stage2_38[81], stage2_38[82], stage2_38[83]},
      {stage2_40[30], stage2_40[31], stage2_40[32], stage2_40[33], stage2_40[34], stage2_40[35]},
      {stage3_42[5],stage3_41[12],stage3_40[19],stage3_39[24],stage3_38[37]}
   );
   gpc606_5 gpc7533 (
      {stage2_38[84], stage2_38[85], stage2_38[86], stage2_38[87], stage2_38[88], stage2_38[89]},
      {stage2_40[36], stage2_40[37], stage2_40[38], stage2_40[39], stage2_40[40], stage2_40[41]},
      {stage3_42[6],stage3_41[13],stage3_40[20],stage3_39[25],stage3_38[38]}
   );
   gpc606_5 gpc7534 (
      {stage2_38[90], stage2_38[91], stage2_38[92], stage2_38[93], stage2_38[94], stage2_38[95]},
      {stage2_40[42], stage2_40[43], stage2_40[44], stage2_40[45], stage2_40[46], stage2_40[47]},
      {stage3_42[7],stage3_41[14],stage3_40[21],stage3_39[26],stage3_38[39]}
   );
   gpc606_5 gpc7535 (
      {stage2_38[96], stage2_38[97], stage2_38[98], stage2_38[99], stage2_38[100], stage2_38[101]},
      {stage2_40[48], stage2_40[49], stage2_40[50], stage2_40[51], stage2_40[52], stage2_40[53]},
      {stage3_42[8],stage3_41[15],stage3_40[22],stage3_39[27],stage3_38[40]}
   );
   gpc606_5 gpc7536 (
      {stage2_38[102], stage2_38[103], stage2_38[104], stage2_38[105], stage2_38[106], stage2_38[107]},
      {stage2_40[54], stage2_40[55], stage2_40[56], stage2_40[57], stage2_40[58], stage2_40[59]},
      {stage3_42[9],stage3_41[16],stage3_40[23],stage3_39[28],stage3_38[41]}
   );
   gpc606_5 gpc7537 (
      {stage2_38[108], stage2_38[109], stage2_38[110], stage2_38[111], stage2_38[112], stage2_38[113]},
      {stage2_40[60], stage2_40[61], stage2_40[62], stage2_40[63], stage2_40[64], stage2_40[65]},
      {stage3_42[10],stage3_41[17],stage3_40[24],stage3_39[29],stage3_38[42]}
   );
   gpc606_5 gpc7538 (
      {stage2_38[114], stage2_38[115], stage2_38[116], stage2_38[117], stage2_38[118], stage2_38[119]},
      {stage2_40[66], stage2_40[67], stage2_40[68], stage2_40[69], stage2_40[70], stage2_40[71]},
      {stage3_42[11],stage3_41[18],stage3_40[25],stage3_39[30],stage3_38[43]}
   );
   gpc615_5 gpc7539 (
      {stage2_38[120], stage2_38[121], stage2_38[122], stage2_38[123], stage2_38[124]},
      {stage2_39[42]},
      {stage2_40[72], stage2_40[73], stage2_40[74], stage2_40[75], stage2_40[76], stage2_40[77]},
      {stage3_42[12],stage3_41[19],stage3_40[26],stage3_39[31],stage3_38[44]}
   );
   gpc615_5 gpc7540 (
      {stage2_39[43], stage2_39[44], stage2_39[45], stage2_39[46], stage2_39[47]},
      {stage2_40[78]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[13],stage3_41[20],stage3_40[27],stage3_39[32]}
   );
   gpc615_5 gpc7541 (
      {stage2_39[48], stage2_39[49], stage2_39[50], stage2_39[51], stage2_39[52]},
      {stage2_40[79]},
      {stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11]},
      {stage3_43[1],stage3_42[14],stage3_41[21],stage3_40[28],stage3_39[33]}
   );
   gpc615_5 gpc7542 (
      {stage2_39[53], stage2_39[54], stage2_39[55], stage2_39[56], stage2_39[57]},
      {stage2_40[80]},
      {stage2_41[12], stage2_41[13], stage2_41[14], stage2_41[15], stage2_41[16], stage2_41[17]},
      {stage3_43[2],stage3_42[15],stage3_41[22],stage3_40[29],stage3_39[34]}
   );
   gpc615_5 gpc7543 (
      {stage2_39[58], stage2_39[59], stage2_39[60], stage2_39[61], stage2_39[62]},
      {stage2_40[81]},
      {stage2_41[18], stage2_41[19], stage2_41[20], stage2_41[21], stage2_41[22], stage2_41[23]},
      {stage3_43[3],stage3_42[16],stage3_41[23],stage3_40[30],stage3_39[35]}
   );
   gpc615_5 gpc7544 (
      {stage2_39[63], stage2_39[64], stage2_39[65], stage2_39[66], stage2_39[67]},
      {stage2_40[82]},
      {stage2_41[24], stage2_41[25], stage2_41[26], stage2_41[27], stage2_41[28], stage2_41[29]},
      {stage3_43[4],stage3_42[17],stage3_41[24],stage3_40[31],stage3_39[36]}
   );
   gpc615_5 gpc7545 (
      {stage2_39[68], stage2_39[69], stage2_39[70], stage2_39[71], stage2_39[72]},
      {stage2_40[83]},
      {stage2_41[30], stage2_41[31], stage2_41[32], stage2_41[33], stage2_41[34], stage2_41[35]},
      {stage3_43[5],stage3_42[18],stage3_41[25],stage3_40[32],stage3_39[37]}
   );
   gpc615_5 gpc7546 (
      {stage2_39[73], stage2_39[74], stage2_39[75], stage2_39[76], stage2_39[77]},
      {stage2_40[84]},
      {stage2_41[36], stage2_41[37], stage2_41[38], stage2_41[39], stage2_41[40], stage2_41[41]},
      {stage3_43[6],stage3_42[19],stage3_41[26],stage3_40[33],stage3_39[38]}
   );
   gpc615_5 gpc7547 (
      {stage2_39[78], stage2_39[79], stage2_39[80], stage2_39[81], stage2_39[82]},
      {stage2_40[85]},
      {stage2_41[42], stage2_41[43], stage2_41[44], stage2_41[45], stage2_41[46], stage2_41[47]},
      {stage3_43[7],stage3_42[20],stage3_41[27],stage3_40[34],stage3_39[39]}
   );
   gpc615_5 gpc7548 (
      {stage2_39[83], stage2_39[84], stage2_39[85], stage2_39[86], stage2_39[87]},
      {stage2_40[86]},
      {stage2_41[48], stage2_41[49], stage2_41[50], stage2_41[51], stage2_41[52], stage2_41[53]},
      {stage3_43[8],stage3_42[21],stage3_41[28],stage3_40[35],stage3_39[40]}
   );
   gpc615_5 gpc7549 (
      {stage2_39[88], stage2_39[89], stage2_39[90], stage2_39[91], stage2_39[92]},
      {stage2_40[87]},
      {stage2_41[54], stage2_41[55], stage2_41[56], stage2_41[57], stage2_41[58], stage2_41[59]},
      {stage3_43[9],stage3_42[22],stage3_41[29],stage3_40[36],stage3_39[41]}
   );
   gpc615_5 gpc7550 (
      {stage2_39[93], stage2_39[94], stage2_39[95], stage2_39[96], stage2_39[97]},
      {stage2_40[88]},
      {stage2_41[60], stage2_41[61], stage2_41[62], stage2_41[63], stage2_41[64], stage2_41[65]},
      {stage3_43[10],stage3_42[23],stage3_41[30],stage3_40[37],stage3_39[42]}
   );
   gpc615_5 gpc7551 (
      {stage2_39[98], stage2_39[99], stage2_39[100], stage2_39[101], stage2_39[102]},
      {stage2_40[89]},
      {stage2_41[66], stage2_41[67], stage2_41[68], stage2_41[69], stage2_41[70], stage2_41[71]},
      {stage3_43[11],stage3_42[24],stage3_41[31],stage3_40[38],stage3_39[43]}
   );
   gpc615_5 gpc7552 (
      {stage2_39[103], stage2_39[104], stage2_39[105], stage2_39[106], stage2_39[107]},
      {stage2_40[90]},
      {stage2_41[72], stage2_41[73], stage2_41[74], stage2_41[75], stage2_41[76], stage2_41[77]},
      {stage3_43[12],stage3_42[25],stage3_41[32],stage3_40[39],stage3_39[44]}
   );
   gpc615_5 gpc7553 (
      {stage2_39[108], stage2_39[109], stage2_39[110], stage2_39[111], stage2_39[112]},
      {stage2_40[91]},
      {stage2_41[78], stage2_41[79], stage2_41[80], stage2_41[81], stage2_41[82], stage2_41[83]},
      {stage3_43[13],stage3_42[26],stage3_41[33],stage3_40[40],stage3_39[45]}
   );
   gpc615_5 gpc7554 (
      {stage2_39[113], stage2_39[114], stage2_39[115], stage2_39[116], stage2_39[117]},
      {stage2_40[92]},
      {stage2_41[84], stage2_41[85], stage2_41[86], stage2_41[87], stage2_41[88], stage2_41[89]},
      {stage3_43[14],stage3_42[27],stage3_41[34],stage3_40[41],stage3_39[46]}
   );
   gpc615_5 gpc7555 (
      {stage2_39[118], stage2_39[119], stage2_39[120], stage2_39[121], stage2_39[122]},
      {stage2_40[93]},
      {stage2_41[90], stage2_41[91], stage2_41[92], stage2_41[93], stage2_41[94], stage2_41[95]},
      {stage3_43[15],stage3_42[28],stage3_41[35],stage3_40[42],stage3_39[47]}
   );
   gpc615_5 gpc7556 (
      {stage2_39[123], stage2_39[124], stage2_39[125], stage2_39[126], stage2_39[127]},
      {stage2_40[94]},
      {stage2_41[96], stage2_41[97], stage2_41[98], stage2_41[99], stage2_41[100], stage2_41[101]},
      {stage3_43[16],stage3_42[29],stage3_41[36],stage3_40[43],stage3_39[48]}
   );
   gpc606_5 gpc7557 (
      {stage2_40[95], stage2_40[96], stage2_40[97], stage2_40[98], stage2_40[99], stage2_40[100]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[17],stage3_42[30],stage3_41[37],stage3_40[44]}
   );
   gpc606_5 gpc7558 (
      {stage2_40[101], stage2_40[102], stage2_40[103], stage2_40[104], stage2_40[105], stage2_40[106]},
      {stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage3_44[1],stage3_43[18],stage3_42[31],stage3_41[38],stage3_40[45]}
   );
   gpc615_5 gpc7559 (
      {stage2_42[12], stage2_42[13], stage2_42[14], stage2_42[15], stage2_42[16]},
      {stage2_43[0]},
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage3_46[0],stage3_45[0],stage3_44[2],stage3_43[19],stage3_42[32]}
   );
   gpc615_5 gpc7560 (
      {stage2_42[17], stage2_42[18], stage2_42[19], stage2_42[20], stage2_42[21]},
      {stage2_43[1]},
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage3_46[1],stage3_45[1],stage3_44[3],stage3_43[20],stage3_42[33]}
   );
   gpc615_5 gpc7561 (
      {stage2_42[22], stage2_42[23], stage2_42[24], stage2_42[25], stage2_42[26]},
      {stage2_43[2]},
      {stage2_44[12], stage2_44[13], stage2_44[14], stage2_44[15], stage2_44[16], stage2_44[17]},
      {stage3_46[2],stage3_45[2],stage3_44[4],stage3_43[21],stage3_42[34]}
   );
   gpc615_5 gpc7562 (
      {stage2_42[27], stage2_42[28], stage2_42[29], stage2_42[30], stage2_42[31]},
      {stage2_43[3]},
      {stage2_44[18], stage2_44[19], stage2_44[20], stage2_44[21], stage2_44[22], stage2_44[23]},
      {stage3_46[3],stage3_45[3],stage3_44[5],stage3_43[22],stage3_42[35]}
   );
   gpc615_5 gpc7563 (
      {stage2_42[32], stage2_42[33], stage2_42[34], stage2_42[35], stage2_42[36]},
      {stage2_43[4]},
      {stage2_44[24], stage2_44[25], stage2_44[26], stage2_44[27], stage2_44[28], stage2_44[29]},
      {stage3_46[4],stage3_45[4],stage3_44[6],stage3_43[23],stage3_42[36]}
   );
   gpc615_5 gpc7564 (
      {stage2_42[37], stage2_42[38], stage2_42[39], stage2_42[40], stage2_42[41]},
      {stage2_43[5]},
      {stage2_44[30], stage2_44[31], stage2_44[32], stage2_44[33], stage2_44[34], stage2_44[35]},
      {stage3_46[5],stage3_45[5],stage3_44[7],stage3_43[24],stage3_42[37]}
   );
   gpc615_5 gpc7565 (
      {stage2_42[42], stage2_42[43], stage2_42[44], stage2_42[45], stage2_42[46]},
      {stage2_43[6]},
      {stage2_44[36], stage2_44[37], stage2_44[38], stage2_44[39], stage2_44[40], stage2_44[41]},
      {stage3_46[6],stage3_45[6],stage3_44[8],stage3_43[25],stage3_42[38]}
   );
   gpc615_5 gpc7566 (
      {stage2_42[47], stage2_42[48], stage2_42[49], stage2_42[50], stage2_42[51]},
      {stage2_43[7]},
      {stage2_44[42], stage2_44[43], stage2_44[44], stage2_44[45], stage2_44[46], stage2_44[47]},
      {stage3_46[7],stage3_45[7],stage3_44[9],stage3_43[26],stage3_42[39]}
   );
   gpc615_5 gpc7567 (
      {stage2_42[52], stage2_42[53], stage2_42[54], stage2_42[55], stage2_42[56]},
      {stage2_43[8]},
      {stage2_44[48], stage2_44[49], stage2_44[50], stage2_44[51], stage2_44[52], stage2_44[53]},
      {stage3_46[8],stage3_45[8],stage3_44[10],stage3_43[27],stage3_42[40]}
   );
   gpc615_5 gpc7568 (
      {stage2_42[57], stage2_42[58], stage2_42[59], stage2_42[60], stage2_42[61]},
      {stage2_43[9]},
      {stage2_44[54], stage2_44[55], stage2_44[56], stage2_44[57], stage2_44[58], stage2_44[59]},
      {stage3_46[9],stage3_45[9],stage3_44[11],stage3_43[28],stage3_42[41]}
   );
   gpc615_5 gpc7569 (
      {stage2_42[62], stage2_42[63], stage2_42[64], stage2_42[65], stage2_42[66]},
      {stage2_43[10]},
      {stage2_44[60], stage2_44[61], stage2_44[62], stage2_44[63], stage2_44[64], stage2_44[65]},
      {stage3_46[10],stage3_45[10],stage3_44[12],stage3_43[29],stage3_42[42]}
   );
   gpc615_5 gpc7570 (
      {stage2_42[67], stage2_42[68], stage2_42[69], stage2_42[70], stage2_42[71]},
      {stage2_43[11]},
      {stage2_44[66], stage2_44[67], stage2_44[68], stage2_44[69], stage2_44[70], stage2_44[71]},
      {stage3_46[11],stage3_45[11],stage3_44[13],stage3_43[30],stage3_42[43]}
   );
   gpc615_5 gpc7571 (
      {stage2_42[72], stage2_42[73], stage2_42[74], stage2_42[75], stage2_42[76]},
      {stage2_43[12]},
      {stage2_44[72], stage2_44[73], stage2_44[74], stage2_44[75], stage2_44[76], stage2_44[77]},
      {stage3_46[12],stage3_45[12],stage3_44[14],stage3_43[31],stage3_42[44]}
   );
   gpc615_5 gpc7572 (
      {stage2_42[77], stage2_42[78], stage2_42[79], stage2_42[80], stage2_42[81]},
      {stage2_43[13]},
      {stage2_44[78], stage2_44[79], stage2_44[80], stage2_44[81], stage2_44[82], stage2_44[83]},
      {stage3_46[13],stage3_45[13],stage3_44[15],stage3_43[32],stage3_42[45]}
   );
   gpc615_5 gpc7573 (
      {stage2_43[14], stage2_43[15], stage2_43[16], stage2_43[17], stage2_43[18]},
      {stage2_44[84]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[14],stage3_45[14],stage3_44[16],stage3_43[33]}
   );
   gpc615_5 gpc7574 (
      {stage2_43[19], stage2_43[20], stage2_43[21], stage2_43[22], stage2_43[23]},
      {stage2_44[85]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[15],stage3_45[15],stage3_44[17],stage3_43[34]}
   );
   gpc615_5 gpc7575 (
      {stage2_43[24], stage2_43[25], stage2_43[26], stage2_43[27], stage2_43[28]},
      {stage2_44[86]},
      {stage2_45[12], stage2_45[13], stage2_45[14], stage2_45[15], stage2_45[16], stage2_45[17]},
      {stage3_47[2],stage3_46[16],stage3_45[16],stage3_44[18],stage3_43[35]}
   );
   gpc615_5 gpc7576 (
      {stage2_43[29], stage2_43[30], stage2_43[31], stage2_43[32], stage2_43[33]},
      {stage2_44[87]},
      {stage2_45[18], stage2_45[19], stage2_45[20], stage2_45[21], stage2_45[22], stage2_45[23]},
      {stage3_47[3],stage3_46[17],stage3_45[17],stage3_44[19],stage3_43[36]}
   );
   gpc615_5 gpc7577 (
      {stage2_43[34], stage2_43[35], stage2_43[36], stage2_43[37], stage2_43[38]},
      {stage2_44[88]},
      {stage2_45[24], stage2_45[25], stage2_45[26], stage2_45[27], stage2_45[28], stage2_45[29]},
      {stage3_47[4],stage3_46[18],stage3_45[18],stage3_44[20],stage3_43[37]}
   );
   gpc615_5 gpc7578 (
      {stage2_43[39], stage2_43[40], stage2_43[41], stage2_43[42], stage2_43[43]},
      {stage2_44[89]},
      {stage2_45[30], stage2_45[31], stage2_45[32], stage2_45[33], stage2_45[34], stage2_45[35]},
      {stage3_47[5],stage3_46[19],stage3_45[19],stage3_44[21],stage3_43[38]}
   );
   gpc615_5 gpc7579 (
      {stage2_43[44], stage2_43[45], stage2_43[46], stage2_43[47], stage2_43[48]},
      {stage2_44[90]},
      {stage2_45[36], stage2_45[37], stage2_45[38], stage2_45[39], stage2_45[40], stage2_45[41]},
      {stage3_47[6],stage3_46[20],stage3_45[20],stage3_44[22],stage3_43[39]}
   );
   gpc615_5 gpc7580 (
      {stage2_43[49], stage2_43[50], stage2_43[51], stage2_43[52], stage2_43[53]},
      {stage2_44[91]},
      {stage2_45[42], stage2_45[43], stage2_45[44], stage2_45[45], stage2_45[46], stage2_45[47]},
      {stage3_47[7],stage3_46[21],stage3_45[21],stage3_44[23],stage3_43[40]}
   );
   gpc615_5 gpc7581 (
      {stage2_43[54], stage2_43[55], stage2_43[56], stage2_43[57], stage2_43[58]},
      {stage2_44[92]},
      {stage2_45[48], stage2_45[49], stage2_45[50], stage2_45[51], stage2_45[52], stage2_45[53]},
      {stage3_47[8],stage3_46[22],stage3_45[22],stage3_44[24],stage3_43[41]}
   );
   gpc615_5 gpc7582 (
      {stage2_43[59], stage2_43[60], stage2_43[61], stage2_43[62], stage2_43[63]},
      {stage2_44[93]},
      {stage2_45[54], stage2_45[55], stage2_45[56], stage2_45[57], stage2_45[58], stage2_45[59]},
      {stage3_47[9],stage3_46[23],stage3_45[23],stage3_44[25],stage3_43[42]}
   );
   gpc615_5 gpc7583 (
      {stage2_43[64], stage2_43[65], stage2_43[66], stage2_43[67], stage2_43[68]},
      {stage2_44[94]},
      {stage2_45[60], stage2_45[61], stage2_45[62], stage2_45[63], stage2_45[64], stage2_45[65]},
      {stage3_47[10],stage3_46[24],stage3_45[24],stage3_44[26],stage3_43[43]}
   );
   gpc615_5 gpc7584 (
      {stage2_43[69], stage2_43[70], stage2_43[71], stage2_43[72], stage2_43[73]},
      {stage2_44[95]},
      {stage2_45[66], stage2_45[67], stage2_45[68], stage2_45[69], stage2_45[70], stage2_45[71]},
      {stage3_47[11],stage3_46[25],stage3_45[25],stage3_44[27],stage3_43[44]}
   );
   gpc615_5 gpc7585 (
      {stage2_43[74], stage2_43[75], stage2_43[76], stage2_43[77], stage2_43[78]},
      {stage2_44[96]},
      {stage2_45[72], stage2_45[73], stage2_45[74], stage2_45[75], stage2_45[76], stage2_45[77]},
      {stage3_47[12],stage3_46[26],stage3_45[26],stage3_44[28],stage3_43[45]}
   );
   gpc606_5 gpc7586 (
      {stage2_44[97], stage2_44[98], stage2_44[99], stage2_44[100], stage2_44[101], stage2_44[102]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[13],stage3_46[27],stage3_45[27],stage3_44[29]}
   );
   gpc606_5 gpc7587 (
      {stage2_44[103], stage2_44[104], stage2_44[105], stage2_44[106], stage2_44[107], stage2_44[108]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[14],stage3_46[28],stage3_45[28],stage3_44[30]}
   );
   gpc606_5 gpc7588 (
      {stage2_45[78], stage2_45[79], stage2_45[80], stage2_45[81], stage2_45[82], stage2_45[83]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[2],stage3_47[15],stage3_46[29],stage3_45[29]}
   );
   gpc606_5 gpc7589 (
      {stage2_45[84], stage2_45[85], stage2_45[86], stage2_45[87], stage2_45[88], stage2_45[89]},
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10], stage2_47[11]},
      {stage3_49[1],stage3_48[3],stage3_47[16],stage3_46[30],stage3_45[30]}
   );
   gpc606_5 gpc7590 (
      {stage2_45[90], stage2_45[91], stage2_45[92], stage2_45[93], stage2_45[94], stage2_45[95]},
      {stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16], stage2_47[17]},
      {stage3_49[2],stage3_48[4],stage3_47[17],stage3_46[31],stage3_45[31]}
   );
   gpc606_5 gpc7591 (
      {stage2_45[96], stage2_45[97], stage2_45[98], stage2_45[99], stage2_45[100], stage2_45[101]},
      {stage2_47[18], stage2_47[19], stage2_47[20], stage2_47[21], stage2_47[22], stage2_47[23]},
      {stage3_49[3],stage3_48[5],stage3_47[18],stage3_46[32],stage3_45[32]}
   );
   gpc606_5 gpc7592 (
      {stage2_45[102], stage2_45[103], stage2_45[104], stage2_45[105], stage2_45[106], stage2_45[107]},
      {stage2_47[24], stage2_47[25], stage2_47[26], stage2_47[27], stage2_47[28], stage2_47[29]},
      {stage3_49[4],stage3_48[6],stage3_47[19],stage3_46[33],stage3_45[33]}
   );
   gpc1163_5 gpc7593 (
      {stage2_46[12], stage2_46[13], stage2_46[14]},
      {stage2_47[30], stage2_47[31], stage2_47[32], stage2_47[33], stage2_47[34], stage2_47[35]},
      {stage2_48[0]},
      {stage2_49[0]},
      {stage3_50[0],stage3_49[5],stage3_48[7],stage3_47[20],stage3_46[34]}
   );
   gpc1163_5 gpc7594 (
      {stage2_46[15], stage2_46[16], stage2_46[17]},
      {stage2_47[36], stage2_47[37], stage2_47[38], stage2_47[39], stage2_47[40], stage2_47[41]},
      {stage2_48[1]},
      {stage2_49[1]},
      {stage3_50[1],stage3_49[6],stage3_48[8],stage3_47[21],stage3_46[35]}
   );
   gpc615_5 gpc7595 (
      {stage2_46[18], stage2_46[19], stage2_46[20], stage2_46[21], stage2_46[22]},
      {stage2_47[42]},
      {stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5], stage2_48[6], stage2_48[7]},
      {stage3_50[2],stage3_49[7],stage3_48[9],stage3_47[22],stage3_46[36]}
   );
   gpc615_5 gpc7596 (
      {stage2_46[23], stage2_46[24], stage2_46[25], stage2_46[26], stage2_46[27]},
      {stage2_47[43]},
      {stage2_48[8], stage2_48[9], stage2_48[10], stage2_48[11], stage2_48[12], stage2_48[13]},
      {stage3_50[3],stage3_49[8],stage3_48[10],stage3_47[23],stage3_46[37]}
   );
   gpc615_5 gpc7597 (
      {stage2_46[28], stage2_46[29], stage2_46[30], stage2_46[31], stage2_46[32]},
      {stage2_47[44]},
      {stage2_48[14], stage2_48[15], stage2_48[16], stage2_48[17], stage2_48[18], stage2_48[19]},
      {stage3_50[4],stage3_49[9],stage3_48[11],stage3_47[24],stage3_46[38]}
   );
   gpc615_5 gpc7598 (
      {stage2_46[33], stage2_46[34], stage2_46[35], stage2_46[36], stage2_46[37]},
      {stage2_47[45]},
      {stage2_48[20], stage2_48[21], stage2_48[22], stage2_48[23], stage2_48[24], stage2_48[25]},
      {stage3_50[5],stage3_49[10],stage3_48[12],stage3_47[25],stage3_46[39]}
   );
   gpc615_5 gpc7599 (
      {stage2_46[38], stage2_46[39], stage2_46[40], stage2_46[41], stage2_46[42]},
      {stage2_47[46]},
      {stage2_48[26], stage2_48[27], stage2_48[28], stage2_48[29], stage2_48[30], stage2_48[31]},
      {stage3_50[6],stage3_49[11],stage3_48[13],stage3_47[26],stage3_46[40]}
   );
   gpc615_5 gpc7600 (
      {stage2_46[43], stage2_46[44], stage2_46[45], stage2_46[46], stage2_46[47]},
      {stage2_47[47]},
      {stage2_48[32], stage2_48[33], stage2_48[34], stage2_48[35], stage2_48[36], stage2_48[37]},
      {stage3_50[7],stage3_49[12],stage3_48[14],stage3_47[27],stage3_46[41]}
   );
   gpc615_5 gpc7601 (
      {stage2_46[48], stage2_46[49], stage2_46[50], stage2_46[51], stage2_46[52]},
      {stage2_47[48]},
      {stage2_48[38], stage2_48[39], stage2_48[40], stage2_48[41], stage2_48[42], stage2_48[43]},
      {stage3_50[8],stage3_49[13],stage3_48[15],stage3_47[28],stage3_46[42]}
   );
   gpc615_5 gpc7602 (
      {stage2_46[53], stage2_46[54], stage2_46[55], stage2_46[56], stage2_46[57]},
      {stage2_47[49]},
      {stage2_48[44], stage2_48[45], stage2_48[46], stage2_48[47], stage2_48[48], stage2_48[49]},
      {stage3_50[9],stage3_49[14],stage3_48[16],stage3_47[29],stage3_46[43]}
   );
   gpc615_5 gpc7603 (
      {stage2_46[58], stage2_46[59], stage2_46[60], stage2_46[61], stage2_46[62]},
      {stage2_47[50]},
      {stage2_48[50], stage2_48[51], stage2_48[52], stage2_48[53], stage2_48[54], stage2_48[55]},
      {stage3_50[10],stage3_49[15],stage3_48[17],stage3_47[30],stage3_46[44]}
   );
   gpc615_5 gpc7604 (
      {stage2_46[63], stage2_46[64], stage2_46[65], stage2_46[66], stage2_46[67]},
      {stage2_47[51]},
      {stage2_48[56], stage2_48[57], stage2_48[58], stage2_48[59], stage2_48[60], stage2_48[61]},
      {stage3_50[11],stage3_49[16],stage3_48[18],stage3_47[31],stage3_46[45]}
   );
   gpc615_5 gpc7605 (
      {stage2_46[68], stage2_46[69], stage2_46[70], stage2_46[71], stage2_46[72]},
      {stage2_47[52]},
      {stage2_48[62], stage2_48[63], stage2_48[64], stage2_48[65], stage2_48[66], stage2_48[67]},
      {stage3_50[12],stage3_49[17],stage3_48[19],stage3_47[32],stage3_46[46]}
   );
   gpc615_5 gpc7606 (
      {stage2_46[73], stage2_46[74], stage2_46[75], stage2_46[76], stage2_46[77]},
      {stage2_47[53]},
      {stage2_48[68], stage2_48[69], stage2_48[70], stage2_48[71], stage2_48[72], stage2_48[73]},
      {stage3_50[13],stage3_49[18],stage3_48[20],stage3_47[33],stage3_46[47]}
   );
   gpc615_5 gpc7607 (
      {stage2_47[54], stage2_47[55], stage2_47[56], stage2_47[57], stage2_47[58]},
      {stage2_48[74]},
      {stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5], stage2_49[6], stage2_49[7]},
      {stage3_51[0],stage3_50[14],stage3_49[19],stage3_48[21],stage3_47[34]}
   );
   gpc615_5 gpc7608 (
      {stage2_47[59], stage2_47[60], stage2_47[61], stage2_47[62], stage2_47[63]},
      {stage2_48[75]},
      {stage2_49[8], stage2_49[9], stage2_49[10], stage2_49[11], stage2_49[12], stage2_49[13]},
      {stage3_51[1],stage3_50[15],stage3_49[20],stage3_48[22],stage3_47[35]}
   );
   gpc615_5 gpc7609 (
      {stage2_47[64], stage2_47[65], stage2_47[66], stage2_47[67], stage2_47[68]},
      {stage2_48[76]},
      {stage2_49[14], stage2_49[15], stage2_49[16], stage2_49[17], stage2_49[18], stage2_49[19]},
      {stage3_51[2],stage3_50[16],stage3_49[21],stage3_48[23],stage3_47[36]}
   );
   gpc615_5 gpc7610 (
      {stage2_47[69], stage2_47[70], stage2_47[71], stage2_47[72], stage2_47[73]},
      {stage2_48[77]},
      {stage2_49[20], stage2_49[21], stage2_49[22], stage2_49[23], stage2_49[24], stage2_49[25]},
      {stage3_51[3],stage3_50[17],stage3_49[22],stage3_48[24],stage3_47[37]}
   );
   gpc615_5 gpc7611 (
      {stage2_47[74], stage2_47[75], stage2_47[76], stage2_47[77], stage2_47[78]},
      {stage2_48[78]},
      {stage2_49[26], stage2_49[27], stage2_49[28], stage2_49[29], stage2_49[30], stage2_49[31]},
      {stage3_51[4],stage3_50[18],stage3_49[23],stage3_48[25],stage3_47[38]}
   );
   gpc615_5 gpc7612 (
      {stage2_47[79], stage2_47[80], stage2_47[81], stage2_47[82], stage2_47[83]},
      {stage2_48[79]},
      {stage2_49[32], stage2_49[33], stage2_49[34], stage2_49[35], stage2_49[36], stage2_49[37]},
      {stage3_51[5],stage3_50[19],stage3_49[24],stage3_48[26],stage3_47[39]}
   );
   gpc615_5 gpc7613 (
      {stage2_47[84], stage2_47[85], stage2_47[86], stage2_47[87], stage2_47[88]},
      {stage2_48[80]},
      {stage2_49[38], stage2_49[39], stage2_49[40], stage2_49[41], stage2_49[42], stage2_49[43]},
      {stage3_51[6],stage3_50[20],stage3_49[25],stage3_48[27],stage3_47[40]}
   );
   gpc615_5 gpc7614 (
      {stage2_47[89], stage2_47[90], stage2_47[91], stage2_47[92], stage2_47[93]},
      {stage2_48[81]},
      {stage2_49[44], stage2_49[45], stage2_49[46], stage2_49[47], stage2_49[48], stage2_49[49]},
      {stage3_51[7],stage3_50[21],stage3_49[26],stage3_48[28],stage3_47[41]}
   );
   gpc615_5 gpc7615 (
      {stage2_47[94], stage2_47[95], stage2_47[96], stage2_47[97], stage2_47[98]},
      {stage2_48[82]},
      {stage2_49[50], stage2_49[51], stage2_49[52], stage2_49[53], stage2_49[54], stage2_49[55]},
      {stage3_51[8],stage3_50[22],stage3_49[27],stage3_48[29],stage3_47[42]}
   );
   gpc615_5 gpc7616 (
      {stage2_47[99], stage2_47[100], stage2_47[101], stage2_47[102], stage2_47[103]},
      {stage2_48[83]},
      {stage2_49[56], stage2_49[57], stage2_49[58], stage2_49[59], stage2_49[60], stage2_49[61]},
      {stage3_51[9],stage3_50[23],stage3_49[28],stage3_48[30],stage3_47[43]}
   );
   gpc606_5 gpc7617 (
      {stage2_48[84], stage2_48[85], stage2_48[86], stage2_48[87], stage2_48[88], stage2_48[89]},
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage3_52[0],stage3_51[10],stage3_50[24],stage3_49[29],stage3_48[31]}
   );
   gpc606_5 gpc7618 (
      {stage2_48[90], stage2_48[91], stage2_48[92], stage2_48[93], stage2_48[94], stage2_48[95]},
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9], stage2_50[10], stage2_50[11]},
      {stage3_52[1],stage3_51[11],stage3_50[25],stage3_49[30],stage3_48[32]}
   );
   gpc606_5 gpc7619 (
      {stage2_48[96], stage2_48[97], stage2_48[98], stage2_48[99], stage2_48[100], stage2_48[101]},
      {stage2_50[12], stage2_50[13], stage2_50[14], stage2_50[15], stage2_50[16], stage2_50[17]},
      {stage3_52[2],stage3_51[12],stage3_50[26],stage3_49[31],stage3_48[33]}
   );
   gpc606_5 gpc7620 (
      {stage2_48[102], stage2_48[103], stage2_48[104], stage2_48[105], stage2_48[106], stage2_48[107]},
      {stage2_50[18], stage2_50[19], stage2_50[20], stage2_50[21], stage2_50[22], stage2_50[23]},
      {stage3_52[3],stage3_51[13],stage3_50[27],stage3_49[32],stage3_48[34]}
   );
   gpc606_5 gpc7621 (
      {stage2_48[108], stage2_48[109], stage2_48[110], stage2_48[111], stage2_48[112], stage2_48[113]},
      {stage2_50[24], stage2_50[25], stage2_50[26], stage2_50[27], stage2_50[28], stage2_50[29]},
      {stage3_52[4],stage3_51[14],stage3_50[28],stage3_49[33],stage3_48[35]}
   );
   gpc606_5 gpc7622 (
      {stage2_48[114], stage2_48[115], stage2_48[116], stage2_48[117], stage2_48[118], stage2_48[119]},
      {stage2_50[30], stage2_50[31], stage2_50[32], stage2_50[33], stage2_50[34], stage2_50[35]},
      {stage3_52[5],stage3_51[15],stage3_50[29],stage3_49[34],stage3_48[36]}
   );
   gpc606_5 gpc7623 (
      {stage2_48[120], stage2_48[121], stage2_48[122], stage2_48[123], stage2_48[124], stage2_48[125]},
      {stage2_50[36], stage2_50[37], stage2_50[38], stage2_50[39], stage2_50[40], stage2_50[41]},
      {stage3_52[6],stage3_51[16],stage3_50[30],stage3_49[35],stage3_48[37]}
   );
   gpc606_5 gpc7624 (
      {stage2_49[62], stage2_49[63], stage2_49[64], stage2_49[65], stage2_49[66], stage2_49[67]},
      {stage2_51[0], stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5]},
      {stage3_53[0],stage3_52[7],stage3_51[17],stage3_50[31],stage3_49[36]}
   );
   gpc606_5 gpc7625 (
      {stage2_49[68], stage2_49[69], stage2_49[70], stage2_49[71], stage2_49[72], stage2_49[73]},
      {stage2_51[6], stage2_51[7], stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11]},
      {stage3_53[1],stage3_52[8],stage3_51[18],stage3_50[32],stage3_49[37]}
   );
   gpc606_5 gpc7626 (
      {stage2_49[74], stage2_49[75], stage2_49[76], stage2_49[77], stage2_49[78], stage2_49[79]},
      {stage2_51[12], stage2_51[13], stage2_51[14], stage2_51[15], stage2_51[16], stage2_51[17]},
      {stage3_53[2],stage3_52[9],stage3_51[19],stage3_50[33],stage3_49[38]}
   );
   gpc606_5 gpc7627 (
      {stage2_49[80], stage2_49[81], stage2_49[82], stage2_49[83], stage2_49[84], stage2_49[85]},
      {stage2_51[18], stage2_51[19], stage2_51[20], stage2_51[21], stage2_51[22], stage2_51[23]},
      {stage3_53[3],stage3_52[10],stage3_51[20],stage3_50[34],stage3_49[39]}
   );
   gpc615_5 gpc7628 (
      {stage2_49[86], stage2_49[87], stage2_49[88], stage2_49[89], stage2_49[90]},
      {stage2_50[42]},
      {stage2_51[24], stage2_51[25], stage2_51[26], stage2_51[27], stage2_51[28], stage2_51[29]},
      {stage3_53[4],stage3_52[11],stage3_51[21],stage3_50[35],stage3_49[40]}
   );
   gpc615_5 gpc7629 (
      {stage2_49[91], stage2_49[92], stage2_49[93], stage2_49[94], stage2_49[95]},
      {stage2_50[43]},
      {stage2_51[30], stage2_51[31], stage2_51[32], stage2_51[33], stage2_51[34], stage2_51[35]},
      {stage3_53[5],stage3_52[12],stage3_51[22],stage3_50[36],stage3_49[41]}
   );
   gpc615_5 gpc7630 (
      {stage2_50[44], stage2_50[45], stage2_50[46], stage2_50[47], stage2_50[48]},
      {stage2_51[36]},
      {stage2_52[0], stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5]},
      {stage3_54[0],stage3_53[6],stage3_52[13],stage3_51[23],stage3_50[37]}
   );
   gpc615_5 gpc7631 (
      {stage2_50[49], stage2_50[50], stage2_50[51], stage2_50[52], stage2_50[53]},
      {stage2_51[37]},
      {stage2_52[6], stage2_52[7], stage2_52[8], stage2_52[9], stage2_52[10], stage2_52[11]},
      {stage3_54[1],stage3_53[7],stage3_52[14],stage3_51[24],stage3_50[38]}
   );
   gpc615_5 gpc7632 (
      {stage2_50[54], stage2_50[55], stage2_50[56], stage2_50[57], stage2_50[58]},
      {stage2_51[38]},
      {stage2_52[12], stage2_52[13], stage2_52[14], stage2_52[15], stage2_52[16], stage2_52[17]},
      {stage3_54[2],stage3_53[8],stage3_52[15],stage3_51[25],stage3_50[39]}
   );
   gpc615_5 gpc7633 (
      {stage2_50[59], stage2_50[60], stage2_50[61], stage2_50[62], stage2_50[63]},
      {stage2_51[39]},
      {stage2_52[18], stage2_52[19], stage2_52[20], stage2_52[21], stage2_52[22], stage2_52[23]},
      {stage3_54[3],stage3_53[9],stage3_52[16],stage3_51[26],stage3_50[40]}
   );
   gpc615_5 gpc7634 (
      {stage2_50[64], stage2_50[65], stage2_50[66], stage2_50[67], stage2_50[68]},
      {stage2_51[40]},
      {stage2_52[24], stage2_52[25], stage2_52[26], stage2_52[27], stage2_52[28], stage2_52[29]},
      {stage3_54[4],stage3_53[10],stage3_52[17],stage3_51[27],stage3_50[41]}
   );
   gpc615_5 gpc7635 (
      {stage2_50[69], stage2_50[70], stage2_50[71], stage2_50[72], stage2_50[73]},
      {stage2_51[41]},
      {stage2_52[30], stage2_52[31], stage2_52[32], stage2_52[33], stage2_52[34], stage2_52[35]},
      {stage3_54[5],stage3_53[11],stage3_52[18],stage3_51[28],stage3_50[42]}
   );
   gpc615_5 gpc7636 (
      {stage2_50[74], stage2_50[75], stage2_50[76], stage2_50[77], stage2_50[78]},
      {stage2_51[42]},
      {stage2_52[36], stage2_52[37], stage2_52[38], stage2_52[39], stage2_52[40], stage2_52[41]},
      {stage3_54[6],stage3_53[12],stage3_52[19],stage3_51[29],stage3_50[43]}
   );
   gpc615_5 gpc7637 (
      {stage2_50[79], stage2_50[80], stage2_50[81], stage2_50[82], stage2_50[83]},
      {stage2_51[43]},
      {stage2_52[42], stage2_52[43], stage2_52[44], stage2_52[45], stage2_52[46], stage2_52[47]},
      {stage3_54[7],stage3_53[13],stage3_52[20],stage3_51[30],stage3_50[44]}
   );
   gpc615_5 gpc7638 (
      {stage2_51[44], stage2_51[45], stage2_51[46], stage2_51[47], stage2_51[48]},
      {stage2_52[48]},
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage3_55[0],stage3_54[8],stage3_53[14],stage3_52[21],stage3_51[31]}
   );
   gpc615_5 gpc7639 (
      {stage2_51[49], stage2_51[50], stage2_51[51], stage2_51[52], stage2_51[53]},
      {stage2_52[49]},
      {stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10], stage2_53[11]},
      {stage3_55[1],stage3_54[9],stage3_53[15],stage3_52[22],stage3_51[32]}
   );
   gpc615_5 gpc7640 (
      {stage2_51[54], stage2_51[55], stage2_51[56], stage2_51[57], stage2_51[58]},
      {stage2_52[50]},
      {stage2_53[12], stage2_53[13], stage2_53[14], stage2_53[15], stage2_53[16], stage2_53[17]},
      {stage3_55[2],stage3_54[10],stage3_53[16],stage3_52[23],stage3_51[33]}
   );
   gpc606_5 gpc7641 (
      {stage2_52[51], stage2_52[52], stage2_52[53], stage2_52[54], stage2_52[55], stage2_52[56]},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage3_56[0],stage3_55[3],stage3_54[11],stage3_53[17],stage3_52[24]}
   );
   gpc606_5 gpc7642 (
      {stage2_52[57], stage2_52[58], stage2_52[59], stage2_52[60], stage2_52[61], stage2_52[62]},
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage3_56[1],stage3_55[4],stage3_54[12],stage3_53[18],stage3_52[25]}
   );
   gpc606_5 gpc7643 (
      {stage2_52[63], stage2_52[64], stage2_52[65], stage2_52[66], stage2_52[67], stage2_52[68]},
      {stage2_54[12], stage2_54[13], stage2_54[14], stage2_54[15], stage2_54[16], stage2_54[17]},
      {stage3_56[2],stage3_55[5],stage3_54[13],stage3_53[19],stage3_52[26]}
   );
   gpc606_5 gpc7644 (
      {stage2_53[18], stage2_53[19], stage2_53[20], stage2_53[21], stage2_53[22], stage2_53[23]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[3],stage3_55[6],stage3_54[14],stage3_53[20]}
   );
   gpc606_5 gpc7645 (
      {stage2_53[24], stage2_53[25], stage2_53[26], stage2_53[27], stage2_53[28], stage2_53[29]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[4],stage3_55[7],stage3_54[15],stage3_53[21]}
   );
   gpc606_5 gpc7646 (
      {stage2_53[30], stage2_53[31], stage2_53[32], stage2_53[33], stage2_53[34], stage2_53[35]},
      {stage2_55[12], stage2_55[13], stage2_55[14], stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage3_57[2],stage3_56[5],stage3_55[8],stage3_54[16],stage3_53[22]}
   );
   gpc606_5 gpc7647 (
      {stage2_53[36], stage2_53[37], stage2_53[38], stage2_53[39], stage2_53[40], stage2_53[41]},
      {stage2_55[18], stage2_55[19], stage2_55[20], stage2_55[21], stage2_55[22], stage2_55[23]},
      {stage3_57[3],stage3_56[6],stage3_55[9],stage3_54[17],stage3_53[23]}
   );
   gpc606_5 gpc7648 (
      {stage2_53[42], stage2_53[43], stage2_53[44], stage2_53[45], stage2_53[46], stage2_53[47]},
      {stage2_55[24], stage2_55[25], stage2_55[26], stage2_55[27], stage2_55[28], stage2_55[29]},
      {stage3_57[4],stage3_56[7],stage3_55[10],stage3_54[18],stage3_53[24]}
   );
   gpc606_5 gpc7649 (
      {stage2_53[48], stage2_53[49], stage2_53[50], stage2_53[51], stage2_53[52], stage2_53[53]},
      {stage2_55[30], stage2_55[31], stage2_55[32], stage2_55[33], stage2_55[34], stage2_55[35]},
      {stage3_57[5],stage3_56[8],stage3_55[11],stage3_54[19],stage3_53[25]}
   );
   gpc615_5 gpc7650 (
      {stage2_53[54], stage2_53[55], stage2_53[56], stage2_53[57], stage2_53[58]},
      {stage2_54[18]},
      {stage2_55[36], stage2_55[37], stage2_55[38], stage2_55[39], stage2_55[40], stage2_55[41]},
      {stage3_57[6],stage3_56[9],stage3_55[12],stage3_54[20],stage3_53[26]}
   );
   gpc615_5 gpc7651 (
      {stage2_53[59], stage2_53[60], stage2_53[61], stage2_53[62], stage2_53[63]},
      {stage2_54[19]},
      {stage2_55[42], stage2_55[43], stage2_55[44], stage2_55[45], stage2_55[46], stage2_55[47]},
      {stage3_57[7],stage3_56[10],stage3_55[13],stage3_54[21],stage3_53[27]}
   );
   gpc615_5 gpc7652 (
      {stage2_53[64], stage2_53[65], stage2_53[66], stage2_53[67], stage2_53[68]},
      {stage2_54[20]},
      {stage2_55[48], stage2_55[49], stage2_55[50], stage2_55[51], stage2_55[52], stage2_55[53]},
      {stage3_57[8],stage3_56[11],stage3_55[14],stage3_54[22],stage3_53[28]}
   );
   gpc615_5 gpc7653 (
      {stage2_54[21], stage2_54[22], stage2_54[23], stage2_54[24], stage2_54[25]},
      {stage2_55[54]},
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5]},
      {stage3_58[0],stage3_57[9],stage3_56[12],stage3_55[15],stage3_54[23]}
   );
   gpc615_5 gpc7654 (
      {stage2_54[26], stage2_54[27], stage2_54[28], stage2_54[29], stage2_54[30]},
      {stage2_55[55]},
      {stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9], stage2_56[10], stage2_56[11]},
      {stage3_58[1],stage3_57[10],stage3_56[13],stage3_55[16],stage3_54[24]}
   );
   gpc615_5 gpc7655 (
      {stage2_54[31], stage2_54[32], stage2_54[33], stage2_54[34], stage2_54[35]},
      {stage2_55[56]},
      {stage2_56[12], stage2_56[13], stage2_56[14], stage2_56[15], stage2_56[16], stage2_56[17]},
      {stage3_58[2],stage3_57[11],stage3_56[14],stage3_55[17],stage3_54[25]}
   );
   gpc615_5 gpc7656 (
      {stage2_54[36], stage2_54[37], stage2_54[38], stage2_54[39], stage2_54[40]},
      {stage2_55[57]},
      {stage2_56[18], stage2_56[19], stage2_56[20], stage2_56[21], stage2_56[22], stage2_56[23]},
      {stage3_58[3],stage3_57[12],stage3_56[15],stage3_55[18],stage3_54[26]}
   );
   gpc615_5 gpc7657 (
      {stage2_54[41], stage2_54[42], stage2_54[43], stage2_54[44], stage2_54[45]},
      {stage2_55[58]},
      {stage2_56[24], stage2_56[25], stage2_56[26], stage2_56[27], stage2_56[28], stage2_56[29]},
      {stage3_58[4],stage3_57[13],stage3_56[16],stage3_55[19],stage3_54[27]}
   );
   gpc615_5 gpc7658 (
      {stage2_54[46], stage2_54[47], stage2_54[48], stage2_54[49], stage2_54[50]},
      {stage2_55[59]},
      {stage2_56[30], stage2_56[31], stage2_56[32], stage2_56[33], stage2_56[34], stage2_56[35]},
      {stage3_58[5],stage3_57[14],stage3_56[17],stage3_55[20],stage3_54[28]}
   );
   gpc615_5 gpc7659 (
      {stage2_54[51], stage2_54[52], stage2_54[53], stage2_54[54], stage2_54[55]},
      {stage2_55[60]},
      {stage2_56[36], stage2_56[37], stage2_56[38], stage2_56[39], stage2_56[40], stage2_56[41]},
      {stage3_58[6],stage3_57[15],stage3_56[18],stage3_55[21],stage3_54[29]}
   );
   gpc615_5 gpc7660 (
      {stage2_54[56], stage2_54[57], stage2_54[58], stage2_54[59], stage2_54[60]},
      {stage2_55[61]},
      {stage2_56[42], stage2_56[43], stage2_56[44], stage2_56[45], stage2_56[46], stage2_56[47]},
      {stage3_58[7],stage3_57[16],stage3_56[19],stage3_55[22],stage3_54[30]}
   );
   gpc615_5 gpc7661 (
      {stage2_54[61], stage2_54[62], stage2_54[63], stage2_54[64], stage2_54[65]},
      {stage2_55[62]},
      {stage2_56[48], stage2_56[49], stage2_56[50], stage2_56[51], stage2_56[52], stage2_56[53]},
      {stage3_58[8],stage3_57[17],stage3_56[20],stage3_55[23],stage3_54[31]}
   );
   gpc615_5 gpc7662 (
      {stage2_54[66], stage2_54[67], stage2_54[68], stage2_54[69], stage2_54[70]},
      {stage2_55[63]},
      {stage2_56[54], stage2_56[55], stage2_56[56], stage2_56[57], stage2_56[58], stage2_56[59]},
      {stage3_58[9],stage3_57[18],stage3_56[21],stage3_55[24],stage3_54[32]}
   );
   gpc615_5 gpc7663 (
      {stage2_54[71], stage2_54[72], stage2_54[73], stage2_54[74], stage2_54[75]},
      {stage2_55[64]},
      {stage2_56[60], stage2_56[61], stage2_56[62], stage2_56[63], stage2_56[64], stage2_56[65]},
      {stage3_58[10],stage3_57[19],stage3_56[22],stage3_55[25],stage3_54[33]}
   );
   gpc615_5 gpc7664 (
      {stage2_54[76], stage2_54[77], stage2_54[78], stage2_54[79], stage2_54[80]},
      {stage2_55[65]},
      {stage2_56[66], stage2_56[67], stage2_56[68], stage2_56[69], stage2_56[70], stage2_56[71]},
      {stage3_58[11],stage3_57[20],stage3_56[23],stage3_55[26],stage3_54[34]}
   );
   gpc615_5 gpc7665 (
      {stage2_54[81], stage2_54[82], stage2_54[83], stage2_54[84], stage2_54[85]},
      {stage2_55[66]},
      {stage2_56[72], stage2_56[73], stage2_56[74], stage2_56[75], stage2_56[76], stage2_56[77]},
      {stage3_58[12],stage3_57[21],stage3_56[24],stage3_55[27],stage3_54[35]}
   );
   gpc615_5 gpc7666 (
      {stage2_54[86], stage2_54[87], stage2_54[88], stage2_54[89], stage2_54[90]},
      {stage2_55[67]},
      {stage2_56[78], stage2_56[79], stage2_56[80], stage2_56[81], stage2_56[82], stage2_56[83]},
      {stage3_58[13],stage3_57[22],stage3_56[25],stage3_55[28],stage3_54[36]}
   );
   gpc615_5 gpc7667 (
      {stage2_54[91], stage2_54[92], stage2_54[93], stage2_54[94], stage2_54[95]},
      {stage2_55[68]},
      {stage2_56[84], stage2_56[85], stage2_56[86], stage2_56[87], stage2_56[88], stage2_56[89]},
      {stage3_58[14],stage3_57[23],stage3_56[26],stage3_55[29],stage3_54[37]}
   );
   gpc615_5 gpc7668 (
      {stage2_54[96], stage2_54[97], stage2_54[98], stage2_54[99], 1'b0},
      {stage2_55[69]},
      {stage2_56[90], stage2_56[91], stage2_56[92], stage2_56[93], stage2_56[94], stage2_56[95]},
      {stage3_58[15],stage3_57[24],stage3_56[27],stage3_55[30],stage3_54[38]}
   );
   gpc615_5 gpc7669 (
      {stage2_56[96], stage2_56[97], stage2_56[98], stage2_56[99], stage2_56[100]},
      {stage2_57[0]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[0],stage3_58[16],stage3_57[25],stage3_56[28]}
   );
   gpc615_5 gpc7670 (
      {stage2_56[101], stage2_56[102], stage2_56[103], stage2_56[104], stage2_56[105]},
      {stage2_57[1]},
      {stage2_58[6], stage2_58[7], stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage3_60[1],stage3_59[1],stage3_58[17],stage3_57[26],stage3_56[29]}
   );
   gpc615_5 gpc7671 (
      {stage2_56[106], stage2_56[107], stage2_56[108], stage2_56[109], stage2_56[110]},
      {stage2_57[2]},
      {stage2_58[12], stage2_58[13], stage2_58[14], stage2_58[15], stage2_58[16], stage2_58[17]},
      {stage3_60[2],stage3_59[2],stage3_58[18],stage3_57[27],stage3_56[30]}
   );
   gpc615_5 gpc7672 (
      {stage2_56[111], stage2_56[112], stage2_56[113], stage2_56[114], 1'b0},
      {stage2_57[3]},
      {stage2_58[18], stage2_58[19], stage2_58[20], stage2_58[21], stage2_58[22], stage2_58[23]},
      {stage3_60[3],stage3_59[3],stage3_58[19],stage3_57[28],stage3_56[31]}
   );
   gpc207_4 gpc7673 (
      {stage2_57[4], stage2_57[5], stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10]},
      {stage2_59[0], stage2_59[1]},
      {stage3_60[4],stage3_59[4],stage3_58[20],stage3_57[29]}
   );
   gpc606_5 gpc7674 (
      {stage2_57[11], stage2_57[12], stage2_57[13], stage2_57[14], stage2_57[15], stage2_57[16]},
      {stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5], stage2_59[6], stage2_59[7]},
      {stage3_61[0],stage3_60[5],stage3_59[5],stage3_58[21],stage3_57[30]}
   );
   gpc606_5 gpc7675 (
      {stage2_57[17], stage2_57[18], stage2_57[19], stage2_57[20], stage2_57[21], stage2_57[22]},
      {stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11], stage2_59[12], stage2_59[13]},
      {stage3_61[1],stage3_60[6],stage3_59[6],stage3_58[22],stage3_57[31]}
   );
   gpc606_5 gpc7676 (
      {stage2_57[23], stage2_57[24], stage2_57[25], stage2_57[26], stage2_57[27], stage2_57[28]},
      {stage2_59[14], stage2_59[15], stage2_59[16], stage2_59[17], stage2_59[18], stage2_59[19]},
      {stage3_61[2],stage3_60[7],stage3_59[7],stage3_58[23],stage3_57[32]}
   );
   gpc615_5 gpc7677 (
      {stage2_57[29], stage2_57[30], stage2_57[31], stage2_57[32], stage2_57[33]},
      {stage2_58[24]},
      {stage2_59[20], stage2_59[21], stage2_59[22], stage2_59[23], stage2_59[24], stage2_59[25]},
      {stage3_61[3],stage3_60[8],stage3_59[8],stage3_58[24],stage3_57[33]}
   );
   gpc615_5 gpc7678 (
      {stage2_57[34], stage2_57[35], stage2_57[36], stage2_57[37], stage2_57[38]},
      {stage2_58[25]},
      {stage2_59[26], stage2_59[27], stage2_59[28], stage2_59[29], stage2_59[30], stage2_59[31]},
      {stage3_61[4],stage3_60[9],stage3_59[9],stage3_58[25],stage3_57[34]}
   );
   gpc615_5 gpc7679 (
      {stage2_57[39], stage2_57[40], stage2_57[41], stage2_57[42], stage2_57[43]},
      {stage2_58[26]},
      {stage2_59[32], stage2_59[33], stage2_59[34], stage2_59[35], stage2_59[36], stage2_59[37]},
      {stage3_61[5],stage3_60[10],stage3_59[10],stage3_58[26],stage3_57[35]}
   );
   gpc615_5 gpc7680 (
      {stage2_57[44], stage2_57[45], stage2_57[46], stage2_57[47], stage2_57[48]},
      {stage2_58[27]},
      {stage2_59[38], stage2_59[39], stage2_59[40], stage2_59[41], stage2_59[42], stage2_59[43]},
      {stage3_61[6],stage3_60[11],stage3_59[11],stage3_58[27],stage3_57[36]}
   );
   gpc615_5 gpc7681 (
      {stage2_58[28], stage2_58[29], stage2_58[30], stage2_58[31], stage2_58[32]},
      {stage2_59[44]},
      {stage2_60[0], stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5]},
      {stage3_62[0],stage3_61[7],stage3_60[12],stage3_59[12],stage3_58[28]}
   );
   gpc615_5 gpc7682 (
      {stage2_58[33], stage2_58[34], stage2_58[35], stage2_58[36], stage2_58[37]},
      {stage2_59[45]},
      {stage2_60[6], stage2_60[7], stage2_60[8], stage2_60[9], stage2_60[10], stage2_60[11]},
      {stage3_62[1],stage3_61[8],stage3_60[13],stage3_59[13],stage3_58[29]}
   );
   gpc615_5 gpc7683 (
      {stage2_58[38], stage2_58[39], stage2_58[40], stage2_58[41], stage2_58[42]},
      {stage2_59[46]},
      {stage2_60[12], stage2_60[13], stage2_60[14], stage2_60[15], stage2_60[16], stage2_60[17]},
      {stage3_62[2],stage3_61[9],stage3_60[14],stage3_59[14],stage3_58[30]}
   );
   gpc615_5 gpc7684 (
      {stage2_58[43], stage2_58[44], stage2_58[45], stage2_58[46], stage2_58[47]},
      {stage2_59[47]},
      {stage2_60[18], stage2_60[19], stage2_60[20], stage2_60[21], stage2_60[22], stage2_60[23]},
      {stage3_62[3],stage3_61[10],stage3_60[15],stage3_59[15],stage3_58[31]}
   );
   gpc615_5 gpc7685 (
      {stage2_58[48], stage2_58[49], stage2_58[50], stage2_58[51], stage2_58[52]},
      {stage2_59[48]},
      {stage2_60[24], stage2_60[25], stage2_60[26], stage2_60[27], stage2_60[28], stage2_60[29]},
      {stage3_62[4],stage3_61[11],stage3_60[16],stage3_59[16],stage3_58[32]}
   );
   gpc615_5 gpc7686 (
      {stage2_58[53], stage2_58[54], stage2_58[55], stage2_58[56], stage2_58[57]},
      {stage2_59[49]},
      {stage2_60[30], stage2_60[31], stage2_60[32], stage2_60[33], stage2_60[34], stage2_60[35]},
      {stage3_62[5],stage3_61[12],stage3_60[17],stage3_59[17],stage3_58[33]}
   );
   gpc615_5 gpc7687 (
      {stage2_59[50], stage2_59[51], stage2_59[52], stage2_59[53], stage2_59[54]},
      {stage2_60[36]},
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage3_63[0],stage3_62[6],stage3_61[13],stage3_60[18],stage3_59[18]}
   );
   gpc615_5 gpc7688 (
      {stage2_59[55], stage2_59[56], stage2_59[57], stage2_59[58], stage2_59[59]},
      {stage2_60[37]},
      {stage2_61[6], stage2_61[7], stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11]},
      {stage3_63[1],stage3_62[7],stage3_61[14],stage3_60[19],stage3_59[19]}
   );
   gpc615_5 gpc7689 (
      {stage2_59[60], stage2_59[61], stage2_59[62], stage2_59[63], stage2_59[64]},
      {stage2_60[38]},
      {stage2_61[12], stage2_61[13], stage2_61[14], stage2_61[15], stage2_61[16], stage2_61[17]},
      {stage3_63[2],stage3_62[8],stage3_61[15],stage3_60[20],stage3_59[20]}
   );
   gpc615_5 gpc7690 (
      {stage2_59[65], stage2_59[66], stage2_59[67], stage2_59[68], stage2_59[69]},
      {stage2_60[39]},
      {stage2_61[18], stage2_61[19], stage2_61[20], stage2_61[21], stage2_61[22], stage2_61[23]},
      {stage3_63[3],stage3_62[9],stage3_61[16],stage3_60[21],stage3_59[21]}
   );
   gpc615_5 gpc7691 (
      {stage2_59[70], stage2_59[71], stage2_59[72], stage2_59[73], stage2_59[74]},
      {stage2_60[40]},
      {stage2_61[24], stage2_61[25], stage2_61[26], stage2_61[27], stage2_61[28], stage2_61[29]},
      {stage3_63[4],stage3_62[10],stage3_61[17],stage3_60[22],stage3_59[22]}
   );
   gpc615_5 gpc7692 (
      {stage2_59[75], stage2_59[76], stage2_59[77], stage2_59[78], stage2_59[79]},
      {stage2_60[41]},
      {stage2_61[30], stage2_61[31], stage2_61[32], stage2_61[33], stage2_61[34], stage2_61[35]},
      {stage3_63[5],stage3_62[11],stage3_61[18],stage3_60[23],stage3_59[23]}
   );
   gpc615_5 gpc7693 (
      {stage2_59[80], stage2_59[81], stage2_59[82], stage2_59[83], stage2_59[84]},
      {stage2_60[42]},
      {stage2_61[36], stage2_61[37], stage2_61[38], stage2_61[39], stage2_61[40], stage2_61[41]},
      {stage3_63[6],stage3_62[12],stage3_61[19],stage3_60[24],stage3_59[24]}
   );
   gpc606_5 gpc7694 (
      {stage2_60[43], stage2_60[44], stage2_60[45], stage2_60[46], stage2_60[47], stage2_60[48]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[7],stage3_62[13],stage3_61[20],stage3_60[25]}
   );
   gpc606_5 gpc7695 (
      {stage2_60[49], stage2_60[50], stage2_60[51], stage2_60[52], stage2_60[53], stage2_60[54]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage3_64[1],stage3_63[8],stage3_62[14],stage3_61[21],stage3_60[26]}
   );
   gpc606_5 gpc7696 (
      {stage2_60[55], stage2_60[56], stage2_60[57], stage2_60[58], stage2_60[59], stage2_60[60]},
      {stage2_62[12], stage2_62[13], stage2_62[14], stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage3_64[2],stage3_63[9],stage3_62[15],stage3_61[22],stage3_60[27]}
   );
   gpc606_5 gpc7697 (
      {stage2_60[61], stage2_60[62], stage2_60[63], stage2_60[64], stage2_60[65], stage2_60[66]},
      {stage2_62[18], stage2_62[19], stage2_62[20], stage2_62[21], stage2_62[22], stage2_62[23]},
      {stage3_64[3],stage3_63[10],stage3_62[16],stage3_61[23],stage3_60[28]}
   );
   gpc606_5 gpc7698 (
      {stage2_60[67], stage2_60[68], stage2_60[69], stage2_60[70], stage2_60[71], stage2_60[72]},
      {stage2_62[24], stage2_62[25], stage2_62[26], stage2_62[27], stage2_62[28], stage2_62[29]},
      {stage3_64[4],stage3_63[11],stage3_62[17],stage3_61[24],stage3_60[29]}
   );
   gpc606_5 gpc7699 (
      {stage2_61[42], stage2_61[43], stage2_61[44], stage2_61[45], stage2_61[46], stage2_61[47]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[5],stage3_63[12],stage3_62[18],stage3_61[25]}
   );
   gpc615_5 gpc7700 (
      {stage2_62[30], stage2_62[31], stage2_62[32], stage2_62[33], stage2_62[34]},
      {stage2_63[6]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[1],stage3_64[6],stage3_63[13],stage3_62[19]}
   );
   gpc615_5 gpc7701 (
      {stage2_62[35], stage2_62[36], stage2_62[37], stage2_62[38], stage2_62[39]},
      {stage2_63[7]},
      {stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9], stage2_64[10], stage2_64[11]},
      {stage3_66[1],stage3_65[2],stage3_64[7],stage3_63[14],stage3_62[20]}
   );
   gpc615_5 gpc7702 (
      {stage2_62[40], stage2_62[41], stage2_62[42], stage2_62[43], stage2_62[44]},
      {stage2_63[8]},
      {stage2_64[12], stage2_64[13], stage2_64[14], stage2_64[15], stage2_64[16], stage2_64[17]},
      {stage3_66[2],stage3_65[3],stage3_64[8],stage3_63[15],stage3_62[21]}
   );
   gpc615_5 gpc7703 (
      {stage2_62[45], stage2_62[46], stage2_62[47], stage2_62[48], stage2_62[49]},
      {stage2_63[9]},
      {stage2_64[18], stage2_64[19], stage2_64[20], stage2_64[21], stage2_64[22], stage2_64[23]},
      {stage3_66[3],stage3_65[4],stage3_64[9],stage3_63[16],stage3_62[22]}
   );
   gpc615_5 gpc7704 (
      {stage2_62[50], stage2_62[51], stage2_62[52], stage2_62[53], stage2_62[54]},
      {stage2_63[10]},
      {stage2_64[24], stage2_64[25], stage2_64[26], stage2_64[27], stage2_64[28], stage2_64[29]},
      {stage3_66[4],stage3_65[5],stage3_64[10],stage3_63[17],stage3_62[23]}
   );
   gpc615_5 gpc7705 (
      {stage2_62[55], stage2_62[56], stage2_62[57], stage2_62[58], stage2_62[59]},
      {stage2_63[11]},
      {stage2_64[30], stage2_64[31], stage2_64[32], stage2_64[33], stage2_64[34], stage2_64[35]},
      {stage3_66[5],stage3_65[6],stage3_64[11],stage3_63[18],stage3_62[24]}
   );
   gpc615_5 gpc7706 (
      {stage2_62[60], stage2_62[61], stage2_62[62], stage2_62[63], stage2_62[64]},
      {stage2_63[12]},
      {stage2_64[36], stage2_64[37], stage2_64[38], stage2_64[39], stage2_64[40], stage2_64[41]},
      {stage3_66[6],stage3_65[7],stage3_64[12],stage3_63[19],stage3_62[25]}
   );
   gpc615_5 gpc7707 (
      {stage2_62[65], stage2_62[66], stage2_62[67], stage2_62[68], stage2_62[69]},
      {stage2_63[13]},
      {stage2_64[42], stage2_64[43], stage2_64[44], stage2_64[45], stage2_64[46], stage2_64[47]},
      {stage3_66[7],stage3_65[8],stage3_64[13],stage3_63[20],stage3_62[26]}
   );
   gpc615_5 gpc7708 (
      {stage2_62[70], stage2_62[71], stage2_62[72], stage2_62[73], stage2_62[74]},
      {stage2_63[14]},
      {stage2_64[48], stage2_64[49], stage2_64[50], stage2_64[51], stage2_64[52], stage2_64[53]},
      {stage3_66[8],stage3_65[9],stage3_64[14],stage3_63[21],stage3_62[27]}
   );
   gpc615_5 gpc7709 (
      {stage2_62[75], stage2_62[76], stage2_62[77], stage2_62[78], stage2_62[79]},
      {stage2_63[15]},
      {stage2_64[54], stage2_64[55], stage2_64[56], stage2_64[57], stage2_64[58], stage2_64[59]},
      {stage3_66[9],stage3_65[10],stage3_64[15],stage3_63[22],stage3_62[28]}
   );
   gpc615_5 gpc7710 (
      {stage2_62[80], stage2_62[81], stage2_62[82], stage2_62[83], stage2_62[84]},
      {stage2_63[16]},
      {stage2_64[60], stage2_64[61], stage2_64[62], stage2_64[63], stage2_64[64], stage2_64[65]},
      {stage3_66[10],stage3_65[11],stage3_64[16],stage3_63[23],stage3_62[29]}
   );
   gpc615_5 gpc7711 (
      {stage2_62[85], stage2_62[86], stage2_62[87], stage2_62[88], stage2_62[89]},
      {stage2_63[17]},
      {stage2_64[66], stage2_64[67], stage2_64[68], stage2_64[69], stage2_64[70], stage2_64[71]},
      {stage3_66[11],stage3_65[12],stage3_64[17],stage3_63[24],stage3_62[30]}
   );
   gpc615_5 gpc7712 (
      {stage2_62[90], stage2_62[91], stage2_62[92], stage2_62[93], stage2_62[94]},
      {stage2_63[18]},
      {stage2_64[72], stage2_64[73], stage2_64[74], stage2_64[75], stage2_64[76], stage2_64[77]},
      {stage3_66[12],stage3_65[13],stage3_64[18],stage3_63[25],stage3_62[31]}
   );
   gpc615_5 gpc7713 (
      {stage2_62[95], stage2_62[96], stage2_62[97], stage2_62[98], stage2_62[99]},
      {stage2_63[19]},
      {stage2_64[78], stage2_64[79], stage2_64[80], stage2_64[81], stage2_64[82], stage2_64[83]},
      {stage3_66[13],stage3_65[14],stage3_64[19],stage3_63[26],stage3_62[32]}
   );
   gpc615_5 gpc7714 (
      {stage2_62[100], stage2_62[101], stage2_62[102], stage2_62[103], stage2_62[104]},
      {stage2_63[20]},
      {stage2_64[84], stage2_64[85], stage2_64[86], stage2_64[87], stage2_64[88], stage2_64[89]},
      {stage3_66[14],stage3_65[15],stage3_64[20],stage3_63[27],stage3_62[33]}
   );
   gpc117_4 gpc7715 (
      {stage2_63[21], stage2_63[22], stage2_63[23], stage2_63[24], stage2_63[25], stage2_63[26], stage2_63[27]},
      {stage2_64[90]},
      {stage2_65[0]},
      {stage3_66[15],stage3_65[16],stage3_64[21],stage3_63[28]}
   );
   gpc117_4 gpc7716 (
      {stage2_63[28], stage2_63[29], stage2_63[30], stage2_63[31], stage2_63[32], stage2_63[33], stage2_63[34]},
      {stage2_64[91]},
      {stage2_65[1]},
      {stage3_66[16],stage3_65[17],stage3_64[22],stage3_63[29]}
   );
   gpc117_4 gpc7717 (
      {stage2_63[35], stage2_63[36], stage2_63[37], stage2_63[38], stage2_63[39], stage2_63[40], stage2_63[41]},
      {stage2_64[92]},
      {stage2_65[2]},
      {stage3_66[17],stage3_65[18],stage3_64[23],stage3_63[30]}
   );
   gpc606_5 gpc7718 (
      {stage2_63[42], stage2_63[43], stage2_63[44], stage2_63[45], stage2_63[46], stage2_63[47]},
      {stage2_65[3], stage2_65[4], stage2_65[5], stage2_65[6], stage2_65[7], stage2_65[8]},
      {stage3_67[0],stage3_66[18],stage3_65[19],stage3_64[24],stage3_63[31]}
   );
   gpc606_5 gpc7719 (
      {stage2_63[48], stage2_63[49], stage2_63[50], stage2_63[51], stage2_63[52], stage2_63[53]},
      {stage2_65[9], stage2_65[10], stage2_65[11], stage2_65[12], stage2_65[13], stage2_65[14]},
      {stage3_67[1],stage3_66[19],stage3_65[20],stage3_64[25],stage3_63[32]}
   );
   gpc606_5 gpc7720 (
      {stage2_63[54], stage2_63[55], stage2_63[56], stage2_63[57], stage2_63[58], stage2_63[59]},
      {stage2_65[15], stage2_65[16], stage2_65[17], stage2_65[18], stage2_65[19], stage2_65[20]},
      {stage3_67[2],stage3_66[20],stage3_65[21],stage3_64[26],stage3_63[33]}
   );
   gpc606_5 gpc7721 (
      {stage2_63[60], stage2_63[61], stage2_63[62], stage2_63[63], stage2_63[64], stage2_63[65]},
      {stage2_65[21], stage2_65[22], stage2_65[23], stage2_65[24], stage2_65[25], stage2_65[26]},
      {stage3_67[3],stage3_66[21],stage3_65[22],stage3_64[27],stage3_63[34]}
   );
   gpc606_5 gpc7722 (
      {stage2_63[66], stage2_63[67], stage2_63[68], stage2_63[69], stage2_63[70], stage2_63[71]},
      {stage2_65[27], stage2_65[28], stage2_65[29], stage2_65[30], stage2_65[31], stage2_65[32]},
      {stage3_67[4],stage3_66[22],stage3_65[23],stage3_64[28],stage3_63[35]}
   );
   gpc606_5 gpc7723 (
      {stage2_63[72], stage2_63[73], stage2_63[74], stage2_63[75], stage2_63[76], stage2_63[77]},
      {stage2_65[33], stage2_65[34], stage2_65[35], stage2_65[36], stage2_65[37], stage2_65[38]},
      {stage3_67[5],stage3_66[23],stage3_65[24],stage3_64[29],stage3_63[36]}
   );
   gpc606_5 gpc7724 (
      {stage2_63[78], stage2_63[79], stage2_63[80], stage2_63[81], stage2_63[82], stage2_63[83]},
      {stage2_65[39], stage2_65[40], stage2_65[41], stage2_65[42], stage2_65[43], stage2_65[44]},
      {stage3_67[6],stage3_66[24],stage3_65[25],stage3_64[30],stage3_63[37]}
   );
   gpc606_5 gpc7725 (
      {stage2_63[84], stage2_63[85], stage2_63[86], stage2_63[87], stage2_63[88], stage2_63[89]},
      {stage2_65[45], stage2_65[46], stage2_65[47], stage2_65[48], stage2_65[49], stage2_65[50]},
      {stage3_67[7],stage3_66[25],stage3_65[26],stage3_64[31],stage3_63[38]}
   );
   gpc606_5 gpc7726 (
      {stage2_64[93], stage2_64[94], stage2_64[95], stage2_64[96], stage2_64[97], stage2_64[98]},
      {stage2_66[0], stage2_66[1], stage2_66[2], stage2_66[3], stage2_66[4], stage2_66[5]},
      {stage3_68[0],stage3_67[8],stage3_66[26],stage3_65[27],stage3_64[32]}
   );
   gpc606_5 gpc7727 (
      {stage2_64[99], stage2_64[100], stage2_64[101], stage2_64[102], stage2_64[103], stage2_64[104]},
      {stage2_66[6], stage2_66[7], stage2_66[8], stage2_66[9], stage2_66[10], stage2_66[11]},
      {stage3_68[1],stage3_67[9],stage3_66[27],stage3_65[28],stage3_64[33]}
   );
   gpc606_5 gpc7728 (
      {stage2_64[105], stage2_64[106], stage2_64[107], stage2_64[108], stage2_64[109], stage2_64[110]},
      {stage2_66[12], stage2_66[13], stage2_66[14], stage2_66[15], stage2_66[16], stage2_66[17]},
      {stage3_68[2],stage3_67[10],stage3_66[28],stage3_65[29],stage3_64[34]}
   );
   gpc606_5 gpc7729 (
      {stage2_64[111], stage2_64[112], stage2_64[113], stage2_64[114], stage2_64[115], stage2_64[116]},
      {stage2_66[18], stage2_66[19], stage2_66[20], stage2_66[21], stage2_66[22], stage2_66[23]},
      {stage3_68[3],stage3_67[11],stage3_66[29],stage3_65[30],stage3_64[35]}
   );
   gpc606_5 gpc7730 (
      {stage2_64[117], stage2_64[118], stage2_64[119], stage2_64[120], stage2_64[121], stage2_64[122]},
      {stage2_66[24], stage2_66[25], stage2_66[26], stage2_66[27], stage2_66[28], stage2_66[29]},
      {stage3_68[4],stage3_67[12],stage3_66[30],stage3_65[31],stage3_64[36]}
   );
   gpc606_5 gpc7731 (
      {stage2_64[123], stage2_64[124], stage2_64[125], stage2_64[126], stage2_64[127], stage2_64[128]},
      {stage2_66[30], stage2_66[31], stage2_66[32], stage2_66[33], stage2_66[34], stage2_66[35]},
      {stage3_68[5],stage3_67[13],stage3_66[31],stage3_65[32],stage3_64[37]}
   );
   gpc1_1 gpc7732 (
      {stage2_0[23]},
      {stage3_0[6]}
   );
   gpc1_1 gpc7733 (
      {stage2_0[24]},
      {stage3_0[7]}
   );
   gpc1_1 gpc7734 (
      {stage2_0[25]},
      {stage3_0[8]}
   );
   gpc1_1 gpc7735 (
      {stage2_0[26]},
      {stage3_0[9]}
   );
   gpc1_1 gpc7736 (
      {stage2_0[27]},
      {stage3_0[10]}
   );
   gpc1_1 gpc7737 (
      {stage2_0[28]},
      {stage3_0[11]}
   );
   gpc1_1 gpc7738 (
      {stage2_0[29]},
      {stage3_0[12]}
   );
   gpc1_1 gpc7739 (
      {stage2_0[30]},
      {stage3_0[13]}
   );
   gpc1_1 gpc7740 (
      {stage2_0[31]},
      {stage3_0[14]}
   );
   gpc1_1 gpc7741 (
      {stage2_0[32]},
      {stage3_0[15]}
   );
   gpc1_1 gpc7742 (
      {stage2_0[33]},
      {stage3_0[16]}
   );
   gpc1_1 gpc7743 (
      {stage2_0[34]},
      {stage3_0[17]}
   );
   gpc1_1 gpc7744 (
      {stage2_0[35]},
      {stage3_0[18]}
   );
   gpc1_1 gpc7745 (
      {stage2_0[36]},
      {stage3_0[19]}
   );
   gpc1_1 gpc7746 (
      {stage2_0[37]},
      {stage3_0[20]}
   );
   gpc1_1 gpc7747 (
      {stage2_1[42]},
      {stage3_1[10]}
   );
   gpc1_1 gpc7748 (
      {stage2_1[43]},
      {stage3_1[11]}
   );
   gpc1_1 gpc7749 (
      {stage2_1[44]},
      {stage3_1[12]}
   );
   gpc1_1 gpc7750 (
      {stage2_1[45]},
      {stage3_1[13]}
   );
   gpc1_1 gpc7751 (
      {stage2_1[46]},
      {stage3_1[14]}
   );
   gpc1_1 gpc7752 (
      {stage2_1[47]},
      {stage3_1[15]}
   );
   gpc1_1 gpc7753 (
      {stage2_1[48]},
      {stage3_1[16]}
   );
   gpc1_1 gpc7754 (
      {stage2_1[49]},
      {stage3_1[17]}
   );
   gpc1_1 gpc7755 (
      {stage2_1[50]},
      {stage3_1[18]}
   );
   gpc1_1 gpc7756 (
      {stage2_1[51]},
      {stage3_1[19]}
   );
   gpc1_1 gpc7757 (
      {stage2_1[52]},
      {stage3_1[20]}
   );
   gpc1_1 gpc7758 (
      {stage2_1[53]},
      {stage3_1[21]}
   );
   gpc1_1 gpc7759 (
      {stage2_2[32]},
      {stage3_2[12]}
   );
   gpc1_1 gpc7760 (
      {stage2_2[33]},
      {stage3_2[13]}
   );
   gpc1_1 gpc7761 (
      {stage2_2[34]},
      {stage3_2[14]}
   );
   gpc1_1 gpc7762 (
      {stage2_2[35]},
      {stage3_2[15]}
   );
   gpc1_1 gpc7763 (
      {stage2_2[36]},
      {stage3_2[16]}
   );
   gpc1_1 gpc7764 (
      {stage2_2[37]},
      {stage3_2[17]}
   );
   gpc1_1 gpc7765 (
      {stage2_2[38]},
      {stage3_2[18]}
   );
   gpc1_1 gpc7766 (
      {stage2_2[39]},
      {stage3_2[19]}
   );
   gpc1_1 gpc7767 (
      {stage2_2[40]},
      {stage3_2[20]}
   );
   gpc1_1 gpc7768 (
      {stage2_2[41]},
      {stage3_2[21]}
   );
   gpc1_1 gpc7769 (
      {stage2_2[42]},
      {stage3_2[22]}
   );
   gpc1_1 gpc7770 (
      {stage2_2[43]},
      {stage3_2[23]}
   );
   gpc1_1 gpc7771 (
      {stage2_2[44]},
      {stage3_2[24]}
   );
   gpc1_1 gpc7772 (
      {stage2_2[45]},
      {stage3_2[25]}
   );
   gpc1_1 gpc7773 (
      {stage2_2[46]},
      {stage3_2[26]}
   );
   gpc1_1 gpc7774 (
      {stage2_2[47]},
      {stage3_2[27]}
   );
   gpc1_1 gpc7775 (
      {stage2_2[48]},
      {stage3_2[28]}
   );
   gpc1_1 gpc7776 (
      {stage2_2[49]},
      {stage3_2[29]}
   );
   gpc1_1 gpc7777 (
      {stage2_2[50]},
      {stage3_2[30]}
   );
   gpc1_1 gpc7778 (
      {stage2_2[51]},
      {stage3_2[31]}
   );
   gpc1_1 gpc7779 (
      {stage2_2[52]},
      {stage3_2[32]}
   );
   gpc1_1 gpc7780 (
      {stage2_2[53]},
      {stage3_2[33]}
   );
   gpc1_1 gpc7781 (
      {stage2_2[54]},
      {stage3_2[34]}
   );
   gpc1_1 gpc7782 (
      {stage2_2[55]},
      {stage3_2[35]}
   );
   gpc1_1 gpc7783 (
      {stage2_2[56]},
      {stage3_2[36]}
   );
   gpc1_1 gpc7784 (
      {stage2_2[57]},
      {stage3_2[37]}
   );
   gpc1_1 gpc7785 (
      {stage2_2[58]},
      {stage3_2[38]}
   );
   gpc1_1 gpc7786 (
      {stage2_2[59]},
      {stage3_2[39]}
   );
   gpc1_1 gpc7787 (
      {stage2_2[60]},
      {stage3_2[40]}
   );
   gpc1_1 gpc7788 (
      {stage2_2[61]},
      {stage3_2[41]}
   );
   gpc1_1 gpc7789 (
      {stage2_2[62]},
      {stage3_2[42]}
   );
   gpc1_1 gpc7790 (
      {stage2_4[29]},
      {stage3_4[29]}
   );
   gpc1_1 gpc7791 (
      {stage2_4[30]},
      {stage3_4[30]}
   );
   gpc1_1 gpc7792 (
      {stage2_4[31]},
      {stage3_4[31]}
   );
   gpc1_1 gpc7793 (
      {stage2_4[32]},
      {stage3_4[32]}
   );
   gpc1_1 gpc7794 (
      {stage2_4[33]},
      {stage3_4[33]}
   );
   gpc1_1 gpc7795 (
      {stage2_4[34]},
      {stage3_4[34]}
   );
   gpc1_1 gpc7796 (
      {stage2_4[35]},
      {stage3_4[35]}
   );
   gpc1_1 gpc7797 (
      {stage2_4[36]},
      {stage3_4[36]}
   );
   gpc1_1 gpc7798 (
      {stage2_4[37]},
      {stage3_4[37]}
   );
   gpc1_1 gpc7799 (
      {stage2_4[38]},
      {stage3_4[38]}
   );
   gpc1_1 gpc7800 (
      {stage2_4[39]},
      {stage3_4[39]}
   );
   gpc1_1 gpc7801 (
      {stage2_4[40]},
      {stage3_4[40]}
   );
   gpc1_1 gpc7802 (
      {stage2_4[41]},
      {stage3_4[41]}
   );
   gpc1_1 gpc7803 (
      {stage2_4[42]},
      {stage3_4[42]}
   );
   gpc1_1 gpc7804 (
      {stage2_4[43]},
      {stage3_4[43]}
   );
   gpc1_1 gpc7805 (
      {stage2_4[44]},
      {stage3_4[44]}
   );
   gpc1_1 gpc7806 (
      {stage2_4[45]},
      {stage3_4[45]}
   );
   gpc1_1 gpc7807 (
      {stage2_4[46]},
      {stage3_4[46]}
   );
   gpc1_1 gpc7808 (
      {stage2_4[47]},
      {stage3_4[47]}
   );
   gpc1_1 gpc7809 (
      {stage2_4[48]},
      {stage3_4[48]}
   );
   gpc1_1 gpc7810 (
      {stage2_4[49]},
      {stage3_4[49]}
   );
   gpc1_1 gpc7811 (
      {stage2_4[50]},
      {stage3_4[50]}
   );
   gpc1_1 gpc7812 (
      {stage2_4[51]},
      {stage3_4[51]}
   );
   gpc1_1 gpc7813 (
      {stage2_4[52]},
      {stage3_4[52]}
   );
   gpc1_1 gpc7814 (
      {stage2_4[53]},
      {stage3_4[53]}
   );
   gpc1_1 gpc7815 (
      {stage2_4[54]},
      {stage3_4[54]}
   );
   gpc1_1 gpc7816 (
      {stage2_4[55]},
      {stage3_4[55]}
   );
   gpc1_1 gpc7817 (
      {stage2_4[56]},
      {stage3_4[56]}
   );
   gpc1_1 gpc7818 (
      {stage2_4[57]},
      {stage3_4[57]}
   );
   gpc1_1 gpc7819 (
      {stage2_4[58]},
      {stage3_4[58]}
   );
   gpc1_1 gpc7820 (
      {stage2_4[59]},
      {stage3_4[59]}
   );
   gpc1_1 gpc7821 (
      {stage2_4[60]},
      {stage3_4[60]}
   );
   gpc1_1 gpc7822 (
      {stage2_4[61]},
      {stage3_4[61]}
   );
   gpc1_1 gpc7823 (
      {stage2_4[62]},
      {stage3_4[62]}
   );
   gpc1_1 gpc7824 (
      {stage2_4[63]},
      {stage3_4[63]}
   );
   gpc1_1 gpc7825 (
      {stage2_4[64]},
      {stage3_4[64]}
   );
   gpc1_1 gpc7826 (
      {stage2_4[65]},
      {stage3_4[65]}
   );
   gpc1_1 gpc7827 (
      {stage2_4[66]},
      {stage3_4[66]}
   );
   gpc1_1 gpc7828 (
      {stage2_4[67]},
      {stage3_4[67]}
   );
   gpc1_1 gpc7829 (
      {stage2_4[68]},
      {stage3_4[68]}
   );
   gpc1_1 gpc7830 (
      {stage2_4[69]},
      {stage3_4[69]}
   );
   gpc1_1 gpc7831 (
      {stage2_4[70]},
      {stage3_4[70]}
   );
   gpc1_1 gpc7832 (
      {stage2_4[71]},
      {stage3_4[71]}
   );
   gpc1_1 gpc7833 (
      {stage2_4[72]},
      {stage3_4[72]}
   );
   gpc1_1 gpc7834 (
      {stage2_4[73]},
      {stage3_4[73]}
   );
   gpc1_1 gpc7835 (
      {stage2_4[74]},
      {stage3_4[74]}
   );
   gpc1_1 gpc7836 (
      {stage2_4[75]},
      {stage3_4[75]}
   );
   gpc1_1 gpc7837 (
      {stage2_4[76]},
      {stage3_4[76]}
   );
   gpc1_1 gpc7838 (
      {stage2_4[77]},
      {stage3_4[77]}
   );
   gpc1_1 gpc7839 (
      {stage2_4[78]},
      {stage3_4[78]}
   );
   gpc1_1 gpc7840 (
      {stage2_4[79]},
      {stage3_4[79]}
   );
   gpc1_1 gpc7841 (
      {stage2_4[80]},
      {stage3_4[80]}
   );
   gpc1_1 gpc7842 (
      {stage2_4[81]},
      {stage3_4[81]}
   );
   gpc1_1 gpc7843 (
      {stage2_4[82]},
      {stage3_4[82]}
   );
   gpc1_1 gpc7844 (
      {stage2_4[83]},
      {stage3_4[83]}
   );
   gpc1_1 gpc7845 (
      {stage2_4[84]},
      {stage3_4[84]}
   );
   gpc1_1 gpc7846 (
      {stage2_4[85]},
      {stage3_4[85]}
   );
   gpc1_1 gpc7847 (
      {stage2_4[86]},
      {stage3_4[86]}
   );
   gpc1_1 gpc7848 (
      {stage2_4[87]},
      {stage3_4[87]}
   );
   gpc1_1 gpc7849 (
      {stage2_4[88]},
      {stage3_4[88]}
   );
   gpc1_1 gpc7850 (
      {stage2_4[89]},
      {stage3_4[89]}
   );
   gpc1_1 gpc7851 (
      {stage2_4[90]},
      {stage3_4[90]}
   );
   gpc1_1 gpc7852 (
      {stage2_4[91]},
      {stage3_4[91]}
   );
   gpc1_1 gpc7853 (
      {stage2_4[92]},
      {stage3_4[92]}
   );
   gpc1_1 gpc7854 (
      {stage2_4[93]},
      {stage3_4[93]}
   );
   gpc1_1 gpc7855 (
      {stage2_4[94]},
      {stage3_4[94]}
   );
   gpc1_1 gpc7856 (
      {stage2_4[95]},
      {stage3_4[95]}
   );
   gpc1_1 gpc7857 (
      {stage2_4[96]},
      {stage3_4[96]}
   );
   gpc1_1 gpc7858 (
      {stage2_4[97]},
      {stage3_4[97]}
   );
   gpc1_1 gpc7859 (
      {stage2_4[98]},
      {stage3_4[98]}
   );
   gpc1_1 gpc7860 (
      {stage2_4[99]},
      {stage3_4[99]}
   );
   gpc1_1 gpc7861 (
      {stage2_4[100]},
      {stage3_4[100]}
   );
   gpc1_1 gpc7862 (
      {stage2_4[101]},
      {stage3_4[101]}
   );
   gpc1_1 gpc7863 (
      {stage2_4[102]},
      {stage3_4[102]}
   );
   gpc1_1 gpc7864 (
      {stage2_4[103]},
      {stage3_4[103]}
   );
   gpc1_1 gpc7865 (
      {stage2_4[104]},
      {stage3_4[104]}
   );
   gpc1_1 gpc7866 (
      {stage2_4[105]},
      {stage3_4[105]}
   );
   gpc1_1 gpc7867 (
      {stage2_4[106]},
      {stage3_4[106]}
   );
   gpc1_1 gpc7868 (
      {stage2_4[107]},
      {stage3_4[107]}
   );
   gpc1_1 gpc7869 (
      {stage2_4[108]},
      {stage3_4[108]}
   );
   gpc1_1 gpc7870 (
      {stage2_4[109]},
      {stage3_4[109]}
   );
   gpc1_1 gpc7871 (
      {stage2_4[110]},
      {stage3_4[110]}
   );
   gpc1_1 gpc7872 (
      {stage2_4[111]},
      {stage3_4[111]}
   );
   gpc1_1 gpc7873 (
      {stage2_5[126]},
      {stage3_5[27]}
   );
   gpc1_1 gpc7874 (
      {stage2_5[127]},
      {stage3_5[28]}
   );
   gpc1_1 gpc7875 (
      {stage2_5[128]},
      {stage3_5[29]}
   );
   gpc1_1 gpc7876 (
      {stage2_5[129]},
      {stage3_5[30]}
   );
   gpc1_1 gpc7877 (
      {stage2_5[130]},
      {stage3_5[31]}
   );
   gpc1_1 gpc7878 (
      {stage2_5[131]},
      {stage3_5[32]}
   );
   gpc1_1 gpc7879 (
      {stage2_5[132]},
      {stage3_5[33]}
   );
   gpc1_1 gpc7880 (
      {stage2_5[133]},
      {stage3_5[34]}
   );
   gpc1_1 gpc7881 (
      {stage2_5[134]},
      {stage3_5[35]}
   );
   gpc1_1 gpc7882 (
      {stage2_5[135]},
      {stage3_5[36]}
   );
   gpc1_1 gpc7883 (
      {stage2_5[136]},
      {stage3_5[37]}
   );
   gpc1_1 gpc7884 (
      {stage2_5[137]},
      {stage3_5[38]}
   );
   gpc1_1 gpc7885 (
      {stage2_5[138]},
      {stage3_5[39]}
   );
   gpc1_1 gpc7886 (
      {stage2_5[139]},
      {stage3_5[40]}
   );
   gpc1_1 gpc7887 (
      {stage2_5[140]},
      {stage3_5[41]}
   );
   gpc1_1 gpc7888 (
      {stage2_5[141]},
      {stage3_5[42]}
   );
   gpc1_1 gpc7889 (
      {stage2_5[142]},
      {stage3_5[43]}
   );
   gpc1_1 gpc7890 (
      {stage2_5[143]},
      {stage3_5[44]}
   );
   gpc1_1 gpc7891 (
      {stage2_5[144]},
      {stage3_5[45]}
   );
   gpc1_1 gpc7892 (
      {stage2_5[145]},
      {stage3_5[46]}
   );
   gpc1_1 gpc7893 (
      {stage2_5[146]},
      {stage3_5[47]}
   );
   gpc1_1 gpc7894 (
      {stage2_5[147]},
      {stage3_5[48]}
   );
   gpc1_1 gpc7895 (
      {stage2_5[148]},
      {stage3_5[49]}
   );
   gpc1_1 gpc7896 (
      {stage2_5[149]},
      {stage3_5[50]}
   );
   gpc1_1 gpc7897 (
      {stage2_5[150]},
      {stage3_5[51]}
   );
   gpc1_1 gpc7898 (
      {stage2_5[151]},
      {stage3_5[52]}
   );
   gpc1_1 gpc7899 (
      {stage2_6[46]},
      {stage3_6[32]}
   );
   gpc1_1 gpc7900 (
      {stage2_6[47]},
      {stage3_6[33]}
   );
   gpc1_1 gpc7901 (
      {stage2_6[48]},
      {stage3_6[34]}
   );
   gpc1_1 gpc7902 (
      {stage2_6[49]},
      {stage3_6[35]}
   );
   gpc1_1 gpc7903 (
      {stage2_6[50]},
      {stage3_6[36]}
   );
   gpc1_1 gpc7904 (
      {stage2_6[51]},
      {stage3_6[37]}
   );
   gpc1_1 gpc7905 (
      {stage2_6[52]},
      {stage3_6[38]}
   );
   gpc1_1 gpc7906 (
      {stage2_6[53]},
      {stage3_6[39]}
   );
   gpc1_1 gpc7907 (
      {stage2_6[54]},
      {stage3_6[40]}
   );
   gpc1_1 gpc7908 (
      {stage2_6[55]},
      {stage3_6[41]}
   );
   gpc1_1 gpc7909 (
      {stage2_6[56]},
      {stage3_6[42]}
   );
   gpc1_1 gpc7910 (
      {stage2_6[57]},
      {stage3_6[43]}
   );
   gpc1_1 gpc7911 (
      {stage2_6[58]},
      {stage3_6[44]}
   );
   gpc1_1 gpc7912 (
      {stage2_6[59]},
      {stage3_6[45]}
   );
   gpc1_1 gpc7913 (
      {stage2_6[60]},
      {stage3_6[46]}
   );
   gpc1_1 gpc7914 (
      {stage2_6[61]},
      {stage3_6[47]}
   );
   gpc1_1 gpc7915 (
      {stage2_6[62]},
      {stage3_6[48]}
   );
   gpc1_1 gpc7916 (
      {stage2_6[63]},
      {stage3_6[49]}
   );
   gpc1_1 gpc7917 (
      {stage2_6[64]},
      {stage3_6[50]}
   );
   gpc1_1 gpc7918 (
      {stage2_6[65]},
      {stage3_6[51]}
   );
   gpc1_1 gpc7919 (
      {stage2_6[66]},
      {stage3_6[52]}
   );
   gpc1_1 gpc7920 (
      {stage2_6[67]},
      {stage3_6[53]}
   );
   gpc1_1 gpc7921 (
      {stage2_6[68]},
      {stage3_6[54]}
   );
   gpc1_1 gpc7922 (
      {stage2_6[69]},
      {stage3_6[55]}
   );
   gpc1_1 gpc7923 (
      {stage2_6[70]},
      {stage3_6[56]}
   );
   gpc1_1 gpc7924 (
      {stage2_6[71]},
      {stage3_6[57]}
   );
   gpc1_1 gpc7925 (
      {stage2_6[72]},
      {stage3_6[58]}
   );
   gpc1_1 gpc7926 (
      {stage2_6[73]},
      {stage3_6[59]}
   );
   gpc1_1 gpc7927 (
      {stage2_6[74]},
      {stage3_6[60]}
   );
   gpc1_1 gpc7928 (
      {stage2_6[75]},
      {stage3_6[61]}
   );
   gpc1_1 gpc7929 (
      {stage2_6[76]},
      {stage3_6[62]}
   );
   gpc1_1 gpc7930 (
      {stage2_6[77]},
      {stage3_6[63]}
   );
   gpc1_1 gpc7931 (
      {stage2_6[78]},
      {stage3_6[64]}
   );
   gpc1_1 gpc7932 (
      {stage2_6[79]},
      {stage3_6[65]}
   );
   gpc1_1 gpc7933 (
      {stage2_6[80]},
      {stage3_6[66]}
   );
   gpc1_1 gpc7934 (
      {stage2_6[81]},
      {stage3_6[67]}
   );
   gpc1_1 gpc7935 (
      {stage2_6[82]},
      {stage3_6[68]}
   );
   gpc1_1 gpc7936 (
      {stage2_6[83]},
      {stage3_6[69]}
   );
   gpc1_1 gpc7937 (
      {stage2_6[84]},
      {stage3_6[70]}
   );
   gpc1_1 gpc7938 (
      {stage2_6[85]},
      {stage3_6[71]}
   );
   gpc1_1 gpc7939 (
      {stage2_6[86]},
      {stage3_6[72]}
   );
   gpc1_1 gpc7940 (
      {stage2_6[87]},
      {stage3_6[73]}
   );
   gpc1_1 gpc7941 (
      {stage2_6[88]},
      {stage3_6[74]}
   );
   gpc1_1 gpc7942 (
      {stage2_6[89]},
      {stage3_6[75]}
   );
   gpc1_1 gpc7943 (
      {stage2_6[90]},
      {stage3_6[76]}
   );
   gpc1_1 gpc7944 (
      {stage2_6[91]},
      {stage3_6[77]}
   );
   gpc1_1 gpc7945 (
      {stage2_7[57]},
      {stage3_7[35]}
   );
   gpc1_1 gpc7946 (
      {stage2_7[58]},
      {stage3_7[36]}
   );
   gpc1_1 gpc7947 (
      {stage2_7[59]},
      {stage3_7[37]}
   );
   gpc1_1 gpc7948 (
      {stage2_7[60]},
      {stage3_7[38]}
   );
   gpc1_1 gpc7949 (
      {stage2_7[61]},
      {stage3_7[39]}
   );
   gpc1_1 gpc7950 (
      {stage2_7[62]},
      {stage3_7[40]}
   );
   gpc1_1 gpc7951 (
      {stage2_7[63]},
      {stage3_7[41]}
   );
   gpc1_1 gpc7952 (
      {stage2_7[64]},
      {stage3_7[42]}
   );
   gpc1_1 gpc7953 (
      {stage2_7[65]},
      {stage3_7[43]}
   );
   gpc1_1 gpc7954 (
      {stage2_7[66]},
      {stage3_7[44]}
   );
   gpc1_1 gpc7955 (
      {stage2_7[67]},
      {stage3_7[45]}
   );
   gpc1_1 gpc7956 (
      {stage2_7[68]},
      {stage3_7[46]}
   );
   gpc1_1 gpc7957 (
      {stage2_7[69]},
      {stage3_7[47]}
   );
   gpc1_1 gpc7958 (
      {stage2_7[70]},
      {stage3_7[48]}
   );
   gpc1_1 gpc7959 (
      {stage2_7[71]},
      {stage3_7[49]}
   );
   gpc1_1 gpc7960 (
      {stage2_7[72]},
      {stage3_7[50]}
   );
   gpc1_1 gpc7961 (
      {stage2_10[117]},
      {stage3_10[53]}
   );
   gpc1_1 gpc7962 (
      {stage2_10[118]},
      {stage3_10[54]}
   );
   gpc1_1 gpc7963 (
      {stage2_10[119]},
      {stage3_10[55]}
   );
   gpc1_1 gpc7964 (
      {stage2_10[120]},
      {stage3_10[56]}
   );
   gpc1_1 gpc7965 (
      {stage2_10[121]},
      {stage3_10[57]}
   );
   gpc1_1 gpc7966 (
      {stage2_10[122]},
      {stage3_10[58]}
   );
   gpc1_1 gpc7967 (
      {stage2_10[123]},
      {stage3_10[59]}
   );
   gpc1_1 gpc7968 (
      {stage2_10[124]},
      {stage3_10[60]}
   );
   gpc1_1 gpc7969 (
      {stage2_10[125]},
      {stage3_10[61]}
   );
   gpc1_1 gpc7970 (
      {stage2_10[126]},
      {stage3_10[62]}
   );
   gpc1_1 gpc7971 (
      {stage2_10[127]},
      {stage3_10[63]}
   );
   gpc1_1 gpc7972 (
      {stage2_10[128]},
      {stage3_10[64]}
   );
   gpc1_1 gpc7973 (
      {stage2_10[129]},
      {stage3_10[65]}
   );
   gpc1_1 gpc7974 (
      {stage2_10[130]},
      {stage3_10[66]}
   );
   gpc1_1 gpc7975 (
      {stage2_10[131]},
      {stage3_10[67]}
   );
   gpc1_1 gpc7976 (
      {stage2_10[132]},
      {stage3_10[68]}
   );
   gpc1_1 gpc7977 (
      {stage2_10[133]},
      {stage3_10[69]}
   );
   gpc1_1 gpc7978 (
      {stage2_10[134]},
      {stage3_10[70]}
   );
   gpc1_1 gpc7979 (
      {stage2_10[135]},
      {stage3_10[71]}
   );
   gpc1_1 gpc7980 (
      {stage2_10[136]},
      {stage3_10[72]}
   );
   gpc1_1 gpc7981 (
      {stage2_10[137]},
      {stage3_10[73]}
   );
   gpc1_1 gpc7982 (
      {stage2_10[138]},
      {stage3_10[74]}
   );
   gpc1_1 gpc7983 (
      {stage2_10[139]},
      {stage3_10[75]}
   );
   gpc1_1 gpc7984 (
      {stage2_10[140]},
      {stage3_10[76]}
   );
   gpc1_1 gpc7985 (
      {stage2_10[141]},
      {stage3_10[77]}
   );
   gpc1_1 gpc7986 (
      {stage2_10[142]},
      {stage3_10[78]}
   );
   gpc1_1 gpc7987 (
      {stage2_10[143]},
      {stage3_10[79]}
   );
   gpc1_1 gpc7988 (
      {stage2_10[144]},
      {stage3_10[80]}
   );
   gpc1_1 gpc7989 (
      {stage2_10[145]},
      {stage3_10[81]}
   );
   gpc1_1 gpc7990 (
      {stage2_10[146]},
      {stage3_10[82]}
   );
   gpc1_1 gpc7991 (
      {stage2_10[147]},
      {stage3_10[83]}
   );
   gpc1_1 gpc7992 (
      {stage2_10[148]},
      {stage3_10[84]}
   );
   gpc1_1 gpc7993 (
      {stage2_10[149]},
      {stage3_10[85]}
   );
   gpc1_1 gpc7994 (
      {stage2_10[150]},
      {stage3_10[86]}
   );
   gpc1_1 gpc7995 (
      {stage2_10[151]},
      {stage3_10[87]}
   );
   gpc1_1 gpc7996 (
      {stage2_10[152]},
      {stage3_10[88]}
   );
   gpc1_1 gpc7997 (
      {stage2_10[153]},
      {stage3_10[89]}
   );
   gpc1_1 gpc7998 (
      {stage2_10[154]},
      {stage3_10[90]}
   );
   gpc1_1 gpc7999 (
      {stage2_10[155]},
      {stage3_10[91]}
   );
   gpc1_1 gpc8000 (
      {stage2_10[156]},
      {stage3_10[92]}
   );
   gpc1_1 gpc8001 (
      {stage2_10[157]},
      {stage3_10[93]}
   );
   gpc1_1 gpc8002 (
      {stage2_10[158]},
      {stage3_10[94]}
   );
   gpc1_1 gpc8003 (
      {stage2_10[159]},
      {stage3_10[95]}
   );
   gpc1_1 gpc8004 (
      {stage2_10[160]},
      {stage3_10[96]}
   );
   gpc1_1 gpc8005 (
      {stage2_10[161]},
      {stage3_10[97]}
   );
   gpc1_1 gpc8006 (
      {stage2_10[162]},
      {stage3_10[98]}
   );
   gpc1_1 gpc8007 (
      {stage2_10[163]},
      {stage3_10[99]}
   );
   gpc1_1 gpc8008 (
      {stage2_11[127]},
      {stage3_11[46]}
   );
   gpc1_1 gpc8009 (
      {stage2_11[128]},
      {stage3_11[47]}
   );
   gpc1_1 gpc8010 (
      {stage2_11[129]},
      {stage3_11[48]}
   );
   gpc1_1 gpc8011 (
      {stage2_11[130]},
      {stage3_11[49]}
   );
   gpc1_1 gpc8012 (
      {stage2_11[131]},
      {stage3_11[50]}
   );
   gpc1_1 gpc8013 (
      {stage2_11[132]},
      {stage3_11[51]}
   );
   gpc1_1 gpc8014 (
      {stage2_11[133]},
      {stage3_11[52]}
   );
   gpc1_1 gpc8015 (
      {stage2_11[134]},
      {stage3_11[53]}
   );
   gpc1_1 gpc8016 (
      {stage2_11[135]},
      {stage3_11[54]}
   );
   gpc1_1 gpc8017 (
      {stage2_11[136]},
      {stage3_11[55]}
   );
   gpc1_1 gpc8018 (
      {stage2_11[137]},
      {stage3_11[56]}
   );
   gpc1_1 gpc8019 (
      {stage2_11[138]},
      {stage3_11[57]}
   );
   gpc1_1 gpc8020 (
      {stage2_12[92]},
      {stage3_12[53]}
   );
   gpc1_1 gpc8021 (
      {stage2_12[93]},
      {stage3_12[54]}
   );
   gpc1_1 gpc8022 (
      {stage2_12[94]},
      {stage3_12[55]}
   );
   gpc1_1 gpc8023 (
      {stage2_12[95]},
      {stage3_12[56]}
   );
   gpc1_1 gpc8024 (
      {stage2_12[96]},
      {stage3_12[57]}
   );
   gpc1_1 gpc8025 (
      {stage2_12[97]},
      {stage3_12[58]}
   );
   gpc1_1 gpc8026 (
      {stage2_12[98]},
      {stage3_12[59]}
   );
   gpc1_1 gpc8027 (
      {stage2_12[99]},
      {stage3_12[60]}
   );
   gpc1_1 gpc8028 (
      {stage2_12[100]},
      {stage3_12[61]}
   );
   gpc1_1 gpc8029 (
      {stage2_12[101]},
      {stage3_12[62]}
   );
   gpc1_1 gpc8030 (
      {stage2_12[102]},
      {stage3_12[63]}
   );
   gpc1_1 gpc8031 (
      {stage2_12[103]},
      {stage3_12[64]}
   );
   gpc1_1 gpc8032 (
      {stage2_12[104]},
      {stage3_12[65]}
   );
   gpc1_1 gpc8033 (
      {stage2_12[105]},
      {stage3_12[66]}
   );
   gpc1_1 gpc8034 (
      {stage2_12[106]},
      {stage3_12[67]}
   );
   gpc1_1 gpc8035 (
      {stage2_13[66]},
      {stage3_13[45]}
   );
   gpc1_1 gpc8036 (
      {stage2_13[67]},
      {stage3_13[46]}
   );
   gpc1_1 gpc8037 (
      {stage2_13[68]},
      {stage3_13[47]}
   );
   gpc1_1 gpc8038 (
      {stage2_13[69]},
      {stage3_13[48]}
   );
   gpc1_1 gpc8039 (
      {stage2_13[70]},
      {stage3_13[49]}
   );
   gpc1_1 gpc8040 (
      {stage2_13[71]},
      {stage3_13[50]}
   );
   gpc1_1 gpc8041 (
      {stage2_13[72]},
      {stage3_13[51]}
   );
   gpc1_1 gpc8042 (
      {stage2_13[73]},
      {stage3_13[52]}
   );
   gpc1_1 gpc8043 (
      {stage2_13[74]},
      {stage3_13[53]}
   );
   gpc1_1 gpc8044 (
      {stage2_13[75]},
      {stage3_13[54]}
   );
   gpc1_1 gpc8045 (
      {stage2_13[76]},
      {stage3_13[55]}
   );
   gpc1_1 gpc8046 (
      {stage2_13[77]},
      {stage3_13[56]}
   );
   gpc1_1 gpc8047 (
      {stage2_15[138]},
      {stage3_15[45]}
   );
   gpc1_1 gpc8048 (
      {stage2_15[139]},
      {stage3_15[46]}
   );
   gpc1_1 gpc8049 (
      {stage2_15[140]},
      {stage3_15[47]}
   );
   gpc1_1 gpc8050 (
      {stage2_16[80]},
      {stage3_16[48]}
   );
   gpc1_1 gpc8051 (
      {stage2_16[81]},
      {stage3_16[49]}
   );
   gpc1_1 gpc8052 (
      {stage2_16[82]},
      {stage3_16[50]}
   );
   gpc1_1 gpc8053 (
      {stage2_18[100]},
      {stage3_18[41]}
   );
   gpc1_1 gpc8054 (
      {stage2_18[101]},
      {stage3_18[42]}
   );
   gpc1_1 gpc8055 (
      {stage2_18[102]},
      {stage3_18[43]}
   );
   gpc1_1 gpc8056 (
      {stage2_18[103]},
      {stage3_18[44]}
   );
   gpc1_1 gpc8057 (
      {stage2_18[104]},
      {stage3_18[45]}
   );
   gpc1_1 gpc8058 (
      {stage2_18[105]},
      {stage3_18[46]}
   );
   gpc1_1 gpc8059 (
      {stage2_18[106]},
      {stage3_18[47]}
   );
   gpc1_1 gpc8060 (
      {stage2_18[107]},
      {stage3_18[48]}
   );
   gpc1_1 gpc8061 (
      {stage2_18[108]},
      {stage3_18[49]}
   );
   gpc1_1 gpc8062 (
      {stage2_18[109]},
      {stage3_18[50]}
   );
   gpc1_1 gpc8063 (
      {stage2_18[110]},
      {stage3_18[51]}
   );
   gpc1_1 gpc8064 (
      {stage2_18[111]},
      {stage3_18[52]}
   );
   gpc1_1 gpc8065 (
      {stage2_18[112]},
      {stage3_18[53]}
   );
   gpc1_1 gpc8066 (
      {stage2_18[113]},
      {stage3_18[54]}
   );
   gpc1_1 gpc8067 (
      {stage2_18[114]},
      {stage3_18[55]}
   );
   gpc1_1 gpc8068 (
      {stage2_18[115]},
      {stage3_18[56]}
   );
   gpc1_1 gpc8069 (
      {stage2_18[116]},
      {stage3_18[57]}
   );
   gpc1_1 gpc8070 (
      {stage2_18[117]},
      {stage3_18[58]}
   );
   gpc1_1 gpc8071 (
      {stage2_18[118]},
      {stage3_18[59]}
   );
   gpc1_1 gpc8072 (
      {stage2_20[45]},
      {stage3_20[35]}
   );
   gpc1_1 gpc8073 (
      {stage2_20[46]},
      {stage3_20[36]}
   );
   gpc1_1 gpc8074 (
      {stage2_20[47]},
      {stage3_20[37]}
   );
   gpc1_1 gpc8075 (
      {stage2_20[48]},
      {stage3_20[38]}
   );
   gpc1_1 gpc8076 (
      {stage2_20[49]},
      {stage3_20[39]}
   );
   gpc1_1 gpc8077 (
      {stage2_20[50]},
      {stage3_20[40]}
   );
   gpc1_1 gpc8078 (
      {stage2_20[51]},
      {stage3_20[41]}
   );
   gpc1_1 gpc8079 (
      {stage2_20[52]},
      {stage3_20[42]}
   );
   gpc1_1 gpc8080 (
      {stage2_20[53]},
      {stage3_20[43]}
   );
   gpc1_1 gpc8081 (
      {stage2_20[54]},
      {stage3_20[44]}
   );
   gpc1_1 gpc8082 (
      {stage2_20[55]},
      {stage3_20[45]}
   );
   gpc1_1 gpc8083 (
      {stage2_20[56]},
      {stage3_20[46]}
   );
   gpc1_1 gpc8084 (
      {stage2_20[57]},
      {stage3_20[47]}
   );
   gpc1_1 gpc8085 (
      {stage2_20[58]},
      {stage3_20[48]}
   );
   gpc1_1 gpc8086 (
      {stage2_20[59]},
      {stage3_20[49]}
   );
   gpc1_1 gpc8087 (
      {stage2_20[60]},
      {stage3_20[50]}
   );
   gpc1_1 gpc8088 (
      {stage2_20[61]},
      {stage3_20[51]}
   );
   gpc1_1 gpc8089 (
      {stage2_20[62]},
      {stage3_20[52]}
   );
   gpc1_1 gpc8090 (
      {stage2_20[63]},
      {stage3_20[53]}
   );
   gpc1_1 gpc8091 (
      {stage2_20[64]},
      {stage3_20[54]}
   );
   gpc1_1 gpc8092 (
      {stage2_20[65]},
      {stage3_20[55]}
   );
   gpc1_1 gpc8093 (
      {stage2_20[66]},
      {stage3_20[56]}
   );
   gpc1_1 gpc8094 (
      {stage2_20[67]},
      {stage3_20[57]}
   );
   gpc1_1 gpc8095 (
      {stage2_20[68]},
      {stage3_20[58]}
   );
   gpc1_1 gpc8096 (
      {stage2_20[69]},
      {stage3_20[59]}
   );
   gpc1_1 gpc8097 (
      {stage2_20[70]},
      {stage3_20[60]}
   );
   gpc1_1 gpc8098 (
      {stage2_20[71]},
      {stage3_20[61]}
   );
   gpc1_1 gpc8099 (
      {stage2_20[72]},
      {stage3_20[62]}
   );
   gpc1_1 gpc8100 (
      {stage2_20[73]},
      {stage3_20[63]}
   );
   gpc1_1 gpc8101 (
      {stage2_20[74]},
      {stage3_20[64]}
   );
   gpc1_1 gpc8102 (
      {stage2_20[75]},
      {stage3_20[65]}
   );
   gpc1_1 gpc8103 (
      {stage2_20[76]},
      {stage3_20[66]}
   );
   gpc1_1 gpc8104 (
      {stage2_20[77]},
      {stage3_20[67]}
   );
   gpc1_1 gpc8105 (
      {stage2_20[78]},
      {stage3_20[68]}
   );
   gpc1_1 gpc8106 (
      {stage2_20[79]},
      {stage3_20[69]}
   );
   gpc1_1 gpc8107 (
      {stage2_20[80]},
      {stage3_20[70]}
   );
   gpc1_1 gpc8108 (
      {stage2_20[81]},
      {stage3_20[71]}
   );
   gpc1_1 gpc8109 (
      {stage2_20[82]},
      {stage3_20[72]}
   );
   gpc1_1 gpc8110 (
      {stage2_20[83]},
      {stage3_20[73]}
   );
   gpc1_1 gpc8111 (
      {stage2_20[84]},
      {stage3_20[74]}
   );
   gpc1_1 gpc8112 (
      {stage2_20[85]},
      {stage3_20[75]}
   );
   gpc1_1 gpc8113 (
      {stage2_20[86]},
      {stage3_20[76]}
   );
   gpc1_1 gpc8114 (
      {stage2_20[87]},
      {stage3_20[77]}
   );
   gpc1_1 gpc8115 (
      {stage2_20[88]},
      {stage3_20[78]}
   );
   gpc1_1 gpc8116 (
      {stage2_20[89]},
      {stage3_20[79]}
   );
   gpc1_1 gpc8117 (
      {stage2_20[90]},
      {stage3_20[80]}
   );
   gpc1_1 gpc8118 (
      {stage2_20[91]},
      {stage3_20[81]}
   );
   gpc1_1 gpc8119 (
      {stage2_20[92]},
      {stage3_20[82]}
   );
   gpc1_1 gpc8120 (
      {stage2_21[120]},
      {stage3_21[31]}
   );
   gpc1_1 gpc8121 (
      {stage2_21[121]},
      {stage3_21[32]}
   );
   gpc1_1 gpc8122 (
      {stage2_21[122]},
      {stage3_21[33]}
   );
   gpc1_1 gpc8123 (
      {stage2_21[123]},
      {stage3_21[34]}
   );
   gpc1_1 gpc8124 (
      {stage2_21[124]},
      {stage3_21[35]}
   );
   gpc1_1 gpc8125 (
      {stage2_21[125]},
      {stage3_21[36]}
   );
   gpc1_1 gpc8126 (
      {stage2_21[126]},
      {stage3_21[37]}
   );
   gpc1_1 gpc8127 (
      {stage2_21[127]},
      {stage3_21[38]}
   );
   gpc1_1 gpc8128 (
      {stage2_22[80]},
      {stage3_22[45]}
   );
   gpc1_1 gpc8129 (
      {stage2_22[81]},
      {stage3_22[46]}
   );
   gpc1_1 gpc8130 (
      {stage2_22[82]},
      {stage3_22[47]}
   );
   gpc1_1 gpc8131 (
      {stage2_22[83]},
      {stage3_22[48]}
   );
   gpc1_1 gpc8132 (
      {stage2_22[84]},
      {stage3_22[49]}
   );
   gpc1_1 gpc8133 (
      {stage2_22[85]},
      {stage3_22[50]}
   );
   gpc1_1 gpc8134 (
      {stage2_22[86]},
      {stage3_22[51]}
   );
   gpc1_1 gpc8135 (
      {stage2_22[87]},
      {stage3_22[52]}
   );
   gpc1_1 gpc8136 (
      {stage2_22[88]},
      {stage3_22[53]}
   );
   gpc1_1 gpc8137 (
      {stage2_22[89]},
      {stage3_22[54]}
   );
   gpc1_1 gpc8138 (
      {stage2_22[90]},
      {stage3_22[55]}
   );
   gpc1_1 gpc8139 (
      {stage2_22[91]},
      {stage3_22[56]}
   );
   gpc1_1 gpc8140 (
      {stage2_22[92]},
      {stage3_22[57]}
   );
   gpc1_1 gpc8141 (
      {stage2_22[93]},
      {stage3_22[58]}
   );
   gpc1_1 gpc8142 (
      {stage2_22[94]},
      {stage3_22[59]}
   );
   gpc1_1 gpc8143 (
      {stage2_22[95]},
      {stage3_22[60]}
   );
   gpc1_1 gpc8144 (
      {stage2_22[96]},
      {stage3_22[61]}
   );
   gpc1_1 gpc8145 (
      {stage2_22[97]},
      {stage3_22[62]}
   );
   gpc1_1 gpc8146 (
      {stage2_22[98]},
      {stage3_22[63]}
   );
   gpc1_1 gpc8147 (
      {stage2_22[99]},
      {stage3_22[64]}
   );
   gpc1_1 gpc8148 (
      {stage2_22[100]},
      {stage3_22[65]}
   );
   gpc1_1 gpc8149 (
      {stage2_22[101]},
      {stage3_22[66]}
   );
   gpc1_1 gpc8150 (
      {stage2_22[102]},
      {stage3_22[67]}
   );
   gpc1_1 gpc8151 (
      {stage2_22[103]},
      {stage3_22[68]}
   );
   gpc1_1 gpc8152 (
      {stage2_22[104]},
      {stage3_22[69]}
   );
   gpc1_1 gpc8153 (
      {stage2_22[105]},
      {stage3_22[70]}
   );
   gpc1_1 gpc8154 (
      {stage2_22[106]},
      {stage3_22[71]}
   );
   gpc1_1 gpc8155 (
      {stage2_22[107]},
      {stage3_22[72]}
   );
   gpc1_1 gpc8156 (
      {stage2_26[83]},
      {stage3_26[47]}
   );
   gpc1_1 gpc8157 (
      {stage2_26[84]},
      {stage3_26[48]}
   );
   gpc1_1 gpc8158 (
      {stage2_27[93]},
      {stage3_27[36]}
   );
   gpc1_1 gpc8159 (
      {stage2_27[94]},
      {stage3_27[37]}
   );
   gpc1_1 gpc8160 (
      {stage2_27[95]},
      {stage3_27[38]}
   );
   gpc1_1 gpc8161 (
      {stage2_27[96]},
      {stage3_27[39]}
   );
   gpc1_1 gpc8162 (
      {stage2_27[97]},
      {stage3_27[40]}
   );
   gpc1_1 gpc8163 (
      {stage2_27[98]},
      {stage3_27[41]}
   );
   gpc1_1 gpc8164 (
      {stage2_27[99]},
      {stage3_27[42]}
   );
   gpc1_1 gpc8165 (
      {stage2_27[100]},
      {stage3_27[43]}
   );
   gpc1_1 gpc8166 (
      {stage2_27[101]},
      {stage3_27[44]}
   );
   gpc1_1 gpc8167 (
      {stage2_27[102]},
      {stage3_27[45]}
   );
   gpc1_1 gpc8168 (
      {stage2_27[103]},
      {stage3_27[46]}
   );
   gpc1_1 gpc8169 (
      {stage2_27[104]},
      {stage3_27[47]}
   );
   gpc1_1 gpc8170 (
      {stage2_27[105]},
      {stage3_27[48]}
   );
   gpc1_1 gpc8171 (
      {stage2_28[69]},
      {stage3_28[34]}
   );
   gpc1_1 gpc8172 (
      {stage2_28[70]},
      {stage3_28[35]}
   );
   gpc1_1 gpc8173 (
      {stage2_28[71]},
      {stage3_28[36]}
   );
   gpc1_1 gpc8174 (
      {stage2_28[72]},
      {stage3_28[37]}
   );
   gpc1_1 gpc8175 (
      {stage2_28[73]},
      {stage3_28[38]}
   );
   gpc1_1 gpc8176 (
      {stage2_28[74]},
      {stage3_28[39]}
   );
   gpc1_1 gpc8177 (
      {stage2_28[75]},
      {stage3_28[40]}
   );
   gpc1_1 gpc8178 (
      {stage2_28[76]},
      {stage3_28[41]}
   );
   gpc1_1 gpc8179 (
      {stage2_28[77]},
      {stage3_28[42]}
   );
   gpc1_1 gpc8180 (
      {stage2_28[78]},
      {stage3_28[43]}
   );
   gpc1_1 gpc8181 (
      {stage2_28[79]},
      {stage3_28[44]}
   );
   gpc1_1 gpc8182 (
      {stage2_28[80]},
      {stage3_28[45]}
   );
   gpc1_1 gpc8183 (
      {stage2_28[81]},
      {stage3_28[46]}
   );
   gpc1_1 gpc8184 (
      {stage2_28[82]},
      {stage3_28[47]}
   );
   gpc1_1 gpc8185 (
      {stage2_28[83]},
      {stage3_28[48]}
   );
   gpc1_1 gpc8186 (
      {stage2_28[84]},
      {stage3_28[49]}
   );
   gpc1_1 gpc8187 (
      {stage2_28[85]},
      {stage3_28[50]}
   );
   gpc1_1 gpc8188 (
      {stage2_28[86]},
      {stage3_28[51]}
   );
   gpc1_1 gpc8189 (
      {stage2_28[87]},
      {stage3_28[52]}
   );
   gpc1_1 gpc8190 (
      {stage2_28[88]},
      {stage3_28[53]}
   );
   gpc1_1 gpc8191 (
      {stage2_28[89]},
      {stage3_28[54]}
   );
   gpc1_1 gpc8192 (
      {stage2_28[90]},
      {stage3_28[55]}
   );
   gpc1_1 gpc8193 (
      {stage2_28[91]},
      {stage3_28[56]}
   );
   gpc1_1 gpc8194 (
      {stage2_30[103]},
      {stage3_30[28]}
   );
   gpc1_1 gpc8195 (
      {stage2_30[104]},
      {stage3_30[29]}
   );
   gpc1_1 gpc8196 (
      {stage2_30[105]},
      {stage3_30[30]}
   );
   gpc1_1 gpc8197 (
      {stage2_30[106]},
      {stage3_30[31]}
   );
   gpc1_1 gpc8198 (
      {stage2_30[107]},
      {stage3_30[32]}
   );
   gpc1_1 gpc8199 (
      {stage2_30[108]},
      {stage3_30[33]}
   );
   gpc1_1 gpc8200 (
      {stage2_30[109]},
      {stage3_30[34]}
   );
   gpc1_1 gpc8201 (
      {stage2_30[110]},
      {stage3_30[35]}
   );
   gpc1_1 gpc8202 (
      {stage2_30[111]},
      {stage3_30[36]}
   );
   gpc1_1 gpc8203 (
      {stage2_30[112]},
      {stage3_30[37]}
   );
   gpc1_1 gpc8204 (
      {stage2_30[113]},
      {stage3_30[38]}
   );
   gpc1_1 gpc8205 (
      {stage2_30[114]},
      {stage3_30[39]}
   );
   gpc1_1 gpc8206 (
      {stage2_30[115]},
      {stage3_30[40]}
   );
   gpc1_1 gpc8207 (
      {stage2_30[116]},
      {stage3_30[41]}
   );
   gpc1_1 gpc8208 (
      {stage2_31[95]},
      {stage3_31[34]}
   );
   gpc1_1 gpc8209 (
      {stage2_31[96]},
      {stage3_31[35]}
   );
   gpc1_1 gpc8210 (
      {stage2_31[97]},
      {stage3_31[36]}
   );
   gpc1_1 gpc8211 (
      {stage2_31[98]},
      {stage3_31[37]}
   );
   gpc1_1 gpc8212 (
      {stage2_32[99]},
      {stage3_32[47]}
   );
   gpc1_1 gpc8213 (
      {stage2_32[100]},
      {stage3_32[48]}
   );
   gpc1_1 gpc8214 (
      {stage2_32[101]},
      {stage3_32[49]}
   );
   gpc1_1 gpc8215 (
      {stage2_32[102]},
      {stage3_32[50]}
   );
   gpc1_1 gpc8216 (
      {stage2_32[103]},
      {stage3_32[51]}
   );
   gpc1_1 gpc8217 (
      {stage2_32[104]},
      {stage3_32[52]}
   );
   gpc1_1 gpc8218 (
      {stage2_32[105]},
      {stage3_32[53]}
   );
   gpc1_1 gpc8219 (
      {stage2_33[72]},
      {stage3_33[42]}
   );
   gpc1_1 gpc8220 (
      {stage2_33[73]},
      {stage3_33[43]}
   );
   gpc1_1 gpc8221 (
      {stage2_33[74]},
      {stage3_33[44]}
   );
   gpc1_1 gpc8222 (
      {stage2_33[75]},
      {stage3_33[45]}
   );
   gpc1_1 gpc8223 (
      {stage2_34[129]},
      {stage3_34[39]}
   );
   gpc1_1 gpc8224 (
      {stage2_34[130]},
      {stage3_34[40]}
   );
   gpc1_1 gpc8225 (
      {stage2_34[131]},
      {stage3_34[41]}
   );
   gpc1_1 gpc8226 (
      {stage2_35[120]},
      {stage3_35[44]}
   );
   gpc1_1 gpc8227 (
      {stage2_35[121]},
      {stage3_35[45]}
   );
   gpc1_1 gpc8228 (
      {stage2_35[122]},
      {stage3_35[46]}
   );
   gpc1_1 gpc8229 (
      {stage2_35[123]},
      {stage3_35[47]}
   );
   gpc1_1 gpc8230 (
      {stage2_35[124]},
      {stage3_35[48]}
   );
   gpc1_1 gpc8231 (
      {stage2_35[125]},
      {stage3_35[49]}
   );
   gpc1_1 gpc8232 (
      {stage2_35[126]},
      {stage3_35[50]}
   );
   gpc1_1 gpc8233 (
      {stage2_35[127]},
      {stage3_35[51]}
   );
   gpc1_1 gpc8234 (
      {stage2_35[128]},
      {stage3_35[52]}
   );
   gpc1_1 gpc8235 (
      {stage2_35[129]},
      {stage3_35[53]}
   );
   gpc1_1 gpc8236 (
      {stage2_35[130]},
      {stage3_35[54]}
   );
   gpc1_1 gpc8237 (
      {stage2_35[131]},
      {stage3_35[55]}
   );
   gpc1_1 gpc8238 (
      {stage2_35[132]},
      {stage3_35[56]}
   );
   gpc1_1 gpc8239 (
      {stage2_36[73]},
      {stage3_36[44]}
   );
   gpc1_1 gpc8240 (
      {stage2_36[74]},
      {stage3_36[45]}
   );
   gpc1_1 gpc8241 (
      {stage2_37[74]},
      {stage3_37[37]}
   );
   gpc1_1 gpc8242 (
      {stage2_37[75]},
      {stage3_37[38]}
   );
   gpc1_1 gpc8243 (
      {stage2_37[76]},
      {stage3_37[39]}
   );
   gpc1_1 gpc8244 (
      {stage2_37[77]},
      {stage3_37[40]}
   );
   gpc1_1 gpc8245 (
      {stage2_37[78]},
      {stage3_37[41]}
   );
   gpc1_1 gpc8246 (
      {stage2_37[79]},
      {stage3_37[42]}
   );
   gpc1_1 gpc8247 (
      {stage2_37[80]},
      {stage3_37[43]}
   );
   gpc1_1 gpc8248 (
      {stage2_37[81]},
      {stage3_37[44]}
   );
   gpc1_1 gpc8249 (
      {stage2_37[82]},
      {stage3_37[45]}
   );
   gpc1_1 gpc8250 (
      {stage2_37[83]},
      {stage3_37[46]}
   );
   gpc1_1 gpc8251 (
      {stage2_37[84]},
      {stage3_37[47]}
   );
   gpc1_1 gpc8252 (
      {stage2_37[85]},
      {stage3_37[48]}
   );
   gpc1_1 gpc8253 (
      {stage2_37[86]},
      {stage3_37[49]}
   );
   gpc1_1 gpc8254 (
      {stage2_37[87]},
      {stage3_37[50]}
   );
   gpc1_1 gpc8255 (
      {stage2_37[88]},
      {stage3_37[51]}
   );
   gpc1_1 gpc8256 (
      {stage2_37[89]},
      {stage3_37[52]}
   );
   gpc1_1 gpc8257 (
      {stage2_38[125]},
      {stage3_38[45]}
   );
   gpc1_1 gpc8258 (
      {stage2_38[126]},
      {stage3_38[46]}
   );
   gpc1_1 gpc8259 (
      {stage2_38[127]},
      {stage3_38[47]}
   );
   gpc1_1 gpc8260 (
      {stage2_38[128]},
      {stage3_38[48]}
   );
   gpc1_1 gpc8261 (
      {stage2_38[129]},
      {stage3_38[49]}
   );
   gpc1_1 gpc8262 (
      {stage2_38[130]},
      {stage3_38[50]}
   );
   gpc1_1 gpc8263 (
      {stage2_38[131]},
      {stage3_38[51]}
   );
   gpc1_1 gpc8264 (
      {stage2_38[132]},
      {stage3_38[52]}
   );
   gpc1_1 gpc8265 (
      {stage2_38[133]},
      {stage3_38[53]}
   );
   gpc1_1 gpc8266 (
      {stage2_38[134]},
      {stage3_38[54]}
   );
   gpc1_1 gpc8267 (
      {stage2_38[135]},
      {stage3_38[55]}
   );
   gpc1_1 gpc8268 (
      {stage2_38[136]},
      {stage3_38[56]}
   );
   gpc1_1 gpc8269 (
      {stage2_38[137]},
      {stage3_38[57]}
   );
   gpc1_1 gpc8270 (
      {stage2_38[138]},
      {stage3_38[58]}
   );
   gpc1_1 gpc8271 (
      {stage2_38[139]},
      {stage3_38[59]}
   );
   gpc1_1 gpc8272 (
      {stage2_39[128]},
      {stage3_39[49]}
   );
   gpc1_1 gpc8273 (
      {stage2_39[129]},
      {stage3_39[50]}
   );
   gpc1_1 gpc8274 (
      {stage2_39[130]},
      {stage3_39[51]}
   );
   gpc1_1 gpc8275 (
      {stage2_39[131]},
      {stage3_39[52]}
   );
   gpc1_1 gpc8276 (
      {stage2_39[132]},
      {stage3_39[53]}
   );
   gpc1_1 gpc8277 (
      {stage2_39[133]},
      {stage3_39[54]}
   );
   gpc1_1 gpc8278 (
      {stage2_39[134]},
      {stage3_39[55]}
   );
   gpc1_1 gpc8279 (
      {stage2_39[135]},
      {stage3_39[56]}
   );
   gpc1_1 gpc8280 (
      {stage2_39[136]},
      {stage3_39[57]}
   );
   gpc1_1 gpc8281 (
      {stage2_40[107]},
      {stage3_40[46]}
   );
   gpc1_1 gpc8282 (
      {stage2_40[108]},
      {stage3_40[47]}
   );
   gpc1_1 gpc8283 (
      {stage2_40[109]},
      {stage3_40[48]}
   );
   gpc1_1 gpc8284 (
      {stage2_40[110]},
      {stage3_40[49]}
   );
   gpc1_1 gpc8285 (
      {stage2_40[111]},
      {stage3_40[50]}
   );
   gpc1_1 gpc8286 (
      {stage2_40[112]},
      {stage3_40[51]}
   );
   gpc1_1 gpc8287 (
      {stage2_41[102]},
      {stage3_41[39]}
   );
   gpc1_1 gpc8288 (
      {stage2_41[103]},
      {stage3_41[40]}
   );
   gpc1_1 gpc8289 (
      {stage2_41[104]},
      {stage3_41[41]}
   );
   gpc1_1 gpc8290 (
      {stage2_41[105]},
      {stage3_41[42]}
   );
   gpc1_1 gpc8291 (
      {stage2_42[82]},
      {stage3_42[46]}
   );
   gpc1_1 gpc8292 (
      {stage2_42[83]},
      {stage3_42[47]}
   );
   gpc1_1 gpc8293 (
      {stage2_42[84]},
      {stage3_42[48]}
   );
   gpc1_1 gpc8294 (
      {stage2_42[85]},
      {stage3_42[49]}
   );
   gpc1_1 gpc8295 (
      {stage2_44[109]},
      {stage3_44[31]}
   );
   gpc1_1 gpc8296 (
      {stage2_44[110]},
      {stage3_44[32]}
   );
   gpc1_1 gpc8297 (
      {stage2_44[111]},
      {stage3_44[33]}
   );
   gpc1_1 gpc8298 (
      {stage2_44[112]},
      {stage3_44[34]}
   );
   gpc1_1 gpc8299 (
      {stage2_44[113]},
      {stage3_44[35]}
   );
   gpc1_1 gpc8300 (
      {stage2_44[114]},
      {stage3_44[36]}
   );
   gpc1_1 gpc8301 (
      {stage2_44[115]},
      {stage3_44[37]}
   );
   gpc1_1 gpc8302 (
      {stage2_44[116]},
      {stage3_44[38]}
   );
   gpc1_1 gpc8303 (
      {stage2_44[117]},
      {stage3_44[39]}
   );
   gpc1_1 gpc8304 (
      {stage2_44[118]},
      {stage3_44[40]}
   );
   gpc1_1 gpc8305 (
      {stage2_45[108]},
      {stage3_45[34]}
   );
   gpc1_1 gpc8306 (
      {stage2_45[109]},
      {stage3_45[35]}
   );
   gpc1_1 gpc8307 (
      {stage2_45[110]},
      {stage3_45[36]}
   );
   gpc1_1 gpc8308 (
      {stage2_45[111]},
      {stage3_45[37]}
   );
   gpc1_1 gpc8309 (
      {stage2_45[112]},
      {stage3_45[38]}
   );
   gpc1_1 gpc8310 (
      {stage2_45[113]},
      {stage3_45[39]}
   );
   gpc1_1 gpc8311 (
      {stage2_45[114]},
      {stage3_45[40]}
   );
   gpc1_1 gpc8312 (
      {stage2_45[115]},
      {stage3_45[41]}
   );
   gpc1_1 gpc8313 (
      {stage2_45[116]},
      {stage3_45[42]}
   );
   gpc1_1 gpc8314 (
      {stage2_45[117]},
      {stage3_45[43]}
   );
   gpc1_1 gpc8315 (
      {stage2_46[78]},
      {stage3_46[48]}
   );
   gpc1_1 gpc8316 (
      {stage2_46[79]},
      {stage3_46[49]}
   );
   gpc1_1 gpc8317 (
      {stage2_46[80]},
      {stage3_46[50]}
   );
   gpc1_1 gpc8318 (
      {stage2_46[81]},
      {stage3_46[51]}
   );
   gpc1_1 gpc8319 (
      {stage2_46[82]},
      {stage3_46[52]}
   );
   gpc1_1 gpc8320 (
      {stage2_46[83]},
      {stage3_46[53]}
   );
   gpc1_1 gpc8321 (
      {stage2_46[84]},
      {stage3_46[54]}
   );
   gpc1_1 gpc8322 (
      {stage2_46[85]},
      {stage3_46[55]}
   );
   gpc1_1 gpc8323 (
      {stage2_46[86]},
      {stage3_46[56]}
   );
   gpc1_1 gpc8324 (
      {stage2_46[87]},
      {stage3_46[57]}
   );
   gpc1_1 gpc8325 (
      {stage2_48[126]},
      {stage3_48[38]}
   );
   gpc1_1 gpc8326 (
      {stage2_48[127]},
      {stage3_48[39]}
   );
   gpc1_1 gpc8327 (
      {stage2_48[128]},
      {stage3_48[40]}
   );
   gpc1_1 gpc8328 (
      {stage2_48[129]},
      {stage3_48[41]}
   );
   gpc1_1 gpc8329 (
      {stage2_50[84]},
      {stage3_50[45]}
   );
   gpc1_1 gpc8330 (
      {stage2_50[85]},
      {stage3_50[46]}
   );
   gpc1_1 gpc8331 (
      {stage2_51[59]},
      {stage3_51[34]}
   );
   gpc1_1 gpc8332 (
      {stage2_51[60]},
      {stage3_51[35]}
   );
   gpc1_1 gpc8333 (
      {stage2_51[61]},
      {stage3_51[36]}
   );
   gpc1_1 gpc8334 (
      {stage2_51[62]},
      {stage3_51[37]}
   );
   gpc1_1 gpc8335 (
      {stage2_51[63]},
      {stage3_51[38]}
   );
   gpc1_1 gpc8336 (
      {stage2_51[64]},
      {stage3_51[39]}
   );
   gpc1_1 gpc8337 (
      {stage2_51[65]},
      {stage3_51[40]}
   );
   gpc1_1 gpc8338 (
      {stage2_51[66]},
      {stage3_51[41]}
   );
   gpc1_1 gpc8339 (
      {stage2_51[67]},
      {stage3_51[42]}
   );
   gpc1_1 gpc8340 (
      {stage2_51[68]},
      {stage3_51[43]}
   );
   gpc1_1 gpc8341 (
      {stage2_51[69]},
      {stage3_51[44]}
   );
   gpc1_1 gpc8342 (
      {stage2_51[70]},
      {stage3_51[45]}
   );
   gpc1_1 gpc8343 (
      {stage2_51[71]},
      {stage3_51[46]}
   );
   gpc1_1 gpc8344 (
      {stage2_51[72]},
      {stage3_51[47]}
   );
   gpc1_1 gpc8345 (
      {stage2_51[73]},
      {stage3_51[48]}
   );
   gpc1_1 gpc8346 (
      {stage2_51[74]},
      {stage3_51[49]}
   );
   gpc1_1 gpc8347 (
      {stage2_51[75]},
      {stage3_51[50]}
   );
   gpc1_1 gpc8348 (
      {stage2_51[76]},
      {stage3_51[51]}
   );
   gpc1_1 gpc8349 (
      {stage2_51[77]},
      {stage3_51[52]}
   );
   gpc1_1 gpc8350 (
      {stage2_51[78]},
      {stage3_51[53]}
   );
   gpc1_1 gpc8351 (
      {stage2_51[79]},
      {stage3_51[54]}
   );
   gpc1_1 gpc8352 (
      {stage2_51[80]},
      {stage3_51[55]}
   );
   gpc1_1 gpc8353 (
      {stage2_51[81]},
      {stage3_51[56]}
   );
   gpc1_1 gpc8354 (
      {stage2_51[82]},
      {stage3_51[57]}
   );
   gpc1_1 gpc8355 (
      {stage2_51[83]},
      {stage3_51[58]}
   );
   gpc1_1 gpc8356 (
      {stage2_51[84]},
      {stage3_51[59]}
   );
   gpc1_1 gpc8357 (
      {stage2_51[85]},
      {stage3_51[60]}
   );
   gpc1_1 gpc8358 (
      {stage2_51[86]},
      {stage3_51[61]}
   );
   gpc1_1 gpc8359 (
      {stage2_51[87]},
      {stage3_51[62]}
   );
   gpc1_1 gpc8360 (
      {stage2_52[69]},
      {stage3_52[27]}
   );
   gpc1_1 gpc8361 (
      {stage2_52[70]},
      {stage3_52[28]}
   );
   gpc1_1 gpc8362 (
      {stage2_52[71]},
      {stage3_52[29]}
   );
   gpc1_1 gpc8363 (
      {stage2_52[72]},
      {stage3_52[30]}
   );
   gpc1_1 gpc8364 (
      {stage2_52[73]},
      {stage3_52[31]}
   );
   gpc1_1 gpc8365 (
      {stage2_52[74]},
      {stage3_52[32]}
   );
   gpc1_1 gpc8366 (
      {stage2_52[75]},
      {stage3_52[33]}
   );
   gpc1_1 gpc8367 (
      {stage2_52[76]},
      {stage3_52[34]}
   );
   gpc1_1 gpc8368 (
      {stage2_52[77]},
      {stage3_52[35]}
   );
   gpc1_1 gpc8369 (
      {stage2_52[78]},
      {stage3_52[36]}
   );
   gpc1_1 gpc8370 (
      {stage2_52[79]},
      {stage3_52[37]}
   );
   gpc1_1 gpc8371 (
      {stage2_52[80]},
      {stage3_52[38]}
   );
   gpc1_1 gpc8372 (
      {stage2_52[81]},
      {stage3_52[39]}
   );
   gpc1_1 gpc8373 (
      {stage2_52[82]},
      {stage3_52[40]}
   );
   gpc1_1 gpc8374 (
      {stage2_52[83]},
      {stage3_52[41]}
   );
   gpc1_1 gpc8375 (
      {stage2_52[84]},
      {stage3_52[42]}
   );
   gpc1_1 gpc8376 (
      {stage2_52[85]},
      {stage3_52[43]}
   );
   gpc1_1 gpc8377 (
      {stage2_52[86]},
      {stage3_52[44]}
   );
   gpc1_1 gpc8378 (
      {stage2_52[87]},
      {stage3_52[45]}
   );
   gpc1_1 gpc8379 (
      {stage2_52[88]},
      {stage3_52[46]}
   );
   gpc1_1 gpc8380 (
      {stage2_52[89]},
      {stage3_52[47]}
   );
   gpc1_1 gpc8381 (
      {stage2_52[90]},
      {stage3_52[48]}
   );
   gpc1_1 gpc8382 (
      {stage2_52[91]},
      {stage3_52[49]}
   );
   gpc1_1 gpc8383 (
      {stage2_52[92]},
      {stage3_52[50]}
   );
   gpc1_1 gpc8384 (
      {stage2_52[93]},
      {stage3_52[51]}
   );
   gpc1_1 gpc8385 (
      {stage2_52[94]},
      {stage3_52[52]}
   );
   gpc1_1 gpc8386 (
      {stage2_52[95]},
      {stage3_52[53]}
   );
   gpc1_1 gpc8387 (
      {stage2_52[96]},
      {stage3_52[54]}
   );
   gpc1_1 gpc8388 (
      {stage2_52[97]},
      {stage3_52[55]}
   );
   gpc1_1 gpc8389 (
      {stage2_52[98]},
      {stage3_52[56]}
   );
   gpc1_1 gpc8390 (
      {stage2_52[99]},
      {stage3_52[57]}
   );
   gpc1_1 gpc8391 (
      {stage2_52[100]},
      {stage3_52[58]}
   );
   gpc1_1 gpc8392 (
      {stage2_52[101]},
      {stage3_52[59]}
   );
   gpc1_1 gpc8393 (
      {stage2_52[102]},
      {stage3_52[60]}
   );
   gpc1_1 gpc8394 (
      {stage2_52[103]},
      {stage3_52[61]}
   );
   gpc1_1 gpc8395 (
      {stage2_52[104]},
      {stage3_52[62]}
   );
   gpc1_1 gpc8396 (
      {stage2_53[69]},
      {stage3_53[29]}
   );
   gpc1_1 gpc8397 (
      {stage2_53[70]},
      {stage3_53[30]}
   );
   gpc1_1 gpc8398 (
      {stage2_53[71]},
      {stage3_53[31]}
   );
   gpc1_1 gpc8399 (
      {stage2_53[72]},
      {stage3_53[32]}
   );
   gpc1_1 gpc8400 (
      {stage2_53[73]},
      {stage3_53[33]}
   );
   gpc1_1 gpc8401 (
      {stage2_53[74]},
      {stage3_53[34]}
   );
   gpc1_1 gpc8402 (
      {stage2_53[75]},
      {stage3_53[35]}
   );
   gpc1_1 gpc8403 (
      {stage2_53[76]},
      {stage3_53[36]}
   );
   gpc1_1 gpc8404 (
      {stage2_53[77]},
      {stage3_53[37]}
   );
   gpc1_1 gpc8405 (
      {stage2_53[78]},
      {stage3_53[38]}
   );
   gpc1_1 gpc8406 (
      {stage2_53[79]},
      {stage3_53[39]}
   );
   gpc1_1 gpc8407 (
      {stage2_53[80]},
      {stage3_53[40]}
   );
   gpc1_1 gpc8408 (
      {stage2_53[81]},
      {stage3_53[41]}
   );
   gpc1_1 gpc8409 (
      {stage2_53[82]},
      {stage3_53[42]}
   );
   gpc1_1 gpc8410 (
      {stage2_53[83]},
      {stage3_53[43]}
   );
   gpc1_1 gpc8411 (
      {stage2_53[84]},
      {stage3_53[44]}
   );
   gpc1_1 gpc8412 (
      {stage2_53[85]},
      {stage3_53[45]}
   );
   gpc1_1 gpc8413 (
      {stage2_53[86]},
      {stage3_53[46]}
   );
   gpc1_1 gpc8414 (
      {stage2_53[87]},
      {stage3_53[47]}
   );
   gpc1_1 gpc8415 (
      {stage2_53[88]},
      {stage3_53[48]}
   );
   gpc1_1 gpc8416 (
      {stage2_53[89]},
      {stage3_53[49]}
   );
   gpc1_1 gpc8417 (
      {stage2_53[90]},
      {stage3_53[50]}
   );
   gpc1_1 gpc8418 (
      {stage2_53[91]},
      {stage3_53[51]}
   );
   gpc1_1 gpc8419 (
      {stage2_53[92]},
      {stage3_53[52]}
   );
   gpc1_1 gpc8420 (
      {stage2_53[93]},
      {stage3_53[53]}
   );
   gpc1_1 gpc8421 (
      {stage2_53[94]},
      {stage3_53[54]}
   );
   gpc1_1 gpc8422 (
      {stage2_53[95]},
      {stage3_53[55]}
   );
   gpc1_1 gpc8423 (
      {stage2_53[96]},
      {stage3_53[56]}
   );
   gpc1_1 gpc8424 (
      {stage2_53[97]},
      {stage3_53[57]}
   );
   gpc1_1 gpc8425 (
      {stage2_53[98]},
      {stage3_53[58]}
   );
   gpc1_1 gpc8426 (
      {stage2_53[99]},
      {stage3_53[59]}
   );
   gpc1_1 gpc8427 (
      {stage2_53[100]},
      {stage3_53[60]}
   );
   gpc1_1 gpc8428 (
      {stage2_53[101]},
      {stage3_53[61]}
   );
   gpc1_1 gpc8429 (
      {stage2_53[102]},
      {stage3_53[62]}
   );
   gpc1_1 gpc8430 (
      {stage2_53[103]},
      {stage3_53[63]}
   );
   gpc1_1 gpc8431 (
      {stage2_53[104]},
      {stage3_53[64]}
   );
   gpc1_1 gpc8432 (
      {stage2_53[105]},
      {stage3_53[65]}
   );
   gpc1_1 gpc8433 (
      {stage2_53[106]},
      {stage3_53[66]}
   );
   gpc1_1 gpc8434 (
      {stage2_53[107]},
      {stage3_53[67]}
   );
   gpc1_1 gpc8435 (
      {stage2_53[108]},
      {stage3_53[68]}
   );
   gpc1_1 gpc8436 (
      {stage2_53[109]},
      {stage3_53[69]}
   );
   gpc1_1 gpc8437 (
      {stage2_53[110]},
      {stage3_53[70]}
   );
   gpc1_1 gpc8438 (
      {stage2_53[111]},
      {stage3_53[71]}
   );
   gpc1_1 gpc8439 (
      {stage2_53[112]},
      {stage3_53[72]}
   );
   gpc1_1 gpc8440 (
      {stage2_53[113]},
      {stage3_53[73]}
   );
   gpc1_1 gpc8441 (
      {stage2_53[114]},
      {stage3_53[74]}
   );
   gpc1_1 gpc8442 (
      {stage2_55[70]},
      {stage3_55[31]}
   );
   gpc1_1 gpc8443 (
      {stage2_55[71]},
      {stage3_55[32]}
   );
   gpc1_1 gpc8444 (
      {stage2_55[72]},
      {stage3_55[33]}
   );
   gpc1_1 gpc8445 (
      {stage2_55[73]},
      {stage3_55[34]}
   );
   gpc1_1 gpc8446 (
      {stage2_55[74]},
      {stage3_55[35]}
   );
   gpc1_1 gpc8447 (
      {stage2_55[75]},
      {stage3_55[36]}
   );
   gpc1_1 gpc8448 (
      {stage2_55[76]},
      {stage3_55[37]}
   );
   gpc1_1 gpc8449 (
      {stage2_55[77]},
      {stage3_55[38]}
   );
   gpc1_1 gpc8450 (
      {stage2_55[78]},
      {stage3_55[39]}
   );
   gpc1_1 gpc8451 (
      {stage2_55[79]},
      {stage3_55[40]}
   );
   gpc1_1 gpc8452 (
      {stage2_55[80]},
      {stage3_55[41]}
   );
   gpc1_1 gpc8453 (
      {stage2_55[81]},
      {stage3_55[42]}
   );
   gpc1_1 gpc8454 (
      {stage2_55[82]},
      {stage3_55[43]}
   );
   gpc1_1 gpc8455 (
      {stage2_55[83]},
      {stage3_55[44]}
   );
   gpc1_1 gpc8456 (
      {stage2_55[84]},
      {stage3_55[45]}
   );
   gpc1_1 gpc8457 (
      {stage2_55[85]},
      {stage3_55[46]}
   );
   gpc1_1 gpc8458 (
      {stage2_55[86]},
      {stage3_55[47]}
   );
   gpc1_1 gpc8459 (
      {stage2_55[87]},
      {stage3_55[48]}
   );
   gpc1_1 gpc8460 (
      {stage2_55[88]},
      {stage3_55[49]}
   );
   gpc1_1 gpc8461 (
      {stage2_55[89]},
      {stage3_55[50]}
   );
   gpc1_1 gpc8462 (
      {stage2_55[90]},
      {stage3_55[51]}
   );
   gpc1_1 gpc8463 (
      {stage2_55[91]},
      {stage3_55[52]}
   );
   gpc1_1 gpc8464 (
      {stage2_55[92]},
      {stage3_55[53]}
   );
   gpc1_1 gpc8465 (
      {stage2_55[93]},
      {stage3_55[54]}
   );
   gpc1_1 gpc8466 (
      {stage2_55[94]},
      {stage3_55[55]}
   );
   gpc1_1 gpc8467 (
      {stage2_55[95]},
      {stage3_55[56]}
   );
   gpc1_1 gpc8468 (
      {stage2_55[96]},
      {stage3_55[57]}
   );
   gpc1_1 gpc8469 (
      {stage2_55[97]},
      {stage3_55[58]}
   );
   gpc1_1 gpc8470 (
      {stage2_55[98]},
      {stage3_55[59]}
   );
   gpc1_1 gpc8471 (
      {stage2_55[99]},
      {stage3_55[60]}
   );
   gpc1_1 gpc8472 (
      {stage2_55[100]},
      {stage3_55[61]}
   );
   gpc1_1 gpc8473 (
      {stage2_55[101]},
      {stage3_55[62]}
   );
   gpc1_1 gpc8474 (
      {stage2_55[102]},
      {stage3_55[63]}
   );
   gpc1_1 gpc8475 (
      {stage2_55[103]},
      {stage3_55[64]}
   );
   gpc1_1 gpc8476 (
      {stage2_55[104]},
      {stage3_55[65]}
   );
   gpc1_1 gpc8477 (
      {stage2_55[105]},
      {stage3_55[66]}
   );
   gpc1_1 gpc8478 (
      {stage2_57[49]},
      {stage3_57[37]}
   );
   gpc1_1 gpc8479 (
      {stage2_57[50]},
      {stage3_57[38]}
   );
   gpc1_1 gpc8480 (
      {stage2_57[51]},
      {stage3_57[39]}
   );
   gpc1_1 gpc8481 (
      {stage2_57[52]},
      {stage3_57[40]}
   );
   gpc1_1 gpc8482 (
      {stage2_57[53]},
      {stage3_57[41]}
   );
   gpc1_1 gpc8483 (
      {stage2_57[54]},
      {stage3_57[42]}
   );
   gpc1_1 gpc8484 (
      {stage2_57[55]},
      {stage3_57[43]}
   );
   gpc1_1 gpc8485 (
      {stage2_57[56]},
      {stage3_57[44]}
   );
   gpc1_1 gpc8486 (
      {stage2_57[57]},
      {stage3_57[45]}
   );
   gpc1_1 gpc8487 (
      {stage2_57[58]},
      {stage3_57[46]}
   );
   gpc1_1 gpc8488 (
      {stage2_57[59]},
      {stage3_57[47]}
   );
   gpc1_1 gpc8489 (
      {stage2_57[60]},
      {stage3_57[48]}
   );
   gpc1_1 gpc8490 (
      {stage2_57[61]},
      {stage3_57[49]}
   );
   gpc1_1 gpc8491 (
      {stage2_57[62]},
      {stage3_57[50]}
   );
   gpc1_1 gpc8492 (
      {stage2_57[63]},
      {stage3_57[51]}
   );
   gpc1_1 gpc8493 (
      {stage2_57[64]},
      {stage3_57[52]}
   );
   gpc1_1 gpc8494 (
      {stage2_57[65]},
      {stage3_57[53]}
   );
   gpc1_1 gpc8495 (
      {stage2_58[58]},
      {stage3_58[34]}
   );
   gpc1_1 gpc8496 (
      {stage2_58[59]},
      {stage3_58[35]}
   );
   gpc1_1 gpc8497 (
      {stage2_58[60]},
      {stage3_58[36]}
   );
   gpc1_1 gpc8498 (
      {stage2_58[61]},
      {stage3_58[37]}
   );
   gpc1_1 gpc8499 (
      {stage2_58[62]},
      {stage3_58[38]}
   );
   gpc1_1 gpc8500 (
      {stage2_58[63]},
      {stage3_58[39]}
   );
   gpc1_1 gpc8501 (
      {stage2_58[64]},
      {stage3_58[40]}
   );
   gpc1_1 gpc8502 (
      {stage2_58[65]},
      {stage3_58[41]}
   );
   gpc1_1 gpc8503 (
      {stage2_58[66]},
      {stage3_58[42]}
   );
   gpc1_1 gpc8504 (
      {stage2_58[67]},
      {stage3_58[43]}
   );
   gpc1_1 gpc8505 (
      {stage2_58[68]},
      {stage3_58[44]}
   );
   gpc1_1 gpc8506 (
      {stage2_58[69]},
      {stage3_58[45]}
   );
   gpc1_1 gpc8507 (
      {stage2_58[70]},
      {stage3_58[46]}
   );
   gpc1_1 gpc8508 (
      {stage2_58[71]},
      {stage3_58[47]}
   );
   gpc1_1 gpc8509 (
      {stage2_58[72]},
      {stage3_58[48]}
   );
   gpc1_1 gpc8510 (
      {stage2_58[73]},
      {stage3_58[49]}
   );
   gpc1_1 gpc8511 (
      {stage2_58[74]},
      {stage3_58[50]}
   );
   gpc1_1 gpc8512 (
      {stage2_58[75]},
      {stage3_58[51]}
   );
   gpc1_1 gpc8513 (
      {stage2_58[76]},
      {stage3_58[52]}
   );
   gpc1_1 gpc8514 (
      {stage2_58[77]},
      {stage3_58[53]}
   );
   gpc1_1 gpc8515 (
      {stage2_58[78]},
      {stage3_58[54]}
   );
   gpc1_1 gpc8516 (
      {stage2_58[79]},
      {stage3_58[55]}
   );
   gpc1_1 gpc8517 (
      {stage2_58[80]},
      {stage3_58[56]}
   );
   gpc1_1 gpc8518 (
      {stage2_58[81]},
      {stage3_58[57]}
   );
   gpc1_1 gpc8519 (
      {stage2_58[82]},
      {stage3_58[58]}
   );
   gpc1_1 gpc8520 (
      {stage2_58[83]},
      {stage3_58[59]}
   );
   gpc1_1 gpc8521 (
      {stage2_58[84]},
      {stage3_58[60]}
   );
   gpc1_1 gpc8522 (
      {stage2_58[85]},
      {stage3_58[61]}
   );
   gpc1_1 gpc8523 (
      {stage2_59[85]},
      {stage3_59[25]}
   );
   gpc1_1 gpc8524 (
      {stage2_59[86]},
      {stage3_59[26]}
   );
   gpc1_1 gpc8525 (
      {stage2_59[87]},
      {stage3_59[27]}
   );
   gpc1_1 gpc8526 (
      {stage2_59[88]},
      {stage3_59[28]}
   );
   gpc1_1 gpc8527 (
      {stage2_59[89]},
      {stage3_59[29]}
   );
   gpc1_1 gpc8528 (
      {stage2_59[90]},
      {stage3_59[30]}
   );
   gpc1_1 gpc8529 (
      {stage2_59[91]},
      {stage3_59[31]}
   );
   gpc1_1 gpc8530 (
      {stage2_59[92]},
      {stage3_59[32]}
   );
   gpc1_1 gpc8531 (
      {stage2_59[93]},
      {stage3_59[33]}
   );
   gpc1_1 gpc8532 (
      {stage2_59[94]},
      {stage3_59[34]}
   );
   gpc1_1 gpc8533 (
      {stage2_59[95]},
      {stage3_59[35]}
   );
   gpc1_1 gpc8534 (
      {stage2_59[96]},
      {stage3_59[36]}
   );
   gpc1_1 gpc8535 (
      {stage2_59[97]},
      {stage3_59[37]}
   );
   gpc1_1 gpc8536 (
      {stage2_59[98]},
      {stage3_59[38]}
   );
   gpc1_1 gpc8537 (
      {stage2_59[99]},
      {stage3_59[39]}
   );
   gpc1_1 gpc8538 (
      {stage2_59[100]},
      {stage3_59[40]}
   );
   gpc1_1 gpc8539 (
      {stage2_59[101]},
      {stage3_59[41]}
   );
   gpc1_1 gpc8540 (
      {stage2_59[102]},
      {stage3_59[42]}
   );
   gpc1_1 gpc8541 (
      {stage2_59[103]},
      {stage3_59[43]}
   );
   gpc1_1 gpc8542 (
      {stage2_59[104]},
      {stage3_59[44]}
   );
   gpc1_1 gpc8543 (
      {stage2_59[105]},
      {stage3_59[45]}
   );
   gpc1_1 gpc8544 (
      {stage2_59[106]},
      {stage3_59[46]}
   );
   gpc1_1 gpc8545 (
      {stage2_59[107]},
      {stage3_59[47]}
   );
   gpc1_1 gpc8546 (
      {stage2_59[108]},
      {stage3_59[48]}
   );
   gpc1_1 gpc8547 (
      {stage2_59[109]},
      {stage3_59[49]}
   );
   gpc1_1 gpc8548 (
      {stage2_60[73]},
      {stage3_60[30]}
   );
   gpc1_1 gpc8549 (
      {stage2_60[74]},
      {stage3_60[31]}
   );
   gpc1_1 gpc8550 (
      {stage2_60[75]},
      {stage3_60[32]}
   );
   gpc1_1 gpc8551 (
      {stage2_60[76]},
      {stage3_60[33]}
   );
   gpc1_1 gpc8552 (
      {stage2_60[77]},
      {stage3_60[34]}
   );
   gpc1_1 gpc8553 (
      {stage2_60[78]},
      {stage3_60[35]}
   );
   gpc1_1 gpc8554 (
      {stage2_60[79]},
      {stage3_60[36]}
   );
   gpc1_1 gpc8555 (
      {stage2_60[80]},
      {stage3_60[37]}
   );
   gpc1_1 gpc8556 (
      {stage2_60[81]},
      {stage3_60[38]}
   );
   gpc1_1 gpc8557 (
      {stage2_60[82]},
      {stage3_60[39]}
   );
   gpc1_1 gpc8558 (
      {stage2_60[83]},
      {stage3_60[40]}
   );
   gpc1_1 gpc8559 (
      {stage2_60[84]},
      {stage3_60[41]}
   );
   gpc1_1 gpc8560 (
      {stage2_61[48]},
      {stage3_61[26]}
   );
   gpc1_1 gpc8561 (
      {stage2_61[49]},
      {stage3_61[27]}
   );
   gpc1_1 gpc8562 (
      {stage2_61[50]},
      {stage3_61[28]}
   );
   gpc1_1 gpc8563 (
      {stage2_61[51]},
      {stage3_61[29]}
   );
   gpc1_1 gpc8564 (
      {stage2_61[52]},
      {stage3_61[30]}
   );
   gpc1_1 gpc8565 (
      {stage2_61[53]},
      {stage3_61[31]}
   );
   gpc1_1 gpc8566 (
      {stage2_61[54]},
      {stage3_61[32]}
   );
   gpc1_1 gpc8567 (
      {stage2_61[55]},
      {stage3_61[33]}
   );
   gpc1_1 gpc8568 (
      {stage2_61[56]},
      {stage3_61[34]}
   );
   gpc1_1 gpc8569 (
      {stage2_61[57]},
      {stage3_61[35]}
   );
   gpc1_1 gpc8570 (
      {stage2_61[58]},
      {stage3_61[36]}
   );
   gpc1_1 gpc8571 (
      {stage2_61[59]},
      {stage3_61[37]}
   );
   gpc1_1 gpc8572 (
      {stage2_61[60]},
      {stage3_61[38]}
   );
   gpc1_1 gpc8573 (
      {stage2_61[61]},
      {stage3_61[39]}
   );
   gpc1_1 gpc8574 (
      {stage2_61[62]},
      {stage3_61[40]}
   );
   gpc1_1 gpc8575 (
      {stage2_61[63]},
      {stage3_61[41]}
   );
   gpc1_1 gpc8576 (
      {stage2_61[64]},
      {stage3_61[42]}
   );
   gpc1_1 gpc8577 (
      {stage2_61[65]},
      {stage3_61[43]}
   );
   gpc1_1 gpc8578 (
      {stage2_61[66]},
      {stage3_61[44]}
   );
   gpc1_1 gpc8579 (
      {stage2_61[67]},
      {stage3_61[45]}
   );
   gpc1_1 gpc8580 (
      {stage2_61[68]},
      {stage3_61[46]}
   );
   gpc1_1 gpc8581 (
      {stage2_61[69]},
      {stage3_61[47]}
   );
   gpc1_1 gpc8582 (
      {stage2_61[70]},
      {stage3_61[48]}
   );
   gpc1_1 gpc8583 (
      {stage2_61[71]},
      {stage3_61[49]}
   );
   gpc1_1 gpc8584 (
      {stage2_61[72]},
      {stage3_61[50]}
   );
   gpc1_1 gpc8585 (
      {stage2_61[73]},
      {stage3_61[51]}
   );
   gpc1_1 gpc8586 (
      {stage2_61[74]},
      {stage3_61[52]}
   );
   gpc1_1 gpc8587 (
      {stage2_63[90]},
      {stage3_63[39]}
   );
   gpc1_1 gpc8588 (
      {stage2_63[91]},
      {stage3_63[40]}
   );
   gpc1_1 gpc8589 (
      {stage2_63[92]},
      {stage3_63[41]}
   );
   gpc1_1 gpc8590 (
      {stage2_63[93]},
      {stage3_63[42]}
   );
   gpc1_1 gpc8591 (
      {stage2_63[94]},
      {stage3_63[43]}
   );
   gpc1_1 gpc8592 (
      {stage2_63[95]},
      {stage3_63[44]}
   );
   gpc1_1 gpc8593 (
      {stage2_63[96]},
      {stage3_63[45]}
   );
   gpc1_1 gpc8594 (
      {stage2_63[97]},
      {stage3_63[46]}
   );
   gpc1_1 gpc8595 (
      {stage2_63[98]},
      {stage3_63[47]}
   );
   gpc1_1 gpc8596 (
      {stage2_64[129]},
      {stage3_64[38]}
   );
   gpc1_1 gpc8597 (
      {stage2_64[130]},
      {stage3_64[39]}
   );
   gpc1_1 gpc8598 (
      {stage2_64[131]},
      {stage3_64[40]}
   );
   gpc1_1 gpc8599 (
      {stage2_64[132]},
      {stage3_64[41]}
   );
   gpc1_1 gpc8600 (
      {stage2_64[133]},
      {stage3_64[42]}
   );
   gpc1_1 gpc8601 (
      {stage2_64[134]},
      {stage3_64[43]}
   );
   gpc1_1 gpc8602 (
      {stage2_64[135]},
      {stage3_64[44]}
   );
   gpc1_1 gpc8603 (
      {stage2_64[136]},
      {stage3_64[45]}
   );
   gpc1_1 gpc8604 (
      {stage2_64[137]},
      {stage3_64[46]}
   );
   gpc1_1 gpc8605 (
      {stage2_64[138]},
      {stage3_64[47]}
   );
   gpc1_1 gpc8606 (
      {stage2_64[139]},
      {stage3_64[48]}
   );
   gpc1_1 gpc8607 (
      {stage2_64[140]},
      {stage3_64[49]}
   );
   gpc1_1 gpc8608 (
      {stage2_64[141]},
      {stage3_64[50]}
   );
   gpc1_1 gpc8609 (
      {stage2_65[51]},
      {stage3_65[33]}
   );
   gpc1_1 gpc8610 (
      {stage2_65[52]},
      {stage3_65[34]}
   );
   gpc1_1 gpc8611 (
      {stage2_65[53]},
      {stage3_65[35]}
   );
   gpc1_1 gpc8612 (
      {stage2_65[54]},
      {stage3_65[36]}
   );
   gpc1_1 gpc8613 (
      {stage2_65[55]},
      {stage3_65[37]}
   );
   gpc1_1 gpc8614 (
      {stage2_66[36]},
      {stage3_66[32]}
   );
   gpc1_1 gpc8615 (
      {stage2_66[37]},
      {stage3_66[33]}
   );
   gpc1_1 gpc8616 (
      {stage2_66[38]},
      {stage3_66[34]}
   );
   gpc1_1 gpc8617 (
      {stage2_66[39]},
      {stage3_66[35]}
   );
   gpc1_1 gpc8618 (
      {stage2_66[40]},
      {stage3_66[36]}
   );
   gpc1_1 gpc8619 (
      {stage2_66[41]},
      {stage3_66[37]}
   );
   gpc615_5 gpc8620 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4]},
      {stage3_1[0]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc8621 (
      {stage3_0[5], stage3_0[6], stage3_0[7], stage3_0[8], stage3_0[9]},
      {stage3_1[1]},
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1],stage4_0[1]}
   );
   gpc615_5 gpc8622 (
      {stage3_0[10], stage3_0[11], stage3_0[12], stage3_0[13], stage3_0[14]},
      {stage3_1[2]},
      {stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15], stage3_2[16], stage3_2[17]},
      {stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2],stage4_0[2]}
   );
   gpc606_5 gpc8623 (
      {stage3_1[3], stage3_1[4], stage3_1[5], stage3_1[6], stage3_1[7], stage3_1[8]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[3],stage4_3[3],stage4_2[3],stage4_1[3]}
   );
   gpc606_5 gpc8624 (
      {stage3_1[9], stage3_1[10], stage3_1[11], stage3_1[12], stage3_1[13], stage3_1[14]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[4],stage4_3[4],stage4_2[4],stage4_1[4]}
   );
   gpc606_5 gpc8625 (
      {stage3_1[15], stage3_1[16], stage3_1[17], stage3_1[18], stage3_1[19], stage3_1[20]},
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17]},
      {stage4_5[2],stage4_4[5],stage4_3[5],stage4_2[5],stage4_1[5]}
   );
   gpc606_5 gpc8626 (
      {stage3_2[18], stage3_2[19], stage3_2[20], stage3_2[21], stage3_2[22], stage3_2[23]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[3],stage4_4[6],stage4_3[6],stage4_2[6]}
   );
   gpc606_5 gpc8627 (
      {stage3_2[24], stage3_2[25], stage3_2[26], stage3_2[27], stage3_2[28], stage3_2[29]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[4],stage4_4[7],stage4_3[7],stage4_2[7]}
   );
   gpc606_5 gpc8628 (
      {stage3_2[30], stage3_2[31], stage3_2[32], stage3_2[33], stage3_2[34], stage3_2[35]},
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage4_6[2],stage4_5[5],stage4_4[8],stage4_3[8],stage4_2[8]}
   );
   gpc606_5 gpc8629 (
      {stage3_2[36], stage3_2[37], stage3_2[38], stage3_2[39], stage3_2[40], stage3_2[41]},
      {stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23]},
      {stage4_6[3],stage4_5[6],stage4_4[9],stage4_3[9],stage4_2[9]}
   );
   gpc615_5 gpc8630 (
      {stage3_3[18], stage3_3[19], stage3_3[20], stage3_3[21], stage3_3[22]},
      {stage3_4[24]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[4],stage4_5[7],stage4_4[10],stage4_3[10]}
   );
   gpc1163_5 gpc8631 (
      {stage3_4[25], stage3_4[26], stage3_4[27]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_6[0]},
      {stage3_7[0]},
      {stage4_8[0],stage4_7[1],stage4_6[5],stage4_5[8],stage4_4[11]}
   );
   gpc1163_5 gpc8632 (
      {stage3_4[28], stage3_4[29], stage3_4[30]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_6[1]},
      {stage3_7[1]},
      {stage4_8[1],stage4_7[2],stage4_6[6],stage4_5[9],stage4_4[12]}
   );
   gpc1163_5 gpc8633 (
      {stage3_4[31], stage3_4[32], stage3_4[33]},
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_6[2]},
      {stage3_7[2]},
      {stage4_8[2],stage4_7[3],stage4_6[7],stage4_5[10],stage4_4[13]}
   );
   gpc1163_5 gpc8634 (
      {stage3_4[34], stage3_4[35], stage3_4[36]},
      {stage3_5[24], stage3_5[25], stage3_5[26], stage3_5[27], stage3_5[28], stage3_5[29]},
      {stage3_6[3]},
      {stage3_7[3]},
      {stage4_8[3],stage4_7[4],stage4_6[8],stage4_5[11],stage4_4[14]}
   );
   gpc1163_5 gpc8635 (
      {stage3_4[37], stage3_4[38], stage3_4[39]},
      {stage3_5[30], stage3_5[31], stage3_5[32], stage3_5[33], stage3_5[34], stage3_5[35]},
      {stage3_6[4]},
      {stage3_7[4]},
      {stage4_8[4],stage4_7[5],stage4_6[9],stage4_5[12],stage4_4[15]}
   );
   gpc1163_5 gpc8636 (
      {stage3_4[40], stage3_4[41], stage3_4[42]},
      {stage3_5[36], stage3_5[37], stage3_5[38], stage3_5[39], stage3_5[40], stage3_5[41]},
      {stage3_6[5]},
      {stage3_7[5]},
      {stage4_8[5],stage4_7[6],stage4_6[10],stage4_5[13],stage4_4[16]}
   );
   gpc606_5 gpc8637 (
      {stage3_4[43], stage3_4[44], stage3_4[45], stage3_4[46], stage3_4[47], stage3_4[48]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[6],stage4_7[7],stage4_6[11],stage4_5[14],stage4_4[17]}
   );
   gpc606_5 gpc8638 (
      {stage3_4[49], stage3_4[50], stage3_4[51], stage3_4[52], stage3_4[53], stage3_4[54]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[7],stage4_7[8],stage4_6[12],stage4_5[15],stage4_4[18]}
   );
   gpc606_5 gpc8639 (
      {stage3_4[55], stage3_4[56], stage3_4[57], stage3_4[58], stage3_4[59], stage3_4[60]},
      {stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage4_8[8],stage4_7[9],stage4_6[13],stage4_5[16],stage4_4[19]}
   );
   gpc606_5 gpc8640 (
      {stage3_4[61], stage3_4[62], stage3_4[63], stage3_4[64], stage3_4[65], stage3_4[66]},
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29]},
      {stage4_8[9],stage4_7[10],stage4_6[14],stage4_5[17],stage4_4[20]}
   );
   gpc606_5 gpc8641 (
      {stage3_4[67], stage3_4[68], stage3_4[69], stage3_4[70], stage3_4[71], stage3_4[72]},
      {stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33], stage3_6[34], stage3_6[35]},
      {stage4_8[10],stage4_7[11],stage4_6[15],stage4_5[18],stage4_4[21]}
   );
   gpc606_5 gpc8642 (
      {stage3_4[73], stage3_4[74], stage3_4[75], stage3_4[76], stage3_4[77], stage3_4[78]},
      {stage3_6[36], stage3_6[37], stage3_6[38], stage3_6[39], stage3_6[40], stage3_6[41]},
      {stage4_8[11],stage4_7[12],stage4_6[16],stage4_5[19],stage4_4[22]}
   );
   gpc606_5 gpc8643 (
      {stage3_4[79], stage3_4[80], stage3_4[81], stage3_4[82], stage3_4[83], stage3_4[84]},
      {stage3_6[42], stage3_6[43], stage3_6[44], stage3_6[45], stage3_6[46], stage3_6[47]},
      {stage4_8[12],stage4_7[13],stage4_6[17],stage4_5[20],stage4_4[23]}
   );
   gpc606_5 gpc8644 (
      {stage3_4[85], stage3_4[86], stage3_4[87], stage3_4[88], stage3_4[89], stage3_4[90]},
      {stage3_6[48], stage3_6[49], stage3_6[50], stage3_6[51], stage3_6[52], stage3_6[53]},
      {stage4_8[13],stage4_7[14],stage4_6[18],stage4_5[21],stage4_4[24]}
   );
   gpc606_5 gpc8645 (
      {stage3_4[91], stage3_4[92], stage3_4[93], stage3_4[94], stage3_4[95], stage3_4[96]},
      {stage3_6[54], stage3_6[55], stage3_6[56], stage3_6[57], stage3_6[58], stage3_6[59]},
      {stage4_8[14],stage4_7[15],stage4_6[19],stage4_5[22],stage4_4[25]}
   );
   gpc606_5 gpc8646 (
      {stage3_4[97], stage3_4[98], stage3_4[99], stage3_4[100], stage3_4[101], stage3_4[102]},
      {stage3_6[60], stage3_6[61], stage3_6[62], stage3_6[63], stage3_6[64], stage3_6[65]},
      {stage4_8[15],stage4_7[16],stage4_6[20],stage4_5[23],stage4_4[26]}
   );
   gpc606_5 gpc8647 (
      {stage3_4[103], stage3_4[104], stage3_4[105], stage3_4[106], stage3_4[107], stage3_4[108]},
      {stage3_6[66], stage3_6[67], stage3_6[68], stage3_6[69], stage3_6[70], stage3_6[71]},
      {stage4_8[16],stage4_7[17],stage4_6[21],stage4_5[24],stage4_4[27]}
   );
   gpc615_5 gpc8648 (
      {stage3_6[72], stage3_6[73], stage3_6[74], stage3_6[75], stage3_6[76]},
      {stage3_7[6]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[17],stage4_7[18],stage4_6[22]}
   );
   gpc615_5 gpc8649 (
      {stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[18],stage4_7[19]}
   );
   gpc615_5 gpc8650 (
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16]},
      {stage3_8[7]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[2],stage4_9[2],stage4_8[19],stage4_7[20]}
   );
   gpc615_5 gpc8651 (
      {stage3_7[17], stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21]},
      {stage3_8[8]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[3],stage4_9[3],stage4_8[20],stage4_7[21]}
   );
   gpc615_5 gpc8652 (
      {stage3_7[22], stage3_7[23], stage3_7[24], stage3_7[25], stage3_7[26]},
      {stage3_8[9]},
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage4_11[3],stage4_10[4],stage4_9[4],stage4_8[21],stage4_7[22]}
   );
   gpc615_5 gpc8653 (
      {stage3_7[27], stage3_7[28], stage3_7[29], stage3_7[30], stage3_7[31]},
      {stage3_8[10]},
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage4_11[4],stage4_10[5],stage4_9[5],stage4_8[22],stage4_7[23]}
   );
   gpc615_5 gpc8654 (
      {stage3_7[32], stage3_7[33], stage3_7[34], stage3_7[35], stage3_7[36]},
      {stage3_8[11]},
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage4_11[5],stage4_10[6],stage4_9[6],stage4_8[23],stage4_7[24]}
   );
   gpc606_5 gpc8655 (
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[6],stage4_10[7],stage4_9[7],stage4_8[24]}
   );
   gpc606_5 gpc8656 (
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22], stage3_8[23]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[7],stage4_10[8],stage4_9[8],stage4_8[25]}
   );
   gpc606_5 gpc8657 (
      {stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27], stage3_8[28], stage3_8[29]},
      {stage3_10[12], stage3_10[13], stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17]},
      {stage4_12[2],stage4_11[8],stage4_10[9],stage4_9[9],stage4_8[26]}
   );
   gpc606_5 gpc8658 (
      {stage3_8[30], stage3_8[31], stage3_8[32], stage3_8[33], stage3_8[34], 1'b0},
      {stage3_10[18], stage3_10[19], stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23]},
      {stage4_12[3],stage4_11[9],stage4_10[10],stage4_9[10],stage4_8[27]}
   );
   gpc606_5 gpc8659 (
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[4],stage4_11[10],stage4_10[11],stage4_9[11]}
   );
   gpc606_5 gpc8660 (
      {stage3_9[42], stage3_9[43], stage3_9[44], stage3_9[45], stage3_9[46], stage3_9[47]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[5],stage4_11[11],stage4_10[12],stage4_9[12]}
   );
   gpc606_5 gpc8661 (
      {stage3_9[48], stage3_9[49], stage3_9[50], stage3_9[51], stage3_9[52], stage3_9[53]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[6],stage4_11[12],stage4_10[13],stage4_9[13]}
   );
   gpc615_5 gpc8662 (
      {stage3_10[24], stage3_10[25], stage3_10[26], stage3_10[27], stage3_10[28]},
      {stage3_11[18]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[3],stage4_12[7],stage4_11[13],stage4_10[14]}
   );
   gpc615_5 gpc8663 (
      {stage3_10[29], stage3_10[30], stage3_10[31], stage3_10[32], stage3_10[33]},
      {stage3_11[19]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[4],stage4_12[8],stage4_11[14],stage4_10[15]}
   );
   gpc615_5 gpc8664 (
      {stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37], stage3_10[38]},
      {stage3_11[20]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[5],stage4_12[9],stage4_11[15],stage4_10[16]}
   );
   gpc615_5 gpc8665 (
      {stage3_10[39], stage3_10[40], stage3_10[41], stage3_10[42], stage3_10[43]},
      {stage3_11[21]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage4_14[3],stage4_13[6],stage4_12[10],stage4_11[16],stage4_10[17]}
   );
   gpc615_5 gpc8666 (
      {stage3_10[44], stage3_10[45], stage3_10[46], stage3_10[47], stage3_10[48]},
      {stage3_11[22]},
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage4_14[4],stage4_13[7],stage4_12[11],stage4_11[17],stage4_10[18]}
   );
   gpc615_5 gpc8667 (
      {stage3_10[49], stage3_10[50], stage3_10[51], stage3_10[52], stage3_10[53]},
      {stage3_11[23]},
      {stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35]},
      {stage4_14[5],stage4_13[8],stage4_12[12],stage4_11[18],stage4_10[19]}
   );
   gpc615_5 gpc8668 (
      {stage3_10[54], stage3_10[55], stage3_10[56], stage3_10[57], stage3_10[58]},
      {stage3_11[24]},
      {stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40], stage3_12[41]},
      {stage4_14[6],stage4_13[9],stage4_12[13],stage4_11[19],stage4_10[20]}
   );
   gpc615_5 gpc8669 (
      {stage3_10[59], stage3_10[60], stage3_10[61], stage3_10[62], stage3_10[63]},
      {stage3_11[25]},
      {stage3_12[42], stage3_12[43], stage3_12[44], stage3_12[45], stage3_12[46], stage3_12[47]},
      {stage4_14[7],stage4_13[10],stage4_12[14],stage4_11[20],stage4_10[21]}
   );
   gpc615_5 gpc8670 (
      {stage3_10[64], stage3_10[65], stage3_10[66], stage3_10[67], stage3_10[68]},
      {stage3_11[26]},
      {stage3_12[48], stage3_12[49], stage3_12[50], stage3_12[51], stage3_12[52], stage3_12[53]},
      {stage4_14[8],stage4_13[11],stage4_12[15],stage4_11[21],stage4_10[22]}
   );
   gpc615_5 gpc8671 (
      {stage3_10[69], stage3_10[70], stage3_10[71], stage3_10[72], stage3_10[73]},
      {stage3_11[27]},
      {stage3_12[54], stage3_12[55], stage3_12[56], stage3_12[57], stage3_12[58], stage3_12[59]},
      {stage4_14[9],stage4_13[12],stage4_12[16],stage4_11[22],stage4_10[23]}
   );
   gpc1325_5 gpc8672 (
      {stage3_10[74], stage3_10[75], stage3_10[76], stage3_10[77], stage3_10[78]},
      {stage3_11[28], stage3_11[29]},
      {stage3_12[60], stage3_12[61], stage3_12[62]},
      {stage3_13[0]},
      {stage4_14[10],stage4_13[13],stage4_12[17],stage4_11[23],stage4_10[24]}
   );
   gpc1325_5 gpc8673 (
      {stage3_10[79], stage3_10[80], stage3_10[81], stage3_10[82], stage3_10[83]},
      {stage3_11[30], stage3_11[31]},
      {stage3_12[63], stage3_12[64], stage3_12[65]},
      {stage3_13[1]},
      {stage4_14[11],stage4_13[14],stage4_12[18],stage4_11[24],stage4_10[25]}
   );
   gpc207_4 gpc8674 (
      {stage3_11[32], stage3_11[33], stage3_11[34], stage3_11[35], stage3_11[36], stage3_11[37], stage3_11[38]},
      {stage3_13[2], stage3_13[3]},
      {stage4_14[12],stage4_13[15],stage4_12[19],stage4_11[25]}
   );
   gpc207_4 gpc8675 (
      {stage3_11[39], stage3_11[40], stage3_11[41], stage3_11[42], stage3_11[43], stage3_11[44], stage3_11[45]},
      {stage3_13[4], stage3_13[5]},
      {stage4_14[13],stage4_13[16],stage4_12[20],stage4_11[26]}
   );
   gpc207_4 gpc8676 (
      {stage3_11[46], stage3_11[47], stage3_11[48], stage3_11[49], stage3_11[50], stage3_11[51], stage3_11[52]},
      {stage3_13[6], stage3_13[7]},
      {stage4_14[14],stage4_13[17],stage4_12[21],stage4_11[27]}
   );
   gpc615_5 gpc8677 (
      {stage3_11[53], stage3_11[54], stage3_11[55], stage3_11[56], stage3_11[57]},
      {stage3_12[66]},
      {stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], stage3_13[13]},
      {stage4_15[0],stage4_14[15],stage4_13[18],stage4_12[22],stage4_11[28]}
   );
   gpc606_5 gpc8678 (
      {stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[0],stage4_15[1],stage4_14[16],stage4_13[19]}
   );
   gpc606_5 gpc8679 (
      {stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24], stage3_13[25]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[1],stage4_15[2],stage4_14[17],stage4_13[20]}
   );
   gpc606_5 gpc8680 (
      {stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30], stage3_13[31]},
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17]},
      {stage4_17[2],stage4_16[2],stage4_15[3],stage4_14[18],stage4_13[21]}
   );
   gpc606_5 gpc8681 (
      {stage3_13[32], stage3_13[33], stage3_13[34], stage3_13[35], stage3_13[36], stage3_13[37]},
      {stage3_15[18], stage3_15[19], stage3_15[20], stage3_15[21], stage3_15[22], stage3_15[23]},
      {stage4_17[3],stage4_16[3],stage4_15[4],stage4_14[19],stage4_13[22]}
   );
   gpc606_5 gpc8682 (
      {stage3_13[38], stage3_13[39], stage3_13[40], stage3_13[41], stage3_13[42], stage3_13[43]},
      {stage3_15[24], stage3_15[25], stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29]},
      {stage4_17[4],stage4_16[4],stage4_15[5],stage4_14[20],stage4_13[23]}
   );
   gpc606_5 gpc8683 (
      {stage3_13[44], stage3_13[45], stage3_13[46], stage3_13[47], stage3_13[48], stage3_13[49]},
      {stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34], stage3_15[35]},
      {stage4_17[5],stage4_16[5],stage4_15[6],stage4_14[21],stage4_13[24]}
   );
   gpc615_5 gpc8684 (
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4]},
      {stage3_15[36]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[6],stage4_16[6],stage4_15[7],stage4_14[22]}
   );
   gpc615_5 gpc8685 (
      {stage3_14[5], stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9]},
      {stage3_15[37]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[7],stage4_16[7],stage4_15[8],stage4_14[23]}
   );
   gpc615_5 gpc8686 (
      {stage3_14[10], stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14]},
      {stage3_15[38]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[8],stage4_16[8],stage4_15[9],stage4_14[24]}
   );
   gpc615_5 gpc8687 (
      {stage3_14[15], stage3_14[16], stage3_14[17], stage3_14[18], stage3_14[19]},
      {stage3_15[39]},
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23]},
      {stage4_18[3],stage4_17[9],stage4_16[9],stage4_15[10],stage4_14[25]}
   );
   gpc615_5 gpc8688 (
      {stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23], stage3_14[24]},
      {stage3_15[40]},
      {stage3_16[24], stage3_16[25], stage3_16[26], stage3_16[27], stage3_16[28], stage3_16[29]},
      {stage4_18[4],stage4_17[10],stage4_16[10],stage4_15[11],stage4_14[26]}
   );
   gpc615_5 gpc8689 (
      {stage3_14[25], stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29]},
      {stage3_15[41]},
      {stage3_16[30], stage3_16[31], stage3_16[32], stage3_16[33], stage3_16[34], stage3_16[35]},
      {stage4_18[5],stage4_17[11],stage4_16[11],stage4_15[12],stage4_14[27]}
   );
   gpc615_5 gpc8690 (
      {stage3_15[42], stage3_15[43], stage3_15[44], stage3_15[45], stage3_15[46]},
      {stage3_16[36]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[6],stage4_17[12],stage4_16[12],stage4_15[13]}
   );
   gpc606_5 gpc8691 (
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[0],stage4_19[1],stage4_18[7],stage4_17[13]}
   );
   gpc606_5 gpc8692 (
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[1],stage4_19[2],stage4_18[8],stage4_17[14]}
   );
   gpc606_5 gpc8693 (
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17]},
      {stage4_21[2],stage4_20[2],stage4_19[3],stage4_18[9],stage4_17[15]}
   );
   gpc606_5 gpc8694 (
      {stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29]},
      {stage3_19[18], stage3_19[19], stage3_19[20], stage3_19[21], stage3_19[22], stage3_19[23]},
      {stage4_21[3],stage4_20[3],stage4_19[4],stage4_18[10],stage4_17[16]}
   );
   gpc606_5 gpc8695 (
      {stage3_17[30], stage3_17[31], stage3_17[32], stage3_17[33], stage3_17[34], stage3_17[35]},
      {stage3_19[24], stage3_19[25], stage3_19[26], stage3_19[27], stage3_19[28], stage3_19[29]},
      {stage4_21[4],stage4_20[4],stage4_19[5],stage4_18[11],stage4_17[17]}
   );
   gpc207_4 gpc8696 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5], stage3_18[6]},
      {stage3_20[0], stage3_20[1]},
      {stage4_21[5],stage4_20[5],stage4_19[6],stage4_18[12]}
   );
   gpc207_4 gpc8697 (
      {stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12], stage3_18[13]},
      {stage3_20[2], stage3_20[3]},
      {stage4_21[6],stage4_20[6],stage4_19[7],stage4_18[13]}
   );
   gpc207_4 gpc8698 (
      {stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17], stage3_18[18], stage3_18[19], stage3_18[20]},
      {stage3_20[4], stage3_20[5]},
      {stage4_21[7],stage4_20[7],stage4_19[8],stage4_18[14]}
   );
   gpc207_4 gpc8699 (
      {stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25], stage3_18[26], stage3_18[27]},
      {stage3_20[6], stage3_20[7]},
      {stage4_21[8],stage4_20[8],stage4_19[9],stage4_18[15]}
   );
   gpc207_4 gpc8700 (
      {stage3_18[28], stage3_18[29], stage3_18[30], stage3_18[31], stage3_18[32], stage3_18[33], stage3_18[34]},
      {stage3_20[8], stage3_20[9]},
      {stage4_21[9],stage4_20[9],stage4_19[10],stage4_18[16]}
   );
   gpc207_4 gpc8701 (
      {stage3_18[35], stage3_18[36], stage3_18[37], stage3_18[38], stage3_18[39], stage3_18[40], stage3_18[41]},
      {stage3_20[10], stage3_20[11]},
      {stage4_21[10],stage4_20[10],stage4_19[11],stage4_18[17]}
   );
   gpc207_4 gpc8702 (
      {stage3_18[42], stage3_18[43], stage3_18[44], stage3_18[45], stage3_18[46], stage3_18[47], stage3_18[48]},
      {stage3_20[12], stage3_20[13]},
      {stage4_21[11],stage4_20[11],stage4_19[12],stage4_18[18]}
   );
   gpc207_4 gpc8703 (
      {stage3_18[49], stage3_18[50], stage3_18[51], stage3_18[52], stage3_18[53], stage3_18[54], stage3_18[55]},
      {stage3_20[14], stage3_20[15]},
      {stage4_21[12],stage4_20[12],stage4_19[13],stage4_18[19]}
   );
   gpc207_4 gpc8704 (
      {stage3_18[56], stage3_18[57], stage3_18[58], stage3_18[59], 1'b0, 1'b0, 1'b0},
      {stage3_20[16], stage3_20[17]},
      {stage4_21[13],stage4_20[13],stage4_19[14],stage4_18[20]}
   );
   gpc615_5 gpc8705 (
      {stage3_19[30], stage3_19[31], stage3_19[32], stage3_19[33], stage3_19[34]},
      {stage3_20[18]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[0],stage4_21[14],stage4_20[14],stage4_19[15]}
   );
   gpc606_5 gpc8706 (
      {stage3_20[19], stage3_20[20], stage3_20[21], stage3_20[22], stage3_20[23], stage3_20[24]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[15],stage4_20[15]}
   );
   gpc606_5 gpc8707 (
      {stage3_20[25], stage3_20[26], stage3_20[27], stage3_20[28], stage3_20[29], stage3_20[30]},
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11]},
      {stage4_24[1],stage4_23[2],stage4_22[2],stage4_21[16],stage4_20[16]}
   );
   gpc606_5 gpc8708 (
      {stage3_20[31], stage3_20[32], stage3_20[33], stage3_20[34], stage3_20[35], stage3_20[36]},
      {stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16], stage3_22[17]},
      {stage4_24[2],stage4_23[3],stage4_22[3],stage4_21[17],stage4_20[17]}
   );
   gpc606_5 gpc8709 (
      {stage3_20[37], stage3_20[38], stage3_20[39], stage3_20[40], stage3_20[41], stage3_20[42]},
      {stage3_22[18], stage3_22[19], stage3_22[20], stage3_22[21], stage3_22[22], stage3_22[23]},
      {stage4_24[3],stage4_23[4],stage4_22[4],stage4_21[18],stage4_20[18]}
   );
   gpc606_5 gpc8710 (
      {stage3_20[43], stage3_20[44], stage3_20[45], stage3_20[46], stage3_20[47], stage3_20[48]},
      {stage3_22[24], stage3_22[25], stage3_22[26], stage3_22[27], stage3_22[28], stage3_22[29]},
      {stage4_24[4],stage4_23[5],stage4_22[5],stage4_21[19],stage4_20[19]}
   );
   gpc606_5 gpc8711 (
      {stage3_20[49], stage3_20[50], stage3_20[51], stage3_20[52], stage3_20[53], stage3_20[54]},
      {stage3_22[30], stage3_22[31], stage3_22[32], stage3_22[33], stage3_22[34], stage3_22[35]},
      {stage4_24[5],stage4_23[6],stage4_22[6],stage4_21[20],stage4_20[20]}
   );
   gpc606_5 gpc8712 (
      {stage3_20[55], stage3_20[56], stage3_20[57], stage3_20[58], stage3_20[59], stage3_20[60]},
      {stage3_22[36], stage3_22[37], stage3_22[38], stage3_22[39], stage3_22[40], stage3_22[41]},
      {stage4_24[6],stage4_23[7],stage4_22[7],stage4_21[21],stage4_20[21]}
   );
   gpc606_5 gpc8713 (
      {stage3_20[61], stage3_20[62], stage3_20[63], stage3_20[64], stage3_20[65], stage3_20[66]},
      {stage3_22[42], stage3_22[43], stage3_22[44], stage3_22[45], stage3_22[46], stage3_22[47]},
      {stage4_24[7],stage4_23[8],stage4_22[8],stage4_21[22],stage4_20[22]}
   );
   gpc606_5 gpc8714 (
      {stage3_20[67], stage3_20[68], stage3_20[69], stage3_20[70], stage3_20[71], stage3_20[72]},
      {stage3_22[48], stage3_22[49], stage3_22[50], stage3_22[51], stage3_22[52], stage3_22[53]},
      {stage4_24[8],stage4_23[9],stage4_22[9],stage4_21[23],stage4_20[23]}
   );
   gpc606_5 gpc8715 (
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[9],stage4_23[10],stage4_22[10],stage4_21[24]}
   );
   gpc606_5 gpc8716 (
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage4_25[1],stage4_24[10],stage4_23[11],stage4_22[11],stage4_21[25]}
   );
   gpc606_5 gpc8717 (
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage3_23[12], stage3_23[13], stage3_23[14], stage3_23[15], stage3_23[16], stage3_23[17]},
      {stage4_25[2],stage4_24[11],stage4_23[12],stage4_22[12],stage4_21[26]}
   );
   gpc606_5 gpc8718 (
      {stage3_21[24], stage3_21[25], stage3_21[26], stage3_21[27], stage3_21[28], stage3_21[29]},
      {stage3_23[18], stage3_23[19], stage3_23[20], stage3_23[21], stage3_23[22], stage3_23[23]},
      {stage4_25[3],stage4_24[12],stage4_23[13],stage4_22[13],stage4_21[27]}
   );
   gpc615_5 gpc8719 (
      {stage3_22[54], stage3_22[55], stage3_22[56], stage3_22[57], stage3_22[58]},
      {stage3_23[24]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[4],stage4_24[13],stage4_23[14],stage4_22[14]}
   );
   gpc615_5 gpc8720 (
      {stage3_22[59], stage3_22[60], stage3_22[61], stage3_22[62], stage3_22[63]},
      {stage3_23[25]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[5],stage4_24[14],stage4_23[15],stage4_22[15]}
   );
   gpc615_5 gpc8721 (
      {stage3_22[64], stage3_22[65], stage3_22[66], stage3_22[67], stage3_22[68]},
      {stage3_23[26]},
      {stage3_24[12], stage3_24[13], stage3_24[14], stage3_24[15], stage3_24[16], stage3_24[17]},
      {stage4_26[2],stage4_25[6],stage4_24[15],stage4_23[16],stage4_22[16]}
   );
   gpc615_5 gpc8722 (
      {stage3_22[69], stage3_22[70], stage3_22[71], stage3_22[72], 1'b0},
      {stage3_23[27]},
      {stage3_24[18], stage3_24[19], stage3_24[20], stage3_24[21], stage3_24[22], stage3_24[23]},
      {stage4_26[3],stage4_25[7],stage4_24[16],stage4_23[17],stage4_22[17]}
   );
   gpc615_5 gpc8723 (
      {stage3_23[28], stage3_23[29], stage3_23[30], stage3_23[31], stage3_23[32]},
      {stage3_24[24]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[4],stage4_25[8],stage4_24[17],stage4_23[18]}
   );
   gpc615_5 gpc8724 (
      {stage3_23[33], stage3_23[34], stage3_23[35], stage3_23[36], stage3_23[37]},
      {stage3_24[25]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[5],stage4_25[9],stage4_24[18],stage4_23[19]}
   );
   gpc615_5 gpc8725 (
      {stage3_23[38], stage3_23[39], stage3_23[40], stage3_23[41], stage3_23[42]},
      {stage3_24[26]},
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage4_27[2],stage4_26[6],stage4_25[10],stage4_24[19],stage4_23[20]}
   );
   gpc606_5 gpc8726 (
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[3],stage4_26[7],stage4_25[11]}
   );
   gpc1163_5 gpc8727 (
      {stage3_26[0], stage3_26[1], stage3_26[2]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage3_28[0]},
      {stage3_29[0]},
      {stage4_30[0],stage4_29[1],stage4_28[1],stage4_27[4],stage4_26[8]}
   );
   gpc1163_5 gpc8728 (
      {stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage3_28[1]},
      {stage3_29[1]},
      {stage4_30[1],stage4_29[2],stage4_28[2],stage4_27[5],stage4_26[9]}
   );
   gpc1163_5 gpc8729 (
      {stage3_26[6], stage3_26[7], stage3_26[8]},
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage3_28[2]},
      {stage3_29[2]},
      {stage4_30[2],stage4_29[3],stage4_28[3],stage4_27[6],stage4_26[10]}
   );
   gpc615_5 gpc8730 (
      {stage3_26[9], stage3_26[10], stage3_26[11], stage3_26[12], stage3_26[13]},
      {stage3_27[24]},
      {stage3_28[3], stage3_28[4], stage3_28[5], stage3_28[6], stage3_28[7], stage3_28[8]},
      {stage4_30[3],stage4_29[4],stage4_28[4],stage4_27[7],stage4_26[11]}
   );
   gpc615_5 gpc8731 (
      {stage3_26[14], stage3_26[15], stage3_26[16], stage3_26[17], stage3_26[18]},
      {stage3_27[25]},
      {stage3_28[9], stage3_28[10], stage3_28[11], stage3_28[12], stage3_28[13], stage3_28[14]},
      {stage4_30[4],stage4_29[5],stage4_28[5],stage4_27[8],stage4_26[12]}
   );
   gpc615_5 gpc8732 (
      {stage3_26[19], stage3_26[20], stage3_26[21], stage3_26[22], stage3_26[23]},
      {stage3_27[26]},
      {stage3_28[15], stage3_28[16], stage3_28[17], stage3_28[18], stage3_28[19], stage3_28[20]},
      {stage4_30[5],stage4_29[6],stage4_28[6],stage4_27[9],stage4_26[13]}
   );
   gpc615_5 gpc8733 (
      {stage3_26[24], stage3_26[25], stage3_26[26], stage3_26[27], stage3_26[28]},
      {stage3_27[27]},
      {stage3_28[21], stage3_28[22], stage3_28[23], stage3_28[24], stage3_28[25], stage3_28[26]},
      {stage4_30[6],stage4_29[7],stage4_28[7],stage4_27[10],stage4_26[14]}
   );
   gpc615_5 gpc8734 (
      {stage3_26[29], stage3_26[30], stage3_26[31], stage3_26[32], stage3_26[33]},
      {stage3_27[28]},
      {stage3_28[27], stage3_28[28], stage3_28[29], stage3_28[30], stage3_28[31], stage3_28[32]},
      {stage4_30[7],stage4_29[8],stage4_28[8],stage4_27[11],stage4_26[15]}
   );
   gpc615_5 gpc8735 (
      {stage3_26[34], stage3_26[35], stage3_26[36], stage3_26[37], stage3_26[38]},
      {stage3_27[29]},
      {stage3_28[33], stage3_28[34], stage3_28[35], stage3_28[36], stage3_28[37], stage3_28[38]},
      {stage4_30[8],stage4_29[9],stage4_28[9],stage4_27[12],stage4_26[16]}
   );
   gpc615_5 gpc8736 (
      {stage3_26[39], stage3_26[40], stage3_26[41], stage3_26[42], stage3_26[43]},
      {stage3_27[30]},
      {stage3_28[39], stage3_28[40], stage3_28[41], stage3_28[42], stage3_28[43], stage3_28[44]},
      {stage4_30[9],stage4_29[10],stage4_28[10],stage4_27[13],stage4_26[17]}
   );
   gpc615_5 gpc8737 (
      {stage3_26[44], stage3_26[45], stage3_26[46], stage3_26[47], stage3_26[48]},
      {stage3_27[31]},
      {stage3_28[45], stage3_28[46], stage3_28[47], stage3_28[48], stage3_28[49], stage3_28[50]},
      {stage4_30[10],stage4_29[11],stage4_28[11],stage4_27[14],stage4_26[18]}
   );
   gpc606_5 gpc8738 (
      {stage3_27[32], stage3_27[33], stage3_27[34], stage3_27[35], stage3_27[36], stage3_27[37]},
      {stage3_29[3], stage3_29[4], stage3_29[5], stage3_29[6], stage3_29[7], stage3_29[8]},
      {stage4_31[0],stage4_30[11],stage4_29[12],stage4_28[12],stage4_27[15]}
   );
   gpc1163_5 gpc8739 (
      {stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[0]},
      {stage3_32[0]},
      {stage4_33[0],stage4_32[0],stage4_31[1],stage4_30[12],stage4_29[13]}
   );
   gpc1163_5 gpc8740 (
      {stage3_29[12], stage3_29[13], stage3_29[14]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage3_31[1]},
      {stage3_32[1]},
      {stage4_33[1],stage4_32[1],stage4_31[2],stage4_30[13],stage4_29[14]}
   );
   gpc1163_5 gpc8741 (
      {stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage3_31[2]},
      {stage3_32[2]},
      {stage4_33[2],stage4_32[2],stage4_31[3],stage4_30[14],stage4_29[15]}
   );
   gpc1163_5 gpc8742 (
      {stage3_29[18], stage3_29[19], stage3_29[20]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage3_31[3]},
      {stage3_32[3]},
      {stage4_33[3],stage4_32[3],stage4_31[4],stage4_30[15],stage4_29[16]}
   );
   gpc1163_5 gpc8743 (
      {stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage3_30[24], stage3_30[25], stage3_30[26], stage3_30[27], stage3_30[28], stage3_30[29]},
      {stage3_31[4]},
      {stage3_32[4]},
      {stage4_33[4],stage4_32[4],stage4_31[5],stage4_30[16],stage4_29[17]}
   );
   gpc606_5 gpc8744 (
      {stage3_29[24], stage3_29[25], stage3_29[26], stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage3_31[5], stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10]},
      {stage4_33[5],stage4_32[5],stage4_31[6],stage4_30[17],stage4_29[18]}
   );
   gpc606_5 gpc8745 (
      {stage3_29[30], stage3_29[31], stage3_29[32], stage3_29[33], stage3_29[34], stage3_29[35]},
      {stage3_31[11], stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16]},
      {stage4_33[6],stage4_32[6],stage4_31[7],stage4_30[18],stage4_29[19]}
   );
   gpc606_5 gpc8746 (
      {stage3_29[36], stage3_29[37], stage3_29[38], stage3_29[39], stage3_29[40], stage3_29[41]},
      {stage3_31[17], stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21], stage3_31[22]},
      {stage4_33[7],stage4_32[7],stage4_31[8],stage4_30[19],stage4_29[20]}
   );
   gpc606_5 gpc8747 (
      {stage3_29[42], stage3_29[43], stage3_29[44], stage3_29[45], stage3_29[46], stage3_29[47]},
      {stage3_31[23], stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27], stage3_31[28]},
      {stage4_33[8],stage4_32[8],stage4_31[9],stage4_30[20],stage4_29[21]}
   );
   gpc615_5 gpc8748 (
      {stage3_31[29], stage3_31[30], stage3_31[31], stage3_31[32], stage3_31[33]},
      {stage3_32[5]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[0],stage4_33[9],stage4_32[9],stage4_31[10]}
   );
   gpc2135_5 gpc8749 (
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10]},
      {stage3_33[6], stage3_33[7], stage3_33[8]},
      {stage3_34[0]},
      {stage3_35[0], stage3_35[1]},
      {stage4_36[0],stage4_35[1],stage4_34[1],stage4_33[10],stage4_32[10]}
   );
   gpc2135_5 gpc8750 (
      {stage3_32[11], stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15]},
      {stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage3_34[1]},
      {stage3_35[2], stage3_35[3]},
      {stage4_36[1],stage4_35[2],stage4_34[2],stage4_33[11],stage4_32[11]}
   );
   gpc615_5 gpc8751 (
      {stage3_32[16], stage3_32[17], stage3_32[18], stage3_32[19], stage3_32[20]},
      {stage3_33[12]},
      {stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5], stage3_34[6], stage3_34[7]},
      {stage4_36[2],stage4_35[3],stage4_34[3],stage4_33[12],stage4_32[12]}
   );
   gpc615_5 gpc8752 (
      {stage3_32[21], stage3_32[22], stage3_32[23], stage3_32[24], stage3_32[25]},
      {stage3_33[13]},
      {stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11], stage3_34[12], stage3_34[13]},
      {stage4_36[3],stage4_35[4],stage4_34[4],stage4_33[13],stage4_32[13]}
   );
   gpc615_5 gpc8753 (
      {stage3_32[26], stage3_32[27], stage3_32[28], stage3_32[29], stage3_32[30]},
      {stage3_33[14]},
      {stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17], stage3_34[18], stage3_34[19]},
      {stage4_36[4],stage4_35[5],stage4_34[5],stage4_33[14],stage4_32[14]}
   );
   gpc615_5 gpc8754 (
      {stage3_32[31], stage3_32[32], stage3_32[33], stage3_32[34], stage3_32[35]},
      {stage3_33[15]},
      {stage3_34[20], stage3_34[21], stage3_34[22], stage3_34[23], stage3_34[24], stage3_34[25]},
      {stage4_36[5],stage4_35[6],stage4_34[6],stage4_33[15],stage4_32[15]}
   );
   gpc615_5 gpc8755 (
      {stage3_32[36], stage3_32[37], stage3_32[38], stage3_32[39], stage3_32[40]},
      {stage3_33[16]},
      {stage3_34[26], stage3_34[27], stage3_34[28], stage3_34[29], stage3_34[30], stage3_34[31]},
      {stage4_36[6],stage4_35[7],stage4_34[7],stage4_33[16],stage4_32[16]}
   );
   gpc117_4 gpc8756 (
      {stage3_33[17], stage3_33[18], stage3_33[19], stage3_33[20], stage3_33[21], stage3_33[22], stage3_33[23]},
      {stage3_34[32]},
      {stage3_35[4]},
      {stage4_36[7],stage4_35[8],stage4_34[8],stage4_33[17]}
   );
   gpc117_4 gpc8757 (
      {stage3_33[24], stage3_33[25], stage3_33[26], stage3_33[27], stage3_33[28], stage3_33[29], stage3_33[30]},
      {stage3_34[33]},
      {stage3_35[5]},
      {stage4_36[8],stage4_35[9],stage4_34[9],stage4_33[18]}
   );
   gpc606_5 gpc8758 (
      {stage3_33[31], stage3_33[32], stage3_33[33], stage3_33[34], stage3_33[35], stage3_33[36]},
      {stage3_35[6], stage3_35[7], stage3_35[8], stage3_35[9], stage3_35[10], stage3_35[11]},
      {stage4_37[0],stage4_36[9],stage4_35[10],stage4_34[10],stage4_33[19]}
   );
   gpc615_5 gpc8759 (
      {stage3_35[12], stage3_35[13], stage3_35[14], stage3_35[15], stage3_35[16]},
      {stage3_36[0]},
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage4_39[0],stage4_38[0],stage4_37[1],stage4_36[10],stage4_35[11]}
   );
   gpc615_5 gpc8760 (
      {stage3_35[17], stage3_35[18], stage3_35[19], stage3_35[20], stage3_35[21]},
      {stage3_36[1]},
      {stage3_37[6], stage3_37[7], stage3_37[8], stage3_37[9], stage3_37[10], stage3_37[11]},
      {stage4_39[1],stage4_38[1],stage4_37[2],stage4_36[11],stage4_35[12]}
   );
   gpc615_5 gpc8761 (
      {stage3_35[22], stage3_35[23], stage3_35[24], stage3_35[25], stage3_35[26]},
      {stage3_36[2]},
      {stage3_37[12], stage3_37[13], stage3_37[14], stage3_37[15], stage3_37[16], stage3_37[17]},
      {stage4_39[2],stage4_38[2],stage4_37[3],stage4_36[12],stage4_35[13]}
   );
   gpc615_5 gpc8762 (
      {stage3_35[27], stage3_35[28], stage3_35[29], stage3_35[30], stage3_35[31]},
      {stage3_36[3]},
      {stage3_37[18], stage3_37[19], stage3_37[20], stage3_37[21], stage3_37[22], stage3_37[23]},
      {stage4_39[3],stage4_38[3],stage4_37[4],stage4_36[13],stage4_35[14]}
   );
   gpc615_5 gpc8763 (
      {stage3_35[32], stage3_35[33], stage3_35[34], stage3_35[35], stage3_35[36]},
      {stage3_36[4]},
      {stage3_37[24], stage3_37[25], stage3_37[26], stage3_37[27], stage3_37[28], stage3_37[29]},
      {stage4_39[4],stage4_38[4],stage4_37[5],stage4_36[14],stage4_35[15]}
   );
   gpc606_5 gpc8764 (
      {stage3_36[5], stage3_36[6], stage3_36[7], stage3_36[8], stage3_36[9], stage3_36[10]},
      {stage3_38[0], stage3_38[1], stage3_38[2], stage3_38[3], stage3_38[4], stage3_38[5]},
      {stage4_40[0],stage4_39[5],stage4_38[5],stage4_37[6],stage4_36[15]}
   );
   gpc606_5 gpc8765 (
      {stage3_36[11], stage3_36[12], stage3_36[13], stage3_36[14], stage3_36[15], stage3_36[16]},
      {stage3_38[6], stage3_38[7], stage3_38[8], stage3_38[9], stage3_38[10], stage3_38[11]},
      {stage4_40[1],stage4_39[6],stage4_38[6],stage4_37[7],stage4_36[16]}
   );
   gpc606_5 gpc8766 (
      {stage3_36[17], stage3_36[18], stage3_36[19], stage3_36[20], stage3_36[21], stage3_36[22]},
      {stage3_38[12], stage3_38[13], stage3_38[14], stage3_38[15], stage3_38[16], stage3_38[17]},
      {stage4_40[2],stage4_39[7],stage4_38[7],stage4_37[8],stage4_36[17]}
   );
   gpc606_5 gpc8767 (
      {stage3_36[23], stage3_36[24], stage3_36[25], stage3_36[26], stage3_36[27], stage3_36[28]},
      {stage3_38[18], stage3_38[19], stage3_38[20], stage3_38[21], stage3_38[22], stage3_38[23]},
      {stage4_40[3],stage4_39[8],stage4_38[8],stage4_37[9],stage4_36[18]}
   );
   gpc606_5 gpc8768 (
      {stage3_37[30], stage3_37[31], stage3_37[32], stage3_37[33], stage3_37[34], stage3_37[35]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[4],stage4_39[9],stage4_38[9],stage4_37[10]}
   );
   gpc606_5 gpc8769 (
      {stage3_37[36], stage3_37[37], stage3_37[38], stage3_37[39], stage3_37[40], stage3_37[41]},
      {stage3_39[6], stage3_39[7], stage3_39[8], stage3_39[9], stage3_39[10], stage3_39[11]},
      {stage4_41[1],stage4_40[5],stage4_39[10],stage4_38[10],stage4_37[11]}
   );
   gpc606_5 gpc8770 (
      {stage3_37[42], stage3_37[43], stage3_37[44], stage3_37[45], stage3_37[46], stage3_37[47]},
      {stage3_39[12], stage3_39[13], stage3_39[14], stage3_39[15], stage3_39[16], stage3_39[17]},
      {stage4_41[2],stage4_40[6],stage4_39[11],stage4_38[11],stage4_37[12]}
   );
   gpc615_5 gpc8771 (
      {stage3_38[24], stage3_38[25], stage3_38[26], stage3_38[27], stage3_38[28]},
      {stage3_39[18]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[3],stage4_40[7],stage4_39[12],stage4_38[12]}
   );
   gpc615_5 gpc8772 (
      {stage3_38[29], stage3_38[30], stage3_38[31], stage3_38[32], stage3_38[33]},
      {stage3_39[19]},
      {stage3_40[6], stage3_40[7], stage3_40[8], stage3_40[9], stage3_40[10], stage3_40[11]},
      {stage4_42[1],stage4_41[4],stage4_40[8],stage4_39[13],stage4_38[13]}
   );
   gpc615_5 gpc8773 (
      {stage3_38[34], stage3_38[35], stage3_38[36], stage3_38[37], stage3_38[38]},
      {stage3_39[20]},
      {stage3_40[12], stage3_40[13], stage3_40[14], stage3_40[15], stage3_40[16], stage3_40[17]},
      {stage4_42[2],stage4_41[5],stage4_40[9],stage4_39[14],stage4_38[14]}
   );
   gpc615_5 gpc8774 (
      {stage3_38[39], stage3_38[40], stage3_38[41], stage3_38[42], stage3_38[43]},
      {stage3_39[21]},
      {stage3_40[18], stage3_40[19], stage3_40[20], stage3_40[21], stage3_40[22], stage3_40[23]},
      {stage4_42[3],stage4_41[6],stage4_40[10],stage4_39[15],stage4_38[15]}
   );
   gpc615_5 gpc8775 (
      {stage3_38[44], stage3_38[45], stage3_38[46], stage3_38[47], stage3_38[48]},
      {stage3_39[22]},
      {stage3_40[24], stage3_40[25], stage3_40[26], stage3_40[27], stage3_40[28], stage3_40[29]},
      {stage4_42[4],stage4_41[7],stage4_40[11],stage4_39[16],stage4_38[16]}
   );
   gpc615_5 gpc8776 (
      {stage3_38[49], stage3_38[50], stage3_38[51], stage3_38[52], stage3_38[53]},
      {stage3_39[23]},
      {stage3_40[30], stage3_40[31], stage3_40[32], stage3_40[33], stage3_40[34], stage3_40[35]},
      {stage4_42[5],stage4_41[8],stage4_40[12],stage4_39[17],stage4_38[17]}
   );
   gpc615_5 gpc8777 (
      {stage3_38[54], stage3_38[55], stage3_38[56], stage3_38[57], stage3_38[58]},
      {stage3_39[24]},
      {stage3_40[36], stage3_40[37], stage3_40[38], stage3_40[39], stage3_40[40], stage3_40[41]},
      {stage4_42[6],stage4_41[9],stage4_40[13],stage4_39[18],stage4_38[18]}
   );
   gpc207_4 gpc8778 (
      {stage3_39[25], stage3_39[26], stage3_39[27], stage3_39[28], stage3_39[29], stage3_39[30], stage3_39[31]},
      {stage3_41[0], stage3_41[1]},
      {stage4_42[7],stage4_41[10],stage4_40[14],stage4_39[19]}
   );
   gpc207_4 gpc8779 (
      {stage3_39[32], stage3_39[33], stage3_39[34], stage3_39[35], stage3_39[36], stage3_39[37], stage3_39[38]},
      {stage3_41[2], stage3_41[3]},
      {stage4_42[8],stage4_41[11],stage4_40[15],stage4_39[20]}
   );
   gpc207_4 gpc8780 (
      {stage3_39[39], stage3_39[40], stage3_39[41], stage3_39[42], stage3_39[43], stage3_39[44], stage3_39[45]},
      {stage3_41[4], stage3_41[5]},
      {stage4_42[9],stage4_41[12],stage4_40[16],stage4_39[21]}
   );
   gpc207_4 gpc8781 (
      {stage3_39[46], stage3_39[47], stage3_39[48], stage3_39[49], stage3_39[50], stage3_39[51], stage3_39[52]},
      {stage3_41[6], stage3_41[7]},
      {stage4_42[10],stage4_41[13],stage4_40[17],stage4_39[22]}
   );
   gpc615_5 gpc8782 (
      {stage3_39[53], stage3_39[54], stage3_39[55], stage3_39[56], stage3_39[57]},
      {stage3_40[42]},
      {stage3_41[8], stage3_41[9], stage3_41[10], stage3_41[11], stage3_41[12], stage3_41[13]},
      {stage4_43[0],stage4_42[11],stage4_41[14],stage4_40[18],stage4_39[23]}
   );
   gpc606_5 gpc8783 (
      {stage3_41[14], stage3_41[15], stage3_41[16], stage3_41[17], stage3_41[18], stage3_41[19]},
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4], stage3_43[5]},
      {stage4_45[0],stage4_44[0],stage4_43[1],stage4_42[12],stage4_41[15]}
   );
   gpc606_5 gpc8784 (
      {stage3_41[20], stage3_41[21], stage3_41[22], stage3_41[23], stage3_41[24], stage3_41[25]},
      {stage3_43[6], stage3_43[7], stage3_43[8], stage3_43[9], stage3_43[10], stage3_43[11]},
      {stage4_45[1],stage4_44[1],stage4_43[2],stage4_42[13],stage4_41[16]}
   );
   gpc606_5 gpc8785 (
      {stage3_41[26], stage3_41[27], stage3_41[28], stage3_41[29], stage3_41[30], stage3_41[31]},
      {stage3_43[12], stage3_43[13], stage3_43[14], stage3_43[15], stage3_43[16], stage3_43[17]},
      {stage4_45[2],stage4_44[2],stage4_43[3],stage4_42[14],stage4_41[17]}
   );
   gpc606_5 gpc8786 (
      {stage3_41[32], stage3_41[33], stage3_41[34], stage3_41[35], stage3_41[36], stage3_41[37]},
      {stage3_43[18], stage3_43[19], stage3_43[20], stage3_43[21], stage3_43[22], stage3_43[23]},
      {stage4_45[3],stage4_44[3],stage4_43[4],stage4_42[15],stage4_41[18]}
   );
   gpc606_5 gpc8787 (
      {stage3_41[38], stage3_41[39], stage3_41[40], stage3_41[41], stage3_41[42], 1'b0},
      {stage3_43[24], stage3_43[25], stage3_43[26], stage3_43[27], stage3_43[28], stage3_43[29]},
      {stage4_45[4],stage4_44[4],stage4_43[5],stage4_42[16],stage4_41[19]}
   );
   gpc207_4 gpc8788 (
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4], stage3_42[5], stage3_42[6]},
      {stage3_44[0], stage3_44[1]},
      {stage4_45[5],stage4_44[5],stage4_43[6],stage4_42[17]}
   );
   gpc207_4 gpc8789 (
      {stage3_42[7], stage3_42[8], stage3_42[9], stage3_42[10], stage3_42[11], stage3_42[12], stage3_42[13]},
      {stage3_44[2], stage3_44[3]},
      {stage4_45[6],stage4_44[6],stage4_43[7],stage4_42[18]}
   );
   gpc207_4 gpc8790 (
      {stage3_42[14], stage3_42[15], stage3_42[16], stage3_42[17], stage3_42[18], stage3_42[19], stage3_42[20]},
      {stage3_44[4], stage3_44[5]},
      {stage4_45[7],stage4_44[7],stage4_43[8],stage4_42[19]}
   );
   gpc207_4 gpc8791 (
      {stage3_42[21], stage3_42[22], stage3_42[23], stage3_42[24], stage3_42[25], stage3_42[26], stage3_42[27]},
      {stage3_44[6], stage3_44[7]},
      {stage4_45[8],stage4_44[8],stage4_43[9],stage4_42[20]}
   );
   gpc606_5 gpc8792 (
      {stage3_42[28], stage3_42[29], stage3_42[30], stage3_42[31], stage3_42[32], stage3_42[33]},
      {stage3_44[8], stage3_44[9], stage3_44[10], stage3_44[11], stage3_44[12], stage3_44[13]},
      {stage4_46[0],stage4_45[9],stage4_44[9],stage4_43[10],stage4_42[21]}
   );
   gpc606_5 gpc8793 (
      {stage3_43[30], stage3_43[31], stage3_43[32], stage3_43[33], stage3_43[34], stage3_43[35]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3], stage3_45[4], stage3_45[5]},
      {stage4_47[0],stage4_46[1],stage4_45[10],stage4_44[10],stage4_43[11]}
   );
   gpc606_5 gpc8794 (
      {stage3_43[36], stage3_43[37], stage3_43[38], stage3_43[39], stage3_43[40], stage3_43[41]},
      {stage3_45[6], stage3_45[7], stage3_45[8], stage3_45[9], stage3_45[10], stage3_45[11]},
      {stage4_47[1],stage4_46[2],stage4_45[11],stage4_44[11],stage4_43[12]}
   );
   gpc615_5 gpc8795 (
      {stage3_43[42], stage3_43[43], stage3_43[44], stage3_43[45], 1'b0},
      {stage3_44[14]},
      {stage3_45[12], stage3_45[13], stage3_45[14], stage3_45[15], stage3_45[16], stage3_45[17]},
      {stage4_47[2],stage4_46[3],stage4_45[12],stage4_44[12],stage4_43[13]}
   );
   gpc606_5 gpc8796 (
      {stage3_44[15], stage3_44[16], stage3_44[17], stage3_44[18], stage3_44[19], stage3_44[20]},
      {stage3_46[0], stage3_46[1], stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5]},
      {stage4_48[0],stage4_47[3],stage4_46[4],stage4_45[13],stage4_44[13]}
   );
   gpc606_5 gpc8797 (
      {stage3_44[21], stage3_44[22], stage3_44[23], stage3_44[24], stage3_44[25], stage3_44[26]},
      {stage3_46[6], stage3_46[7], stage3_46[8], stage3_46[9], stage3_46[10], stage3_46[11]},
      {stage4_48[1],stage4_47[4],stage4_46[5],stage4_45[14],stage4_44[14]}
   );
   gpc615_5 gpc8798 (
      {stage3_44[27], stage3_44[28], stage3_44[29], stage3_44[30], stage3_44[31]},
      {stage3_45[18]},
      {stage3_46[12], stage3_46[13], stage3_46[14], stage3_46[15], stage3_46[16], stage3_46[17]},
      {stage4_48[2],stage4_47[5],stage4_46[6],stage4_45[15],stage4_44[15]}
   );
   gpc135_4 gpc8799 (
      {stage3_45[19], stage3_45[20], stage3_45[21], stage3_45[22], stage3_45[23]},
      {stage3_46[18], stage3_46[19], stage3_46[20]},
      {stage3_47[0]},
      {stage4_48[3],stage4_47[6],stage4_46[7],stage4_45[16]}
   );
   gpc135_4 gpc8800 (
      {stage3_45[24], stage3_45[25], stage3_45[26], stage3_45[27], stage3_45[28]},
      {stage3_46[21], stage3_46[22], stage3_46[23]},
      {stage3_47[1]},
      {stage4_48[4],stage4_47[7],stage4_46[8],stage4_45[17]}
   );
   gpc135_4 gpc8801 (
      {stage3_45[29], stage3_45[30], stage3_45[31], stage3_45[32], stage3_45[33]},
      {stage3_46[24], stage3_46[25], stage3_46[26]},
      {stage3_47[2]},
      {stage4_48[5],stage4_47[8],stage4_46[9],stage4_45[18]}
   );
   gpc615_5 gpc8802 (
      {stage3_46[27], stage3_46[28], stage3_46[29], stage3_46[30], stage3_46[31]},
      {stage3_47[3]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[0],stage4_48[6],stage4_47[9],stage4_46[10]}
   );
   gpc615_5 gpc8803 (
      {stage3_46[32], stage3_46[33], stage3_46[34], stage3_46[35], stage3_46[36]},
      {stage3_47[4]},
      {stage3_48[6], stage3_48[7], stage3_48[8], stage3_48[9], stage3_48[10], stage3_48[11]},
      {stage4_50[1],stage4_49[1],stage4_48[7],stage4_47[10],stage4_46[11]}
   );
   gpc615_5 gpc8804 (
      {stage3_46[37], stage3_46[38], stage3_46[39], stage3_46[40], stage3_46[41]},
      {stage3_47[5]},
      {stage3_48[12], stage3_48[13], stage3_48[14], stage3_48[15], stage3_48[16], stage3_48[17]},
      {stage4_50[2],stage4_49[2],stage4_48[8],stage4_47[11],stage4_46[12]}
   );
   gpc615_5 gpc8805 (
      {stage3_46[42], stage3_46[43], stage3_46[44], stage3_46[45], stage3_46[46]},
      {stage3_47[6]},
      {stage3_48[18], stage3_48[19], stage3_48[20], stage3_48[21], stage3_48[22], stage3_48[23]},
      {stage4_50[3],stage4_49[3],stage4_48[9],stage4_47[12],stage4_46[13]}
   );
   gpc615_5 gpc8806 (
      {stage3_46[47], stage3_46[48], stage3_46[49], stage3_46[50], stage3_46[51]},
      {stage3_47[7]},
      {stage3_48[24], stage3_48[25], stage3_48[26], stage3_48[27], stage3_48[28], stage3_48[29]},
      {stage4_50[4],stage4_49[4],stage4_48[10],stage4_47[13],stage4_46[14]}
   );
   gpc615_5 gpc8807 (
      {stage3_46[52], stage3_46[53], stage3_46[54], stage3_46[55], stage3_46[56]},
      {stage3_47[8]},
      {stage3_48[30], stage3_48[31], stage3_48[32], stage3_48[33], stage3_48[34], stage3_48[35]},
      {stage4_50[5],stage4_49[5],stage4_48[11],stage4_47[14],stage4_46[15]}
   );
   gpc606_5 gpc8808 (
      {stage3_47[9], stage3_47[10], stage3_47[11], stage3_47[12], stage3_47[13], stage3_47[14]},
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5]},
      {stage4_51[0],stage4_50[6],stage4_49[6],stage4_48[12],stage4_47[15]}
   );
   gpc606_5 gpc8809 (
      {stage3_47[15], stage3_47[16], stage3_47[17], stage3_47[18], stage3_47[19], stage3_47[20]},
      {stage3_49[6], stage3_49[7], stage3_49[8], stage3_49[9], stage3_49[10], stage3_49[11]},
      {stage4_51[1],stage4_50[7],stage4_49[7],stage4_48[13],stage4_47[16]}
   );
   gpc606_5 gpc8810 (
      {stage3_47[21], stage3_47[22], stage3_47[23], stage3_47[24], stage3_47[25], stage3_47[26]},
      {stage3_49[12], stage3_49[13], stage3_49[14], stage3_49[15], stage3_49[16], stage3_49[17]},
      {stage4_51[2],stage4_50[8],stage4_49[8],stage4_48[14],stage4_47[17]}
   );
   gpc606_5 gpc8811 (
      {stage3_47[27], stage3_47[28], stage3_47[29], stage3_47[30], stage3_47[31], stage3_47[32]},
      {stage3_49[18], stage3_49[19], stage3_49[20], stage3_49[21], stage3_49[22], stage3_49[23]},
      {stage4_51[3],stage4_50[9],stage4_49[9],stage4_48[15],stage4_47[18]}
   );
   gpc606_5 gpc8812 (
      {stage3_47[33], stage3_47[34], stage3_47[35], stage3_47[36], stage3_47[37], stage3_47[38]},
      {stage3_49[24], stage3_49[25], stage3_49[26], stage3_49[27], stage3_49[28], stage3_49[29]},
      {stage4_51[4],stage4_50[10],stage4_49[10],stage4_48[16],stage4_47[19]}
   );
   gpc615_5 gpc8813 (
      {stage3_47[39], stage3_47[40], stage3_47[41], stage3_47[42], stage3_47[43]},
      {stage3_48[36]},
      {stage3_49[30], stage3_49[31], stage3_49[32], stage3_49[33], stage3_49[34], stage3_49[35]},
      {stage4_51[5],stage4_50[11],stage4_49[11],stage4_48[17],stage4_47[20]}
   );
   gpc606_5 gpc8814 (
      {stage3_49[36], stage3_49[37], stage3_49[38], stage3_49[39], stage3_49[40], stage3_49[41]},
      {stage3_51[0], stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5]},
      {stage4_53[0],stage4_52[0],stage4_51[6],stage4_50[12],stage4_49[12]}
   );
   gpc117_4 gpc8815 (
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5], stage3_50[6]},
      {stage3_51[6]},
      {stage3_52[0]},
      {stage4_53[1],stage4_52[1],stage4_51[7],stage4_50[13]}
   );
   gpc117_4 gpc8816 (
      {stage3_50[7], stage3_50[8], stage3_50[9], stage3_50[10], stage3_50[11], stage3_50[12], stage3_50[13]},
      {stage3_51[7]},
      {stage3_52[1]},
      {stage4_53[2],stage4_52[2],stage4_51[8],stage4_50[14]}
   );
   gpc615_5 gpc8817 (
      {stage3_50[14], stage3_50[15], stage3_50[16], stage3_50[17], stage3_50[18]},
      {stage3_51[8]},
      {stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5], stage3_52[6], stage3_52[7]},
      {stage4_54[0],stage4_53[3],stage4_52[3],stage4_51[9],stage4_50[15]}
   );
   gpc615_5 gpc8818 (
      {stage3_50[19], stage3_50[20], stage3_50[21], stage3_50[22], stage3_50[23]},
      {stage3_51[9]},
      {stage3_52[8], stage3_52[9], stage3_52[10], stage3_52[11], stage3_52[12], stage3_52[13]},
      {stage4_54[1],stage4_53[4],stage4_52[4],stage4_51[10],stage4_50[16]}
   );
   gpc615_5 gpc8819 (
      {stage3_50[24], stage3_50[25], stage3_50[26], stage3_50[27], stage3_50[28]},
      {stage3_51[10]},
      {stage3_52[14], stage3_52[15], stage3_52[16], stage3_52[17], stage3_52[18], stage3_52[19]},
      {stage4_54[2],stage4_53[5],stage4_52[5],stage4_51[11],stage4_50[17]}
   );
   gpc615_5 gpc8820 (
      {stage3_50[29], stage3_50[30], stage3_50[31], stage3_50[32], stage3_50[33]},
      {stage3_51[11]},
      {stage3_52[20], stage3_52[21], stage3_52[22], stage3_52[23], stage3_52[24], stage3_52[25]},
      {stage4_54[3],stage4_53[6],stage4_52[6],stage4_51[12],stage4_50[18]}
   );
   gpc615_5 gpc8821 (
      {stage3_50[34], stage3_50[35], stage3_50[36], stage3_50[37], stage3_50[38]},
      {stage3_51[12]},
      {stage3_52[26], stage3_52[27], stage3_52[28], stage3_52[29], stage3_52[30], stage3_52[31]},
      {stage4_54[4],stage4_53[7],stage4_52[7],stage4_51[13],stage4_50[19]}
   );
   gpc615_5 gpc8822 (
      {stage3_50[39], stage3_50[40], stage3_50[41], stage3_50[42], stage3_50[43]},
      {stage3_51[13]},
      {stage3_52[32], stage3_52[33], stage3_52[34], stage3_52[35], stage3_52[36], stage3_52[37]},
      {stage4_54[5],stage4_53[8],stage4_52[8],stage4_51[14],stage4_50[20]}
   );
   gpc615_5 gpc8823 (
      {stage3_50[44], stage3_50[45], stage3_50[46], 1'b0, 1'b0},
      {stage3_51[14]},
      {stage3_52[38], stage3_52[39], stage3_52[40], stage3_52[41], stage3_52[42], stage3_52[43]},
      {stage4_54[6],stage4_53[9],stage4_52[9],stage4_51[15],stage4_50[21]}
   );
   gpc2135_5 gpc8824 (
      {stage3_51[15], stage3_51[16], stage3_51[17], stage3_51[18], stage3_51[19]},
      {stage3_52[44], stage3_52[45], stage3_52[46]},
      {stage3_53[0]},
      {stage3_54[0], stage3_54[1]},
      {stage4_55[0],stage4_54[7],stage4_53[10],stage4_52[10],stage4_51[16]}
   );
   gpc2135_5 gpc8825 (
      {stage3_51[20], stage3_51[21], stage3_51[22], stage3_51[23], stage3_51[24]},
      {stage3_52[47], stage3_52[48], stage3_52[49]},
      {stage3_53[1]},
      {stage3_54[2], stage3_54[3]},
      {stage4_55[1],stage4_54[8],stage4_53[11],stage4_52[11],stage4_51[17]}
   );
   gpc2135_5 gpc8826 (
      {stage3_51[25], stage3_51[26], stage3_51[27], stage3_51[28], stage3_51[29]},
      {stage3_52[50], stage3_52[51], stage3_52[52]},
      {stage3_53[2]},
      {stage3_54[4], stage3_54[5]},
      {stage4_55[2],stage4_54[9],stage4_53[12],stage4_52[12],stage4_51[18]}
   );
   gpc2135_5 gpc8827 (
      {stage3_51[30], stage3_51[31], stage3_51[32], stage3_51[33], stage3_51[34]},
      {stage3_52[53], stage3_52[54], stage3_52[55]},
      {stage3_53[3]},
      {stage3_54[6], stage3_54[7]},
      {stage4_55[3],stage4_54[10],stage4_53[13],stage4_52[13],stage4_51[19]}
   );
   gpc2135_5 gpc8828 (
      {stage3_51[35], stage3_51[36], stage3_51[37], stage3_51[38], stage3_51[39]},
      {stage3_52[56], stage3_52[57], stage3_52[58]},
      {stage3_53[4]},
      {stage3_54[8], stage3_54[9]},
      {stage4_55[4],stage4_54[11],stage4_53[14],stage4_52[14],stage4_51[20]}
   );
   gpc615_5 gpc8829 (
      {stage3_51[40], stage3_51[41], stage3_51[42], stage3_51[43], stage3_51[44]},
      {stage3_52[59]},
      {stage3_53[5], stage3_53[6], stage3_53[7], stage3_53[8], stage3_53[9], stage3_53[10]},
      {stage4_55[5],stage4_54[12],stage4_53[15],stage4_52[15],stage4_51[21]}
   );
   gpc615_5 gpc8830 (
      {stage3_51[45], stage3_51[46], stage3_51[47], stage3_51[48], stage3_51[49]},
      {stage3_52[60]},
      {stage3_53[11], stage3_53[12], stage3_53[13], stage3_53[14], stage3_53[15], stage3_53[16]},
      {stage4_55[6],stage4_54[13],stage4_53[16],stage4_52[16],stage4_51[22]}
   );
   gpc606_5 gpc8831 (
      {stage3_53[17], stage3_53[18], stage3_53[19], stage3_53[20], stage3_53[21], stage3_53[22]},
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3], stage3_55[4], stage3_55[5]},
      {stage4_57[0],stage4_56[0],stage4_55[7],stage4_54[14],stage4_53[17]}
   );
   gpc606_5 gpc8832 (
      {stage3_53[23], stage3_53[24], stage3_53[25], stage3_53[26], stage3_53[27], stage3_53[28]},
      {stage3_55[6], stage3_55[7], stage3_55[8], stage3_55[9], stage3_55[10], stage3_55[11]},
      {stage4_57[1],stage4_56[1],stage4_55[8],stage4_54[15],stage4_53[18]}
   );
   gpc606_5 gpc8833 (
      {stage3_53[29], stage3_53[30], stage3_53[31], stage3_53[32], stage3_53[33], stage3_53[34]},
      {stage3_55[12], stage3_55[13], stage3_55[14], stage3_55[15], stage3_55[16], stage3_55[17]},
      {stage4_57[2],stage4_56[2],stage4_55[9],stage4_54[16],stage4_53[19]}
   );
   gpc615_5 gpc8834 (
      {stage3_53[35], stage3_53[36], stage3_53[37], stage3_53[38], stage3_53[39]},
      {stage3_54[10]},
      {stage3_55[18], stage3_55[19], stage3_55[20], stage3_55[21], stage3_55[22], stage3_55[23]},
      {stage4_57[3],stage4_56[3],stage4_55[10],stage4_54[17],stage4_53[20]}
   );
   gpc615_5 gpc8835 (
      {stage3_53[40], stage3_53[41], stage3_53[42], stage3_53[43], stage3_53[44]},
      {stage3_54[11]},
      {stage3_55[24], stage3_55[25], stage3_55[26], stage3_55[27], stage3_55[28], stage3_55[29]},
      {stage4_57[4],stage4_56[4],stage4_55[11],stage4_54[18],stage4_53[21]}
   );
   gpc615_5 gpc8836 (
      {stage3_53[45], stage3_53[46], stage3_53[47], stage3_53[48], stage3_53[49]},
      {stage3_54[12]},
      {stage3_55[30], stage3_55[31], stage3_55[32], stage3_55[33], stage3_55[34], stage3_55[35]},
      {stage4_57[5],stage4_56[5],stage4_55[12],stage4_54[19],stage4_53[22]}
   );
   gpc615_5 gpc8837 (
      {stage3_53[50], stage3_53[51], stage3_53[52], stage3_53[53], stage3_53[54]},
      {stage3_54[13]},
      {stage3_55[36], stage3_55[37], stage3_55[38], stage3_55[39], stage3_55[40], stage3_55[41]},
      {stage4_57[6],stage4_56[6],stage4_55[13],stage4_54[20],stage4_53[23]}
   );
   gpc615_5 gpc8838 (
      {stage3_54[14], stage3_54[15], stage3_54[16], stage3_54[17], stage3_54[18]},
      {stage3_55[42]},
      {stage3_56[0], stage3_56[1], stage3_56[2], stage3_56[3], stage3_56[4], stage3_56[5]},
      {stage4_58[0],stage4_57[7],stage4_56[7],stage4_55[14],stage4_54[21]}
   );
   gpc615_5 gpc8839 (
      {stage3_54[19], stage3_54[20], stage3_54[21], stage3_54[22], stage3_54[23]},
      {stage3_55[43]},
      {stage3_56[6], stage3_56[7], stage3_56[8], stage3_56[9], stage3_56[10], stage3_56[11]},
      {stage4_58[1],stage4_57[8],stage4_56[8],stage4_55[15],stage4_54[22]}
   );
   gpc615_5 gpc8840 (
      {stage3_54[24], stage3_54[25], stage3_54[26], stage3_54[27], stage3_54[28]},
      {stage3_55[44]},
      {stage3_56[12], stage3_56[13], stage3_56[14], stage3_56[15], stage3_56[16], stage3_56[17]},
      {stage4_58[2],stage4_57[9],stage4_56[9],stage4_55[16],stage4_54[23]}
   );
   gpc615_5 gpc8841 (
      {stage3_54[29], stage3_54[30], stage3_54[31], stage3_54[32], stage3_54[33]},
      {stage3_55[45]},
      {stage3_56[18], stage3_56[19], stage3_56[20], stage3_56[21], stage3_56[22], stage3_56[23]},
      {stage4_58[3],stage4_57[10],stage4_56[10],stage4_55[17],stage4_54[24]}
   );
   gpc615_5 gpc8842 (
      {stage3_54[34], stage3_54[35], stage3_54[36], stage3_54[37], stage3_54[38]},
      {stage3_55[46]},
      {stage3_56[24], stage3_56[25], stage3_56[26], stage3_56[27], stage3_56[28], stage3_56[29]},
      {stage4_58[4],stage4_57[11],stage4_56[11],stage4_55[18],stage4_54[25]}
   );
   gpc1163_5 gpc8843 (
      {stage3_57[0], stage3_57[1], stage3_57[2]},
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4], stage3_58[5]},
      {stage3_59[0]},
      {stage3_60[0]},
      {stage4_61[0],stage4_60[0],stage4_59[0],stage4_58[5],stage4_57[12]}
   );
   gpc1163_5 gpc8844 (
      {stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage3_58[6], stage3_58[7], stage3_58[8], stage3_58[9], stage3_58[10], stage3_58[11]},
      {stage3_59[1]},
      {stage3_60[1]},
      {stage4_61[1],stage4_60[1],stage4_59[1],stage4_58[6],stage4_57[13]}
   );
   gpc1163_5 gpc8845 (
      {stage3_57[6], stage3_57[7], stage3_57[8]},
      {stage3_58[12], stage3_58[13], stage3_58[14], stage3_58[15], stage3_58[16], stage3_58[17]},
      {stage3_59[2]},
      {stage3_60[2]},
      {stage4_61[2],stage4_60[2],stage4_59[2],stage4_58[7],stage4_57[14]}
   );
   gpc1163_5 gpc8846 (
      {stage3_57[9], stage3_57[10], stage3_57[11]},
      {stage3_58[18], stage3_58[19], stage3_58[20], stage3_58[21], stage3_58[22], stage3_58[23]},
      {stage3_59[3]},
      {stage3_60[3]},
      {stage4_61[3],stage4_60[3],stage4_59[3],stage4_58[8],stage4_57[15]}
   );
   gpc1163_5 gpc8847 (
      {stage3_57[12], stage3_57[13], stage3_57[14]},
      {stage3_58[24], stage3_58[25], stage3_58[26], stage3_58[27], stage3_58[28], stage3_58[29]},
      {stage3_59[4]},
      {stage3_60[4]},
      {stage4_61[4],stage4_60[4],stage4_59[4],stage4_58[9],stage4_57[16]}
   );
   gpc1163_5 gpc8848 (
      {stage3_57[15], stage3_57[16], stage3_57[17]},
      {stage3_58[30], stage3_58[31], stage3_58[32], stage3_58[33], stage3_58[34], stage3_58[35]},
      {stage3_59[5]},
      {stage3_60[5]},
      {stage4_61[5],stage4_60[5],stage4_59[5],stage4_58[10],stage4_57[17]}
   );
   gpc1163_5 gpc8849 (
      {stage3_57[18], stage3_57[19], stage3_57[20]},
      {stage3_58[36], stage3_58[37], stage3_58[38], stage3_58[39], stage3_58[40], stage3_58[41]},
      {stage3_59[6]},
      {stage3_60[6]},
      {stage4_61[6],stage4_60[6],stage4_59[6],stage4_58[11],stage4_57[18]}
   );
   gpc1163_5 gpc8850 (
      {stage3_57[21], stage3_57[22], stage3_57[23]},
      {stage3_58[42], stage3_58[43], stage3_58[44], stage3_58[45], stage3_58[46], stage3_58[47]},
      {stage3_59[7]},
      {stage3_60[7]},
      {stage4_61[7],stage4_60[7],stage4_59[7],stage4_58[12],stage4_57[19]}
   );
   gpc1163_5 gpc8851 (
      {stage3_57[24], stage3_57[25], stage3_57[26]},
      {stage3_58[48], stage3_58[49], stage3_58[50], stage3_58[51], stage3_58[52], stage3_58[53]},
      {stage3_59[8]},
      {stage3_60[8]},
      {stage4_61[8],stage4_60[8],stage4_59[8],stage4_58[13],stage4_57[20]}
   );
   gpc606_5 gpc8852 (
      {stage3_57[27], stage3_57[28], stage3_57[29], stage3_57[30], stage3_57[31], stage3_57[32]},
      {stage3_59[9], stage3_59[10], stage3_59[11], stage3_59[12], stage3_59[13], stage3_59[14]},
      {stage4_61[9],stage4_60[9],stage4_59[9],stage4_58[14],stage4_57[21]}
   );
   gpc606_5 gpc8853 (
      {stage3_57[33], stage3_57[34], stage3_57[35], stage3_57[36], stage3_57[37], stage3_57[38]},
      {stage3_59[15], stage3_59[16], stage3_59[17], stage3_59[18], stage3_59[19], stage3_59[20]},
      {stage4_61[10],stage4_60[10],stage4_59[10],stage4_58[15],stage4_57[22]}
   );
   gpc615_5 gpc8854 (
      {stage3_57[39], stage3_57[40], stage3_57[41], stage3_57[42], stage3_57[43]},
      {stage3_58[54]},
      {stage3_59[21], stage3_59[22], stage3_59[23], stage3_59[24], stage3_59[25], stage3_59[26]},
      {stage4_61[11],stage4_60[11],stage4_59[11],stage4_58[16],stage4_57[23]}
   );
   gpc615_5 gpc8855 (
      {stage3_57[44], stage3_57[45], stage3_57[46], stage3_57[47], stage3_57[48]},
      {stage3_58[55]},
      {stage3_59[27], stage3_59[28], stage3_59[29], stage3_59[30], stage3_59[31], stage3_59[32]},
      {stage4_61[12],stage4_60[12],stage4_59[12],stage4_58[17],stage4_57[24]}
   );
   gpc615_5 gpc8856 (
      {stage3_57[49], stage3_57[50], stage3_57[51], stage3_57[52], stage3_57[53]},
      {stage3_58[56]},
      {stage3_59[33], stage3_59[34], stage3_59[35], stage3_59[36], stage3_59[37], stage3_59[38]},
      {stage4_61[13],stage4_60[13],stage4_59[13],stage4_58[18],stage4_57[25]}
   );
   gpc615_5 gpc8857 (
      {stage3_59[39], stage3_59[40], stage3_59[41], stage3_59[42], stage3_59[43]},
      {stage3_60[9]},
      {stage3_61[0], stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5]},
      {stage4_63[0],stage4_62[0],stage4_61[14],stage4_60[14],stage4_59[14]}
   );
   gpc606_5 gpc8858 (
      {stage3_60[10], stage3_60[11], stage3_60[12], stage3_60[13], stage3_60[14], stage3_60[15]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], stage3_62[5]},
      {stage4_64[0],stage4_63[1],stage4_62[1],stage4_61[15],stage4_60[15]}
   );
   gpc606_5 gpc8859 (
      {stage3_60[16], stage3_60[17], stage3_60[18], stage3_60[19], stage3_60[20], stage3_60[21]},
      {stage3_62[6], stage3_62[7], stage3_62[8], stage3_62[9], stage3_62[10], stage3_62[11]},
      {stage4_64[1],stage4_63[2],stage4_62[2],stage4_61[16],stage4_60[16]}
   );
   gpc606_5 gpc8860 (
      {stage3_60[22], stage3_60[23], stage3_60[24], stage3_60[25], stage3_60[26], stage3_60[27]},
      {stage3_62[12], stage3_62[13], stage3_62[14], stage3_62[15], stage3_62[16], stage3_62[17]},
      {stage4_64[2],stage4_63[3],stage4_62[3],stage4_61[17],stage4_60[17]}
   );
   gpc606_5 gpc8861 (
      {stage3_60[28], stage3_60[29], stage3_60[30], stage3_60[31], stage3_60[32], stage3_60[33]},
      {stage3_62[18], stage3_62[19], stage3_62[20], stage3_62[21], stage3_62[22], stage3_62[23]},
      {stage4_64[3],stage4_63[4],stage4_62[4],stage4_61[18],stage4_60[18]}
   );
   gpc606_5 gpc8862 (
      {stage3_60[34], stage3_60[35], stage3_60[36], stage3_60[37], stage3_60[38], stage3_60[39]},
      {stage3_62[24], stage3_62[25], stage3_62[26], stage3_62[27], stage3_62[28], stage3_62[29]},
      {stage4_64[4],stage4_63[5],stage4_62[5],stage4_61[19],stage4_60[19]}
   );
   gpc606_5 gpc8863 (
      {stage3_61[6], stage3_61[7], stage3_61[8], stage3_61[9], stage3_61[10], stage3_61[11]},
      {stage3_63[0], stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5]},
      {stage4_65[0],stage4_64[5],stage4_63[6],stage4_62[6],stage4_61[20]}
   );
   gpc606_5 gpc8864 (
      {stage3_61[12], stage3_61[13], stage3_61[14], stage3_61[15], stage3_61[16], stage3_61[17]},
      {stage3_63[6], stage3_63[7], stage3_63[8], stage3_63[9], stage3_63[10], stage3_63[11]},
      {stage4_65[1],stage4_64[6],stage4_63[7],stage4_62[7],stage4_61[21]}
   );
   gpc606_5 gpc8865 (
      {stage3_61[18], stage3_61[19], stage3_61[20], stage3_61[21], stage3_61[22], stage3_61[23]},
      {stage3_63[12], stage3_63[13], stage3_63[14], stage3_63[15], stage3_63[16], stage3_63[17]},
      {stage4_65[2],stage4_64[7],stage4_63[8],stage4_62[8],stage4_61[22]}
   );
   gpc606_5 gpc8866 (
      {stage3_61[24], stage3_61[25], stage3_61[26], stage3_61[27], stage3_61[28], stage3_61[29]},
      {stage3_63[18], stage3_63[19], stage3_63[20], stage3_63[21], stage3_63[22], stage3_63[23]},
      {stage4_65[3],stage4_64[8],stage4_63[9],stage4_62[9],stage4_61[23]}
   );
   gpc606_5 gpc8867 (
      {stage3_61[30], stage3_61[31], stage3_61[32], stage3_61[33], stage3_61[34], stage3_61[35]},
      {stage3_63[24], stage3_63[25], stage3_63[26], stage3_63[27], stage3_63[28], stage3_63[29]},
      {stage4_65[4],stage4_64[9],stage4_63[10],stage4_62[10],stage4_61[24]}
   );
   gpc606_5 gpc8868 (
      {stage3_61[36], stage3_61[37], stage3_61[38], stage3_61[39], stage3_61[40], stage3_61[41]},
      {stage3_63[30], stage3_63[31], stage3_63[32], stage3_63[33], stage3_63[34], stage3_63[35]},
      {stage4_65[5],stage4_64[10],stage4_63[11],stage4_62[11],stage4_61[25]}
   );
   gpc606_5 gpc8869 (
      {stage3_61[42], stage3_61[43], stage3_61[44], stage3_61[45], stage3_61[46], stage3_61[47]},
      {stage3_63[36], stage3_63[37], stage3_63[38], stage3_63[39], stage3_63[40], stage3_63[41]},
      {stage4_65[6],stage4_64[11],stage4_63[12],stage4_62[12],stage4_61[26]}
   );
   gpc606_5 gpc8870 (
      {stage3_63[42], stage3_63[43], stage3_63[44], stage3_63[45], stage3_63[46], stage3_63[47]},
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5]},
      {stage4_67[0],stage4_66[0],stage4_65[7],stage4_64[12],stage4_63[13]}
   );
   gpc606_5 gpc8871 (
      {stage3_64[0], stage3_64[1], stage3_64[2], stage3_64[3], stage3_64[4], stage3_64[5]},
      {stage3_66[0], stage3_66[1], stage3_66[2], stage3_66[3], stage3_66[4], stage3_66[5]},
      {stage4_68[0],stage4_67[1],stage4_66[1],stage4_65[8],stage4_64[13]}
   );
   gpc606_5 gpc8872 (
      {stage3_64[6], stage3_64[7], stage3_64[8], stage3_64[9], stage3_64[10], stage3_64[11]},
      {stage3_66[6], stage3_66[7], stage3_66[8], stage3_66[9], stage3_66[10], stage3_66[11]},
      {stage4_68[1],stage4_67[2],stage4_66[2],stage4_65[9],stage4_64[14]}
   );
   gpc606_5 gpc8873 (
      {stage3_64[12], stage3_64[13], stage3_64[14], stage3_64[15], stage3_64[16], stage3_64[17]},
      {stage3_66[12], stage3_66[13], stage3_66[14], stage3_66[15], stage3_66[16], stage3_66[17]},
      {stage4_68[2],stage4_67[3],stage4_66[3],stage4_65[10],stage4_64[15]}
   );
   gpc606_5 gpc8874 (
      {stage3_64[18], stage3_64[19], stage3_64[20], stage3_64[21], stage3_64[22], stage3_64[23]},
      {stage3_66[18], stage3_66[19], stage3_66[20], stage3_66[21], stage3_66[22], stage3_66[23]},
      {stage4_68[3],stage4_67[4],stage4_66[4],stage4_65[11],stage4_64[16]}
   );
   gpc606_5 gpc8875 (
      {stage3_64[24], stage3_64[25], stage3_64[26], stage3_64[27], stage3_64[28], stage3_64[29]},
      {stage3_66[24], stage3_66[25], stage3_66[26], stage3_66[27], stage3_66[28], stage3_66[29]},
      {stage4_68[4],stage4_67[5],stage4_66[5],stage4_65[12],stage4_64[17]}
   );
   gpc606_5 gpc8876 (
      {stage3_64[30], stage3_64[31], stage3_64[32], stage3_64[33], stage3_64[34], stage3_64[35]},
      {stage3_66[30], stage3_66[31], stage3_66[32], stage3_66[33], stage3_66[34], stage3_66[35]},
      {stage4_68[5],stage4_67[6],stage4_66[6],stage4_65[13],stage4_64[18]}
   );
   gpc606_5 gpc8877 (
      {stage3_65[6], stage3_65[7], stage3_65[8], stage3_65[9], stage3_65[10], stage3_65[11]},
      {stage3_67[0], stage3_67[1], stage3_67[2], stage3_67[3], stage3_67[4], stage3_67[5]},
      {stage4_69[0],stage4_68[6],stage4_67[7],stage4_66[7],stage4_65[14]}
   );
   gpc606_5 gpc8878 (
      {stage3_65[12], stage3_65[13], stage3_65[14], stage3_65[15], stage3_65[16], stage3_65[17]},
      {stage3_67[6], stage3_67[7], stage3_67[8], stage3_67[9], stage3_67[10], stage3_67[11]},
      {stage4_69[1],stage4_68[7],stage4_67[8],stage4_66[8],stage4_65[15]}
   );
   gpc1_1 gpc8879 (
      {stage3_0[15]},
      {stage4_0[3]}
   );
   gpc1_1 gpc8880 (
      {stage3_0[16]},
      {stage4_0[4]}
   );
   gpc1_1 gpc8881 (
      {stage3_0[17]},
      {stage4_0[5]}
   );
   gpc1_1 gpc8882 (
      {stage3_0[18]},
      {stage4_0[6]}
   );
   gpc1_1 gpc8883 (
      {stage3_0[19]},
      {stage4_0[7]}
   );
   gpc1_1 gpc8884 (
      {stage3_0[20]},
      {stage4_0[8]}
   );
   gpc1_1 gpc8885 (
      {stage3_1[21]},
      {stage4_1[6]}
   );
   gpc1_1 gpc8886 (
      {stage3_2[42]},
      {stage4_2[10]}
   );
   gpc1_1 gpc8887 (
      {stage3_3[23]},
      {stage4_3[11]}
   );
   gpc1_1 gpc8888 (
      {stage3_3[24]},
      {stage4_3[12]}
   );
   gpc1_1 gpc8889 (
      {stage3_3[25]},
      {stage4_3[13]}
   );
   gpc1_1 gpc8890 (
      {stage3_3[26]},
      {stage4_3[14]}
   );
   gpc1_1 gpc8891 (
      {stage3_3[27]},
      {stage4_3[15]}
   );
   gpc1_1 gpc8892 (
      {stage3_3[28]},
      {stage4_3[16]}
   );
   gpc1_1 gpc8893 (
      {stage3_4[109]},
      {stage4_4[28]}
   );
   gpc1_1 gpc8894 (
      {stage3_4[110]},
      {stage4_4[29]}
   );
   gpc1_1 gpc8895 (
      {stage3_4[111]},
      {stage4_4[30]}
   );
   gpc1_1 gpc8896 (
      {stage3_5[42]},
      {stage4_5[25]}
   );
   gpc1_1 gpc8897 (
      {stage3_5[43]},
      {stage4_5[26]}
   );
   gpc1_1 gpc8898 (
      {stage3_5[44]},
      {stage4_5[27]}
   );
   gpc1_1 gpc8899 (
      {stage3_5[45]},
      {stage4_5[28]}
   );
   gpc1_1 gpc8900 (
      {stage3_5[46]},
      {stage4_5[29]}
   );
   gpc1_1 gpc8901 (
      {stage3_5[47]},
      {stage4_5[30]}
   );
   gpc1_1 gpc8902 (
      {stage3_5[48]},
      {stage4_5[31]}
   );
   gpc1_1 gpc8903 (
      {stage3_5[49]},
      {stage4_5[32]}
   );
   gpc1_1 gpc8904 (
      {stage3_5[50]},
      {stage4_5[33]}
   );
   gpc1_1 gpc8905 (
      {stage3_5[51]},
      {stage4_5[34]}
   );
   gpc1_1 gpc8906 (
      {stage3_5[52]},
      {stage4_5[35]}
   );
   gpc1_1 gpc8907 (
      {stage3_6[77]},
      {stage4_6[23]}
   );
   gpc1_1 gpc8908 (
      {stage3_7[37]},
      {stage4_7[25]}
   );
   gpc1_1 gpc8909 (
      {stage3_7[38]},
      {stage4_7[26]}
   );
   gpc1_1 gpc8910 (
      {stage3_7[39]},
      {stage4_7[27]}
   );
   gpc1_1 gpc8911 (
      {stage3_7[40]},
      {stage4_7[28]}
   );
   gpc1_1 gpc8912 (
      {stage3_7[41]},
      {stage4_7[29]}
   );
   gpc1_1 gpc8913 (
      {stage3_7[42]},
      {stage4_7[30]}
   );
   gpc1_1 gpc8914 (
      {stage3_7[43]},
      {stage4_7[31]}
   );
   gpc1_1 gpc8915 (
      {stage3_7[44]},
      {stage4_7[32]}
   );
   gpc1_1 gpc8916 (
      {stage3_7[45]},
      {stage4_7[33]}
   );
   gpc1_1 gpc8917 (
      {stage3_7[46]},
      {stage4_7[34]}
   );
   gpc1_1 gpc8918 (
      {stage3_7[47]},
      {stage4_7[35]}
   );
   gpc1_1 gpc8919 (
      {stage3_7[48]},
      {stage4_7[36]}
   );
   gpc1_1 gpc8920 (
      {stage3_7[49]},
      {stage4_7[37]}
   );
   gpc1_1 gpc8921 (
      {stage3_7[50]},
      {stage4_7[38]}
   );
   gpc1_1 gpc8922 (
      {stage3_10[84]},
      {stage4_10[26]}
   );
   gpc1_1 gpc8923 (
      {stage3_10[85]},
      {stage4_10[27]}
   );
   gpc1_1 gpc8924 (
      {stage3_10[86]},
      {stage4_10[28]}
   );
   gpc1_1 gpc8925 (
      {stage3_10[87]},
      {stage4_10[29]}
   );
   gpc1_1 gpc8926 (
      {stage3_10[88]},
      {stage4_10[30]}
   );
   gpc1_1 gpc8927 (
      {stage3_10[89]},
      {stage4_10[31]}
   );
   gpc1_1 gpc8928 (
      {stage3_10[90]},
      {stage4_10[32]}
   );
   gpc1_1 gpc8929 (
      {stage3_10[91]},
      {stage4_10[33]}
   );
   gpc1_1 gpc8930 (
      {stage3_10[92]},
      {stage4_10[34]}
   );
   gpc1_1 gpc8931 (
      {stage3_10[93]},
      {stage4_10[35]}
   );
   gpc1_1 gpc8932 (
      {stage3_10[94]},
      {stage4_10[36]}
   );
   gpc1_1 gpc8933 (
      {stage3_10[95]},
      {stage4_10[37]}
   );
   gpc1_1 gpc8934 (
      {stage3_10[96]},
      {stage4_10[38]}
   );
   gpc1_1 gpc8935 (
      {stage3_10[97]},
      {stage4_10[39]}
   );
   gpc1_1 gpc8936 (
      {stage3_10[98]},
      {stage4_10[40]}
   );
   gpc1_1 gpc8937 (
      {stage3_10[99]},
      {stage4_10[41]}
   );
   gpc1_1 gpc8938 (
      {stage3_12[67]},
      {stage4_12[23]}
   );
   gpc1_1 gpc8939 (
      {stage3_13[50]},
      {stage4_13[25]}
   );
   gpc1_1 gpc8940 (
      {stage3_13[51]},
      {stage4_13[26]}
   );
   gpc1_1 gpc8941 (
      {stage3_13[52]},
      {stage4_13[27]}
   );
   gpc1_1 gpc8942 (
      {stage3_13[53]},
      {stage4_13[28]}
   );
   gpc1_1 gpc8943 (
      {stage3_13[54]},
      {stage4_13[29]}
   );
   gpc1_1 gpc8944 (
      {stage3_13[55]},
      {stage4_13[30]}
   );
   gpc1_1 gpc8945 (
      {stage3_13[56]},
      {stage4_13[31]}
   );
   gpc1_1 gpc8946 (
      {stage3_14[30]},
      {stage4_14[28]}
   );
   gpc1_1 gpc8947 (
      {stage3_14[31]},
      {stage4_14[29]}
   );
   gpc1_1 gpc8948 (
      {stage3_15[47]},
      {stage4_15[14]}
   );
   gpc1_1 gpc8949 (
      {stage3_16[37]},
      {stage4_16[13]}
   );
   gpc1_1 gpc8950 (
      {stage3_16[38]},
      {stage4_16[14]}
   );
   gpc1_1 gpc8951 (
      {stage3_16[39]},
      {stage4_16[15]}
   );
   gpc1_1 gpc8952 (
      {stage3_16[40]},
      {stage4_16[16]}
   );
   gpc1_1 gpc8953 (
      {stage3_16[41]},
      {stage4_16[17]}
   );
   gpc1_1 gpc8954 (
      {stage3_16[42]},
      {stage4_16[18]}
   );
   gpc1_1 gpc8955 (
      {stage3_16[43]},
      {stage4_16[19]}
   );
   gpc1_1 gpc8956 (
      {stage3_16[44]},
      {stage4_16[20]}
   );
   gpc1_1 gpc8957 (
      {stage3_16[45]},
      {stage4_16[21]}
   );
   gpc1_1 gpc8958 (
      {stage3_16[46]},
      {stage4_16[22]}
   );
   gpc1_1 gpc8959 (
      {stage3_16[47]},
      {stage4_16[23]}
   );
   gpc1_1 gpc8960 (
      {stage3_16[48]},
      {stage4_16[24]}
   );
   gpc1_1 gpc8961 (
      {stage3_16[49]},
      {stage4_16[25]}
   );
   gpc1_1 gpc8962 (
      {stage3_16[50]},
      {stage4_16[26]}
   );
   gpc1_1 gpc8963 (
      {stage3_19[35]},
      {stage4_19[16]}
   );
   gpc1_1 gpc8964 (
      {stage3_19[36]},
      {stage4_19[17]}
   );
   gpc1_1 gpc8965 (
      {stage3_19[37]},
      {stage4_19[18]}
   );
   gpc1_1 gpc8966 (
      {stage3_19[38]},
      {stage4_19[19]}
   );
   gpc1_1 gpc8967 (
      {stage3_19[39]},
      {stage4_19[20]}
   );
   gpc1_1 gpc8968 (
      {stage3_19[40]},
      {stage4_19[21]}
   );
   gpc1_1 gpc8969 (
      {stage3_19[41]},
      {stage4_19[22]}
   );
   gpc1_1 gpc8970 (
      {stage3_19[42]},
      {stage4_19[23]}
   );
   gpc1_1 gpc8971 (
      {stage3_19[43]},
      {stage4_19[24]}
   );
   gpc1_1 gpc8972 (
      {stage3_19[44]},
      {stage4_19[25]}
   );
   gpc1_1 gpc8973 (
      {stage3_19[45]},
      {stage4_19[26]}
   );
   gpc1_1 gpc8974 (
      {stage3_19[46]},
      {stage4_19[27]}
   );
   gpc1_1 gpc8975 (
      {stage3_19[47]},
      {stage4_19[28]}
   );
   gpc1_1 gpc8976 (
      {stage3_20[73]},
      {stage4_20[24]}
   );
   gpc1_1 gpc8977 (
      {stage3_20[74]},
      {stage4_20[25]}
   );
   gpc1_1 gpc8978 (
      {stage3_20[75]},
      {stage4_20[26]}
   );
   gpc1_1 gpc8979 (
      {stage3_20[76]},
      {stage4_20[27]}
   );
   gpc1_1 gpc8980 (
      {stage3_20[77]},
      {stage4_20[28]}
   );
   gpc1_1 gpc8981 (
      {stage3_20[78]},
      {stage4_20[29]}
   );
   gpc1_1 gpc8982 (
      {stage3_20[79]},
      {stage4_20[30]}
   );
   gpc1_1 gpc8983 (
      {stage3_20[80]},
      {stage4_20[31]}
   );
   gpc1_1 gpc8984 (
      {stage3_20[81]},
      {stage4_20[32]}
   );
   gpc1_1 gpc8985 (
      {stage3_20[82]},
      {stage4_20[33]}
   );
   gpc1_1 gpc8986 (
      {stage3_21[30]},
      {stage4_21[28]}
   );
   gpc1_1 gpc8987 (
      {stage3_21[31]},
      {stage4_21[29]}
   );
   gpc1_1 gpc8988 (
      {stage3_21[32]},
      {stage4_21[30]}
   );
   gpc1_1 gpc8989 (
      {stage3_21[33]},
      {stage4_21[31]}
   );
   gpc1_1 gpc8990 (
      {stage3_21[34]},
      {stage4_21[32]}
   );
   gpc1_1 gpc8991 (
      {stage3_21[35]},
      {stage4_21[33]}
   );
   gpc1_1 gpc8992 (
      {stage3_21[36]},
      {stage4_21[34]}
   );
   gpc1_1 gpc8993 (
      {stage3_21[37]},
      {stage4_21[35]}
   );
   gpc1_1 gpc8994 (
      {stage3_21[38]},
      {stage4_21[36]}
   );
   gpc1_1 gpc8995 (
      {stage3_24[27]},
      {stage4_24[20]}
   );
   gpc1_1 gpc8996 (
      {stage3_24[28]},
      {stage4_24[21]}
   );
   gpc1_1 gpc8997 (
      {stage3_25[24]},
      {stage4_25[12]}
   );
   gpc1_1 gpc8998 (
      {stage3_25[25]},
      {stage4_25[13]}
   );
   gpc1_1 gpc8999 (
      {stage3_25[26]},
      {stage4_25[14]}
   );
   gpc1_1 gpc9000 (
      {stage3_25[27]},
      {stage4_25[15]}
   );
   gpc1_1 gpc9001 (
      {stage3_25[28]},
      {stage4_25[16]}
   );
   gpc1_1 gpc9002 (
      {stage3_25[29]},
      {stage4_25[17]}
   );
   gpc1_1 gpc9003 (
      {stage3_25[30]},
      {stage4_25[18]}
   );
   gpc1_1 gpc9004 (
      {stage3_25[31]},
      {stage4_25[19]}
   );
   gpc1_1 gpc9005 (
      {stage3_25[32]},
      {stage4_25[20]}
   );
   gpc1_1 gpc9006 (
      {stage3_27[38]},
      {stage4_27[16]}
   );
   gpc1_1 gpc9007 (
      {stage3_27[39]},
      {stage4_27[17]}
   );
   gpc1_1 gpc9008 (
      {stage3_27[40]},
      {stage4_27[18]}
   );
   gpc1_1 gpc9009 (
      {stage3_27[41]},
      {stage4_27[19]}
   );
   gpc1_1 gpc9010 (
      {stage3_27[42]},
      {stage4_27[20]}
   );
   gpc1_1 gpc9011 (
      {stage3_27[43]},
      {stage4_27[21]}
   );
   gpc1_1 gpc9012 (
      {stage3_27[44]},
      {stage4_27[22]}
   );
   gpc1_1 gpc9013 (
      {stage3_27[45]},
      {stage4_27[23]}
   );
   gpc1_1 gpc9014 (
      {stage3_27[46]},
      {stage4_27[24]}
   );
   gpc1_1 gpc9015 (
      {stage3_27[47]},
      {stage4_27[25]}
   );
   gpc1_1 gpc9016 (
      {stage3_27[48]},
      {stage4_27[26]}
   );
   gpc1_1 gpc9017 (
      {stage3_28[51]},
      {stage4_28[13]}
   );
   gpc1_1 gpc9018 (
      {stage3_28[52]},
      {stage4_28[14]}
   );
   gpc1_1 gpc9019 (
      {stage3_28[53]},
      {stage4_28[15]}
   );
   gpc1_1 gpc9020 (
      {stage3_28[54]},
      {stage4_28[16]}
   );
   gpc1_1 gpc9021 (
      {stage3_28[55]},
      {stage4_28[17]}
   );
   gpc1_1 gpc9022 (
      {stage3_28[56]},
      {stage4_28[18]}
   );
   gpc1_1 gpc9023 (
      {stage3_30[30]},
      {stage4_30[21]}
   );
   gpc1_1 gpc9024 (
      {stage3_30[31]},
      {stage4_30[22]}
   );
   gpc1_1 gpc9025 (
      {stage3_30[32]},
      {stage4_30[23]}
   );
   gpc1_1 gpc9026 (
      {stage3_30[33]},
      {stage4_30[24]}
   );
   gpc1_1 gpc9027 (
      {stage3_30[34]},
      {stage4_30[25]}
   );
   gpc1_1 gpc9028 (
      {stage3_30[35]},
      {stage4_30[26]}
   );
   gpc1_1 gpc9029 (
      {stage3_30[36]},
      {stage4_30[27]}
   );
   gpc1_1 gpc9030 (
      {stage3_30[37]},
      {stage4_30[28]}
   );
   gpc1_1 gpc9031 (
      {stage3_30[38]},
      {stage4_30[29]}
   );
   gpc1_1 gpc9032 (
      {stage3_30[39]},
      {stage4_30[30]}
   );
   gpc1_1 gpc9033 (
      {stage3_30[40]},
      {stage4_30[31]}
   );
   gpc1_1 gpc9034 (
      {stage3_30[41]},
      {stage4_30[32]}
   );
   gpc1_1 gpc9035 (
      {stage3_31[34]},
      {stage4_31[11]}
   );
   gpc1_1 gpc9036 (
      {stage3_31[35]},
      {stage4_31[12]}
   );
   gpc1_1 gpc9037 (
      {stage3_31[36]},
      {stage4_31[13]}
   );
   gpc1_1 gpc9038 (
      {stage3_31[37]},
      {stage4_31[14]}
   );
   gpc1_1 gpc9039 (
      {stage3_32[41]},
      {stage4_32[17]}
   );
   gpc1_1 gpc9040 (
      {stage3_32[42]},
      {stage4_32[18]}
   );
   gpc1_1 gpc9041 (
      {stage3_32[43]},
      {stage4_32[19]}
   );
   gpc1_1 gpc9042 (
      {stage3_32[44]},
      {stage4_32[20]}
   );
   gpc1_1 gpc9043 (
      {stage3_32[45]},
      {stage4_32[21]}
   );
   gpc1_1 gpc9044 (
      {stage3_32[46]},
      {stage4_32[22]}
   );
   gpc1_1 gpc9045 (
      {stage3_32[47]},
      {stage4_32[23]}
   );
   gpc1_1 gpc9046 (
      {stage3_32[48]},
      {stage4_32[24]}
   );
   gpc1_1 gpc9047 (
      {stage3_32[49]},
      {stage4_32[25]}
   );
   gpc1_1 gpc9048 (
      {stage3_32[50]},
      {stage4_32[26]}
   );
   gpc1_1 gpc9049 (
      {stage3_32[51]},
      {stage4_32[27]}
   );
   gpc1_1 gpc9050 (
      {stage3_32[52]},
      {stage4_32[28]}
   );
   gpc1_1 gpc9051 (
      {stage3_32[53]},
      {stage4_32[29]}
   );
   gpc1_1 gpc9052 (
      {stage3_33[37]},
      {stage4_33[20]}
   );
   gpc1_1 gpc9053 (
      {stage3_33[38]},
      {stage4_33[21]}
   );
   gpc1_1 gpc9054 (
      {stage3_33[39]},
      {stage4_33[22]}
   );
   gpc1_1 gpc9055 (
      {stage3_33[40]},
      {stage4_33[23]}
   );
   gpc1_1 gpc9056 (
      {stage3_33[41]},
      {stage4_33[24]}
   );
   gpc1_1 gpc9057 (
      {stage3_33[42]},
      {stage4_33[25]}
   );
   gpc1_1 gpc9058 (
      {stage3_33[43]},
      {stage4_33[26]}
   );
   gpc1_1 gpc9059 (
      {stage3_33[44]},
      {stage4_33[27]}
   );
   gpc1_1 gpc9060 (
      {stage3_33[45]},
      {stage4_33[28]}
   );
   gpc1_1 gpc9061 (
      {stage3_34[34]},
      {stage4_34[11]}
   );
   gpc1_1 gpc9062 (
      {stage3_34[35]},
      {stage4_34[12]}
   );
   gpc1_1 gpc9063 (
      {stage3_34[36]},
      {stage4_34[13]}
   );
   gpc1_1 gpc9064 (
      {stage3_34[37]},
      {stage4_34[14]}
   );
   gpc1_1 gpc9065 (
      {stage3_34[38]},
      {stage4_34[15]}
   );
   gpc1_1 gpc9066 (
      {stage3_34[39]},
      {stage4_34[16]}
   );
   gpc1_1 gpc9067 (
      {stage3_34[40]},
      {stage4_34[17]}
   );
   gpc1_1 gpc9068 (
      {stage3_34[41]},
      {stage4_34[18]}
   );
   gpc1_1 gpc9069 (
      {stage3_35[37]},
      {stage4_35[16]}
   );
   gpc1_1 gpc9070 (
      {stage3_35[38]},
      {stage4_35[17]}
   );
   gpc1_1 gpc9071 (
      {stage3_35[39]},
      {stage4_35[18]}
   );
   gpc1_1 gpc9072 (
      {stage3_35[40]},
      {stage4_35[19]}
   );
   gpc1_1 gpc9073 (
      {stage3_35[41]},
      {stage4_35[20]}
   );
   gpc1_1 gpc9074 (
      {stage3_35[42]},
      {stage4_35[21]}
   );
   gpc1_1 gpc9075 (
      {stage3_35[43]},
      {stage4_35[22]}
   );
   gpc1_1 gpc9076 (
      {stage3_35[44]},
      {stage4_35[23]}
   );
   gpc1_1 gpc9077 (
      {stage3_35[45]},
      {stage4_35[24]}
   );
   gpc1_1 gpc9078 (
      {stage3_35[46]},
      {stage4_35[25]}
   );
   gpc1_1 gpc9079 (
      {stage3_35[47]},
      {stage4_35[26]}
   );
   gpc1_1 gpc9080 (
      {stage3_35[48]},
      {stage4_35[27]}
   );
   gpc1_1 gpc9081 (
      {stage3_35[49]},
      {stage4_35[28]}
   );
   gpc1_1 gpc9082 (
      {stage3_35[50]},
      {stage4_35[29]}
   );
   gpc1_1 gpc9083 (
      {stage3_35[51]},
      {stage4_35[30]}
   );
   gpc1_1 gpc9084 (
      {stage3_35[52]},
      {stage4_35[31]}
   );
   gpc1_1 gpc9085 (
      {stage3_35[53]},
      {stage4_35[32]}
   );
   gpc1_1 gpc9086 (
      {stage3_35[54]},
      {stage4_35[33]}
   );
   gpc1_1 gpc9087 (
      {stage3_35[55]},
      {stage4_35[34]}
   );
   gpc1_1 gpc9088 (
      {stage3_35[56]},
      {stage4_35[35]}
   );
   gpc1_1 gpc9089 (
      {stage3_36[29]},
      {stage4_36[19]}
   );
   gpc1_1 gpc9090 (
      {stage3_36[30]},
      {stage4_36[20]}
   );
   gpc1_1 gpc9091 (
      {stage3_36[31]},
      {stage4_36[21]}
   );
   gpc1_1 gpc9092 (
      {stage3_36[32]},
      {stage4_36[22]}
   );
   gpc1_1 gpc9093 (
      {stage3_36[33]},
      {stage4_36[23]}
   );
   gpc1_1 gpc9094 (
      {stage3_36[34]},
      {stage4_36[24]}
   );
   gpc1_1 gpc9095 (
      {stage3_36[35]},
      {stage4_36[25]}
   );
   gpc1_1 gpc9096 (
      {stage3_36[36]},
      {stage4_36[26]}
   );
   gpc1_1 gpc9097 (
      {stage3_36[37]},
      {stage4_36[27]}
   );
   gpc1_1 gpc9098 (
      {stage3_36[38]},
      {stage4_36[28]}
   );
   gpc1_1 gpc9099 (
      {stage3_36[39]},
      {stage4_36[29]}
   );
   gpc1_1 gpc9100 (
      {stage3_36[40]},
      {stage4_36[30]}
   );
   gpc1_1 gpc9101 (
      {stage3_36[41]},
      {stage4_36[31]}
   );
   gpc1_1 gpc9102 (
      {stage3_36[42]},
      {stage4_36[32]}
   );
   gpc1_1 gpc9103 (
      {stage3_36[43]},
      {stage4_36[33]}
   );
   gpc1_1 gpc9104 (
      {stage3_36[44]},
      {stage4_36[34]}
   );
   gpc1_1 gpc9105 (
      {stage3_36[45]},
      {stage4_36[35]}
   );
   gpc1_1 gpc9106 (
      {stage3_37[48]},
      {stage4_37[13]}
   );
   gpc1_1 gpc9107 (
      {stage3_37[49]},
      {stage4_37[14]}
   );
   gpc1_1 gpc9108 (
      {stage3_37[50]},
      {stage4_37[15]}
   );
   gpc1_1 gpc9109 (
      {stage3_37[51]},
      {stage4_37[16]}
   );
   gpc1_1 gpc9110 (
      {stage3_37[52]},
      {stage4_37[17]}
   );
   gpc1_1 gpc9111 (
      {stage3_38[59]},
      {stage4_38[19]}
   );
   gpc1_1 gpc9112 (
      {stage3_40[43]},
      {stage4_40[19]}
   );
   gpc1_1 gpc9113 (
      {stage3_40[44]},
      {stage4_40[20]}
   );
   gpc1_1 gpc9114 (
      {stage3_40[45]},
      {stage4_40[21]}
   );
   gpc1_1 gpc9115 (
      {stage3_40[46]},
      {stage4_40[22]}
   );
   gpc1_1 gpc9116 (
      {stage3_40[47]},
      {stage4_40[23]}
   );
   gpc1_1 gpc9117 (
      {stage3_40[48]},
      {stage4_40[24]}
   );
   gpc1_1 gpc9118 (
      {stage3_40[49]},
      {stage4_40[25]}
   );
   gpc1_1 gpc9119 (
      {stage3_40[50]},
      {stage4_40[26]}
   );
   gpc1_1 gpc9120 (
      {stage3_40[51]},
      {stage4_40[27]}
   );
   gpc1_1 gpc9121 (
      {stage3_42[34]},
      {stage4_42[22]}
   );
   gpc1_1 gpc9122 (
      {stage3_42[35]},
      {stage4_42[23]}
   );
   gpc1_1 gpc9123 (
      {stage3_42[36]},
      {stage4_42[24]}
   );
   gpc1_1 gpc9124 (
      {stage3_42[37]},
      {stage4_42[25]}
   );
   gpc1_1 gpc9125 (
      {stage3_42[38]},
      {stage4_42[26]}
   );
   gpc1_1 gpc9126 (
      {stage3_42[39]},
      {stage4_42[27]}
   );
   gpc1_1 gpc9127 (
      {stage3_42[40]},
      {stage4_42[28]}
   );
   gpc1_1 gpc9128 (
      {stage3_42[41]},
      {stage4_42[29]}
   );
   gpc1_1 gpc9129 (
      {stage3_42[42]},
      {stage4_42[30]}
   );
   gpc1_1 gpc9130 (
      {stage3_42[43]},
      {stage4_42[31]}
   );
   gpc1_1 gpc9131 (
      {stage3_42[44]},
      {stage4_42[32]}
   );
   gpc1_1 gpc9132 (
      {stage3_42[45]},
      {stage4_42[33]}
   );
   gpc1_1 gpc9133 (
      {stage3_42[46]},
      {stage4_42[34]}
   );
   gpc1_1 gpc9134 (
      {stage3_42[47]},
      {stage4_42[35]}
   );
   gpc1_1 gpc9135 (
      {stage3_42[48]},
      {stage4_42[36]}
   );
   gpc1_1 gpc9136 (
      {stage3_42[49]},
      {stage4_42[37]}
   );
   gpc1_1 gpc9137 (
      {stage3_44[32]},
      {stage4_44[16]}
   );
   gpc1_1 gpc9138 (
      {stage3_44[33]},
      {stage4_44[17]}
   );
   gpc1_1 gpc9139 (
      {stage3_44[34]},
      {stage4_44[18]}
   );
   gpc1_1 gpc9140 (
      {stage3_44[35]},
      {stage4_44[19]}
   );
   gpc1_1 gpc9141 (
      {stage3_44[36]},
      {stage4_44[20]}
   );
   gpc1_1 gpc9142 (
      {stage3_44[37]},
      {stage4_44[21]}
   );
   gpc1_1 gpc9143 (
      {stage3_44[38]},
      {stage4_44[22]}
   );
   gpc1_1 gpc9144 (
      {stage3_44[39]},
      {stage4_44[23]}
   );
   gpc1_1 gpc9145 (
      {stage3_44[40]},
      {stage4_44[24]}
   );
   gpc1_1 gpc9146 (
      {stage3_45[34]},
      {stage4_45[19]}
   );
   gpc1_1 gpc9147 (
      {stage3_45[35]},
      {stage4_45[20]}
   );
   gpc1_1 gpc9148 (
      {stage3_45[36]},
      {stage4_45[21]}
   );
   gpc1_1 gpc9149 (
      {stage3_45[37]},
      {stage4_45[22]}
   );
   gpc1_1 gpc9150 (
      {stage3_45[38]},
      {stage4_45[23]}
   );
   gpc1_1 gpc9151 (
      {stage3_45[39]},
      {stage4_45[24]}
   );
   gpc1_1 gpc9152 (
      {stage3_45[40]},
      {stage4_45[25]}
   );
   gpc1_1 gpc9153 (
      {stage3_45[41]},
      {stage4_45[26]}
   );
   gpc1_1 gpc9154 (
      {stage3_45[42]},
      {stage4_45[27]}
   );
   gpc1_1 gpc9155 (
      {stage3_45[43]},
      {stage4_45[28]}
   );
   gpc1_1 gpc9156 (
      {stage3_46[57]},
      {stage4_46[16]}
   );
   gpc1_1 gpc9157 (
      {stage3_48[37]},
      {stage4_48[18]}
   );
   gpc1_1 gpc9158 (
      {stage3_48[38]},
      {stage4_48[19]}
   );
   gpc1_1 gpc9159 (
      {stage3_48[39]},
      {stage4_48[20]}
   );
   gpc1_1 gpc9160 (
      {stage3_48[40]},
      {stage4_48[21]}
   );
   gpc1_1 gpc9161 (
      {stage3_48[41]},
      {stage4_48[22]}
   );
   gpc1_1 gpc9162 (
      {stage3_51[50]},
      {stage4_51[23]}
   );
   gpc1_1 gpc9163 (
      {stage3_51[51]},
      {stage4_51[24]}
   );
   gpc1_1 gpc9164 (
      {stage3_51[52]},
      {stage4_51[25]}
   );
   gpc1_1 gpc9165 (
      {stage3_51[53]},
      {stage4_51[26]}
   );
   gpc1_1 gpc9166 (
      {stage3_51[54]},
      {stage4_51[27]}
   );
   gpc1_1 gpc9167 (
      {stage3_51[55]},
      {stage4_51[28]}
   );
   gpc1_1 gpc9168 (
      {stage3_51[56]},
      {stage4_51[29]}
   );
   gpc1_1 gpc9169 (
      {stage3_51[57]},
      {stage4_51[30]}
   );
   gpc1_1 gpc9170 (
      {stage3_51[58]},
      {stage4_51[31]}
   );
   gpc1_1 gpc9171 (
      {stage3_51[59]},
      {stage4_51[32]}
   );
   gpc1_1 gpc9172 (
      {stage3_51[60]},
      {stage4_51[33]}
   );
   gpc1_1 gpc9173 (
      {stage3_51[61]},
      {stage4_51[34]}
   );
   gpc1_1 gpc9174 (
      {stage3_51[62]},
      {stage4_51[35]}
   );
   gpc1_1 gpc9175 (
      {stage3_52[61]},
      {stage4_52[17]}
   );
   gpc1_1 gpc9176 (
      {stage3_52[62]},
      {stage4_52[18]}
   );
   gpc1_1 gpc9177 (
      {stage3_53[55]},
      {stage4_53[24]}
   );
   gpc1_1 gpc9178 (
      {stage3_53[56]},
      {stage4_53[25]}
   );
   gpc1_1 gpc9179 (
      {stage3_53[57]},
      {stage4_53[26]}
   );
   gpc1_1 gpc9180 (
      {stage3_53[58]},
      {stage4_53[27]}
   );
   gpc1_1 gpc9181 (
      {stage3_53[59]},
      {stage4_53[28]}
   );
   gpc1_1 gpc9182 (
      {stage3_53[60]},
      {stage4_53[29]}
   );
   gpc1_1 gpc9183 (
      {stage3_53[61]},
      {stage4_53[30]}
   );
   gpc1_1 gpc9184 (
      {stage3_53[62]},
      {stage4_53[31]}
   );
   gpc1_1 gpc9185 (
      {stage3_53[63]},
      {stage4_53[32]}
   );
   gpc1_1 gpc9186 (
      {stage3_53[64]},
      {stage4_53[33]}
   );
   gpc1_1 gpc9187 (
      {stage3_53[65]},
      {stage4_53[34]}
   );
   gpc1_1 gpc9188 (
      {stage3_53[66]},
      {stage4_53[35]}
   );
   gpc1_1 gpc9189 (
      {stage3_53[67]},
      {stage4_53[36]}
   );
   gpc1_1 gpc9190 (
      {stage3_53[68]},
      {stage4_53[37]}
   );
   gpc1_1 gpc9191 (
      {stage3_53[69]},
      {stage4_53[38]}
   );
   gpc1_1 gpc9192 (
      {stage3_53[70]},
      {stage4_53[39]}
   );
   gpc1_1 gpc9193 (
      {stage3_53[71]},
      {stage4_53[40]}
   );
   gpc1_1 gpc9194 (
      {stage3_53[72]},
      {stage4_53[41]}
   );
   gpc1_1 gpc9195 (
      {stage3_53[73]},
      {stage4_53[42]}
   );
   gpc1_1 gpc9196 (
      {stage3_53[74]},
      {stage4_53[43]}
   );
   gpc1_1 gpc9197 (
      {stage3_55[47]},
      {stage4_55[19]}
   );
   gpc1_1 gpc9198 (
      {stage3_55[48]},
      {stage4_55[20]}
   );
   gpc1_1 gpc9199 (
      {stage3_55[49]},
      {stage4_55[21]}
   );
   gpc1_1 gpc9200 (
      {stage3_55[50]},
      {stage4_55[22]}
   );
   gpc1_1 gpc9201 (
      {stage3_55[51]},
      {stage4_55[23]}
   );
   gpc1_1 gpc9202 (
      {stage3_55[52]},
      {stage4_55[24]}
   );
   gpc1_1 gpc9203 (
      {stage3_55[53]},
      {stage4_55[25]}
   );
   gpc1_1 gpc9204 (
      {stage3_55[54]},
      {stage4_55[26]}
   );
   gpc1_1 gpc9205 (
      {stage3_55[55]},
      {stage4_55[27]}
   );
   gpc1_1 gpc9206 (
      {stage3_55[56]},
      {stage4_55[28]}
   );
   gpc1_1 gpc9207 (
      {stage3_55[57]},
      {stage4_55[29]}
   );
   gpc1_1 gpc9208 (
      {stage3_55[58]},
      {stage4_55[30]}
   );
   gpc1_1 gpc9209 (
      {stage3_55[59]},
      {stage4_55[31]}
   );
   gpc1_1 gpc9210 (
      {stage3_55[60]},
      {stage4_55[32]}
   );
   gpc1_1 gpc9211 (
      {stage3_55[61]},
      {stage4_55[33]}
   );
   gpc1_1 gpc9212 (
      {stage3_55[62]},
      {stage4_55[34]}
   );
   gpc1_1 gpc9213 (
      {stage3_55[63]},
      {stage4_55[35]}
   );
   gpc1_1 gpc9214 (
      {stage3_55[64]},
      {stage4_55[36]}
   );
   gpc1_1 gpc9215 (
      {stage3_55[65]},
      {stage4_55[37]}
   );
   gpc1_1 gpc9216 (
      {stage3_55[66]},
      {stage4_55[38]}
   );
   gpc1_1 gpc9217 (
      {stage3_56[30]},
      {stage4_56[12]}
   );
   gpc1_1 gpc9218 (
      {stage3_56[31]},
      {stage4_56[13]}
   );
   gpc1_1 gpc9219 (
      {stage3_58[57]},
      {stage4_58[19]}
   );
   gpc1_1 gpc9220 (
      {stage3_58[58]},
      {stage4_58[20]}
   );
   gpc1_1 gpc9221 (
      {stage3_58[59]},
      {stage4_58[21]}
   );
   gpc1_1 gpc9222 (
      {stage3_58[60]},
      {stage4_58[22]}
   );
   gpc1_1 gpc9223 (
      {stage3_58[61]},
      {stage4_58[23]}
   );
   gpc1_1 gpc9224 (
      {stage3_59[44]},
      {stage4_59[15]}
   );
   gpc1_1 gpc9225 (
      {stage3_59[45]},
      {stage4_59[16]}
   );
   gpc1_1 gpc9226 (
      {stage3_59[46]},
      {stage4_59[17]}
   );
   gpc1_1 gpc9227 (
      {stage3_59[47]},
      {stage4_59[18]}
   );
   gpc1_1 gpc9228 (
      {stage3_59[48]},
      {stage4_59[19]}
   );
   gpc1_1 gpc9229 (
      {stage3_59[49]},
      {stage4_59[20]}
   );
   gpc1_1 gpc9230 (
      {stage3_60[40]},
      {stage4_60[20]}
   );
   gpc1_1 gpc9231 (
      {stage3_60[41]},
      {stage4_60[21]}
   );
   gpc1_1 gpc9232 (
      {stage3_61[48]},
      {stage4_61[27]}
   );
   gpc1_1 gpc9233 (
      {stage3_61[49]},
      {stage4_61[28]}
   );
   gpc1_1 gpc9234 (
      {stage3_61[50]},
      {stage4_61[29]}
   );
   gpc1_1 gpc9235 (
      {stage3_61[51]},
      {stage4_61[30]}
   );
   gpc1_1 gpc9236 (
      {stage3_61[52]},
      {stage4_61[31]}
   );
   gpc1_1 gpc9237 (
      {stage3_62[30]},
      {stage4_62[13]}
   );
   gpc1_1 gpc9238 (
      {stage3_62[31]},
      {stage4_62[14]}
   );
   gpc1_1 gpc9239 (
      {stage3_62[32]},
      {stage4_62[15]}
   );
   gpc1_1 gpc9240 (
      {stage3_62[33]},
      {stage4_62[16]}
   );
   gpc1_1 gpc9241 (
      {stage3_64[36]},
      {stage4_64[19]}
   );
   gpc1_1 gpc9242 (
      {stage3_64[37]},
      {stage4_64[20]}
   );
   gpc1_1 gpc9243 (
      {stage3_64[38]},
      {stage4_64[21]}
   );
   gpc1_1 gpc9244 (
      {stage3_64[39]},
      {stage4_64[22]}
   );
   gpc1_1 gpc9245 (
      {stage3_64[40]},
      {stage4_64[23]}
   );
   gpc1_1 gpc9246 (
      {stage3_64[41]},
      {stage4_64[24]}
   );
   gpc1_1 gpc9247 (
      {stage3_64[42]},
      {stage4_64[25]}
   );
   gpc1_1 gpc9248 (
      {stage3_64[43]},
      {stage4_64[26]}
   );
   gpc1_1 gpc9249 (
      {stage3_64[44]},
      {stage4_64[27]}
   );
   gpc1_1 gpc9250 (
      {stage3_64[45]},
      {stage4_64[28]}
   );
   gpc1_1 gpc9251 (
      {stage3_64[46]},
      {stage4_64[29]}
   );
   gpc1_1 gpc9252 (
      {stage3_64[47]},
      {stage4_64[30]}
   );
   gpc1_1 gpc9253 (
      {stage3_64[48]},
      {stage4_64[31]}
   );
   gpc1_1 gpc9254 (
      {stage3_64[49]},
      {stage4_64[32]}
   );
   gpc1_1 gpc9255 (
      {stage3_64[50]},
      {stage4_64[33]}
   );
   gpc1_1 gpc9256 (
      {stage3_65[18]},
      {stage4_65[16]}
   );
   gpc1_1 gpc9257 (
      {stage3_65[19]},
      {stage4_65[17]}
   );
   gpc1_1 gpc9258 (
      {stage3_65[20]},
      {stage4_65[18]}
   );
   gpc1_1 gpc9259 (
      {stage3_65[21]},
      {stage4_65[19]}
   );
   gpc1_1 gpc9260 (
      {stage3_65[22]},
      {stage4_65[20]}
   );
   gpc1_1 gpc9261 (
      {stage3_65[23]},
      {stage4_65[21]}
   );
   gpc1_1 gpc9262 (
      {stage3_65[24]},
      {stage4_65[22]}
   );
   gpc1_1 gpc9263 (
      {stage3_65[25]},
      {stage4_65[23]}
   );
   gpc1_1 gpc9264 (
      {stage3_65[26]},
      {stage4_65[24]}
   );
   gpc1_1 gpc9265 (
      {stage3_65[27]},
      {stage4_65[25]}
   );
   gpc1_1 gpc9266 (
      {stage3_65[28]},
      {stage4_65[26]}
   );
   gpc1_1 gpc9267 (
      {stage3_65[29]},
      {stage4_65[27]}
   );
   gpc1_1 gpc9268 (
      {stage3_65[30]},
      {stage4_65[28]}
   );
   gpc1_1 gpc9269 (
      {stage3_65[31]},
      {stage4_65[29]}
   );
   gpc1_1 gpc9270 (
      {stage3_65[32]},
      {stage4_65[30]}
   );
   gpc1_1 gpc9271 (
      {stage3_65[33]},
      {stage4_65[31]}
   );
   gpc1_1 gpc9272 (
      {stage3_65[34]},
      {stage4_65[32]}
   );
   gpc1_1 gpc9273 (
      {stage3_65[35]},
      {stage4_65[33]}
   );
   gpc1_1 gpc9274 (
      {stage3_65[36]},
      {stage4_65[34]}
   );
   gpc1_1 gpc9275 (
      {stage3_65[37]},
      {stage4_65[35]}
   );
   gpc1_1 gpc9276 (
      {stage3_66[36]},
      {stage4_66[9]}
   );
   gpc1_1 gpc9277 (
      {stage3_66[37]},
      {stage4_66[10]}
   );
   gpc1_1 gpc9278 (
      {stage3_67[12]},
      {stage4_67[9]}
   );
   gpc1_1 gpc9279 (
      {stage3_67[13]},
      {stage4_67[10]}
   );
   gpc1_1 gpc9280 (
      {stage3_68[0]},
      {stage4_68[8]}
   );
   gpc1_1 gpc9281 (
      {stage3_68[1]},
      {stage4_68[9]}
   );
   gpc1_1 gpc9282 (
      {stage3_68[2]},
      {stage4_68[10]}
   );
   gpc1_1 gpc9283 (
      {stage3_68[3]},
      {stage4_68[11]}
   );
   gpc1_1 gpc9284 (
      {stage3_68[4]},
      {stage4_68[12]}
   );
   gpc1_1 gpc9285 (
      {stage3_68[5]},
      {stage4_68[13]}
   );
   gpc615_5 gpc9286 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4]},
      {stage4_1[0]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc606_5 gpc9287 (
      {stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5], stage4_1[6]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc1163_5 gpc9288 (
      {stage4_2[6], stage4_2[7], stage4_2[8]},
      {stage4_3[6], stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage4_4[0]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[1],stage5_4[2],stage5_3[2],stage5_2[2]}
   );
   gpc1163_5 gpc9289 (
      {stage4_4[1], stage4_4[2], stage4_4[3]},
      {stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6]},
      {stage4_6[0]},
      {stage4_7[0]},
      {stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[2],stage5_4[3]}
   );
   gpc606_5 gpc9290 (
      {stage4_4[4], stage4_4[5], stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9]},
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5], stage4_6[6]},
      {stage5_8[1],stage5_7[1],stage5_6[2],stage5_5[3],stage5_4[4]}
   );
   gpc606_5 gpc9291 (
      {stage4_4[10], stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15]},
      {stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11], stage4_6[12]},
      {stage5_8[2],stage5_7[2],stage5_6[3],stage5_5[4],stage5_4[5]}
   );
   gpc606_5 gpc9292 (
      {stage4_4[16], stage4_4[17], stage4_4[18], stage4_4[19], stage4_4[20], stage4_4[21]},
      {stage4_6[13], stage4_6[14], stage4_6[15], stage4_6[16], stage4_6[17], stage4_6[18]},
      {stage5_8[3],stage5_7[3],stage5_6[4],stage5_5[5],stage5_4[6]}
   );
   gpc606_5 gpc9293 (
      {stage4_4[22], stage4_4[23], stage4_4[24], stage4_4[25], stage4_4[26], stage4_4[27]},
      {stage4_6[19], stage4_6[20], stage4_6[21], stage4_6[22], stage4_6[23], 1'b0},
      {stage5_8[4],stage5_7[4],stage5_6[5],stage5_5[6],stage5_4[7]}
   );
   gpc606_5 gpc9294 (
      {stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11], stage4_5[12]},
      {stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5], stage4_7[6]},
      {stage5_9[0],stage5_8[5],stage5_7[5],stage5_6[6],stage5_5[7]}
   );
   gpc606_5 gpc9295 (
      {stage4_5[13], stage4_5[14], stage4_5[15], stage4_5[16], stage4_5[17], stage4_5[18]},
      {stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11], stage4_7[12]},
      {stage5_9[1],stage5_8[6],stage5_7[6],stage5_6[7],stage5_5[8]}
   );
   gpc606_5 gpc9296 (
      {stage4_5[19], stage4_5[20], stage4_5[21], stage4_5[22], stage4_5[23], stage4_5[24]},
      {stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16], stage4_7[17], stage4_7[18]},
      {stage5_9[2],stage5_8[7],stage5_7[7],stage5_6[8],stage5_5[9]}
   );
   gpc606_5 gpc9297 (
      {stage4_5[25], stage4_5[26], stage4_5[27], stage4_5[28], stage4_5[29], stage4_5[30]},
      {stage4_7[19], stage4_7[20], stage4_7[21], stage4_7[22], stage4_7[23], stage4_7[24]},
      {stage5_9[3],stage5_8[8],stage5_7[8],stage5_6[9],stage5_5[10]}
   );
   gpc207_4 gpc9298 (
      {stage4_7[25], stage4_7[26], stage4_7[27], stage4_7[28], stage4_7[29], stage4_7[30], stage4_7[31]},
      {stage4_9[0], stage4_9[1]},
      {stage5_10[0],stage5_9[4],stage5_8[9],stage5_7[9]}
   );
   gpc207_4 gpc9299 (
      {stage4_7[32], stage4_7[33], stage4_7[34], stage4_7[35], stage4_7[36], stage4_7[37], stage4_7[38]},
      {stage4_9[2], stage4_9[3]},
      {stage5_10[1],stage5_9[5],stage5_8[10],stage5_7[10]}
   );
   gpc135_4 gpc9300 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[4], stage4_9[5], stage4_9[6]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[2],stage5_9[6],stage5_8[11]}
   );
   gpc117_4 gpc9301 (
      {stage4_8[5], stage4_8[6], stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11]},
      {stage4_9[7]},
      {stage4_10[1]},
      {stage5_11[1],stage5_10[3],stage5_9[7],stage5_8[12]}
   );
   gpc606_5 gpc9302 (
      {stage4_8[12], stage4_8[13], stage4_8[14], stage4_8[15], stage4_8[16], stage4_8[17]},
      {stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage5_12[0],stage5_11[2],stage5_10[4],stage5_9[8],stage5_8[13]}
   );
   gpc606_5 gpc9303 (
      {stage4_8[18], stage4_8[19], stage4_8[20], stage4_8[21], stage4_8[22], stage4_8[23]},
      {stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11], stage4_10[12], stage4_10[13]},
      {stage5_12[1],stage5_11[3],stage5_10[5],stage5_9[9],stage5_8[14]}
   );
   gpc606_5 gpc9304 (
      {stage4_9[8], stage4_9[9], stage4_9[10], stage4_9[11], stage4_9[12], stage4_9[13]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[2],stage5_11[4],stage5_10[6],stage5_9[10]}
   );
   gpc2135_5 gpc9305 (
      {stage4_10[14], stage4_10[15], stage4_10[16], stage4_10[17], stage4_10[18]},
      {stage4_11[6], stage4_11[7], stage4_11[8]},
      {stage4_12[0]},
      {stage4_13[0], stage4_13[1]},
      {stage5_14[0],stage5_13[1],stage5_12[3],stage5_11[5],stage5_10[7]}
   );
   gpc606_5 gpc9306 (
      {stage4_10[19], stage4_10[20], stage4_10[21], stage4_10[22], stage4_10[23], stage4_10[24]},
      {stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6]},
      {stage5_14[1],stage5_13[2],stage5_12[4],stage5_11[6],stage5_10[8]}
   );
   gpc606_5 gpc9307 (
      {stage4_10[25], stage4_10[26], stage4_10[27], stage4_10[28], stage4_10[29], stage4_10[30]},
      {stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11], stage4_12[12]},
      {stage5_14[2],stage5_13[3],stage5_12[5],stage5_11[7],stage5_10[9]}
   );
   gpc615_5 gpc9308 (
      {stage4_11[9], stage4_11[10], stage4_11[11], stage4_11[12], stage4_11[13]},
      {stage4_12[13]},
      {stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6], stage4_13[7]},
      {stage5_15[0],stage5_14[3],stage5_13[4],stage5_12[6],stage5_11[8]}
   );
   gpc615_5 gpc9309 (
      {stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17], stage4_11[18]},
      {stage4_12[14]},
      {stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12], stage4_13[13]},
      {stage5_15[1],stage5_14[4],stage5_13[5],stage5_12[7],stage5_11[9]}
   );
   gpc615_5 gpc9310 (
      {stage4_11[19], stage4_11[20], stage4_11[21], stage4_11[22], stage4_11[23]},
      {stage4_12[15]},
      {stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18], stage4_13[19]},
      {stage5_15[2],stage5_14[5],stage5_13[6],stage5_12[8],stage5_11[10]}
   );
   gpc623_5 gpc9311 (
      {stage4_11[24], stage4_11[25], stage4_11[26]},
      {stage4_12[16], stage4_12[17]},
      {stage4_13[20], stage4_13[21], stage4_13[22], stage4_13[23], stage4_13[24], stage4_13[25]},
      {stage5_15[3],stage5_14[6],stage5_13[7],stage5_12[9],stage5_11[11]}
   );
   gpc606_5 gpc9312 (
      {stage4_12[18], stage4_12[19], stage4_12[20], stage4_12[21], stage4_12[22], stage4_12[23]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[4],stage5_14[7],stage5_13[8],stage5_12[10]}
   );
   gpc615_5 gpc9313 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[0]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[5],stage5_14[8]}
   );
   gpc615_5 gpc9314 (
      {stage4_14[11], stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15]},
      {stage4_15[1]},
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11]},
      {stage5_18[1],stage5_17[1],stage5_16[2],stage5_15[6],stage5_14[9]}
   );
   gpc615_5 gpc9315 (
      {stage4_14[16], stage4_14[17], stage4_14[18], stage4_14[19], stage4_14[20]},
      {stage4_15[2]},
      {stage4_16[12], stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17]},
      {stage5_18[2],stage5_17[2],stage5_16[3],stage5_15[7],stage5_14[10]}
   );
   gpc615_5 gpc9316 (
      {stage4_14[21], stage4_14[22], stage4_14[23], stage4_14[24], stage4_14[25]},
      {stage4_15[3]},
      {stage4_16[18], stage4_16[19], stage4_16[20], stage4_16[21], stage4_16[22], stage4_16[23]},
      {stage5_18[3],stage5_17[3],stage5_16[4],stage5_15[8],stage5_14[11]}
   );
   gpc615_5 gpc9317 (
      {stage4_15[4], stage4_15[5], stage4_15[6], stage4_15[7], stage4_15[8]},
      {stage4_16[24]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[4],stage5_17[4],stage5_16[5],stage5_15[9]}
   );
   gpc615_5 gpc9318 (
      {stage4_15[9], stage4_15[10], stage4_15[11], stage4_15[12], stage4_15[13]},
      {stage4_16[25]},
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage5_19[1],stage5_18[5],stage5_17[5],stage5_16[6],stage5_15[10]}
   );
   gpc615_5 gpc9319 (
      {stage4_15[14], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage4_16[26]},
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17]},
      {stage5_19[2],stage5_18[6],stage5_17[6],stage5_16[7],stage5_15[11]}
   );
   gpc615_5 gpc9320 (
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4]},
      {stage4_19[0]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[0],stage5_20[0],stage5_19[3],stage5_18[7]}
   );
   gpc615_5 gpc9321 (
      {stage4_18[5], stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9]},
      {stage4_19[1]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], stage4_20[11]},
      {stage5_22[1],stage5_21[1],stage5_20[1],stage5_19[4],stage5_18[8]}
   );
   gpc615_5 gpc9322 (
      {stage4_18[10], stage4_18[11], stage4_18[12], stage4_18[13], stage4_18[14]},
      {stage4_19[2]},
      {stage4_20[12], stage4_20[13], stage4_20[14], stage4_20[15], stage4_20[16], stage4_20[17]},
      {stage5_22[2],stage5_21[2],stage5_20[2],stage5_19[5],stage5_18[9]}
   );
   gpc615_5 gpc9323 (
      {stage4_18[15], stage4_18[16], stage4_18[17], stage4_18[18], stage4_18[19]},
      {stage4_19[3]},
      {stage4_20[18], stage4_20[19], stage4_20[20], stage4_20[21], stage4_20[22], stage4_20[23]},
      {stage5_22[3],stage5_21[3],stage5_20[3],stage5_19[6],stage5_18[10]}
   );
   gpc615_5 gpc9324 (
      {stage4_19[4], stage4_19[5], stage4_19[6], stage4_19[7], stage4_19[8]},
      {stage4_20[24]},
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5]},
      {stage5_23[0],stage5_22[4],stage5_21[4],stage5_20[4],stage5_19[7]}
   );
   gpc615_5 gpc9325 (
      {stage4_19[9], stage4_19[10], stage4_19[11], stage4_19[12], stage4_19[13]},
      {stage4_20[25]},
      {stage4_21[6], stage4_21[7], stage4_21[8], stage4_21[9], stage4_21[10], stage4_21[11]},
      {stage5_23[1],stage5_22[5],stage5_21[5],stage5_20[5],stage5_19[8]}
   );
   gpc615_5 gpc9326 (
      {stage4_19[14], stage4_19[15], stage4_19[16], stage4_19[17], stage4_19[18]},
      {stage4_20[26]},
      {stage4_21[12], stage4_21[13], stage4_21[14], stage4_21[15], stage4_21[16], stage4_21[17]},
      {stage5_23[2],stage5_22[6],stage5_21[6],stage5_20[6],stage5_19[9]}
   );
   gpc615_5 gpc9327 (
      {stage4_19[19], stage4_19[20], stage4_19[21], stage4_19[22], stage4_19[23]},
      {stage4_20[27]},
      {stage4_21[18], stage4_21[19], stage4_21[20], stage4_21[21], stage4_21[22], stage4_21[23]},
      {stage5_23[3],stage5_22[7],stage5_21[7],stage5_20[7],stage5_19[10]}
   );
   gpc606_5 gpc9328 (
      {stage4_21[24], stage4_21[25], stage4_21[26], stage4_21[27], stage4_21[28], stage4_21[29]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage5_25[0],stage5_24[0],stage5_23[4],stage5_22[8],stage5_21[8]}
   );
   gpc606_5 gpc9329 (
      {stage4_21[30], stage4_21[31], stage4_21[32], stage4_21[33], stage4_21[34], stage4_21[35]},
      {stage4_23[6], stage4_23[7], stage4_23[8], stage4_23[9], stage4_23[10], stage4_23[11]},
      {stage5_25[1],stage5_24[1],stage5_23[5],stage5_22[9],stage5_21[9]}
   );
   gpc1163_5 gpc9330 (
      {stage4_22[0], stage4_22[1], stage4_22[2]},
      {stage4_23[12], stage4_23[13], stage4_23[14], stage4_23[15], stage4_23[16], stage4_23[17]},
      {stage4_24[0]},
      {stage4_25[0]},
      {stage5_26[0],stage5_25[2],stage5_24[2],stage5_23[6],stage5_22[10]}
   );
   gpc615_5 gpc9331 (
      {stage4_22[3], stage4_22[4], stage4_22[5], stage4_22[6], stage4_22[7]},
      {stage4_23[18]},
      {stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5], stage4_24[6]},
      {stage5_26[1],stage5_25[3],stage5_24[3],stage5_23[7],stage5_22[11]}
   );
   gpc615_5 gpc9332 (
      {stage4_22[8], stage4_22[9], stage4_22[10], stage4_22[11], stage4_22[12]},
      {stage4_23[19]},
      {stage4_24[7], stage4_24[8], stage4_24[9], stage4_24[10], stage4_24[11], stage4_24[12]},
      {stage5_26[2],stage5_25[4],stage5_24[4],stage5_23[8],stage5_22[12]}
   );
   gpc615_5 gpc9333 (
      {stage4_22[13], stage4_22[14], stage4_22[15], stage4_22[16], stage4_22[17]},
      {stage4_23[20]},
      {stage4_24[13], stage4_24[14], stage4_24[15], stage4_24[16], stage4_24[17], stage4_24[18]},
      {stage5_26[3],stage5_25[5],stage5_24[5],stage5_23[9],stage5_22[13]}
   );
   gpc606_5 gpc9334 (
      {stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5], stage4_25[6]},
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage5_29[0],stage5_28[0],stage5_27[0],stage5_26[4],stage5_25[6]}
   );
   gpc606_5 gpc9335 (
      {stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11], stage4_25[12]},
      {stage4_27[6], stage4_27[7], stage4_27[8], stage4_27[9], stage4_27[10], stage4_27[11]},
      {stage5_29[1],stage5_28[1],stage5_27[1],stage5_26[5],stage5_25[7]}
   );
   gpc606_5 gpc9336 (
      {stage4_25[13], stage4_25[14], stage4_25[15], stage4_25[16], stage4_25[17], stage4_25[18]},
      {stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16], stage4_27[17]},
      {stage5_29[2],stage5_28[2],stage5_27[2],stage5_26[6],stage5_25[8]}
   );
   gpc623_5 gpc9337 (
      {stage4_25[19], stage4_25[20], 1'b0},
      {stage4_26[0], stage4_26[1]},
      {stage4_27[18], stage4_27[19], stage4_27[20], stage4_27[21], stage4_27[22], stage4_27[23]},
      {stage5_29[3],stage5_28[3],stage5_27[3],stage5_26[7],stage5_25[9]}
   );
   gpc2135_5 gpc9338 (
      {stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5], stage4_26[6]},
      {stage4_27[24], stage4_27[25], stage4_27[26]},
      {stage4_28[0]},
      {stage4_29[0], stage4_29[1]},
      {stage5_30[0],stage5_29[4],stage5_28[4],stage5_27[4],stage5_26[8]}
   );
   gpc117_4 gpc9339 (
      {stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10], stage4_26[11], stage4_26[12], stage4_26[13]},
      {1'b0},
      {stage4_28[1]},
      {stage5_29[5],stage5_28[5],stage5_27[5],stage5_26[9]}
   );
   gpc606_5 gpc9340 (
      {stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5], stage4_28[6], stage4_28[7]},
      {stage4_30[0], stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5]},
      {stage5_32[0],stage5_31[0],stage5_30[1],stage5_29[6],stage5_28[6]}
   );
   gpc615_5 gpc9341 (
      {stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11], stage4_28[12]},
      {stage4_29[2]},
      {stage4_30[6], stage4_30[7], stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11]},
      {stage5_32[1],stage5_31[1],stage5_30[2],stage5_29[7],stage5_28[7]}
   );
   gpc615_5 gpc9342 (
      {stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16], stage4_28[17]},
      {stage4_29[3]},
      {stage4_30[12], stage4_30[13], stage4_30[14], stage4_30[15], stage4_30[16], stage4_30[17]},
      {stage5_32[2],stage5_31[2],stage5_30[3],stage5_29[8],stage5_28[8]}
   );
   gpc117_4 gpc9343 (
      {stage4_29[4], stage4_29[5], stage4_29[6], stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10]},
      {stage4_30[18]},
      {stage4_31[0]},
      {stage5_32[3],stage5_31[3],stage5_30[4],stage5_29[9]}
   );
   gpc117_4 gpc9344 (
      {stage4_29[11], stage4_29[12], stage4_29[13], stage4_29[14], stage4_29[15], stage4_29[16], stage4_29[17]},
      {stage4_30[19]},
      {stage4_31[1]},
      {stage5_32[4],stage5_31[4],stage5_30[5],stage5_29[10]}
   );
   gpc615_5 gpc9345 (
      {stage4_30[20], stage4_30[21], stage4_30[22], stage4_30[23], stage4_30[24]},
      {stage4_31[2]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[0],stage5_32[5],stage5_31[5],stage5_30[6]}
   );
   gpc615_5 gpc9346 (
      {stage4_30[25], stage4_30[26], stage4_30[27], stage4_30[28], stage4_30[29]},
      {stage4_31[3]},
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11]},
      {stage5_34[1],stage5_33[1],stage5_32[6],stage5_31[6],stage5_30[7]}
   );
   gpc615_5 gpc9347 (
      {stage4_30[30], stage4_30[31], stage4_30[32], 1'b0, 1'b0},
      {stage4_31[4]},
      {stage4_32[12], stage4_32[13], stage4_32[14], stage4_32[15], stage4_32[16], stage4_32[17]},
      {stage5_34[2],stage5_33[2],stage5_32[7],stage5_31[7],stage5_30[8]}
   );
   gpc615_5 gpc9348 (
      {stage4_31[5], stage4_31[6], stage4_31[7], stage4_31[8], stage4_31[9]},
      {stage4_32[18]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[3],stage5_33[3],stage5_32[8],stage5_31[8]}
   );
   gpc615_5 gpc9349 (
      {stage4_31[10], stage4_31[11], stage4_31[12], stage4_31[13], stage4_31[14]},
      {stage4_32[19]},
      {stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage5_35[1],stage5_34[4],stage5_33[4],stage5_32[9],stage5_31[9]}
   );
   gpc606_5 gpc9350 (
      {stage4_33[12], stage4_33[13], stage4_33[14], stage4_33[15], stage4_33[16], stage4_33[17]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[0],stage5_35[2],stage5_34[5],stage5_33[5]}
   );
   gpc606_5 gpc9351 (
      {stage4_33[18], stage4_33[19], stage4_33[20], stage4_33[21], stage4_33[22], stage4_33[23]},
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10], stage4_35[11]},
      {stage5_37[1],stage5_36[1],stage5_35[3],stage5_34[6],stage5_33[6]}
   );
   gpc135_4 gpc9352 (
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4]},
      {stage4_35[12], stage4_35[13], stage4_35[14]},
      {stage4_36[0]},
      {stage5_37[2],stage5_36[2],stage5_35[4],stage5_34[7]}
   );
   gpc615_5 gpc9353 (
      {stage4_34[5], stage4_34[6], stage4_34[7], stage4_34[8], stage4_34[9]},
      {stage4_35[15]},
      {stage4_36[1], stage4_36[2], stage4_36[3], stage4_36[4], stage4_36[5], stage4_36[6]},
      {stage5_38[0],stage5_37[3],stage5_36[3],stage5_35[5],stage5_34[8]}
   );
   gpc615_5 gpc9354 (
      {stage4_34[10], stage4_34[11], stage4_34[12], stage4_34[13], stage4_34[14]},
      {stage4_35[16]},
      {stage4_36[7], stage4_36[8], stage4_36[9], stage4_36[10], stage4_36[11], stage4_36[12]},
      {stage5_38[1],stage5_37[4],stage5_36[4],stage5_35[6],stage5_34[9]}
   );
   gpc615_5 gpc9355 (
      {stage4_35[17], stage4_35[18], stage4_35[19], stage4_35[20], stage4_35[21]},
      {stage4_36[13]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage5_39[0],stage5_38[2],stage5_37[5],stage5_36[5],stage5_35[7]}
   );
   gpc615_5 gpc9356 (
      {stage4_35[22], stage4_35[23], stage4_35[24], stage4_35[25], stage4_35[26]},
      {stage4_36[14]},
      {stage4_37[6], stage4_37[7], stage4_37[8], stage4_37[9], stage4_37[10], stage4_37[11]},
      {stage5_39[1],stage5_38[3],stage5_37[6],stage5_36[6],stage5_35[8]}
   );
   gpc615_5 gpc9357 (
      {stage4_35[27], stage4_35[28], stage4_35[29], stage4_35[30], stage4_35[31]},
      {stage4_36[15]},
      {stage4_37[12], stage4_37[13], stage4_37[14], stage4_37[15], stage4_37[16], stage4_37[17]},
      {stage5_39[2],stage5_38[4],stage5_37[7],stage5_36[7],stage5_35[9]}
   );
   gpc606_5 gpc9358 (
      {stage4_36[16], stage4_36[17], stage4_36[18], stage4_36[19], stage4_36[20], stage4_36[21]},
      {stage4_38[0], stage4_38[1], stage4_38[2], stage4_38[3], stage4_38[4], stage4_38[5]},
      {stage5_40[0],stage5_39[3],stage5_38[5],stage5_37[8],stage5_36[8]}
   );
   gpc606_5 gpc9359 (
      {stage4_36[22], stage4_36[23], stage4_36[24], stage4_36[25], stage4_36[26], stage4_36[27]},
      {stage4_38[6], stage4_38[7], stage4_38[8], stage4_38[9], stage4_38[10], stage4_38[11]},
      {stage5_40[1],stage5_39[4],stage5_38[6],stage5_37[9],stage5_36[9]}
   );
   gpc606_5 gpc9360 (
      {stage4_36[28], stage4_36[29], stage4_36[30], stage4_36[31], stage4_36[32], stage4_36[33]},
      {stage4_38[12], stage4_38[13], stage4_38[14], stage4_38[15], stage4_38[16], stage4_38[17]},
      {stage5_40[2],stage5_39[5],stage5_38[7],stage5_37[10],stage5_36[10]}
   );
   gpc117_4 gpc9361 (
      {stage4_39[0], stage4_39[1], stage4_39[2], stage4_39[3], stage4_39[4], stage4_39[5], stage4_39[6]},
      {stage4_40[0]},
      {stage4_41[0]},
      {stage5_42[0],stage5_41[0],stage5_40[3],stage5_39[6]}
   );
   gpc117_4 gpc9362 (
      {stage4_39[7], stage4_39[8], stage4_39[9], stage4_39[10], stage4_39[11], stage4_39[12], stage4_39[13]},
      {stage4_40[1]},
      {stage4_41[1]},
      {stage5_42[1],stage5_41[1],stage5_40[4],stage5_39[7]}
   );
   gpc615_5 gpc9363 (
      {stage4_39[14], stage4_39[15], stage4_39[16], stage4_39[17], stage4_39[18]},
      {stage4_40[2]},
      {stage4_41[2], stage4_41[3], stage4_41[4], stage4_41[5], stage4_41[6], stage4_41[7]},
      {stage5_43[0],stage5_42[2],stage5_41[2],stage5_40[5],stage5_39[8]}
   );
   gpc615_5 gpc9364 (
      {stage4_39[19], stage4_39[20], stage4_39[21], stage4_39[22], stage4_39[23]},
      {stage4_40[3]},
      {stage4_41[8], stage4_41[9], stage4_41[10], stage4_41[11], stage4_41[12], stage4_41[13]},
      {stage5_43[1],stage5_42[3],stage5_41[3],stage5_40[6],stage5_39[9]}
   );
   gpc606_5 gpc9365 (
      {stage4_40[4], stage4_40[5], stage4_40[6], stage4_40[7], stage4_40[8], stage4_40[9]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3], stage4_42[4], stage4_42[5]},
      {stage5_44[0],stage5_43[2],stage5_42[4],stage5_41[4],stage5_40[7]}
   );
   gpc606_5 gpc9366 (
      {stage4_40[10], stage4_40[11], stage4_40[12], stage4_40[13], stage4_40[14], stage4_40[15]},
      {stage4_42[6], stage4_42[7], stage4_42[8], stage4_42[9], stage4_42[10], stage4_42[11]},
      {stage5_44[1],stage5_43[3],stage5_42[5],stage5_41[5],stage5_40[8]}
   );
   gpc606_5 gpc9367 (
      {stage4_40[16], stage4_40[17], stage4_40[18], stage4_40[19], stage4_40[20], stage4_40[21]},
      {stage4_42[12], stage4_42[13], stage4_42[14], stage4_42[15], stage4_42[16], stage4_42[17]},
      {stage5_44[2],stage5_43[4],stage5_42[6],stage5_41[6],stage5_40[9]}
   );
   gpc606_5 gpc9368 (
      {stage4_40[22], stage4_40[23], stage4_40[24], stage4_40[25], stage4_40[26], stage4_40[27]},
      {stage4_42[18], stage4_42[19], stage4_42[20], stage4_42[21], stage4_42[22], stage4_42[23]},
      {stage5_44[3],stage5_43[5],stage5_42[7],stage5_41[7],stage5_40[10]}
   );
   gpc606_5 gpc9369 (
      {stage4_41[14], stage4_41[15], stage4_41[16], stage4_41[17], stage4_41[18], stage4_41[19]},
      {stage4_43[0], stage4_43[1], stage4_43[2], stage4_43[3], stage4_43[4], stage4_43[5]},
      {stage5_45[0],stage5_44[4],stage5_43[6],stage5_42[8],stage5_41[8]}
   );
   gpc615_5 gpc9370 (
      {stage4_42[24], stage4_42[25], stage4_42[26], stage4_42[27], stage4_42[28]},
      {stage4_43[6]},
      {stage4_44[0], stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage5_46[0],stage5_45[1],stage5_44[5],stage5_43[7],stage5_42[9]}
   );
   gpc615_5 gpc9371 (
      {stage4_43[7], stage4_43[8], stage4_43[9], stage4_43[10], stage4_43[11]},
      {stage4_44[6]},
      {stage4_45[0], stage4_45[1], stage4_45[2], stage4_45[3], stage4_45[4], stage4_45[5]},
      {stage5_47[0],stage5_46[1],stage5_45[2],stage5_44[6],stage5_43[8]}
   );
   gpc135_4 gpc9372 (
      {stage4_44[7], stage4_44[8], stage4_44[9], stage4_44[10], stage4_44[11]},
      {stage4_45[6], stage4_45[7], stage4_45[8]},
      {stage4_46[0]},
      {stage5_47[1],stage5_46[2],stage5_45[3],stage5_44[7]}
   );
   gpc135_4 gpc9373 (
      {stage4_44[12], stage4_44[13], stage4_44[14], stage4_44[15], stage4_44[16]},
      {stage4_45[9], stage4_45[10], stage4_45[11]},
      {stage4_46[1]},
      {stage5_47[2],stage5_46[3],stage5_45[4],stage5_44[8]}
   );
   gpc135_4 gpc9374 (
      {stage4_44[17], stage4_44[18], stage4_44[19], stage4_44[20], stage4_44[21]},
      {stage4_45[12], stage4_45[13], stage4_45[14]},
      {stage4_46[2]},
      {stage5_47[3],stage5_46[4],stage5_45[5],stage5_44[9]}
   );
   gpc606_5 gpc9375 (
      {stage4_45[15], stage4_45[16], stage4_45[17], stage4_45[18], stage4_45[19], stage4_45[20]},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3], stage4_47[4], stage4_47[5]},
      {stage5_49[0],stage5_48[0],stage5_47[4],stage5_46[5],stage5_45[6]}
   );
   gpc615_5 gpc9376 (
      {stage4_46[3], stage4_46[4], stage4_46[5], stage4_46[6], stage4_46[7]},
      {stage4_47[6]},
      {stage4_48[0], stage4_48[1], stage4_48[2], stage4_48[3], stage4_48[4], stage4_48[5]},
      {stage5_50[0],stage5_49[1],stage5_48[1],stage5_47[5],stage5_46[6]}
   );
   gpc615_5 gpc9377 (
      {stage4_46[8], stage4_46[9], stage4_46[10], stage4_46[11], stage4_46[12]},
      {stage4_47[7]},
      {stage4_48[6], stage4_48[7], stage4_48[8], stage4_48[9], stage4_48[10], stage4_48[11]},
      {stage5_50[1],stage5_49[2],stage5_48[2],stage5_47[6],stage5_46[7]}
   );
   gpc615_5 gpc9378 (
      {stage4_47[8], stage4_47[9], stage4_47[10], stage4_47[11], stage4_47[12]},
      {stage4_48[12]},
      {stage4_49[0], stage4_49[1], stage4_49[2], stage4_49[3], stage4_49[4], stage4_49[5]},
      {stage5_51[0],stage5_50[2],stage5_49[3],stage5_48[3],stage5_47[7]}
   );
   gpc615_5 gpc9379 (
      {stage4_47[13], stage4_47[14], stage4_47[15], stage4_47[16], stage4_47[17]},
      {stage4_48[13]},
      {stage4_49[6], stage4_49[7], stage4_49[8], stage4_49[9], stage4_49[10], stage4_49[11]},
      {stage5_51[1],stage5_50[3],stage5_49[4],stage5_48[4],stage5_47[8]}
   );
   gpc7_3 gpc9380 (
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3], stage4_50[4], stage4_50[5], stage4_50[6]},
      {stage5_52[0],stage5_51[2],stage5_50[4]}
   );
   gpc615_5 gpc9381 (
      {stage4_50[7], stage4_50[8], stage4_50[9], stage4_50[10], stage4_50[11]},
      {stage4_51[0]},
      {stage4_52[0], stage4_52[1], stage4_52[2], stage4_52[3], stage4_52[4], stage4_52[5]},
      {stage5_54[0],stage5_53[0],stage5_52[1],stage5_51[3],stage5_50[5]}
   );
   gpc615_5 gpc9382 (
      {stage4_50[12], stage4_50[13], stage4_50[14], stage4_50[15], stage4_50[16]},
      {stage4_51[1]},
      {stage4_52[6], stage4_52[7], stage4_52[8], stage4_52[9], stage4_52[10], stage4_52[11]},
      {stage5_54[1],stage5_53[1],stage5_52[2],stage5_51[4],stage5_50[6]}
   );
   gpc615_5 gpc9383 (
      {stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5], stage4_51[6]},
      {stage4_52[12]},
      {stage4_53[0], stage4_53[1], stage4_53[2], stage4_53[3], stage4_53[4], stage4_53[5]},
      {stage5_55[0],stage5_54[2],stage5_53[2],stage5_52[3],stage5_51[5]}
   );
   gpc615_5 gpc9384 (
      {stage4_51[7], stage4_51[8], stage4_51[9], stage4_51[10], stage4_51[11]},
      {stage4_52[13]},
      {stage4_53[6], stage4_53[7], stage4_53[8], stage4_53[9], stage4_53[10], stage4_53[11]},
      {stage5_55[1],stage5_54[3],stage5_53[3],stage5_52[4],stage5_51[6]}
   );
   gpc615_5 gpc9385 (
      {stage4_51[12], stage4_51[13], stage4_51[14], stage4_51[15], stage4_51[16]},
      {stage4_52[14]},
      {stage4_53[12], stage4_53[13], stage4_53[14], stage4_53[15], stage4_53[16], stage4_53[17]},
      {stage5_55[2],stage5_54[4],stage5_53[4],stage5_52[5],stage5_51[7]}
   );
   gpc615_5 gpc9386 (
      {stage4_51[17], stage4_51[18], stage4_51[19], stage4_51[20], stage4_51[21]},
      {stage4_52[15]},
      {stage4_53[18], stage4_53[19], stage4_53[20], stage4_53[21], stage4_53[22], stage4_53[23]},
      {stage5_55[3],stage5_54[5],stage5_53[5],stage5_52[6],stage5_51[8]}
   );
   gpc615_5 gpc9387 (
      {stage4_51[22], stage4_51[23], stage4_51[24], stage4_51[25], stage4_51[26]},
      {stage4_52[16]},
      {stage4_53[24], stage4_53[25], stage4_53[26], stage4_53[27], stage4_53[28], stage4_53[29]},
      {stage5_55[4],stage5_54[6],stage5_53[6],stage5_52[7],stage5_51[9]}
   );
   gpc615_5 gpc9388 (
      {stage4_53[30], stage4_53[31], stage4_53[32], stage4_53[33], stage4_53[34]},
      {stage4_54[0]},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5]},
      {stage5_57[0],stage5_56[0],stage5_55[5],stage5_54[7],stage5_53[7]}
   );
   gpc615_5 gpc9389 (
      {stage4_53[35], stage4_53[36], stage4_53[37], stage4_53[38], stage4_53[39]},
      {stage4_54[1]},
      {stage4_55[6], stage4_55[7], stage4_55[8], stage4_55[9], stage4_55[10], stage4_55[11]},
      {stage5_57[1],stage5_56[1],stage5_55[6],stage5_54[8],stage5_53[8]}
   );
   gpc2135_5 gpc9390 (
      {stage4_54[2], stage4_54[3], stage4_54[4], stage4_54[5], stage4_54[6]},
      {stage4_55[12], stage4_55[13], stage4_55[14]},
      {stage4_56[0]},
      {stage4_57[0], stage4_57[1]},
      {stage5_58[0],stage5_57[2],stage5_56[2],stage5_55[7],stage5_54[9]}
   );
   gpc2135_5 gpc9391 (
      {stage4_54[7], stage4_54[8], stage4_54[9], stage4_54[10], stage4_54[11]},
      {stage4_55[15], stage4_55[16], stage4_55[17]},
      {stage4_56[1]},
      {stage4_57[2], stage4_57[3]},
      {stage5_58[1],stage5_57[3],stage5_56[3],stage5_55[8],stage5_54[10]}
   );
   gpc2135_5 gpc9392 (
      {stage4_54[12], stage4_54[13], stage4_54[14], stage4_54[15], stage4_54[16]},
      {stage4_55[18], stage4_55[19], stage4_55[20]},
      {stage4_56[2]},
      {stage4_57[4], stage4_57[5]},
      {stage5_58[2],stage5_57[4],stage5_56[4],stage5_55[9],stage5_54[11]}
   );
   gpc2135_5 gpc9393 (
      {stage4_54[17], stage4_54[18], stage4_54[19], stage4_54[20], stage4_54[21]},
      {stage4_55[21], stage4_55[22], stage4_55[23]},
      {stage4_56[3]},
      {stage4_57[6], stage4_57[7]},
      {stage5_58[3],stage5_57[5],stage5_56[5],stage5_55[10],stage5_54[12]}
   );
   gpc615_5 gpc9394 (
      {stage4_55[24], stage4_55[25], stage4_55[26], stage4_55[27], stage4_55[28]},
      {stage4_56[4]},
      {stage4_57[8], stage4_57[9], stage4_57[10], stage4_57[11], stage4_57[12], stage4_57[13]},
      {stage5_59[0],stage5_58[4],stage5_57[6],stage5_56[6],stage5_55[11]}
   );
   gpc606_5 gpc9395 (
      {stage4_56[5], stage4_56[6], stage4_56[7], stage4_56[8], stage4_56[9], stage4_56[10]},
      {stage4_58[0], stage4_58[1], stage4_58[2], stage4_58[3], stage4_58[4], stage4_58[5]},
      {stage5_60[0],stage5_59[1],stage5_58[5],stage5_57[7],stage5_56[7]}
   );
   gpc623_5 gpc9396 (
      {stage4_56[11], stage4_56[12], stage4_56[13]},
      {stage4_57[14], stage4_57[15]},
      {stage4_58[6], stage4_58[7], stage4_58[8], stage4_58[9], stage4_58[10], stage4_58[11]},
      {stage5_60[1],stage5_59[2],stage5_58[6],stage5_57[8],stage5_56[8]}
   );
   gpc606_5 gpc9397 (
      {stage4_57[16], stage4_57[17], stage4_57[18], stage4_57[19], stage4_57[20], stage4_57[21]},
      {stage4_59[0], stage4_59[1], stage4_59[2], stage4_59[3], stage4_59[4], stage4_59[5]},
      {stage5_61[0],stage5_60[2],stage5_59[3],stage5_58[7],stage5_57[9]}
   );
   gpc615_5 gpc9398 (
      {stage4_58[12], stage4_58[13], stage4_58[14], stage4_58[15], stage4_58[16]},
      {stage4_59[6]},
      {stage4_60[0], stage4_60[1], stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5]},
      {stage5_62[0],stage5_61[1],stage5_60[3],stage5_59[4],stage5_58[8]}
   );
   gpc615_5 gpc9399 (
      {stage4_59[7], stage4_59[8], stage4_59[9], stage4_59[10], stage4_59[11]},
      {stage4_60[6]},
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage5_63[0],stage5_62[1],stage5_61[2],stage5_60[4],stage5_59[5]}
   );
   gpc615_5 gpc9400 (
      {stage4_59[12], stage4_59[13], stage4_59[14], stage4_59[15], stage4_59[16]},
      {stage4_60[7]},
      {stage4_61[6], stage4_61[7], stage4_61[8], stage4_61[9], stage4_61[10], stage4_61[11]},
      {stage5_63[1],stage5_62[2],stage5_61[3],stage5_60[5],stage5_59[6]}
   );
   gpc615_5 gpc9401 (
      {stage4_59[17], stage4_59[18], stage4_59[19], stage4_59[20], 1'b0},
      {stage4_60[8]},
      {stage4_61[12], stage4_61[13], stage4_61[14], stage4_61[15], stage4_61[16], stage4_61[17]},
      {stage5_63[2],stage5_62[3],stage5_61[4],stage5_60[6],stage5_59[7]}
   );
   gpc606_5 gpc9402 (
      {stage4_60[9], stage4_60[10], stage4_60[11], stage4_60[12], stage4_60[13], stage4_60[14]},
      {stage4_62[0], stage4_62[1], stage4_62[2], stage4_62[3], stage4_62[4], stage4_62[5]},
      {stage5_64[0],stage5_63[3],stage5_62[4],stage5_61[5],stage5_60[7]}
   );
   gpc615_5 gpc9403 (
      {stage4_61[18], stage4_61[19], stage4_61[20], stage4_61[21], stage4_61[22]},
      {stage4_62[6]},
      {stage4_63[0], stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4], stage4_63[5]},
      {stage5_65[0],stage5_64[1],stage5_63[4],stage5_62[5],stage5_61[6]}
   );
   gpc615_5 gpc9404 (
      {stage4_62[7], stage4_62[8], stage4_62[9], stage4_62[10], stage4_62[11]},
      {stage4_63[6]},
      {stage4_64[0], stage4_64[1], stage4_64[2], stage4_64[3], stage4_64[4], stage4_64[5]},
      {stage5_66[0],stage5_65[1],stage5_64[2],stage5_63[5],stage5_62[6]}
   );
   gpc615_5 gpc9405 (
      {stage4_63[7], stage4_63[8], stage4_63[9], stage4_63[10], stage4_63[11]},
      {stage4_64[6]},
      {stage4_65[0], stage4_65[1], stage4_65[2], stage4_65[3], stage4_65[4], stage4_65[5]},
      {stage5_67[0],stage5_66[1],stage5_65[2],stage5_64[3],stage5_63[6]}
   );
   gpc2135_5 gpc9406 (
      {stage4_64[7], stage4_64[8], stage4_64[9], stage4_64[10], stage4_64[11]},
      {stage4_65[6], stage4_65[7], stage4_65[8]},
      {stage4_66[0]},
      {stage4_67[0], stage4_67[1]},
      {stage5_68[0],stage5_67[1],stage5_66[2],stage5_65[3],stage5_64[4]}
   );
   gpc2135_5 gpc9407 (
      {stage4_64[12], stage4_64[13], stage4_64[14], stage4_64[15], stage4_64[16]},
      {stage4_65[9], stage4_65[10], stage4_65[11]},
      {stage4_66[1]},
      {stage4_67[2], stage4_67[3]},
      {stage5_68[1],stage5_67[2],stage5_66[3],stage5_65[4],stage5_64[5]}
   );
   gpc1163_5 gpc9408 (
      {stage4_64[17], stage4_64[18], stage4_64[19]},
      {stage4_65[12], stage4_65[13], stage4_65[14], stage4_65[15], stage4_65[16], stage4_65[17]},
      {stage4_66[2]},
      {stage4_67[4]},
      {stage5_68[2],stage5_67[3],stage5_66[4],stage5_65[5],stage5_64[6]}
   );
   gpc1163_5 gpc9409 (
      {stage4_64[20], stage4_64[21], stage4_64[22]},
      {stage4_65[18], stage4_65[19], stage4_65[20], stage4_65[21], stage4_65[22], stage4_65[23]},
      {stage4_66[3]},
      {stage4_67[5]},
      {stage5_68[3],stage5_67[4],stage5_66[5],stage5_65[6],stage5_64[7]}
   );
   gpc1325_5 gpc9410 (
      {stage4_64[23], stage4_64[24], stage4_64[25], stage4_64[26], stage4_64[27]},
      {stage4_65[24], stage4_65[25]},
      {stage4_66[4], stage4_66[5], stage4_66[6]},
      {stage4_67[6]},
      {stage5_68[4],stage5_67[5],stage5_66[6],stage5_65[7],stage5_64[8]}
   );
   gpc606_5 gpc9411 (
      {stage4_66[7], stage4_66[8], stage4_66[9], stage4_66[10], 1'b0, 1'b0},
      {stage4_68[0], stage4_68[1], stage4_68[2], stage4_68[3], stage4_68[4], stage4_68[5]},
      {stage5_70[0],stage5_69[0],stage5_68[5],stage5_67[6],stage5_66[7]}
   );
   gpc1_1 gpc9412 (
      {stage4_0[5]},
      {stage5_0[1]}
   );
   gpc1_1 gpc9413 (
      {stage4_0[6]},
      {stage5_0[2]}
   );
   gpc1_1 gpc9414 (
      {stage4_0[7]},
      {stage5_0[3]}
   );
   gpc1_1 gpc9415 (
      {stage4_0[8]},
      {stage5_0[4]}
   );
   gpc1_1 gpc9416 (
      {stage4_2[9]},
      {stage5_2[3]}
   );
   gpc1_1 gpc9417 (
      {stage4_2[10]},
      {stage5_2[4]}
   );
   gpc1_1 gpc9418 (
      {stage4_3[12]},
      {stage5_3[3]}
   );
   gpc1_1 gpc9419 (
      {stage4_3[13]},
      {stage5_3[4]}
   );
   gpc1_1 gpc9420 (
      {stage4_3[14]},
      {stage5_3[5]}
   );
   gpc1_1 gpc9421 (
      {stage4_3[15]},
      {stage5_3[6]}
   );
   gpc1_1 gpc9422 (
      {stage4_3[16]},
      {stage5_3[7]}
   );
   gpc1_1 gpc9423 (
      {stage4_4[28]},
      {stage5_4[8]}
   );
   gpc1_1 gpc9424 (
      {stage4_4[29]},
      {stage5_4[9]}
   );
   gpc1_1 gpc9425 (
      {stage4_4[30]},
      {stage5_4[10]}
   );
   gpc1_1 gpc9426 (
      {stage4_5[31]},
      {stage5_5[11]}
   );
   gpc1_1 gpc9427 (
      {stage4_5[32]},
      {stage5_5[12]}
   );
   gpc1_1 gpc9428 (
      {stage4_5[33]},
      {stage5_5[13]}
   );
   gpc1_1 gpc9429 (
      {stage4_5[34]},
      {stage5_5[14]}
   );
   gpc1_1 gpc9430 (
      {stage4_5[35]},
      {stage5_5[15]}
   );
   gpc1_1 gpc9431 (
      {stage4_8[24]},
      {stage5_8[15]}
   );
   gpc1_1 gpc9432 (
      {stage4_8[25]},
      {stage5_8[16]}
   );
   gpc1_1 gpc9433 (
      {stage4_8[26]},
      {stage5_8[17]}
   );
   gpc1_1 gpc9434 (
      {stage4_8[27]},
      {stage5_8[18]}
   );
   gpc1_1 gpc9435 (
      {stage4_10[31]},
      {stage5_10[10]}
   );
   gpc1_1 gpc9436 (
      {stage4_10[32]},
      {stage5_10[11]}
   );
   gpc1_1 gpc9437 (
      {stage4_10[33]},
      {stage5_10[12]}
   );
   gpc1_1 gpc9438 (
      {stage4_10[34]},
      {stage5_10[13]}
   );
   gpc1_1 gpc9439 (
      {stage4_10[35]},
      {stage5_10[14]}
   );
   gpc1_1 gpc9440 (
      {stage4_10[36]},
      {stage5_10[15]}
   );
   gpc1_1 gpc9441 (
      {stage4_10[37]},
      {stage5_10[16]}
   );
   gpc1_1 gpc9442 (
      {stage4_10[38]},
      {stage5_10[17]}
   );
   gpc1_1 gpc9443 (
      {stage4_10[39]},
      {stage5_10[18]}
   );
   gpc1_1 gpc9444 (
      {stage4_10[40]},
      {stage5_10[19]}
   );
   gpc1_1 gpc9445 (
      {stage4_10[41]},
      {stage5_10[20]}
   );
   gpc1_1 gpc9446 (
      {stage4_11[27]},
      {stage5_11[12]}
   );
   gpc1_1 gpc9447 (
      {stage4_11[28]},
      {stage5_11[13]}
   );
   gpc1_1 gpc9448 (
      {stage4_13[26]},
      {stage5_13[9]}
   );
   gpc1_1 gpc9449 (
      {stage4_13[27]},
      {stage5_13[10]}
   );
   gpc1_1 gpc9450 (
      {stage4_13[28]},
      {stage5_13[11]}
   );
   gpc1_1 gpc9451 (
      {stage4_13[29]},
      {stage5_13[12]}
   );
   gpc1_1 gpc9452 (
      {stage4_13[30]},
      {stage5_13[13]}
   );
   gpc1_1 gpc9453 (
      {stage4_13[31]},
      {stage5_13[14]}
   );
   gpc1_1 gpc9454 (
      {stage4_14[26]},
      {stage5_14[12]}
   );
   gpc1_1 gpc9455 (
      {stage4_14[27]},
      {stage5_14[13]}
   );
   gpc1_1 gpc9456 (
      {stage4_14[28]},
      {stage5_14[14]}
   );
   gpc1_1 gpc9457 (
      {stage4_14[29]},
      {stage5_14[15]}
   );
   gpc1_1 gpc9458 (
      {stage4_18[20]},
      {stage5_18[11]}
   );
   gpc1_1 gpc9459 (
      {stage4_19[24]},
      {stage5_19[11]}
   );
   gpc1_1 gpc9460 (
      {stage4_19[25]},
      {stage5_19[12]}
   );
   gpc1_1 gpc9461 (
      {stage4_19[26]},
      {stage5_19[13]}
   );
   gpc1_1 gpc9462 (
      {stage4_19[27]},
      {stage5_19[14]}
   );
   gpc1_1 gpc9463 (
      {stage4_19[28]},
      {stage5_19[15]}
   );
   gpc1_1 gpc9464 (
      {stage4_20[28]},
      {stage5_20[8]}
   );
   gpc1_1 gpc9465 (
      {stage4_20[29]},
      {stage5_20[9]}
   );
   gpc1_1 gpc9466 (
      {stage4_20[30]},
      {stage5_20[10]}
   );
   gpc1_1 gpc9467 (
      {stage4_20[31]},
      {stage5_20[11]}
   );
   gpc1_1 gpc9468 (
      {stage4_20[32]},
      {stage5_20[12]}
   );
   gpc1_1 gpc9469 (
      {stage4_20[33]},
      {stage5_20[13]}
   );
   gpc1_1 gpc9470 (
      {stage4_21[36]},
      {stage5_21[10]}
   );
   gpc1_1 gpc9471 (
      {stage4_24[19]},
      {stage5_24[6]}
   );
   gpc1_1 gpc9472 (
      {stage4_24[20]},
      {stage5_24[7]}
   );
   gpc1_1 gpc9473 (
      {stage4_24[21]},
      {stage5_24[8]}
   );
   gpc1_1 gpc9474 (
      {stage4_26[14]},
      {stage5_26[10]}
   );
   gpc1_1 gpc9475 (
      {stage4_26[15]},
      {stage5_26[11]}
   );
   gpc1_1 gpc9476 (
      {stage4_26[16]},
      {stage5_26[12]}
   );
   gpc1_1 gpc9477 (
      {stage4_26[17]},
      {stage5_26[13]}
   );
   gpc1_1 gpc9478 (
      {stage4_26[18]},
      {stage5_26[14]}
   );
   gpc1_1 gpc9479 (
      {stage4_28[18]},
      {stage5_28[9]}
   );
   gpc1_1 gpc9480 (
      {stage4_29[18]},
      {stage5_29[11]}
   );
   gpc1_1 gpc9481 (
      {stage4_29[19]},
      {stage5_29[12]}
   );
   gpc1_1 gpc9482 (
      {stage4_29[20]},
      {stage5_29[13]}
   );
   gpc1_1 gpc9483 (
      {stage4_29[21]},
      {stage5_29[14]}
   );
   gpc1_1 gpc9484 (
      {stage4_32[20]},
      {stage5_32[10]}
   );
   gpc1_1 gpc9485 (
      {stage4_32[21]},
      {stage5_32[11]}
   );
   gpc1_1 gpc9486 (
      {stage4_32[22]},
      {stage5_32[12]}
   );
   gpc1_1 gpc9487 (
      {stage4_32[23]},
      {stage5_32[13]}
   );
   gpc1_1 gpc9488 (
      {stage4_32[24]},
      {stage5_32[14]}
   );
   gpc1_1 gpc9489 (
      {stage4_32[25]},
      {stage5_32[15]}
   );
   gpc1_1 gpc9490 (
      {stage4_32[26]},
      {stage5_32[16]}
   );
   gpc1_1 gpc9491 (
      {stage4_32[27]},
      {stage5_32[17]}
   );
   gpc1_1 gpc9492 (
      {stage4_32[28]},
      {stage5_32[18]}
   );
   gpc1_1 gpc9493 (
      {stage4_32[29]},
      {stage5_32[19]}
   );
   gpc1_1 gpc9494 (
      {stage4_33[24]},
      {stage5_33[7]}
   );
   gpc1_1 gpc9495 (
      {stage4_33[25]},
      {stage5_33[8]}
   );
   gpc1_1 gpc9496 (
      {stage4_33[26]},
      {stage5_33[9]}
   );
   gpc1_1 gpc9497 (
      {stage4_33[27]},
      {stage5_33[10]}
   );
   gpc1_1 gpc9498 (
      {stage4_33[28]},
      {stage5_33[11]}
   );
   gpc1_1 gpc9499 (
      {stage4_34[15]},
      {stage5_34[10]}
   );
   gpc1_1 gpc9500 (
      {stage4_34[16]},
      {stage5_34[11]}
   );
   gpc1_1 gpc9501 (
      {stage4_34[17]},
      {stage5_34[12]}
   );
   gpc1_1 gpc9502 (
      {stage4_34[18]},
      {stage5_34[13]}
   );
   gpc1_1 gpc9503 (
      {stage4_35[32]},
      {stage5_35[10]}
   );
   gpc1_1 gpc9504 (
      {stage4_35[33]},
      {stage5_35[11]}
   );
   gpc1_1 gpc9505 (
      {stage4_35[34]},
      {stage5_35[12]}
   );
   gpc1_1 gpc9506 (
      {stage4_35[35]},
      {stage5_35[13]}
   );
   gpc1_1 gpc9507 (
      {stage4_36[34]},
      {stage5_36[11]}
   );
   gpc1_1 gpc9508 (
      {stage4_36[35]},
      {stage5_36[12]}
   );
   gpc1_1 gpc9509 (
      {stage4_38[18]},
      {stage5_38[8]}
   );
   gpc1_1 gpc9510 (
      {stage4_38[19]},
      {stage5_38[9]}
   );
   gpc1_1 gpc9511 (
      {stage4_42[29]},
      {stage5_42[10]}
   );
   gpc1_1 gpc9512 (
      {stage4_42[30]},
      {stage5_42[11]}
   );
   gpc1_1 gpc9513 (
      {stage4_42[31]},
      {stage5_42[12]}
   );
   gpc1_1 gpc9514 (
      {stage4_42[32]},
      {stage5_42[13]}
   );
   gpc1_1 gpc9515 (
      {stage4_42[33]},
      {stage5_42[14]}
   );
   gpc1_1 gpc9516 (
      {stage4_42[34]},
      {stage5_42[15]}
   );
   gpc1_1 gpc9517 (
      {stage4_42[35]},
      {stage5_42[16]}
   );
   gpc1_1 gpc9518 (
      {stage4_42[36]},
      {stage5_42[17]}
   );
   gpc1_1 gpc9519 (
      {stage4_42[37]},
      {stage5_42[18]}
   );
   gpc1_1 gpc9520 (
      {stage4_43[12]},
      {stage5_43[9]}
   );
   gpc1_1 gpc9521 (
      {stage4_43[13]},
      {stage5_43[10]}
   );
   gpc1_1 gpc9522 (
      {stage4_44[22]},
      {stage5_44[10]}
   );
   gpc1_1 gpc9523 (
      {stage4_44[23]},
      {stage5_44[11]}
   );
   gpc1_1 gpc9524 (
      {stage4_44[24]},
      {stage5_44[12]}
   );
   gpc1_1 gpc9525 (
      {stage4_45[21]},
      {stage5_45[7]}
   );
   gpc1_1 gpc9526 (
      {stage4_45[22]},
      {stage5_45[8]}
   );
   gpc1_1 gpc9527 (
      {stage4_45[23]},
      {stage5_45[9]}
   );
   gpc1_1 gpc9528 (
      {stage4_45[24]},
      {stage5_45[10]}
   );
   gpc1_1 gpc9529 (
      {stage4_45[25]},
      {stage5_45[11]}
   );
   gpc1_1 gpc9530 (
      {stage4_45[26]},
      {stage5_45[12]}
   );
   gpc1_1 gpc9531 (
      {stage4_45[27]},
      {stage5_45[13]}
   );
   gpc1_1 gpc9532 (
      {stage4_45[28]},
      {stage5_45[14]}
   );
   gpc1_1 gpc9533 (
      {stage4_46[13]},
      {stage5_46[8]}
   );
   gpc1_1 gpc9534 (
      {stage4_46[14]},
      {stage5_46[9]}
   );
   gpc1_1 gpc9535 (
      {stage4_46[15]},
      {stage5_46[10]}
   );
   gpc1_1 gpc9536 (
      {stage4_46[16]},
      {stage5_46[11]}
   );
   gpc1_1 gpc9537 (
      {stage4_47[18]},
      {stage5_47[9]}
   );
   gpc1_1 gpc9538 (
      {stage4_47[19]},
      {stage5_47[10]}
   );
   gpc1_1 gpc9539 (
      {stage4_47[20]},
      {stage5_47[11]}
   );
   gpc1_1 gpc9540 (
      {stage4_48[14]},
      {stage5_48[5]}
   );
   gpc1_1 gpc9541 (
      {stage4_48[15]},
      {stage5_48[6]}
   );
   gpc1_1 gpc9542 (
      {stage4_48[16]},
      {stage5_48[7]}
   );
   gpc1_1 gpc9543 (
      {stage4_48[17]},
      {stage5_48[8]}
   );
   gpc1_1 gpc9544 (
      {stage4_48[18]},
      {stage5_48[9]}
   );
   gpc1_1 gpc9545 (
      {stage4_48[19]},
      {stage5_48[10]}
   );
   gpc1_1 gpc9546 (
      {stage4_48[20]},
      {stage5_48[11]}
   );
   gpc1_1 gpc9547 (
      {stage4_48[21]},
      {stage5_48[12]}
   );
   gpc1_1 gpc9548 (
      {stage4_48[22]},
      {stage5_48[13]}
   );
   gpc1_1 gpc9549 (
      {stage4_49[12]},
      {stage5_49[5]}
   );
   gpc1_1 gpc9550 (
      {stage4_50[17]},
      {stage5_50[7]}
   );
   gpc1_1 gpc9551 (
      {stage4_50[18]},
      {stage5_50[8]}
   );
   gpc1_1 gpc9552 (
      {stage4_50[19]},
      {stage5_50[9]}
   );
   gpc1_1 gpc9553 (
      {stage4_50[20]},
      {stage5_50[10]}
   );
   gpc1_1 gpc9554 (
      {stage4_50[21]},
      {stage5_50[11]}
   );
   gpc1_1 gpc9555 (
      {stage4_51[27]},
      {stage5_51[10]}
   );
   gpc1_1 gpc9556 (
      {stage4_51[28]},
      {stage5_51[11]}
   );
   gpc1_1 gpc9557 (
      {stage4_51[29]},
      {stage5_51[12]}
   );
   gpc1_1 gpc9558 (
      {stage4_51[30]},
      {stage5_51[13]}
   );
   gpc1_1 gpc9559 (
      {stage4_51[31]},
      {stage5_51[14]}
   );
   gpc1_1 gpc9560 (
      {stage4_51[32]},
      {stage5_51[15]}
   );
   gpc1_1 gpc9561 (
      {stage4_51[33]},
      {stage5_51[16]}
   );
   gpc1_1 gpc9562 (
      {stage4_51[34]},
      {stage5_51[17]}
   );
   gpc1_1 gpc9563 (
      {stage4_51[35]},
      {stage5_51[18]}
   );
   gpc1_1 gpc9564 (
      {stage4_52[17]},
      {stage5_52[8]}
   );
   gpc1_1 gpc9565 (
      {stage4_52[18]},
      {stage5_52[9]}
   );
   gpc1_1 gpc9566 (
      {stage4_53[40]},
      {stage5_53[9]}
   );
   gpc1_1 gpc9567 (
      {stage4_53[41]},
      {stage5_53[10]}
   );
   gpc1_1 gpc9568 (
      {stage4_53[42]},
      {stage5_53[11]}
   );
   gpc1_1 gpc9569 (
      {stage4_53[43]},
      {stage5_53[12]}
   );
   gpc1_1 gpc9570 (
      {stage4_54[22]},
      {stage5_54[13]}
   );
   gpc1_1 gpc9571 (
      {stage4_54[23]},
      {stage5_54[14]}
   );
   gpc1_1 gpc9572 (
      {stage4_54[24]},
      {stage5_54[15]}
   );
   gpc1_1 gpc9573 (
      {stage4_54[25]},
      {stage5_54[16]}
   );
   gpc1_1 gpc9574 (
      {stage4_55[29]},
      {stage5_55[12]}
   );
   gpc1_1 gpc9575 (
      {stage4_55[30]},
      {stage5_55[13]}
   );
   gpc1_1 gpc9576 (
      {stage4_55[31]},
      {stage5_55[14]}
   );
   gpc1_1 gpc9577 (
      {stage4_55[32]},
      {stage5_55[15]}
   );
   gpc1_1 gpc9578 (
      {stage4_55[33]},
      {stage5_55[16]}
   );
   gpc1_1 gpc9579 (
      {stage4_55[34]},
      {stage5_55[17]}
   );
   gpc1_1 gpc9580 (
      {stage4_55[35]},
      {stage5_55[18]}
   );
   gpc1_1 gpc9581 (
      {stage4_55[36]},
      {stage5_55[19]}
   );
   gpc1_1 gpc9582 (
      {stage4_55[37]},
      {stage5_55[20]}
   );
   gpc1_1 gpc9583 (
      {stage4_55[38]},
      {stage5_55[21]}
   );
   gpc1_1 gpc9584 (
      {stage4_57[22]},
      {stage5_57[10]}
   );
   gpc1_1 gpc9585 (
      {stage4_57[23]},
      {stage5_57[11]}
   );
   gpc1_1 gpc9586 (
      {stage4_57[24]},
      {stage5_57[12]}
   );
   gpc1_1 gpc9587 (
      {stage4_57[25]},
      {stage5_57[13]}
   );
   gpc1_1 gpc9588 (
      {stage4_58[17]},
      {stage5_58[9]}
   );
   gpc1_1 gpc9589 (
      {stage4_58[18]},
      {stage5_58[10]}
   );
   gpc1_1 gpc9590 (
      {stage4_58[19]},
      {stage5_58[11]}
   );
   gpc1_1 gpc9591 (
      {stage4_58[20]},
      {stage5_58[12]}
   );
   gpc1_1 gpc9592 (
      {stage4_58[21]},
      {stage5_58[13]}
   );
   gpc1_1 gpc9593 (
      {stage4_58[22]},
      {stage5_58[14]}
   );
   gpc1_1 gpc9594 (
      {stage4_58[23]},
      {stage5_58[15]}
   );
   gpc1_1 gpc9595 (
      {stage4_60[15]},
      {stage5_60[8]}
   );
   gpc1_1 gpc9596 (
      {stage4_60[16]},
      {stage5_60[9]}
   );
   gpc1_1 gpc9597 (
      {stage4_60[17]},
      {stage5_60[10]}
   );
   gpc1_1 gpc9598 (
      {stage4_60[18]},
      {stage5_60[11]}
   );
   gpc1_1 gpc9599 (
      {stage4_60[19]},
      {stage5_60[12]}
   );
   gpc1_1 gpc9600 (
      {stage4_60[20]},
      {stage5_60[13]}
   );
   gpc1_1 gpc9601 (
      {stage4_60[21]},
      {stage5_60[14]}
   );
   gpc1_1 gpc9602 (
      {stage4_61[23]},
      {stage5_61[7]}
   );
   gpc1_1 gpc9603 (
      {stage4_61[24]},
      {stage5_61[8]}
   );
   gpc1_1 gpc9604 (
      {stage4_61[25]},
      {stage5_61[9]}
   );
   gpc1_1 gpc9605 (
      {stage4_61[26]},
      {stage5_61[10]}
   );
   gpc1_1 gpc9606 (
      {stage4_61[27]},
      {stage5_61[11]}
   );
   gpc1_1 gpc9607 (
      {stage4_61[28]},
      {stage5_61[12]}
   );
   gpc1_1 gpc9608 (
      {stage4_61[29]},
      {stage5_61[13]}
   );
   gpc1_1 gpc9609 (
      {stage4_61[30]},
      {stage5_61[14]}
   );
   gpc1_1 gpc9610 (
      {stage4_61[31]},
      {stage5_61[15]}
   );
   gpc1_1 gpc9611 (
      {stage4_62[12]},
      {stage5_62[7]}
   );
   gpc1_1 gpc9612 (
      {stage4_62[13]},
      {stage5_62[8]}
   );
   gpc1_1 gpc9613 (
      {stage4_62[14]},
      {stage5_62[9]}
   );
   gpc1_1 gpc9614 (
      {stage4_62[15]},
      {stage5_62[10]}
   );
   gpc1_1 gpc9615 (
      {stage4_62[16]},
      {stage5_62[11]}
   );
   gpc1_1 gpc9616 (
      {stage4_63[12]},
      {stage5_63[7]}
   );
   gpc1_1 gpc9617 (
      {stage4_63[13]},
      {stage5_63[8]}
   );
   gpc1_1 gpc9618 (
      {stage4_64[28]},
      {stage5_64[9]}
   );
   gpc1_1 gpc9619 (
      {stage4_64[29]},
      {stage5_64[10]}
   );
   gpc1_1 gpc9620 (
      {stage4_64[30]},
      {stage5_64[11]}
   );
   gpc1_1 gpc9621 (
      {stage4_64[31]},
      {stage5_64[12]}
   );
   gpc1_1 gpc9622 (
      {stage4_64[32]},
      {stage5_64[13]}
   );
   gpc1_1 gpc9623 (
      {stage4_64[33]},
      {stage5_64[14]}
   );
   gpc1_1 gpc9624 (
      {stage4_65[26]},
      {stage5_65[8]}
   );
   gpc1_1 gpc9625 (
      {stage4_65[27]},
      {stage5_65[9]}
   );
   gpc1_1 gpc9626 (
      {stage4_65[28]},
      {stage5_65[10]}
   );
   gpc1_1 gpc9627 (
      {stage4_65[29]},
      {stage5_65[11]}
   );
   gpc1_1 gpc9628 (
      {stage4_65[30]},
      {stage5_65[12]}
   );
   gpc1_1 gpc9629 (
      {stage4_65[31]},
      {stage5_65[13]}
   );
   gpc1_1 gpc9630 (
      {stage4_65[32]},
      {stage5_65[14]}
   );
   gpc1_1 gpc9631 (
      {stage4_65[33]},
      {stage5_65[15]}
   );
   gpc1_1 gpc9632 (
      {stage4_65[34]},
      {stage5_65[16]}
   );
   gpc1_1 gpc9633 (
      {stage4_65[35]},
      {stage5_65[17]}
   );
   gpc1_1 gpc9634 (
      {stage4_67[7]},
      {stage5_67[7]}
   );
   gpc1_1 gpc9635 (
      {stage4_67[8]},
      {stage5_67[8]}
   );
   gpc1_1 gpc9636 (
      {stage4_67[9]},
      {stage5_67[9]}
   );
   gpc1_1 gpc9637 (
      {stage4_67[10]},
      {stage5_67[10]}
   );
   gpc1_1 gpc9638 (
      {stage4_68[6]},
      {stage5_68[6]}
   );
   gpc1_1 gpc9639 (
      {stage4_68[7]},
      {stage5_68[7]}
   );
   gpc1_1 gpc9640 (
      {stage4_68[8]},
      {stage5_68[8]}
   );
   gpc1_1 gpc9641 (
      {stage4_68[9]},
      {stage5_68[9]}
   );
   gpc1_1 gpc9642 (
      {stage4_68[10]},
      {stage5_68[10]}
   );
   gpc1_1 gpc9643 (
      {stage4_68[11]},
      {stage5_68[11]}
   );
   gpc1_1 gpc9644 (
      {stage4_68[12]},
      {stage5_68[12]}
   );
   gpc1_1 gpc9645 (
      {stage4_68[13]},
      {stage5_68[13]}
   );
   gpc1_1 gpc9646 (
      {stage4_69[0]},
      {stage5_69[1]}
   );
   gpc1_1 gpc9647 (
      {stage4_69[1]},
      {stage5_69[2]}
   );
   gpc615_5 gpc9648 (
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0]}
   );
   gpc615_5 gpc9649 (
      {stage5_3[5], stage5_3[6], stage5_3[7], 1'b0, 1'b0},
      {stage5_4[1]},
      {stage5_5[6], stage5_5[7], stage5_5[8], stage5_5[9], stage5_5[10], stage5_5[11]},
      {stage6_7[1],stage6_6[1],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc606_5 gpc9650 (
      {stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6], stage5_4[7]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5]},
      {stage6_8[0],stage6_7[2],stage6_6[2],stage6_5[2],stage6_4[2]}
   );
   gpc606_5 gpc9651 (
      {stage5_5[12], stage5_5[13], stage5_5[14], stage5_5[15], 1'b0, 1'b0},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage6_9[0],stage6_8[1],stage6_7[3],stage6_6[3],stage6_5[3]}
   );
   gpc615_5 gpc9652 (
      {stage5_7[6], stage5_7[7], stage5_7[8], stage5_7[9], stage5_7[10]},
      {stage5_8[0]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[2],stage6_7[4]}
   );
   gpc606_5 gpc9653 (
      {stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5], stage5_8[6]},
      {stage5_10[0], stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage6_12[0],stage6_11[1],stage6_10[1],stage6_9[2],stage6_8[3]}
   );
   gpc606_5 gpc9654 (
      {stage5_8[7], stage5_8[8], stage5_8[9], stage5_8[10], stage5_8[11], stage5_8[12]},
      {stage5_10[6], stage5_10[7], stage5_10[8], stage5_10[9], stage5_10[10], stage5_10[11]},
      {stage6_12[1],stage6_11[2],stage6_10[2],stage6_9[3],stage6_8[4]}
   );
   gpc606_5 gpc9655 (
      {stage5_8[13], stage5_8[14], stage5_8[15], stage5_8[16], stage5_8[17], stage5_8[18]},
      {stage5_10[12], stage5_10[13], stage5_10[14], stage5_10[15], stage5_10[16], stage5_10[17]},
      {stage6_12[2],stage6_11[3],stage6_10[3],stage6_9[4],stage6_8[5]}
   );
   gpc615_5 gpc9656 (
      {stage5_10[18], stage5_10[19], stage5_10[20], 1'b0, 1'b0},
      {stage5_11[0]},
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5]},
      {stage6_14[0],stage6_13[0],stage6_12[3],stage6_11[4],stage6_10[4]}
   );
   gpc1406_5 gpc9657 (
      {stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[0]},
      {stage6_15[0],stage6_14[1],stage6_13[1],stage6_12[4],stage6_11[5]}
   );
   gpc7_3 gpc9658 (
      {stage5_11[7], stage5_11[8], stage5_11[9], stage5_11[10], stage5_11[11], stage5_11[12], stage5_11[13]},
      {stage6_13[2],stage6_12[5],stage6_11[6]}
   );
   gpc606_5 gpc9659 (
      {stage5_12[6], stage5_12[7], stage5_12[8], stage5_12[9], stage5_12[10], 1'b0},
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5], stage5_14[6]},
      {stage6_16[0],stage6_15[1],stage6_14[2],stage6_13[3],stage6_12[6]}
   );
   gpc606_5 gpc9660 (
      {stage5_13[4], stage5_13[5], stage5_13[6], stage5_13[7], stage5_13[8], stage5_13[9]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage6_17[0],stage6_16[1],stage6_15[2],stage6_14[3],stage6_13[4]}
   );
   gpc1343_5 gpc9661 (
      {stage5_14[7], stage5_14[8], stage5_14[9]},
      {stage5_15[6], stage5_15[7], stage5_15[8], stage5_15[9]},
      {stage5_16[0], stage5_16[1], stage5_16[2]},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[1],stage6_16[2],stage6_15[3],stage6_14[4]}
   );
   gpc615_5 gpc9662 (
      {stage5_14[10], stage5_14[11], stage5_14[12], stage5_14[13], stage5_14[14]},
      {stage5_15[10]},
      {stage5_16[3], stage5_16[4], stage5_16[5], stage5_16[6], stage5_16[7], 1'b0},
      {stage6_18[1],stage6_17[2],stage6_16[3],stage6_15[4],stage6_14[5]}
   );
   gpc615_5 gpc9663 (
      {stage5_14[15], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage5_15[11]},
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage6_18[2],stage6_17[3],stage6_16[4],stage6_15[5],stage6_14[6]}
   );
   gpc606_5 gpc9664 (
      {stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5], stage5_17[6]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[3],stage6_17[4]}
   );
   gpc117_4 gpc9665 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5], stage5_18[6]},
      {stage5_19[6]},
      {stage5_20[0]},
      {stage6_21[1],stage6_20[1],stage6_19[1],stage6_18[4]}
   );
   gpc615_5 gpc9666 (
      {stage5_18[7], stage5_18[8], stage5_18[9], stage5_18[10], stage5_18[11]},
      {stage5_19[7]},
      {stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5], stage5_20[6]},
      {stage6_22[0],stage6_21[2],stage6_20[2],stage6_19[2],stage6_18[5]}
   );
   gpc615_5 gpc9667 (
      {stage5_19[8], stage5_19[9], stage5_19[10], stage5_19[11], stage5_19[12]},
      {stage5_20[7]},
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5]},
      {stage6_23[0],stage6_22[1],stage6_21[3],stage6_20[3],stage6_19[3]}
   );
   gpc615_5 gpc9668 (
      {stage5_19[13], stage5_19[14], stage5_19[15], 1'b0, 1'b0},
      {stage5_20[8]},
      {stage5_21[6], stage5_21[7], stage5_21[8], stage5_21[9], stage5_21[10], 1'b0},
      {stage6_23[1],stage6_22[2],stage6_21[4],stage6_20[4],stage6_19[4]}
   );
   gpc606_5 gpc9669 (
      {stage5_20[9], stage5_20[10], stage5_20[11], stage5_20[12], stage5_20[13], 1'b0},
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4], stage5_22[5]},
      {stage6_24[0],stage6_23[2],stage6_22[3],stage6_21[5],stage6_20[5]}
   );
   gpc15_3 gpc9670 (
      {stage5_22[6], stage5_22[7], stage5_22[8], stage5_22[9], stage5_22[10]},
      {stage5_23[0]},
      {stage6_24[1],stage6_23[3],stage6_22[4]}
   );
   gpc15_3 gpc9671 (
      {stage5_22[11], stage5_22[12], stage5_22[13], 1'b0, 1'b0},
      {stage5_23[1]},
      {stage6_24[2],stage6_23[4],stage6_22[5]}
   );
   gpc615_5 gpc9672 (
      {stage5_23[2], stage5_23[3], stage5_23[4], stage5_23[5], stage5_23[6]},
      {stage5_24[0]},
      {stage5_25[0], stage5_25[1], stage5_25[2], stage5_25[3], stage5_25[4], stage5_25[5]},
      {stage6_27[0],stage6_26[0],stage6_25[0],stage6_24[3],stage6_23[5]}
   );
   gpc615_5 gpc9673 (
      {stage5_23[7], stage5_23[8], stage5_23[9], 1'b0, 1'b0},
      {stage5_24[1]},
      {stage5_25[6], stage5_25[7], stage5_25[8], stage5_25[9], 1'b0, 1'b0},
      {stage6_27[1],stage6_26[1],stage6_25[1],stage6_24[4],stage6_23[6]}
   );
   gpc606_5 gpc9674 (
      {stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], stage5_24[6], stage5_24[7]},
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5]},
      {stage6_28[0],stage6_27[2],stage6_26[2],stage6_25[2],stage6_24[5]}
   );
   gpc615_5 gpc9675 (
      {stage5_26[6], stage5_26[7], stage5_26[8], stage5_26[9], stage5_26[10]},
      {stage5_27[0]},
      {stage5_28[0], stage5_28[1], stage5_28[2], stage5_28[3], stage5_28[4], stage5_28[5]},
      {stage6_30[0],stage6_29[0],stage6_28[1],stage6_27[3],stage6_26[3]}
   );
   gpc615_5 gpc9676 (
      {stage5_27[1], stage5_27[2], stage5_27[3], stage5_27[4], stage5_27[5]},
      {stage5_28[6]},
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage6_31[0],stage6_30[1],stage6_29[1],stage6_28[2],stage6_27[4]}
   );
   gpc606_5 gpc9677 (
      {stage5_29[6], stage5_29[7], stage5_29[8], stage5_29[9], stage5_29[10], stage5_29[11]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[0],stage6_31[1],stage6_30[2],stage6_29[2]}
   );
   gpc615_5 gpc9678 (
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4]},
      {stage5_31[6]},
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4], stage5_32[5]},
      {stage6_34[0],stage6_33[1],stage6_32[1],stage6_31[2],stage6_30[3]}
   );
   gpc615_5 gpc9679 (
      {stage5_30[5], stage5_30[6], stage5_30[7], stage5_30[8], 1'b0},
      {stage5_31[7]},
      {stage5_32[6], stage5_32[7], stage5_32[8], stage5_32[9], stage5_32[10], stage5_32[11]},
      {stage6_34[1],stage6_33[2],stage6_32[2],stage6_31[3],stage6_30[4]}
   );
   gpc606_5 gpc9680 (
      {stage5_32[12], stage5_32[13], stage5_32[14], stage5_32[15], stage5_32[16], stage5_32[17]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], stage5_34[4], stage5_34[5]},
      {stage6_36[0],stage6_35[0],stage6_34[2],stage6_33[3],stage6_32[3]}
   );
   gpc606_5 gpc9681 (
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage6_37[0],stage6_36[1],stage6_35[1],stage6_34[3],stage6_33[4]}
   );
   gpc606_5 gpc9682 (
      {stage5_33[6], stage5_33[7], stage5_33[8], stage5_33[9], stage5_33[10], stage5_33[11]},
      {stage5_35[6], stage5_35[7], stage5_35[8], stage5_35[9], stage5_35[10], stage5_35[11]},
      {stage6_37[1],stage6_36[2],stage6_35[2],stage6_34[4],stage6_33[5]}
   );
   gpc615_5 gpc9683 (
      {stage5_34[6], stage5_34[7], stage5_34[8], stage5_34[9], stage5_34[10]},
      {stage5_35[12]},
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3], stage5_36[4], stage5_36[5]},
      {stage6_38[0],stage6_37[2],stage6_36[3],stage6_35[3],stage6_34[5]}
   );
   gpc606_5 gpc9684 (
      {stage5_36[6], stage5_36[7], stage5_36[8], stage5_36[9], stage5_36[10], stage5_36[11]},
      {stage5_38[0], stage5_38[1], stage5_38[2], stage5_38[3], stage5_38[4], stage5_38[5]},
      {stage6_40[0],stage6_39[0],stage6_38[1],stage6_37[3],stage6_36[4]}
   );
   gpc2135_5 gpc9685 (
      {stage5_37[0], stage5_37[1], stage5_37[2], stage5_37[3], stage5_37[4]},
      {stage5_38[6], stage5_38[7], stage5_38[8]},
      {stage5_39[0]},
      {stage5_40[0], stage5_40[1]},
      {stage6_41[0],stage6_40[1],stage6_39[1],stage6_38[2],stage6_37[4]}
   );
   gpc606_5 gpc9686 (
      {stage5_37[5], stage5_37[6], stage5_37[7], stage5_37[8], stage5_37[9], stage5_37[10]},
      {stage5_39[1], stage5_39[2], stage5_39[3], stage5_39[4], stage5_39[5], stage5_39[6]},
      {stage6_41[1],stage6_40[2],stage6_39[2],stage6_38[3],stage6_37[5]}
   );
   gpc23_3 gpc9687 (
      {stage5_39[7], stage5_39[8], stage5_39[9]},
      {stage5_40[2], stage5_40[3]},
      {stage6_41[2],stage6_40[3],stage6_39[3]}
   );
   gpc606_5 gpc9688 (
      {stage5_40[4], stage5_40[5], stage5_40[6], stage5_40[7], stage5_40[8], stage5_40[9]},
      {stage5_42[0], stage5_42[1], stage5_42[2], stage5_42[3], stage5_42[4], stage5_42[5]},
      {stage6_44[0],stage6_43[0],stage6_42[0],stage6_41[3],stage6_40[4]}
   );
   gpc606_5 gpc9689 (
      {stage5_41[0], stage5_41[1], stage5_41[2], stage5_41[3], stage5_41[4], stage5_41[5]},
      {stage5_43[0], stage5_43[1], stage5_43[2], stage5_43[3], stage5_43[4], stage5_43[5]},
      {stage6_45[0],stage6_44[1],stage6_43[1],stage6_42[1],stage6_41[4]}
   );
   gpc615_5 gpc9690 (
      {stage5_42[6], stage5_42[7], stage5_42[8], stage5_42[9], stage5_42[10]},
      {stage5_43[6]},
      {stage5_44[0], stage5_44[1], stage5_44[2], stage5_44[3], stage5_44[4], stage5_44[5]},
      {stage6_46[0],stage6_45[1],stage6_44[2],stage6_43[2],stage6_42[2]}
   );
   gpc615_5 gpc9691 (
      {stage5_42[11], stage5_42[12], stage5_42[13], stage5_42[14], stage5_42[15]},
      {stage5_43[7]},
      {stage5_44[6], stage5_44[7], stage5_44[8], stage5_44[9], stage5_44[10], stage5_44[11]},
      {stage6_46[1],stage6_45[2],stage6_44[3],stage6_43[3],stage6_42[3]}
   );
   gpc1163_5 gpc9692 (
      {stage5_45[0], stage5_45[1], stage5_45[2]},
      {stage5_46[0], stage5_46[1], stage5_46[2], stage5_46[3], stage5_46[4], stage5_46[5]},
      {stage5_47[0]},
      {stage5_48[0]},
      {stage6_49[0],stage6_48[0],stage6_47[0],stage6_46[2],stage6_45[3]}
   );
   gpc1163_5 gpc9693 (
      {stage5_45[3], stage5_45[4], stage5_45[5]},
      {stage5_46[6], stage5_46[7], stage5_46[8], stage5_46[9], stage5_46[10], stage5_46[11]},
      {stage5_47[1]},
      {stage5_48[1]},
      {stage6_49[1],stage6_48[1],stage6_47[1],stage6_46[3],stage6_45[4]}
   );
   gpc606_5 gpc9694 (
      {stage5_45[6], stage5_45[7], stage5_45[8], stage5_45[9], stage5_45[10], stage5_45[11]},
      {stage5_47[2], stage5_47[3], stage5_47[4], stage5_47[5], stage5_47[6], stage5_47[7]},
      {stage6_49[2],stage6_48[2],stage6_47[2],stage6_46[4],stage6_45[5]}
   );
   gpc606_5 gpc9695 (
      {stage5_48[2], stage5_48[3], stage5_48[4], stage5_48[5], stage5_48[6], stage5_48[7]},
      {stage5_50[0], stage5_50[1], stage5_50[2], stage5_50[3], stage5_50[4], stage5_50[5]},
      {stage6_52[0],stage6_51[0],stage6_50[0],stage6_49[3],stage6_48[3]}
   );
   gpc606_5 gpc9696 (
      {stage5_48[8], stage5_48[9], stage5_48[10], stage5_48[11], stage5_48[12], stage5_48[13]},
      {stage5_50[6], stage5_50[7], stage5_50[8], stage5_50[9], stage5_50[10], stage5_50[11]},
      {stage6_52[1],stage6_51[1],stage6_50[1],stage6_49[4],stage6_48[4]}
   );
   gpc606_5 gpc9697 (
      {stage5_49[0], stage5_49[1], stage5_49[2], stage5_49[3], stage5_49[4], stage5_49[5]},
      {stage5_51[0], stage5_51[1], stage5_51[2], stage5_51[3], stage5_51[4], stage5_51[5]},
      {stage6_53[0],stage6_52[2],stage6_51[2],stage6_50[2],stage6_49[5]}
   );
   gpc7_3 gpc9698 (
      {stage5_51[6], stage5_51[7], stage5_51[8], stage5_51[9], stage5_51[10], stage5_51[11], stage5_51[12]},
      {stage6_53[1],stage6_52[3],stage6_51[3]}
   );
   gpc623_5 gpc9699 (
      {stage5_51[13], stage5_51[14], stage5_51[15]},
      {stage5_52[0], stage5_52[1]},
      {stage5_53[0], stage5_53[1], stage5_53[2], stage5_53[3], stage5_53[4], stage5_53[5]},
      {stage6_55[0],stage6_54[0],stage6_53[2],stage6_52[4],stage6_51[4]}
   );
   gpc117_4 gpc9700 (
      {stage5_52[2], stage5_52[3], stage5_52[4], stage5_52[5], stage5_52[6], stage5_52[7], stage5_52[8]},
      {stage5_53[6]},
      {stage5_54[0]},
      {stage6_55[1],stage6_54[1],stage6_53[3],stage6_52[5]}
   );
   gpc117_4 gpc9701 (
      {stage5_53[7], stage5_53[8], stage5_53[9], stage5_53[10], stage5_53[11], stage5_53[12], 1'b0},
      {stage5_54[1]},
      {stage5_55[0]},
      {stage6_56[0],stage6_55[2],stage6_54[2],stage6_53[4]}
   );
   gpc135_4 gpc9702 (
      {stage5_54[2], stage5_54[3], stage5_54[4], stage5_54[5], stage5_54[6]},
      {stage5_55[1], stage5_55[2], stage5_55[3]},
      {stage5_56[0]},
      {stage6_57[0],stage6_56[1],stage6_55[3],stage6_54[3]}
   );
   gpc135_4 gpc9703 (
      {stage5_54[7], stage5_54[8], stage5_54[9], stage5_54[10], stage5_54[11]},
      {stage5_55[4], stage5_55[5], stage5_55[6]},
      {stage5_56[1]},
      {stage6_57[1],stage6_56[2],stage6_55[4],stage6_54[4]}
   );
   gpc135_4 gpc9704 (
      {stage5_54[12], stage5_54[13], stage5_54[14], stage5_54[15], stage5_54[16]},
      {stage5_55[7], stage5_55[8], stage5_55[9]},
      {stage5_56[2]},
      {stage6_57[2],stage6_56[3],stage6_55[5],stage6_54[5]}
   );
   gpc615_5 gpc9705 (
      {stage5_55[10], stage5_55[11], stage5_55[12], stage5_55[13], stage5_55[14]},
      {stage5_56[3]},
      {stage5_57[0], stage5_57[1], stage5_57[2], stage5_57[3], stage5_57[4], stage5_57[5]},
      {stage6_59[0],stage6_58[0],stage6_57[3],stage6_56[4],stage6_55[6]}
   );
   gpc615_5 gpc9706 (
      {stage5_55[15], stage5_55[16], stage5_55[17], stage5_55[18], stage5_55[19]},
      {stage5_56[4]},
      {stage5_57[6], stage5_57[7], stage5_57[8], stage5_57[9], stage5_57[10], stage5_57[11]},
      {stage6_59[1],stage6_58[1],stage6_57[4],stage6_56[5],stage6_55[7]}
   );
   gpc2135_5 gpc9707 (
      {stage5_58[0], stage5_58[1], stage5_58[2], stage5_58[3], stage5_58[4]},
      {stage5_59[0], stage5_59[1], stage5_59[2]},
      {stage5_60[0]},
      {stage5_61[0], stage5_61[1]},
      {stage6_62[0],stage6_61[0],stage6_60[0],stage6_59[2],stage6_58[2]}
   );
   gpc2135_5 gpc9708 (
      {stage5_58[5], stage5_58[6], stage5_58[7], stage5_58[8], stage5_58[9]},
      {stage5_59[3], stage5_59[4], stage5_59[5]},
      {stage5_60[1]},
      {stage5_61[2], stage5_61[3]},
      {stage6_62[1],stage6_61[1],stage6_60[1],stage6_59[3],stage6_58[3]}
   );
   gpc2135_5 gpc9709 (
      {stage5_58[10], stage5_58[11], stage5_58[12], stage5_58[13], stage5_58[14]},
      {stage5_59[6], stage5_59[7], 1'b0},
      {stage5_60[2]},
      {stage5_61[4], stage5_61[5]},
      {stage6_62[2],stage6_61[2],stage6_60[2],stage6_59[4],stage6_58[4]}
   );
   gpc606_5 gpc9710 (
      {stage5_60[3], stage5_60[4], stage5_60[5], stage5_60[6], stage5_60[7], stage5_60[8]},
      {stage5_62[0], stage5_62[1], stage5_62[2], stage5_62[3], stage5_62[4], stage5_62[5]},
      {stage6_64[0],stage6_63[0],stage6_62[3],stage6_61[3],stage6_60[3]}
   );
   gpc606_5 gpc9711 (
      {stage5_60[9], stage5_60[10], stage5_60[11], stage5_60[12], stage5_60[13], stage5_60[14]},
      {stage5_62[6], stage5_62[7], stage5_62[8], stage5_62[9], stage5_62[10], stage5_62[11]},
      {stage6_64[1],stage6_63[1],stage6_62[4],stage6_61[4],stage6_60[4]}
   );
   gpc207_4 gpc9712 (
      {stage5_61[6], stage5_61[7], stage5_61[8], stage5_61[9], stage5_61[10], stage5_61[11], stage5_61[12]},
      {stage5_63[0], stage5_63[1]},
      {stage6_64[2],stage6_63[2],stage6_62[5],stage6_61[5]}
   );
   gpc606_5 gpc9713 (
      {stage5_63[2], stage5_63[3], stage5_63[4], stage5_63[5], stage5_63[6], stage5_63[7]},
      {stage5_65[0], stage5_65[1], stage5_65[2], stage5_65[3], stage5_65[4], stage5_65[5]},
      {stage6_67[0],stage6_66[0],stage6_65[0],stage6_64[3],stage6_63[3]}
   );
   gpc1406_5 gpc9714 (
      {stage5_64[0], stage5_64[1], stage5_64[2], stage5_64[3], stage5_64[4], stage5_64[5]},
      {stage5_66[0], stage5_66[1], stage5_66[2], stage5_66[3]},
      {stage5_67[0]},
      {stage6_68[0],stage6_67[1],stage6_66[1],stage6_65[1],stage6_64[4]}
   );
   gpc1406_5 gpc9715 (
      {stage5_64[6], stage5_64[7], stage5_64[8], stage5_64[9], stage5_64[10], stage5_64[11]},
      {stage5_66[4], stage5_66[5], stage5_66[6], stage5_66[7]},
      {stage5_67[1]},
      {stage6_68[1],stage6_67[2],stage6_66[2],stage6_65[2],stage6_64[5]}
   );
   gpc1406_5 gpc9716 (
      {stage5_65[6], stage5_65[7], stage5_65[8], stage5_65[9], stage5_65[10], stage5_65[11]},
      {stage5_67[2], stage5_67[3], stage5_67[4], stage5_67[5]},
      {stage5_68[0]},
      {stage6_69[0],stage6_68[2],stage6_67[3],stage6_66[3],stage6_65[3]}
   );
   gpc606_5 gpc9717 (
      {stage5_65[12], stage5_65[13], stage5_65[14], stage5_65[15], stage5_65[16], stage5_65[17]},
      {stage5_67[6], stage5_67[7], stage5_67[8], stage5_67[9], stage5_67[10], 1'b0},
      {stage6_69[1],stage6_68[3],stage6_67[4],stage6_66[4],stage6_65[4]}
   );
   gpc1_1 gpc9718 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc9719 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc9720 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc9721 (
      {stage5_0[3]},
      {stage6_0[3]}
   );
   gpc1_1 gpc9722 (
      {stage5_0[4]},
      {stage6_0[4]}
   );
   gpc1_1 gpc9723 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc9724 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc9725 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc9726 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc9727 (
      {stage5_2[2]},
      {stage6_2[2]}
   );
   gpc1_1 gpc9728 (
      {stage5_2[3]},
      {stage6_2[3]}
   );
   gpc1_1 gpc9729 (
      {stage5_2[4]},
      {stage6_2[4]}
   );
   gpc1_1 gpc9730 (
      {stage5_4[8]},
      {stage6_4[3]}
   );
   gpc1_1 gpc9731 (
      {stage5_4[9]},
      {stage6_4[4]}
   );
   gpc1_1 gpc9732 (
      {stage5_4[10]},
      {stage6_4[5]}
   );
   gpc1_1 gpc9733 (
      {stage5_6[6]},
      {stage6_6[4]}
   );
   gpc1_1 gpc9734 (
      {stage5_6[7]},
      {stage6_6[5]}
   );
   gpc1_1 gpc9735 (
      {stage5_6[8]},
      {stage6_6[6]}
   );
   gpc1_1 gpc9736 (
      {stage5_6[9]},
      {stage6_6[7]}
   );
   gpc1_1 gpc9737 (
      {stage5_9[6]},
      {stage6_9[5]}
   );
   gpc1_1 gpc9738 (
      {stage5_9[7]},
      {stage6_9[6]}
   );
   gpc1_1 gpc9739 (
      {stage5_9[8]},
      {stage6_9[7]}
   );
   gpc1_1 gpc9740 (
      {stage5_9[9]},
      {stage6_9[8]}
   );
   gpc1_1 gpc9741 (
      {stage5_9[10]},
      {stage6_9[9]}
   );
   gpc1_1 gpc9742 (
      {stage5_13[10]},
      {stage6_13[5]}
   );
   gpc1_1 gpc9743 (
      {stage5_13[11]},
      {stage6_13[6]}
   );
   gpc1_1 gpc9744 (
      {stage5_13[12]},
      {stage6_13[7]}
   );
   gpc1_1 gpc9745 (
      {stage5_13[13]},
      {stage6_13[8]}
   );
   gpc1_1 gpc9746 (
      {stage5_13[14]},
      {stage6_13[9]}
   );
   gpc1_1 gpc9747 (
      {stage5_24[8]},
      {stage6_24[6]}
   );
   gpc1_1 gpc9748 (
      {stage5_26[11]},
      {stage6_26[4]}
   );
   gpc1_1 gpc9749 (
      {stage5_26[12]},
      {stage6_26[5]}
   );
   gpc1_1 gpc9750 (
      {stage5_26[13]},
      {stage6_26[6]}
   );
   gpc1_1 gpc9751 (
      {stage5_26[14]},
      {stage6_26[7]}
   );
   gpc1_1 gpc9752 (
      {stage5_28[7]},
      {stage6_28[3]}
   );
   gpc1_1 gpc9753 (
      {stage5_28[8]},
      {stage6_28[4]}
   );
   gpc1_1 gpc9754 (
      {stage5_28[9]},
      {stage6_28[5]}
   );
   gpc1_1 gpc9755 (
      {stage5_29[12]},
      {stage6_29[3]}
   );
   gpc1_1 gpc9756 (
      {stage5_29[13]},
      {stage6_29[4]}
   );
   gpc1_1 gpc9757 (
      {stage5_29[14]},
      {stage6_29[5]}
   );
   gpc1_1 gpc9758 (
      {stage5_31[8]},
      {stage6_31[4]}
   );
   gpc1_1 gpc9759 (
      {stage5_31[9]},
      {stage6_31[5]}
   );
   gpc1_1 gpc9760 (
      {stage5_32[18]},
      {stage6_32[4]}
   );
   gpc1_1 gpc9761 (
      {stage5_32[19]},
      {stage6_32[5]}
   );
   gpc1_1 gpc9762 (
      {stage5_34[11]},
      {stage6_34[6]}
   );
   gpc1_1 gpc9763 (
      {stage5_34[12]},
      {stage6_34[7]}
   );
   gpc1_1 gpc9764 (
      {stage5_34[13]},
      {stage6_34[8]}
   );
   gpc1_1 gpc9765 (
      {stage5_35[13]},
      {stage6_35[4]}
   );
   gpc1_1 gpc9766 (
      {stage5_36[12]},
      {stage6_36[5]}
   );
   gpc1_1 gpc9767 (
      {stage5_38[9]},
      {stage6_38[4]}
   );
   gpc1_1 gpc9768 (
      {stage5_40[10]},
      {stage6_40[5]}
   );
   gpc1_1 gpc9769 (
      {stage5_41[6]},
      {stage6_41[5]}
   );
   gpc1_1 gpc9770 (
      {stage5_41[7]},
      {stage6_41[6]}
   );
   gpc1_1 gpc9771 (
      {stage5_41[8]},
      {stage6_41[7]}
   );
   gpc1_1 gpc9772 (
      {stage5_42[16]},
      {stage6_42[4]}
   );
   gpc1_1 gpc9773 (
      {stage5_42[17]},
      {stage6_42[5]}
   );
   gpc1_1 gpc9774 (
      {stage5_42[18]},
      {stage6_42[6]}
   );
   gpc1_1 gpc9775 (
      {stage5_43[8]},
      {stage6_43[4]}
   );
   gpc1_1 gpc9776 (
      {stage5_43[9]},
      {stage6_43[5]}
   );
   gpc1_1 gpc9777 (
      {stage5_43[10]},
      {stage6_43[6]}
   );
   gpc1_1 gpc9778 (
      {stage5_44[12]},
      {stage6_44[4]}
   );
   gpc1_1 gpc9779 (
      {stage5_45[12]},
      {stage6_45[6]}
   );
   gpc1_1 gpc9780 (
      {stage5_45[13]},
      {stage6_45[7]}
   );
   gpc1_1 gpc9781 (
      {stage5_45[14]},
      {stage6_45[8]}
   );
   gpc1_1 gpc9782 (
      {stage5_47[8]},
      {stage6_47[3]}
   );
   gpc1_1 gpc9783 (
      {stage5_47[9]},
      {stage6_47[4]}
   );
   gpc1_1 gpc9784 (
      {stage5_47[10]},
      {stage6_47[5]}
   );
   gpc1_1 gpc9785 (
      {stage5_47[11]},
      {stage6_47[6]}
   );
   gpc1_1 gpc9786 (
      {stage5_51[16]},
      {stage6_51[5]}
   );
   gpc1_1 gpc9787 (
      {stage5_51[17]},
      {stage6_51[6]}
   );
   gpc1_1 gpc9788 (
      {stage5_51[18]},
      {stage6_51[7]}
   );
   gpc1_1 gpc9789 (
      {stage5_52[9]},
      {stage6_52[6]}
   );
   gpc1_1 gpc9790 (
      {stage5_55[20]},
      {stage6_55[8]}
   );
   gpc1_1 gpc9791 (
      {stage5_55[21]},
      {stage6_55[9]}
   );
   gpc1_1 gpc9792 (
      {stage5_56[5]},
      {stage6_56[6]}
   );
   gpc1_1 gpc9793 (
      {stage5_56[6]},
      {stage6_56[7]}
   );
   gpc1_1 gpc9794 (
      {stage5_56[7]},
      {stage6_56[8]}
   );
   gpc1_1 gpc9795 (
      {stage5_56[8]},
      {stage6_56[9]}
   );
   gpc1_1 gpc9796 (
      {stage5_57[12]},
      {stage6_57[5]}
   );
   gpc1_1 gpc9797 (
      {stage5_57[13]},
      {stage6_57[6]}
   );
   gpc1_1 gpc9798 (
      {stage5_58[15]},
      {stage6_58[5]}
   );
   gpc1_1 gpc9799 (
      {stage5_61[13]},
      {stage6_61[6]}
   );
   gpc1_1 gpc9800 (
      {stage5_61[14]},
      {stage6_61[7]}
   );
   gpc1_1 gpc9801 (
      {stage5_61[15]},
      {stage6_61[8]}
   );
   gpc1_1 gpc9802 (
      {stage5_63[8]},
      {stage6_63[4]}
   );
   gpc1_1 gpc9803 (
      {stage5_64[12]},
      {stage6_64[6]}
   );
   gpc1_1 gpc9804 (
      {stage5_64[13]},
      {stage6_64[7]}
   );
   gpc1_1 gpc9805 (
      {stage5_64[14]},
      {stage6_64[8]}
   );
   gpc1_1 gpc9806 (
      {stage5_68[1]},
      {stage6_68[4]}
   );
   gpc1_1 gpc9807 (
      {stage5_68[2]},
      {stage6_68[5]}
   );
   gpc1_1 gpc9808 (
      {stage5_68[3]},
      {stage6_68[6]}
   );
   gpc1_1 gpc9809 (
      {stage5_68[4]},
      {stage6_68[7]}
   );
   gpc1_1 gpc9810 (
      {stage5_68[5]},
      {stage6_68[8]}
   );
   gpc1_1 gpc9811 (
      {stage5_68[6]},
      {stage6_68[9]}
   );
   gpc1_1 gpc9812 (
      {stage5_68[7]},
      {stage6_68[10]}
   );
   gpc1_1 gpc9813 (
      {stage5_68[8]},
      {stage6_68[11]}
   );
   gpc1_1 gpc9814 (
      {stage5_68[9]},
      {stage6_68[12]}
   );
   gpc1_1 gpc9815 (
      {stage5_68[10]},
      {stage6_68[13]}
   );
   gpc1_1 gpc9816 (
      {stage5_68[11]},
      {stage6_68[14]}
   );
   gpc1_1 gpc9817 (
      {stage5_68[12]},
      {stage6_68[15]}
   );
   gpc1_1 gpc9818 (
      {stage5_68[13]},
      {stage6_68[16]}
   );
   gpc1_1 gpc9819 (
      {stage5_69[0]},
      {stage6_69[2]}
   );
   gpc1_1 gpc9820 (
      {stage5_69[1]},
      {stage6_69[3]}
   );
   gpc1_1 gpc9821 (
      {stage5_69[2]},
      {stage6_69[4]}
   );
   gpc1_1 gpc9822 (
      {stage5_70[0]},
      {stage6_70[0]}
   );
   gpc1406_5 gpc9823 (
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3], stage6_4[4], stage6_4[5]},
      {stage6_6[0], stage6_6[1], stage6_6[2], stage6_6[3]},
      {stage6_7[0]},
      {stage7_8[0],stage7_7[0],stage7_6[0],stage7_5[0],stage7_4[0]}
   );
   gpc2135_5 gpc9824 (
      {stage6_5[0], stage6_5[1], stage6_5[2], stage6_5[3], 1'b0},
      {stage6_6[4], stage6_6[5], stage6_6[6]},
      {stage6_7[1]},
      {stage6_8[0], stage6_8[1]},
      {stage7_9[0],stage7_8[1],stage7_7[1],stage7_6[1],stage7_5[1]}
   );
   gpc623_5 gpc9825 (
      {stage6_7[2], stage6_7[3], stage6_7[4]},
      {stage6_8[2], stage6_8[3]},
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4], stage6_9[5]},
      {stage7_11[0],stage7_10[0],stage7_9[1],stage7_8[2],stage7_7[2]}
   );
   gpc615_5 gpc9826 (
      {stage6_10[0], stage6_10[1], stage6_10[2], stage6_10[3], stage6_10[4]},
      {stage6_11[0]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage7_14[0],stage7_13[0],stage7_12[0],stage7_11[1],stage7_10[1]}
   );
   gpc615_5 gpc9827 (
      {stage6_11[1], stage6_11[2], stage6_11[3], stage6_11[4], stage6_11[5]},
      {stage6_12[6]},
      {stage6_13[0], stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5]},
      {stage7_15[0],stage7_14[1],stage7_13[1],stage7_12[1],stage7_11[2]}
   );
   gpc7_3 gpc9828 (
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], stage6_14[5], stage6_14[6]},
      {stage7_16[0],stage7_15[1],stage7_14[2]}
   );
   gpc623_5 gpc9829 (
      {stage6_15[0], stage6_15[1], stage6_15[2]},
      {stage6_16[0], stage6_16[1]},
      {stage6_17[0], stage6_17[1], stage6_17[2], stage6_17[3], stage6_17[4], 1'b0},
      {stage7_19[0],stage7_18[0],stage7_17[0],stage7_16[1],stage7_15[2]}
   );
   gpc606_5 gpc9830 (
      {stage6_16[2], stage6_16[3], stage6_16[4], 1'b0, 1'b0, 1'b0},
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage7_20[0],stage7_19[1],stage7_18[1],stage7_17[1],stage7_16[2]}
   );
   gpc15_3 gpc9831 (
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4]},
      {stage6_21[0]},
      {stage7_22[0],stage7_21[0],stage7_20[1]}
   );
   gpc207_4 gpc9832 (
      {stage6_23[0], stage6_23[1], stage6_23[2], stage6_23[3], stage6_23[4], stage6_23[5], stage6_23[6]},
      {stage6_25[0], stage6_25[1]},
      {stage7_26[0],stage7_25[0],stage7_24[0],stage7_23[0]}
   );
   gpc15_3 gpc9833 (
      {stage6_24[0], stage6_24[1], stage6_24[2], stage6_24[3], stage6_24[4]},
      {stage6_25[2]},
      {stage7_26[1],stage7_25[1],stage7_24[1]}
   );
   gpc615_5 gpc9834 (
      {stage6_26[0], stage6_26[1], stage6_26[2], stage6_26[3], stage6_26[4]},
      {stage6_27[0]},
      {stage6_28[0], stage6_28[1], stage6_28[2], stage6_28[3], stage6_28[4], stage6_28[5]},
      {stage7_30[0],stage7_29[0],stage7_28[0],stage7_27[0],stage7_26[2]}
   );
   gpc3_2 gpc9835 (
      {stage6_29[0], stage6_29[1], stage6_29[2]},
      {stage7_30[1],stage7_29[1]}
   );
   gpc615_5 gpc9836 (
      {stage6_31[0], stage6_31[1], stage6_31[2], stage6_31[3], stage6_31[4]},
      {stage6_32[0]},
      {stage6_33[0], stage6_33[1], stage6_33[2], stage6_33[3], stage6_33[4], stage6_33[5]},
      {stage7_35[0],stage7_34[0],stage7_33[0],stage7_32[0],stage7_31[0]}
   );
   gpc615_5 gpc9837 (
      {stage6_34[0], stage6_34[1], stage6_34[2], stage6_34[3], stage6_34[4]},
      {stage6_35[0]},
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3], stage6_36[4], stage6_36[5]},
      {stage7_38[0],stage7_37[0],stage7_36[0],stage7_35[1],stage7_34[1]}
   );
   gpc606_5 gpc9838 (
      {stage6_37[0], stage6_37[1], stage6_37[2], stage6_37[3], stage6_37[4], stage6_37[5]},
      {stage6_39[0], stage6_39[1], stage6_39[2], stage6_39[3], 1'b0, 1'b0},
      {stage7_41[0],stage7_40[0],stage7_39[0],stage7_38[1],stage7_37[1]}
   );
   gpc15_3 gpc9839 (
      {stage6_41[0], stage6_41[1], stage6_41[2], stage6_41[3], stage6_41[4]},
      {stage6_42[0]},
      {stage7_43[0],stage7_42[0],stage7_41[1]}
   );
   gpc615_5 gpc9840 (
      {stage6_42[1], stage6_42[2], stage6_42[3], stage6_42[4], stage6_42[5]},
      {stage6_43[0]},
      {stage6_44[0], stage6_44[1], stage6_44[2], stage6_44[3], stage6_44[4], 1'b0},
      {stage7_46[0],stage7_45[0],stage7_44[0],stage7_43[1],stage7_42[1]}
   );
   gpc615_5 gpc9841 (
      {stage6_43[1], stage6_43[2], stage6_43[3], stage6_43[4], stage6_43[5]},
      {1'b0},
      {stage6_45[0], stage6_45[1], stage6_45[2], stage6_45[3], stage6_45[4], stage6_45[5]},
      {stage7_47[0],stage7_46[1],stage7_45[1],stage7_44[1],stage7_43[2]}
   );
   gpc615_5 gpc9842 (
      {stage6_46[0], stage6_46[1], stage6_46[2], stage6_46[3], stage6_46[4]},
      {stage6_47[0]},
      {stage6_48[0], stage6_48[1], stage6_48[2], stage6_48[3], stage6_48[4], 1'b0},
      {stage7_50[0],stage7_49[0],stage7_48[0],stage7_47[1],stage7_46[2]}
   );
   gpc606_5 gpc9843 (
      {stage6_49[0], stage6_49[1], stage6_49[2], stage6_49[3], stage6_49[4], stage6_49[5]},
      {stage6_51[0], stage6_51[1], stage6_51[2], stage6_51[3], stage6_51[4], stage6_51[5]},
      {stage7_53[0],stage7_52[0],stage7_51[0],stage7_50[1],stage7_49[1]}
   );
   gpc3_2 gpc9844 (
      {stage6_50[0], stage6_50[1], stage6_50[2]},
      {stage7_51[1],stage7_50[2]}
   );
   gpc615_5 gpc9845 (
      {stage6_52[0], stage6_52[1], stage6_52[2], stage6_52[3], stage6_52[4]},
      {stage6_53[0]},
      {stage6_54[0], stage6_54[1], stage6_54[2], stage6_54[3], stage6_54[4], stage6_54[5]},
      {stage7_56[0],stage7_55[0],stage7_54[0],stage7_53[1],stage7_52[1]}
   );
   gpc615_5 gpc9846 (
      {stage6_55[0], stage6_55[1], stage6_55[2], stage6_55[3], stage6_55[4]},
      {stage6_56[0]},
      {stage6_57[0], stage6_57[1], stage6_57[2], stage6_57[3], stage6_57[4], stage6_57[5]},
      {stage7_59[0],stage7_58[0],stage7_57[0],stage7_56[1],stage7_55[1]}
   );
   gpc615_5 gpc9847 (
      {stage6_56[1], stage6_56[2], stage6_56[3], stage6_56[4], stage6_56[5]},
      {stage6_57[6]},
      {stage6_58[0], stage6_58[1], stage6_58[2], stage6_58[3], stage6_58[4], stage6_58[5]},
      {stage7_60[0],stage7_59[1],stage7_58[1],stage7_57[1],stage7_56[2]}
   );
   gpc135_4 gpc9848 (
      {stage6_61[0], stage6_61[1], stage6_61[2], stage6_61[3], stage6_61[4]},
      {stage6_62[0], stage6_62[1], stage6_62[2]},
      {stage6_63[0]},
      {stage7_64[0],stage7_63[0],stage7_62[0],stage7_61[0]}
   );
   gpc135_4 gpc9849 (
      {stage6_61[5], stage6_61[6], stage6_61[7], stage6_61[8], 1'b0},
      {stage6_62[3], stage6_62[4], stage6_62[5]},
      {stage6_63[1]},
      {stage7_64[1],stage7_63[1],stage7_62[1],stage7_61[1]}
   );
   gpc223_4 gpc9850 (
      {stage6_63[2], stage6_63[3], stage6_63[4]},
      {stage6_64[0], stage6_64[1]},
      {stage6_65[0], stage6_65[1]},
      {stage7_66[0],stage7_65[0],stage7_64[2],stage7_63[2]}
   );
   gpc7_3 gpc9851 (
      {stage6_64[2], stage6_64[3], stage6_64[4], stage6_64[5], stage6_64[6], stage6_64[7], stage6_64[8]},
      {stage7_66[1],stage7_65[1],stage7_64[3]}
   );
   gpc3_2 gpc9852 (
      {stage6_65[2], stage6_65[3], stage6_65[4]},
      {stage7_66[2],stage7_65[2]}
   );
   gpc1163_5 gpc9853 (
      {stage6_66[0], stage6_66[1], stage6_66[2]},
      {stage6_67[0], stage6_67[1], stage6_67[2], stage6_67[3], stage6_67[4], 1'b0},
      {stage6_68[0]},
      {stage6_69[0]},
      {stage7_70[0],stage7_69[0],stage7_68[0],stage7_67[0],stage7_66[3]}
   );
   gpc117_4 gpc9854 (
      {stage6_68[1], stage6_68[2], stage6_68[3], stage6_68[4], stage6_68[5], stage6_68[6], stage6_68[7]},
      {stage6_69[1]},
      {stage6_70[0]},
      {stage7_71[0],stage7_70[1],stage7_69[1],stage7_68[1]}
   );
   gpc117_4 gpc9855 (
      {stage6_68[8], stage6_68[9], stage6_68[10], stage6_68[11], stage6_68[12], stage6_68[13], stage6_68[14]},
      {stage6_69[2]},
      {1'b0},
      {stage7_71[1],stage7_70[2],stage7_69[2],stage7_68[2]}
   );
   gpc1_1 gpc9856 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc9857 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc9858 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc9859 (
      {stage6_0[3]},
      {stage7_0[3]}
   );
   gpc1_1 gpc9860 (
      {stage6_0[4]},
      {stage7_0[4]}
   );
   gpc1_1 gpc9861 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc9862 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc9863 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc9864 (
      {stage6_2[1]},
      {stage7_2[1]}
   );
   gpc1_1 gpc9865 (
      {stage6_2[2]},
      {stage7_2[2]}
   );
   gpc1_1 gpc9866 (
      {stage6_2[3]},
      {stage7_2[3]}
   );
   gpc1_1 gpc9867 (
      {stage6_2[4]},
      {stage7_2[4]}
   );
   gpc1_1 gpc9868 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc9869 (
      {stage6_3[1]},
      {stage7_3[1]}
   );
   gpc1_1 gpc9870 (
      {stage6_6[7]},
      {stage7_6[2]}
   );
   gpc1_1 gpc9871 (
      {stage6_8[4]},
      {stage7_8[3]}
   );
   gpc1_1 gpc9872 (
      {stage6_8[5]},
      {stage7_8[4]}
   );
   gpc1_1 gpc9873 (
      {stage6_9[6]},
      {stage7_9[2]}
   );
   gpc1_1 gpc9874 (
      {stage6_9[7]},
      {stage7_9[3]}
   );
   gpc1_1 gpc9875 (
      {stage6_9[8]},
      {stage7_9[4]}
   );
   gpc1_1 gpc9876 (
      {stage6_9[9]},
      {stage7_9[5]}
   );
   gpc1_1 gpc9877 (
      {stage6_11[6]},
      {stage7_11[3]}
   );
   gpc1_1 gpc9878 (
      {stage6_13[6]},
      {stage7_13[2]}
   );
   gpc1_1 gpc9879 (
      {stage6_13[7]},
      {stage7_13[3]}
   );
   gpc1_1 gpc9880 (
      {stage6_13[8]},
      {stage7_13[4]}
   );
   gpc1_1 gpc9881 (
      {stage6_13[9]},
      {stage7_13[5]}
   );
   gpc1_1 gpc9882 (
      {stage6_15[3]},
      {stage7_15[3]}
   );
   gpc1_1 gpc9883 (
      {stage6_15[4]},
      {stage7_15[4]}
   );
   gpc1_1 gpc9884 (
      {stage6_15[5]},
      {stage7_15[5]}
   );
   gpc1_1 gpc9885 (
      {stage6_19[0]},
      {stage7_19[2]}
   );
   gpc1_1 gpc9886 (
      {stage6_19[1]},
      {stage7_19[3]}
   );
   gpc1_1 gpc9887 (
      {stage6_19[2]},
      {stage7_19[4]}
   );
   gpc1_1 gpc9888 (
      {stage6_19[3]},
      {stage7_19[5]}
   );
   gpc1_1 gpc9889 (
      {stage6_19[4]},
      {stage7_19[6]}
   );
   gpc1_1 gpc9890 (
      {stage6_20[5]},
      {stage7_20[2]}
   );
   gpc1_1 gpc9891 (
      {stage6_21[1]},
      {stage7_21[1]}
   );
   gpc1_1 gpc9892 (
      {stage6_21[2]},
      {stage7_21[2]}
   );
   gpc1_1 gpc9893 (
      {stage6_21[3]},
      {stage7_21[3]}
   );
   gpc1_1 gpc9894 (
      {stage6_21[4]},
      {stage7_21[4]}
   );
   gpc1_1 gpc9895 (
      {stage6_21[5]},
      {stage7_21[5]}
   );
   gpc1_1 gpc9896 (
      {stage6_22[0]},
      {stage7_22[1]}
   );
   gpc1_1 gpc9897 (
      {stage6_22[1]},
      {stage7_22[2]}
   );
   gpc1_1 gpc9898 (
      {stage6_22[2]},
      {stage7_22[3]}
   );
   gpc1_1 gpc9899 (
      {stage6_22[3]},
      {stage7_22[4]}
   );
   gpc1_1 gpc9900 (
      {stage6_22[4]},
      {stage7_22[5]}
   );
   gpc1_1 gpc9901 (
      {stage6_22[5]},
      {stage7_22[6]}
   );
   gpc1_1 gpc9902 (
      {stage6_24[5]},
      {stage7_24[2]}
   );
   gpc1_1 gpc9903 (
      {stage6_24[6]},
      {stage7_24[3]}
   );
   gpc1_1 gpc9904 (
      {stage6_26[5]},
      {stage7_26[3]}
   );
   gpc1_1 gpc9905 (
      {stage6_26[6]},
      {stage7_26[4]}
   );
   gpc1_1 gpc9906 (
      {stage6_26[7]},
      {stage7_26[5]}
   );
   gpc1_1 gpc9907 (
      {stage6_27[1]},
      {stage7_27[1]}
   );
   gpc1_1 gpc9908 (
      {stage6_27[2]},
      {stage7_27[2]}
   );
   gpc1_1 gpc9909 (
      {stage6_27[3]},
      {stage7_27[3]}
   );
   gpc1_1 gpc9910 (
      {stage6_27[4]},
      {stage7_27[4]}
   );
   gpc1_1 gpc9911 (
      {stage6_29[3]},
      {stage7_29[2]}
   );
   gpc1_1 gpc9912 (
      {stage6_29[4]},
      {stage7_29[3]}
   );
   gpc1_1 gpc9913 (
      {stage6_29[5]},
      {stage7_29[4]}
   );
   gpc1_1 gpc9914 (
      {stage6_30[0]},
      {stage7_30[2]}
   );
   gpc1_1 gpc9915 (
      {stage6_30[1]},
      {stage7_30[3]}
   );
   gpc1_1 gpc9916 (
      {stage6_30[2]},
      {stage7_30[4]}
   );
   gpc1_1 gpc9917 (
      {stage6_30[3]},
      {stage7_30[5]}
   );
   gpc1_1 gpc9918 (
      {stage6_30[4]},
      {stage7_30[6]}
   );
   gpc1_1 gpc9919 (
      {stage6_31[5]},
      {stage7_31[1]}
   );
   gpc1_1 gpc9920 (
      {stage6_32[1]},
      {stage7_32[1]}
   );
   gpc1_1 gpc9921 (
      {stage6_32[2]},
      {stage7_32[2]}
   );
   gpc1_1 gpc9922 (
      {stage6_32[3]},
      {stage7_32[3]}
   );
   gpc1_1 gpc9923 (
      {stage6_32[4]},
      {stage7_32[4]}
   );
   gpc1_1 gpc9924 (
      {stage6_32[5]},
      {stage7_32[5]}
   );
   gpc1_1 gpc9925 (
      {stage6_34[5]},
      {stage7_34[2]}
   );
   gpc1_1 gpc9926 (
      {stage6_34[6]},
      {stage7_34[3]}
   );
   gpc1_1 gpc9927 (
      {stage6_34[7]},
      {stage7_34[4]}
   );
   gpc1_1 gpc9928 (
      {stage6_34[8]},
      {stage7_34[5]}
   );
   gpc1_1 gpc9929 (
      {stage6_35[1]},
      {stage7_35[2]}
   );
   gpc1_1 gpc9930 (
      {stage6_35[2]},
      {stage7_35[3]}
   );
   gpc1_1 gpc9931 (
      {stage6_35[3]},
      {stage7_35[4]}
   );
   gpc1_1 gpc9932 (
      {stage6_35[4]},
      {stage7_35[5]}
   );
   gpc1_1 gpc9933 (
      {stage6_38[0]},
      {stage7_38[2]}
   );
   gpc1_1 gpc9934 (
      {stage6_38[1]},
      {stage7_38[3]}
   );
   gpc1_1 gpc9935 (
      {stage6_38[2]},
      {stage7_38[4]}
   );
   gpc1_1 gpc9936 (
      {stage6_38[3]},
      {stage7_38[5]}
   );
   gpc1_1 gpc9937 (
      {stage6_38[4]},
      {stage7_38[6]}
   );
   gpc1_1 gpc9938 (
      {stage6_40[0]},
      {stage7_40[1]}
   );
   gpc1_1 gpc9939 (
      {stage6_40[1]},
      {stage7_40[2]}
   );
   gpc1_1 gpc9940 (
      {stage6_40[2]},
      {stage7_40[3]}
   );
   gpc1_1 gpc9941 (
      {stage6_40[3]},
      {stage7_40[4]}
   );
   gpc1_1 gpc9942 (
      {stage6_40[4]},
      {stage7_40[5]}
   );
   gpc1_1 gpc9943 (
      {stage6_40[5]},
      {stage7_40[6]}
   );
   gpc1_1 gpc9944 (
      {stage6_41[5]},
      {stage7_41[2]}
   );
   gpc1_1 gpc9945 (
      {stage6_41[6]},
      {stage7_41[3]}
   );
   gpc1_1 gpc9946 (
      {stage6_41[7]},
      {stage7_41[4]}
   );
   gpc1_1 gpc9947 (
      {stage6_42[6]},
      {stage7_42[2]}
   );
   gpc1_1 gpc9948 (
      {stage6_43[6]},
      {stage7_43[3]}
   );
   gpc1_1 gpc9949 (
      {stage6_45[6]},
      {stage7_45[2]}
   );
   gpc1_1 gpc9950 (
      {stage6_45[7]},
      {stage7_45[3]}
   );
   gpc1_1 gpc9951 (
      {stage6_45[8]},
      {stage7_45[4]}
   );
   gpc1_1 gpc9952 (
      {stage6_47[1]},
      {stage7_47[2]}
   );
   gpc1_1 gpc9953 (
      {stage6_47[2]},
      {stage7_47[3]}
   );
   gpc1_1 gpc9954 (
      {stage6_47[3]},
      {stage7_47[4]}
   );
   gpc1_1 gpc9955 (
      {stage6_47[4]},
      {stage7_47[5]}
   );
   gpc1_1 gpc9956 (
      {stage6_47[5]},
      {stage7_47[6]}
   );
   gpc1_1 gpc9957 (
      {stage6_47[6]},
      {stage7_47[7]}
   );
   gpc1_1 gpc9958 (
      {stage6_51[6]},
      {stage7_51[2]}
   );
   gpc1_1 gpc9959 (
      {stage6_51[7]},
      {stage7_51[3]}
   );
   gpc1_1 gpc9960 (
      {stage6_52[5]},
      {stage7_52[2]}
   );
   gpc1_1 gpc9961 (
      {stage6_52[6]},
      {stage7_52[3]}
   );
   gpc1_1 gpc9962 (
      {stage6_53[1]},
      {stage7_53[2]}
   );
   gpc1_1 gpc9963 (
      {stage6_53[2]},
      {stage7_53[3]}
   );
   gpc1_1 gpc9964 (
      {stage6_53[3]},
      {stage7_53[4]}
   );
   gpc1_1 gpc9965 (
      {stage6_53[4]},
      {stage7_53[5]}
   );
   gpc1_1 gpc9966 (
      {stage6_55[5]},
      {stage7_55[2]}
   );
   gpc1_1 gpc9967 (
      {stage6_55[6]},
      {stage7_55[3]}
   );
   gpc1_1 gpc9968 (
      {stage6_55[7]},
      {stage7_55[4]}
   );
   gpc1_1 gpc9969 (
      {stage6_55[8]},
      {stage7_55[5]}
   );
   gpc1_1 gpc9970 (
      {stage6_55[9]},
      {stage7_55[6]}
   );
   gpc1_1 gpc9971 (
      {stage6_56[6]},
      {stage7_56[3]}
   );
   gpc1_1 gpc9972 (
      {stage6_56[7]},
      {stage7_56[4]}
   );
   gpc1_1 gpc9973 (
      {stage6_56[8]},
      {stage7_56[5]}
   );
   gpc1_1 gpc9974 (
      {stage6_56[9]},
      {stage7_56[6]}
   );
   gpc1_1 gpc9975 (
      {stage6_59[0]},
      {stage7_59[2]}
   );
   gpc1_1 gpc9976 (
      {stage6_59[1]},
      {stage7_59[3]}
   );
   gpc1_1 gpc9977 (
      {stage6_59[2]},
      {stage7_59[4]}
   );
   gpc1_1 gpc9978 (
      {stage6_59[3]},
      {stage7_59[5]}
   );
   gpc1_1 gpc9979 (
      {stage6_59[4]},
      {stage7_59[6]}
   );
   gpc1_1 gpc9980 (
      {stage6_60[0]},
      {stage7_60[1]}
   );
   gpc1_1 gpc9981 (
      {stage6_60[1]},
      {stage7_60[2]}
   );
   gpc1_1 gpc9982 (
      {stage6_60[2]},
      {stage7_60[3]}
   );
   gpc1_1 gpc9983 (
      {stage6_60[3]},
      {stage7_60[4]}
   );
   gpc1_1 gpc9984 (
      {stage6_60[4]},
      {stage7_60[5]}
   );
   gpc1_1 gpc9985 (
      {stage6_66[3]},
      {stage7_66[4]}
   );
   gpc1_1 gpc9986 (
      {stage6_66[4]},
      {stage7_66[5]}
   );
   gpc1_1 gpc9987 (
      {stage6_68[15]},
      {stage7_68[3]}
   );
   gpc1_1 gpc9988 (
      {stage6_68[16]},
      {stage7_68[4]}
   );
   gpc1_1 gpc9989 (
      {stage6_69[3]},
      {stage7_69[3]}
   );
   gpc1_1 gpc9990 (
      {stage6_69[4]},
      {stage7_69[4]}
   );
   gpc1415_5 gpc9991 (
      {stage7_0[0], stage7_0[1], stage7_0[2], stage7_0[3], stage7_0[4]},
      {stage7_1[0]},
      {stage7_2[0], stage7_2[1], stage7_2[2], stage7_2[3]},
      {stage7_3[0]},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc3_2 gpc9992 (
      {stage7_6[0], stage7_6[1], stage7_6[2]},
      {stage8_7[0],stage8_6[0]}
   );
   gpc3_2 gpc9993 (
      {stage7_7[0], stage7_7[1], stage7_7[2]},
      {stage8_8[0],stage8_7[1]}
   );
   gpc215_4 gpc9994 (
      {stage7_8[0], stage7_8[1], stage7_8[2], stage7_8[3], stage7_8[4]},
      {stage7_9[0]},
      {stage7_10[0], stage7_10[1]},
      {stage8_11[0],stage8_10[0],stage8_9[0],stage8_8[1]}
   );
   gpc1415_5 gpc9995 (
      {stage7_9[1], stage7_9[2], stage7_9[3], stage7_9[4], stage7_9[5]},
      {1'b0},
      {stage7_11[0], stage7_11[1], stage7_11[2], stage7_11[3]},
      {stage7_12[0]},
      {stage8_13[0],stage8_12[0],stage8_11[1],stage8_10[1],stage8_9[1]}
   );
   gpc207_4 gpc9996 (
      {stage7_13[0], stage7_13[1], stage7_13[2], stage7_13[3], stage7_13[4], stage7_13[5], 1'b0},
      {stage7_15[0], stage7_15[1]},
      {stage8_16[0],stage8_15[0],stage8_14[0],stage8_13[1]}
   );
   gpc1343_5 gpc9997 (
      {stage7_14[0], stage7_14[1], stage7_14[2]},
      {stage7_15[2], stage7_15[3], stage7_15[4], stage7_15[5]},
      {stage7_16[0], stage7_16[1], stage7_16[2]},
      {stage7_17[0]},
      {stage8_18[0],stage8_17[0],stage8_16[1],stage8_15[1],stage8_14[1]}
   );
   gpc623_5 gpc9998 (
      {stage7_17[1], 1'b0, 1'b0},
      {stage7_18[0], stage7_18[1]},
      {stage7_19[0], stage7_19[1], stage7_19[2], stage7_19[3], stage7_19[4], stage7_19[5]},
      {stage8_21[0],stage8_20[0],stage8_19[0],stage8_18[1],stage8_17[1]}
   );
   gpc1163_5 gpc9999 (
      {stage7_20[0], stage7_20[1], stage7_20[2]},
      {stage7_21[0], stage7_21[1], stage7_21[2], stage7_21[3], stage7_21[4], stage7_21[5]},
      {stage7_22[0]},
      {stage7_23[0]},
      {stage8_24[0],stage8_23[0],stage8_22[0],stage8_21[1],stage8_20[1]}
   );
   gpc1406_5 gpc10000 (
      {stage7_22[1], stage7_22[2], stage7_22[3], stage7_22[4], stage7_22[5], stage7_22[6]},
      {stage7_24[0], stage7_24[1], stage7_24[2], stage7_24[3]},
      {stage7_25[0]},
      {stage8_26[0],stage8_25[0],stage8_24[1],stage8_23[1],stage8_22[1]}
   );
   gpc7_3 gpc10001 (
      {stage7_26[0], stage7_26[1], stage7_26[2], stage7_26[3], stage7_26[4], stage7_26[5], 1'b0},
      {stage8_28[0],stage8_27[0],stage8_26[1]}
   );
   gpc15_3 gpc10002 (
      {stage7_27[0], stage7_27[1], stage7_27[2], stage7_27[3], stage7_27[4]},
      {stage7_28[0]},
      {stage8_29[0],stage8_28[1],stage8_27[1]}
   );
   gpc135_4 gpc10003 (
      {stage7_29[0], stage7_29[1], stage7_29[2], stage7_29[3], stage7_29[4]},
      {stage7_30[0], stage7_30[1], stage7_30[2]},
      {stage7_31[0]},
      {stage8_32[0],stage8_31[0],stage8_30[0],stage8_29[1]}
   );
   gpc615_5 gpc10004 (
      {stage7_30[3], stage7_30[4], stage7_30[5], stage7_30[6], 1'b0},
      {stage7_31[1]},
      {stage7_32[0], stage7_32[1], stage7_32[2], stage7_32[3], stage7_32[4], stage7_32[5]},
      {stage8_34[0],stage8_33[0],stage8_32[1],stage8_31[1],stage8_30[1]}
   );
   gpc7_3 gpc10005 (
      {stage7_34[0], stage7_34[1], stage7_34[2], stage7_34[3], stage7_34[4], stage7_34[5], 1'b0},
      {stage8_36[0],stage8_35[0],stage8_34[1]}
   );
   gpc117_4 gpc10006 (
      {stage7_35[0], stage7_35[1], stage7_35[2], stage7_35[3], stage7_35[4], stage7_35[5], 1'b0},
      {stage7_36[0]},
      {stage7_37[0]},
      {stage8_38[0],stage8_37[0],stage8_36[1],stage8_35[1]}
   );
   gpc7_3 gpc10007 (
      {stage7_38[0], stage7_38[1], stage7_38[2], stage7_38[3], stage7_38[4], stage7_38[5], stage7_38[6]},
      {stage8_40[0],stage8_39[0],stage8_38[1]}
   );
   gpc207_4 gpc10008 (
      {stage7_40[0], stage7_40[1], stage7_40[2], stage7_40[3], stage7_40[4], stage7_40[5], stage7_40[6]},
      {stage7_42[0], stage7_42[1]},
      {stage8_43[0],stage8_42[0],stage8_41[0],stage8_40[1]}
   );
   gpc1415_5 gpc10009 (
      {stage7_41[0], stage7_41[1], stage7_41[2], stage7_41[3], stage7_41[4]},
      {stage7_42[2]},
      {stage7_43[0], stage7_43[1], stage7_43[2], stage7_43[3]},
      {stage7_44[0]},
      {stage8_45[0],stage8_44[0],stage8_43[1],stage8_42[1],stage8_41[1]}
   );
   gpc2135_5 gpc10010 (
      {stage7_45[0], stage7_45[1], stage7_45[2], stage7_45[3], stage7_45[4]},
      {stage7_46[0], stage7_46[1], stage7_46[2]},
      {stage7_47[0]},
      {stage7_48[0], 1'b0},
      {stage8_49[0],stage8_48[0],stage8_47[0],stage8_46[0],stage8_45[1]}
   );
   gpc207_4 gpc10011 (
      {stage7_47[1], stage7_47[2], stage7_47[3], stage7_47[4], stage7_47[5], stage7_47[6], stage7_47[7]},
      {stage7_49[0], stage7_49[1]},
      {stage8_50[0],stage8_49[1],stage8_48[1],stage8_47[1]}
   );
   gpc3_2 gpc10012 (
      {stage7_50[0], stage7_50[1], stage7_50[2]},
      {stage8_51[0],stage8_50[1]}
   );
   gpc615_5 gpc10013 (
      {stage7_51[0], stage7_51[1], stage7_51[2], stage7_51[3], 1'b0},
      {stage7_52[0]},
      {stage7_53[0], stage7_53[1], stage7_53[2], stage7_53[3], stage7_53[4], stage7_53[5]},
      {stage8_55[0],stage8_54[0],stage8_53[0],stage8_52[0],stage8_51[1]}
   );
   gpc3_2 gpc10014 (
      {stage7_52[1], stage7_52[2], stage7_52[3]},
      {stage8_53[1],stage8_52[1]}
   );
   gpc207_4 gpc10015 (
      {stage7_55[0], stage7_55[1], stage7_55[2], stage7_55[3], stage7_55[4], stage7_55[5], stage7_55[6]},
      {stage7_57[0], stage7_57[1]},
      {stage8_58[0],stage8_57[0],stage8_56[0],stage8_55[1]}
   );
   gpc207_4 gpc10016 (
      {stage7_56[0], stage7_56[1], stage7_56[2], stage7_56[3], stage7_56[4], stage7_56[5], stage7_56[6]},
      {stage7_58[0], stage7_58[1]},
      {stage8_59[0],stage8_58[1],stage8_57[1],stage8_56[1]}
   );
   gpc117_4 gpc10017 (
      {stage7_59[0], stage7_59[1], stage7_59[2], stage7_59[3], stage7_59[4], stage7_59[5], stage7_59[6]},
      {stage7_60[0]},
      {stage7_61[0]},
      {stage8_62[0],stage8_61[0],stage8_60[0],stage8_59[1]}
   );
   gpc215_4 gpc10018 (
      {stage7_60[1], stage7_60[2], stage7_60[3], stage7_60[4], stage7_60[5]},
      {stage7_61[1]},
      {stage7_62[0], stage7_62[1]},
      {stage8_63[0],stage8_62[1],stage8_61[1],stage8_60[1]}
   );
   gpc3_2 gpc10019 (
      {stage7_63[0], stage7_63[1], stage7_63[2]},
      {stage8_64[0],stage8_63[1]}
   );
   gpc606_5 gpc10020 (
      {stage7_64[0], stage7_64[1], stage7_64[2], stage7_64[3], 1'b0, 1'b0},
      {stage7_66[0], stage7_66[1], stage7_66[2], stage7_66[3], stage7_66[4], stage7_66[5]},
      {stage8_68[0],stage8_67[0],stage8_66[0],stage8_65[0],stage8_64[1]}
   );
   gpc3_2 gpc10021 (
      {stage7_65[0], stage7_65[1], stage7_65[2]},
      {stage8_66[1],stage8_65[1]}
   );
   gpc615_5 gpc10022 (
      {stage7_68[0], stage7_68[1], stage7_68[2], stage7_68[3], stage7_68[4]},
      {stage7_69[0]},
      {stage7_70[0], stage7_70[1], stage7_70[2], 1'b0, 1'b0, 1'b0},
      {stage8_72[0],stage8_71[0],stage8_70[0],stage8_69[0],stage8_68[1]}
   );
   gpc606_5 gpc10023 (
      {stage7_69[1], stage7_69[2], stage7_69[3], stage7_69[4], 1'b0, 1'b0},
      {stage7_71[0], stage7_71[1], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage8_72[1],stage8_71[1],stage8_70[1],stage8_69[1]}
   );
   gpc1_1 gpc10024 (
      {stage7_1[1]},
      {stage8_1[1]}
   );
   gpc1_1 gpc10025 (
      {stage7_2[4]},
      {stage8_2[1]}
   );
   gpc1_1 gpc10026 (
      {stage7_3[1]},
      {stage8_3[1]}
   );
   gpc1_1 gpc10027 (
      {stage7_4[0]},
      {stage8_4[1]}
   );
   gpc1_1 gpc10028 (
      {stage7_5[0]},
      {stage8_5[0]}
   );
   gpc1_1 gpc10029 (
      {stage7_5[1]},
      {stage8_5[1]}
   );
   gpc1_1 gpc10030 (
      {stage7_12[1]},
      {stage8_12[1]}
   );
   gpc1_1 gpc10031 (
      {stage7_19[6]},
      {stage8_19[1]}
   );
   gpc1_1 gpc10032 (
      {stage7_25[1]},
      {stage8_25[1]}
   );
   gpc1_1 gpc10033 (
      {stage7_33[0]},
      {stage8_33[1]}
   );
   gpc1_1 gpc10034 (
      {stage7_37[1]},
      {stage8_37[1]}
   );
   gpc1_1 gpc10035 (
      {stage7_39[0]},
      {stage8_39[1]}
   );
   gpc1_1 gpc10036 (
      {stage7_44[1]},
      {stage8_44[1]}
   );
   gpc1_1 gpc10037 (
      {stage7_54[0]},
      {stage8_54[1]}
   );
   gpc1_1 gpc10038 (
      {stage7_67[0]},
      {stage8_67[1]}
   );
endmodule

module testbench();
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    reg [485:0] src16;
    reg [485:0] src17;
    reg [485:0] src18;
    reg [485:0] src19;
    reg [485:0] src20;
    reg [485:0] src21;
    reg [485:0] src22;
    reg [485:0] src23;
    reg [485:0] src24;
    reg [485:0] src25;
    reg [485:0] src26;
    reg [485:0] src27;
    reg [485:0] src28;
    reg [485:0] src29;
    reg [485:0] src30;
    reg [485:0] src31;
    reg [485:0] src32;
    reg [485:0] src33;
    reg [485:0] src34;
    reg [485:0] src35;
    reg [485:0] src36;
    reg [485:0] src37;
    reg [485:0] src38;
    reg [485:0] src39;
    reg [485:0] src40;
    reg [485:0] src41;
    reg [485:0] src42;
    reg [485:0] src43;
    reg [485:0] src44;
    reg [485:0] src45;
    reg [485:0] src46;
    reg [485:0] src47;
    reg [485:0] src48;
    reg [485:0] src49;
    reg [485:0] src50;
    reg [485:0] src51;
    reg [485:0] src52;
    reg [485:0] src53;
    reg [485:0] src54;
    reg [485:0] src55;
    reg [485:0] src56;
    reg [485:0] src57;
    reg [485:0] src58;
    reg [485:0] src59;
    reg [485:0] src60;
    reg [485:0] src61;
    reg [485:0] src62;
    reg [485:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [0:0] dst70;
    wire [0:0] dst71;
    wire [0:0] dst72;
    wire [72:0] srcsum;
    wire [72:0] dstsum;
    wire test;
    compressor_CLA486_64 compressor_CLA486_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69),
        .dst70(dst70),
        .dst71(dst71),
        .dst72(dst72));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255] + src16[256] + src16[257] + src16[258] + src16[259] + src16[260] + src16[261] + src16[262] + src16[263] + src16[264] + src16[265] + src16[266] + src16[267] + src16[268] + src16[269] + src16[270] + src16[271] + src16[272] + src16[273] + src16[274] + src16[275] + src16[276] + src16[277] + src16[278] + src16[279] + src16[280] + src16[281] + src16[282] + src16[283] + src16[284] + src16[285] + src16[286] + src16[287] + src16[288] + src16[289] + src16[290] + src16[291] + src16[292] + src16[293] + src16[294] + src16[295] + src16[296] + src16[297] + src16[298] + src16[299] + src16[300] + src16[301] + src16[302] + src16[303] + src16[304] + src16[305] + src16[306] + src16[307] + src16[308] + src16[309] + src16[310] + src16[311] + src16[312] + src16[313] + src16[314] + src16[315] + src16[316] + src16[317] + src16[318] + src16[319] + src16[320] + src16[321] + src16[322] + src16[323] + src16[324] + src16[325] + src16[326] + src16[327] + src16[328] + src16[329] + src16[330] + src16[331] + src16[332] + src16[333] + src16[334] + src16[335] + src16[336] + src16[337] + src16[338] + src16[339] + src16[340] + src16[341] + src16[342] + src16[343] + src16[344] + src16[345] + src16[346] + src16[347] + src16[348] + src16[349] + src16[350] + src16[351] + src16[352] + src16[353] + src16[354] + src16[355] + src16[356] + src16[357] + src16[358] + src16[359] + src16[360] + src16[361] + src16[362] + src16[363] + src16[364] + src16[365] + src16[366] + src16[367] + src16[368] + src16[369] + src16[370] + src16[371] + src16[372] + src16[373] + src16[374] + src16[375] + src16[376] + src16[377] + src16[378] + src16[379] + src16[380] + src16[381] + src16[382] + src16[383] + src16[384] + src16[385] + src16[386] + src16[387] + src16[388] + src16[389] + src16[390] + src16[391] + src16[392] + src16[393] + src16[394] + src16[395] + src16[396] + src16[397] + src16[398] + src16[399] + src16[400] + src16[401] + src16[402] + src16[403] + src16[404] + src16[405] + src16[406] + src16[407] + src16[408] + src16[409] + src16[410] + src16[411] + src16[412] + src16[413] + src16[414] + src16[415] + src16[416] + src16[417] + src16[418] + src16[419] + src16[420] + src16[421] + src16[422] + src16[423] + src16[424] + src16[425] + src16[426] + src16[427] + src16[428] + src16[429] + src16[430] + src16[431] + src16[432] + src16[433] + src16[434] + src16[435] + src16[436] + src16[437] + src16[438] + src16[439] + src16[440] + src16[441] + src16[442] + src16[443] + src16[444] + src16[445] + src16[446] + src16[447] + src16[448] + src16[449] + src16[450] + src16[451] + src16[452] + src16[453] + src16[454] + src16[455] + src16[456] + src16[457] + src16[458] + src16[459] + src16[460] + src16[461] + src16[462] + src16[463] + src16[464] + src16[465] + src16[466] + src16[467] + src16[468] + src16[469] + src16[470] + src16[471] + src16[472] + src16[473] + src16[474] + src16[475] + src16[476] + src16[477] + src16[478] + src16[479] + src16[480] + src16[481] + src16[482] + src16[483] + src16[484] + src16[485])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255] + src17[256] + src17[257] + src17[258] + src17[259] + src17[260] + src17[261] + src17[262] + src17[263] + src17[264] + src17[265] + src17[266] + src17[267] + src17[268] + src17[269] + src17[270] + src17[271] + src17[272] + src17[273] + src17[274] + src17[275] + src17[276] + src17[277] + src17[278] + src17[279] + src17[280] + src17[281] + src17[282] + src17[283] + src17[284] + src17[285] + src17[286] + src17[287] + src17[288] + src17[289] + src17[290] + src17[291] + src17[292] + src17[293] + src17[294] + src17[295] + src17[296] + src17[297] + src17[298] + src17[299] + src17[300] + src17[301] + src17[302] + src17[303] + src17[304] + src17[305] + src17[306] + src17[307] + src17[308] + src17[309] + src17[310] + src17[311] + src17[312] + src17[313] + src17[314] + src17[315] + src17[316] + src17[317] + src17[318] + src17[319] + src17[320] + src17[321] + src17[322] + src17[323] + src17[324] + src17[325] + src17[326] + src17[327] + src17[328] + src17[329] + src17[330] + src17[331] + src17[332] + src17[333] + src17[334] + src17[335] + src17[336] + src17[337] + src17[338] + src17[339] + src17[340] + src17[341] + src17[342] + src17[343] + src17[344] + src17[345] + src17[346] + src17[347] + src17[348] + src17[349] + src17[350] + src17[351] + src17[352] + src17[353] + src17[354] + src17[355] + src17[356] + src17[357] + src17[358] + src17[359] + src17[360] + src17[361] + src17[362] + src17[363] + src17[364] + src17[365] + src17[366] + src17[367] + src17[368] + src17[369] + src17[370] + src17[371] + src17[372] + src17[373] + src17[374] + src17[375] + src17[376] + src17[377] + src17[378] + src17[379] + src17[380] + src17[381] + src17[382] + src17[383] + src17[384] + src17[385] + src17[386] + src17[387] + src17[388] + src17[389] + src17[390] + src17[391] + src17[392] + src17[393] + src17[394] + src17[395] + src17[396] + src17[397] + src17[398] + src17[399] + src17[400] + src17[401] + src17[402] + src17[403] + src17[404] + src17[405] + src17[406] + src17[407] + src17[408] + src17[409] + src17[410] + src17[411] + src17[412] + src17[413] + src17[414] + src17[415] + src17[416] + src17[417] + src17[418] + src17[419] + src17[420] + src17[421] + src17[422] + src17[423] + src17[424] + src17[425] + src17[426] + src17[427] + src17[428] + src17[429] + src17[430] + src17[431] + src17[432] + src17[433] + src17[434] + src17[435] + src17[436] + src17[437] + src17[438] + src17[439] + src17[440] + src17[441] + src17[442] + src17[443] + src17[444] + src17[445] + src17[446] + src17[447] + src17[448] + src17[449] + src17[450] + src17[451] + src17[452] + src17[453] + src17[454] + src17[455] + src17[456] + src17[457] + src17[458] + src17[459] + src17[460] + src17[461] + src17[462] + src17[463] + src17[464] + src17[465] + src17[466] + src17[467] + src17[468] + src17[469] + src17[470] + src17[471] + src17[472] + src17[473] + src17[474] + src17[475] + src17[476] + src17[477] + src17[478] + src17[479] + src17[480] + src17[481] + src17[482] + src17[483] + src17[484] + src17[485])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255] + src18[256] + src18[257] + src18[258] + src18[259] + src18[260] + src18[261] + src18[262] + src18[263] + src18[264] + src18[265] + src18[266] + src18[267] + src18[268] + src18[269] + src18[270] + src18[271] + src18[272] + src18[273] + src18[274] + src18[275] + src18[276] + src18[277] + src18[278] + src18[279] + src18[280] + src18[281] + src18[282] + src18[283] + src18[284] + src18[285] + src18[286] + src18[287] + src18[288] + src18[289] + src18[290] + src18[291] + src18[292] + src18[293] + src18[294] + src18[295] + src18[296] + src18[297] + src18[298] + src18[299] + src18[300] + src18[301] + src18[302] + src18[303] + src18[304] + src18[305] + src18[306] + src18[307] + src18[308] + src18[309] + src18[310] + src18[311] + src18[312] + src18[313] + src18[314] + src18[315] + src18[316] + src18[317] + src18[318] + src18[319] + src18[320] + src18[321] + src18[322] + src18[323] + src18[324] + src18[325] + src18[326] + src18[327] + src18[328] + src18[329] + src18[330] + src18[331] + src18[332] + src18[333] + src18[334] + src18[335] + src18[336] + src18[337] + src18[338] + src18[339] + src18[340] + src18[341] + src18[342] + src18[343] + src18[344] + src18[345] + src18[346] + src18[347] + src18[348] + src18[349] + src18[350] + src18[351] + src18[352] + src18[353] + src18[354] + src18[355] + src18[356] + src18[357] + src18[358] + src18[359] + src18[360] + src18[361] + src18[362] + src18[363] + src18[364] + src18[365] + src18[366] + src18[367] + src18[368] + src18[369] + src18[370] + src18[371] + src18[372] + src18[373] + src18[374] + src18[375] + src18[376] + src18[377] + src18[378] + src18[379] + src18[380] + src18[381] + src18[382] + src18[383] + src18[384] + src18[385] + src18[386] + src18[387] + src18[388] + src18[389] + src18[390] + src18[391] + src18[392] + src18[393] + src18[394] + src18[395] + src18[396] + src18[397] + src18[398] + src18[399] + src18[400] + src18[401] + src18[402] + src18[403] + src18[404] + src18[405] + src18[406] + src18[407] + src18[408] + src18[409] + src18[410] + src18[411] + src18[412] + src18[413] + src18[414] + src18[415] + src18[416] + src18[417] + src18[418] + src18[419] + src18[420] + src18[421] + src18[422] + src18[423] + src18[424] + src18[425] + src18[426] + src18[427] + src18[428] + src18[429] + src18[430] + src18[431] + src18[432] + src18[433] + src18[434] + src18[435] + src18[436] + src18[437] + src18[438] + src18[439] + src18[440] + src18[441] + src18[442] + src18[443] + src18[444] + src18[445] + src18[446] + src18[447] + src18[448] + src18[449] + src18[450] + src18[451] + src18[452] + src18[453] + src18[454] + src18[455] + src18[456] + src18[457] + src18[458] + src18[459] + src18[460] + src18[461] + src18[462] + src18[463] + src18[464] + src18[465] + src18[466] + src18[467] + src18[468] + src18[469] + src18[470] + src18[471] + src18[472] + src18[473] + src18[474] + src18[475] + src18[476] + src18[477] + src18[478] + src18[479] + src18[480] + src18[481] + src18[482] + src18[483] + src18[484] + src18[485])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255] + src19[256] + src19[257] + src19[258] + src19[259] + src19[260] + src19[261] + src19[262] + src19[263] + src19[264] + src19[265] + src19[266] + src19[267] + src19[268] + src19[269] + src19[270] + src19[271] + src19[272] + src19[273] + src19[274] + src19[275] + src19[276] + src19[277] + src19[278] + src19[279] + src19[280] + src19[281] + src19[282] + src19[283] + src19[284] + src19[285] + src19[286] + src19[287] + src19[288] + src19[289] + src19[290] + src19[291] + src19[292] + src19[293] + src19[294] + src19[295] + src19[296] + src19[297] + src19[298] + src19[299] + src19[300] + src19[301] + src19[302] + src19[303] + src19[304] + src19[305] + src19[306] + src19[307] + src19[308] + src19[309] + src19[310] + src19[311] + src19[312] + src19[313] + src19[314] + src19[315] + src19[316] + src19[317] + src19[318] + src19[319] + src19[320] + src19[321] + src19[322] + src19[323] + src19[324] + src19[325] + src19[326] + src19[327] + src19[328] + src19[329] + src19[330] + src19[331] + src19[332] + src19[333] + src19[334] + src19[335] + src19[336] + src19[337] + src19[338] + src19[339] + src19[340] + src19[341] + src19[342] + src19[343] + src19[344] + src19[345] + src19[346] + src19[347] + src19[348] + src19[349] + src19[350] + src19[351] + src19[352] + src19[353] + src19[354] + src19[355] + src19[356] + src19[357] + src19[358] + src19[359] + src19[360] + src19[361] + src19[362] + src19[363] + src19[364] + src19[365] + src19[366] + src19[367] + src19[368] + src19[369] + src19[370] + src19[371] + src19[372] + src19[373] + src19[374] + src19[375] + src19[376] + src19[377] + src19[378] + src19[379] + src19[380] + src19[381] + src19[382] + src19[383] + src19[384] + src19[385] + src19[386] + src19[387] + src19[388] + src19[389] + src19[390] + src19[391] + src19[392] + src19[393] + src19[394] + src19[395] + src19[396] + src19[397] + src19[398] + src19[399] + src19[400] + src19[401] + src19[402] + src19[403] + src19[404] + src19[405] + src19[406] + src19[407] + src19[408] + src19[409] + src19[410] + src19[411] + src19[412] + src19[413] + src19[414] + src19[415] + src19[416] + src19[417] + src19[418] + src19[419] + src19[420] + src19[421] + src19[422] + src19[423] + src19[424] + src19[425] + src19[426] + src19[427] + src19[428] + src19[429] + src19[430] + src19[431] + src19[432] + src19[433] + src19[434] + src19[435] + src19[436] + src19[437] + src19[438] + src19[439] + src19[440] + src19[441] + src19[442] + src19[443] + src19[444] + src19[445] + src19[446] + src19[447] + src19[448] + src19[449] + src19[450] + src19[451] + src19[452] + src19[453] + src19[454] + src19[455] + src19[456] + src19[457] + src19[458] + src19[459] + src19[460] + src19[461] + src19[462] + src19[463] + src19[464] + src19[465] + src19[466] + src19[467] + src19[468] + src19[469] + src19[470] + src19[471] + src19[472] + src19[473] + src19[474] + src19[475] + src19[476] + src19[477] + src19[478] + src19[479] + src19[480] + src19[481] + src19[482] + src19[483] + src19[484] + src19[485])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255] + src20[256] + src20[257] + src20[258] + src20[259] + src20[260] + src20[261] + src20[262] + src20[263] + src20[264] + src20[265] + src20[266] + src20[267] + src20[268] + src20[269] + src20[270] + src20[271] + src20[272] + src20[273] + src20[274] + src20[275] + src20[276] + src20[277] + src20[278] + src20[279] + src20[280] + src20[281] + src20[282] + src20[283] + src20[284] + src20[285] + src20[286] + src20[287] + src20[288] + src20[289] + src20[290] + src20[291] + src20[292] + src20[293] + src20[294] + src20[295] + src20[296] + src20[297] + src20[298] + src20[299] + src20[300] + src20[301] + src20[302] + src20[303] + src20[304] + src20[305] + src20[306] + src20[307] + src20[308] + src20[309] + src20[310] + src20[311] + src20[312] + src20[313] + src20[314] + src20[315] + src20[316] + src20[317] + src20[318] + src20[319] + src20[320] + src20[321] + src20[322] + src20[323] + src20[324] + src20[325] + src20[326] + src20[327] + src20[328] + src20[329] + src20[330] + src20[331] + src20[332] + src20[333] + src20[334] + src20[335] + src20[336] + src20[337] + src20[338] + src20[339] + src20[340] + src20[341] + src20[342] + src20[343] + src20[344] + src20[345] + src20[346] + src20[347] + src20[348] + src20[349] + src20[350] + src20[351] + src20[352] + src20[353] + src20[354] + src20[355] + src20[356] + src20[357] + src20[358] + src20[359] + src20[360] + src20[361] + src20[362] + src20[363] + src20[364] + src20[365] + src20[366] + src20[367] + src20[368] + src20[369] + src20[370] + src20[371] + src20[372] + src20[373] + src20[374] + src20[375] + src20[376] + src20[377] + src20[378] + src20[379] + src20[380] + src20[381] + src20[382] + src20[383] + src20[384] + src20[385] + src20[386] + src20[387] + src20[388] + src20[389] + src20[390] + src20[391] + src20[392] + src20[393] + src20[394] + src20[395] + src20[396] + src20[397] + src20[398] + src20[399] + src20[400] + src20[401] + src20[402] + src20[403] + src20[404] + src20[405] + src20[406] + src20[407] + src20[408] + src20[409] + src20[410] + src20[411] + src20[412] + src20[413] + src20[414] + src20[415] + src20[416] + src20[417] + src20[418] + src20[419] + src20[420] + src20[421] + src20[422] + src20[423] + src20[424] + src20[425] + src20[426] + src20[427] + src20[428] + src20[429] + src20[430] + src20[431] + src20[432] + src20[433] + src20[434] + src20[435] + src20[436] + src20[437] + src20[438] + src20[439] + src20[440] + src20[441] + src20[442] + src20[443] + src20[444] + src20[445] + src20[446] + src20[447] + src20[448] + src20[449] + src20[450] + src20[451] + src20[452] + src20[453] + src20[454] + src20[455] + src20[456] + src20[457] + src20[458] + src20[459] + src20[460] + src20[461] + src20[462] + src20[463] + src20[464] + src20[465] + src20[466] + src20[467] + src20[468] + src20[469] + src20[470] + src20[471] + src20[472] + src20[473] + src20[474] + src20[475] + src20[476] + src20[477] + src20[478] + src20[479] + src20[480] + src20[481] + src20[482] + src20[483] + src20[484] + src20[485])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255] + src21[256] + src21[257] + src21[258] + src21[259] + src21[260] + src21[261] + src21[262] + src21[263] + src21[264] + src21[265] + src21[266] + src21[267] + src21[268] + src21[269] + src21[270] + src21[271] + src21[272] + src21[273] + src21[274] + src21[275] + src21[276] + src21[277] + src21[278] + src21[279] + src21[280] + src21[281] + src21[282] + src21[283] + src21[284] + src21[285] + src21[286] + src21[287] + src21[288] + src21[289] + src21[290] + src21[291] + src21[292] + src21[293] + src21[294] + src21[295] + src21[296] + src21[297] + src21[298] + src21[299] + src21[300] + src21[301] + src21[302] + src21[303] + src21[304] + src21[305] + src21[306] + src21[307] + src21[308] + src21[309] + src21[310] + src21[311] + src21[312] + src21[313] + src21[314] + src21[315] + src21[316] + src21[317] + src21[318] + src21[319] + src21[320] + src21[321] + src21[322] + src21[323] + src21[324] + src21[325] + src21[326] + src21[327] + src21[328] + src21[329] + src21[330] + src21[331] + src21[332] + src21[333] + src21[334] + src21[335] + src21[336] + src21[337] + src21[338] + src21[339] + src21[340] + src21[341] + src21[342] + src21[343] + src21[344] + src21[345] + src21[346] + src21[347] + src21[348] + src21[349] + src21[350] + src21[351] + src21[352] + src21[353] + src21[354] + src21[355] + src21[356] + src21[357] + src21[358] + src21[359] + src21[360] + src21[361] + src21[362] + src21[363] + src21[364] + src21[365] + src21[366] + src21[367] + src21[368] + src21[369] + src21[370] + src21[371] + src21[372] + src21[373] + src21[374] + src21[375] + src21[376] + src21[377] + src21[378] + src21[379] + src21[380] + src21[381] + src21[382] + src21[383] + src21[384] + src21[385] + src21[386] + src21[387] + src21[388] + src21[389] + src21[390] + src21[391] + src21[392] + src21[393] + src21[394] + src21[395] + src21[396] + src21[397] + src21[398] + src21[399] + src21[400] + src21[401] + src21[402] + src21[403] + src21[404] + src21[405] + src21[406] + src21[407] + src21[408] + src21[409] + src21[410] + src21[411] + src21[412] + src21[413] + src21[414] + src21[415] + src21[416] + src21[417] + src21[418] + src21[419] + src21[420] + src21[421] + src21[422] + src21[423] + src21[424] + src21[425] + src21[426] + src21[427] + src21[428] + src21[429] + src21[430] + src21[431] + src21[432] + src21[433] + src21[434] + src21[435] + src21[436] + src21[437] + src21[438] + src21[439] + src21[440] + src21[441] + src21[442] + src21[443] + src21[444] + src21[445] + src21[446] + src21[447] + src21[448] + src21[449] + src21[450] + src21[451] + src21[452] + src21[453] + src21[454] + src21[455] + src21[456] + src21[457] + src21[458] + src21[459] + src21[460] + src21[461] + src21[462] + src21[463] + src21[464] + src21[465] + src21[466] + src21[467] + src21[468] + src21[469] + src21[470] + src21[471] + src21[472] + src21[473] + src21[474] + src21[475] + src21[476] + src21[477] + src21[478] + src21[479] + src21[480] + src21[481] + src21[482] + src21[483] + src21[484] + src21[485])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255] + src22[256] + src22[257] + src22[258] + src22[259] + src22[260] + src22[261] + src22[262] + src22[263] + src22[264] + src22[265] + src22[266] + src22[267] + src22[268] + src22[269] + src22[270] + src22[271] + src22[272] + src22[273] + src22[274] + src22[275] + src22[276] + src22[277] + src22[278] + src22[279] + src22[280] + src22[281] + src22[282] + src22[283] + src22[284] + src22[285] + src22[286] + src22[287] + src22[288] + src22[289] + src22[290] + src22[291] + src22[292] + src22[293] + src22[294] + src22[295] + src22[296] + src22[297] + src22[298] + src22[299] + src22[300] + src22[301] + src22[302] + src22[303] + src22[304] + src22[305] + src22[306] + src22[307] + src22[308] + src22[309] + src22[310] + src22[311] + src22[312] + src22[313] + src22[314] + src22[315] + src22[316] + src22[317] + src22[318] + src22[319] + src22[320] + src22[321] + src22[322] + src22[323] + src22[324] + src22[325] + src22[326] + src22[327] + src22[328] + src22[329] + src22[330] + src22[331] + src22[332] + src22[333] + src22[334] + src22[335] + src22[336] + src22[337] + src22[338] + src22[339] + src22[340] + src22[341] + src22[342] + src22[343] + src22[344] + src22[345] + src22[346] + src22[347] + src22[348] + src22[349] + src22[350] + src22[351] + src22[352] + src22[353] + src22[354] + src22[355] + src22[356] + src22[357] + src22[358] + src22[359] + src22[360] + src22[361] + src22[362] + src22[363] + src22[364] + src22[365] + src22[366] + src22[367] + src22[368] + src22[369] + src22[370] + src22[371] + src22[372] + src22[373] + src22[374] + src22[375] + src22[376] + src22[377] + src22[378] + src22[379] + src22[380] + src22[381] + src22[382] + src22[383] + src22[384] + src22[385] + src22[386] + src22[387] + src22[388] + src22[389] + src22[390] + src22[391] + src22[392] + src22[393] + src22[394] + src22[395] + src22[396] + src22[397] + src22[398] + src22[399] + src22[400] + src22[401] + src22[402] + src22[403] + src22[404] + src22[405] + src22[406] + src22[407] + src22[408] + src22[409] + src22[410] + src22[411] + src22[412] + src22[413] + src22[414] + src22[415] + src22[416] + src22[417] + src22[418] + src22[419] + src22[420] + src22[421] + src22[422] + src22[423] + src22[424] + src22[425] + src22[426] + src22[427] + src22[428] + src22[429] + src22[430] + src22[431] + src22[432] + src22[433] + src22[434] + src22[435] + src22[436] + src22[437] + src22[438] + src22[439] + src22[440] + src22[441] + src22[442] + src22[443] + src22[444] + src22[445] + src22[446] + src22[447] + src22[448] + src22[449] + src22[450] + src22[451] + src22[452] + src22[453] + src22[454] + src22[455] + src22[456] + src22[457] + src22[458] + src22[459] + src22[460] + src22[461] + src22[462] + src22[463] + src22[464] + src22[465] + src22[466] + src22[467] + src22[468] + src22[469] + src22[470] + src22[471] + src22[472] + src22[473] + src22[474] + src22[475] + src22[476] + src22[477] + src22[478] + src22[479] + src22[480] + src22[481] + src22[482] + src22[483] + src22[484] + src22[485])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255] + src23[256] + src23[257] + src23[258] + src23[259] + src23[260] + src23[261] + src23[262] + src23[263] + src23[264] + src23[265] + src23[266] + src23[267] + src23[268] + src23[269] + src23[270] + src23[271] + src23[272] + src23[273] + src23[274] + src23[275] + src23[276] + src23[277] + src23[278] + src23[279] + src23[280] + src23[281] + src23[282] + src23[283] + src23[284] + src23[285] + src23[286] + src23[287] + src23[288] + src23[289] + src23[290] + src23[291] + src23[292] + src23[293] + src23[294] + src23[295] + src23[296] + src23[297] + src23[298] + src23[299] + src23[300] + src23[301] + src23[302] + src23[303] + src23[304] + src23[305] + src23[306] + src23[307] + src23[308] + src23[309] + src23[310] + src23[311] + src23[312] + src23[313] + src23[314] + src23[315] + src23[316] + src23[317] + src23[318] + src23[319] + src23[320] + src23[321] + src23[322] + src23[323] + src23[324] + src23[325] + src23[326] + src23[327] + src23[328] + src23[329] + src23[330] + src23[331] + src23[332] + src23[333] + src23[334] + src23[335] + src23[336] + src23[337] + src23[338] + src23[339] + src23[340] + src23[341] + src23[342] + src23[343] + src23[344] + src23[345] + src23[346] + src23[347] + src23[348] + src23[349] + src23[350] + src23[351] + src23[352] + src23[353] + src23[354] + src23[355] + src23[356] + src23[357] + src23[358] + src23[359] + src23[360] + src23[361] + src23[362] + src23[363] + src23[364] + src23[365] + src23[366] + src23[367] + src23[368] + src23[369] + src23[370] + src23[371] + src23[372] + src23[373] + src23[374] + src23[375] + src23[376] + src23[377] + src23[378] + src23[379] + src23[380] + src23[381] + src23[382] + src23[383] + src23[384] + src23[385] + src23[386] + src23[387] + src23[388] + src23[389] + src23[390] + src23[391] + src23[392] + src23[393] + src23[394] + src23[395] + src23[396] + src23[397] + src23[398] + src23[399] + src23[400] + src23[401] + src23[402] + src23[403] + src23[404] + src23[405] + src23[406] + src23[407] + src23[408] + src23[409] + src23[410] + src23[411] + src23[412] + src23[413] + src23[414] + src23[415] + src23[416] + src23[417] + src23[418] + src23[419] + src23[420] + src23[421] + src23[422] + src23[423] + src23[424] + src23[425] + src23[426] + src23[427] + src23[428] + src23[429] + src23[430] + src23[431] + src23[432] + src23[433] + src23[434] + src23[435] + src23[436] + src23[437] + src23[438] + src23[439] + src23[440] + src23[441] + src23[442] + src23[443] + src23[444] + src23[445] + src23[446] + src23[447] + src23[448] + src23[449] + src23[450] + src23[451] + src23[452] + src23[453] + src23[454] + src23[455] + src23[456] + src23[457] + src23[458] + src23[459] + src23[460] + src23[461] + src23[462] + src23[463] + src23[464] + src23[465] + src23[466] + src23[467] + src23[468] + src23[469] + src23[470] + src23[471] + src23[472] + src23[473] + src23[474] + src23[475] + src23[476] + src23[477] + src23[478] + src23[479] + src23[480] + src23[481] + src23[482] + src23[483] + src23[484] + src23[485])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255] + src24[256] + src24[257] + src24[258] + src24[259] + src24[260] + src24[261] + src24[262] + src24[263] + src24[264] + src24[265] + src24[266] + src24[267] + src24[268] + src24[269] + src24[270] + src24[271] + src24[272] + src24[273] + src24[274] + src24[275] + src24[276] + src24[277] + src24[278] + src24[279] + src24[280] + src24[281] + src24[282] + src24[283] + src24[284] + src24[285] + src24[286] + src24[287] + src24[288] + src24[289] + src24[290] + src24[291] + src24[292] + src24[293] + src24[294] + src24[295] + src24[296] + src24[297] + src24[298] + src24[299] + src24[300] + src24[301] + src24[302] + src24[303] + src24[304] + src24[305] + src24[306] + src24[307] + src24[308] + src24[309] + src24[310] + src24[311] + src24[312] + src24[313] + src24[314] + src24[315] + src24[316] + src24[317] + src24[318] + src24[319] + src24[320] + src24[321] + src24[322] + src24[323] + src24[324] + src24[325] + src24[326] + src24[327] + src24[328] + src24[329] + src24[330] + src24[331] + src24[332] + src24[333] + src24[334] + src24[335] + src24[336] + src24[337] + src24[338] + src24[339] + src24[340] + src24[341] + src24[342] + src24[343] + src24[344] + src24[345] + src24[346] + src24[347] + src24[348] + src24[349] + src24[350] + src24[351] + src24[352] + src24[353] + src24[354] + src24[355] + src24[356] + src24[357] + src24[358] + src24[359] + src24[360] + src24[361] + src24[362] + src24[363] + src24[364] + src24[365] + src24[366] + src24[367] + src24[368] + src24[369] + src24[370] + src24[371] + src24[372] + src24[373] + src24[374] + src24[375] + src24[376] + src24[377] + src24[378] + src24[379] + src24[380] + src24[381] + src24[382] + src24[383] + src24[384] + src24[385] + src24[386] + src24[387] + src24[388] + src24[389] + src24[390] + src24[391] + src24[392] + src24[393] + src24[394] + src24[395] + src24[396] + src24[397] + src24[398] + src24[399] + src24[400] + src24[401] + src24[402] + src24[403] + src24[404] + src24[405] + src24[406] + src24[407] + src24[408] + src24[409] + src24[410] + src24[411] + src24[412] + src24[413] + src24[414] + src24[415] + src24[416] + src24[417] + src24[418] + src24[419] + src24[420] + src24[421] + src24[422] + src24[423] + src24[424] + src24[425] + src24[426] + src24[427] + src24[428] + src24[429] + src24[430] + src24[431] + src24[432] + src24[433] + src24[434] + src24[435] + src24[436] + src24[437] + src24[438] + src24[439] + src24[440] + src24[441] + src24[442] + src24[443] + src24[444] + src24[445] + src24[446] + src24[447] + src24[448] + src24[449] + src24[450] + src24[451] + src24[452] + src24[453] + src24[454] + src24[455] + src24[456] + src24[457] + src24[458] + src24[459] + src24[460] + src24[461] + src24[462] + src24[463] + src24[464] + src24[465] + src24[466] + src24[467] + src24[468] + src24[469] + src24[470] + src24[471] + src24[472] + src24[473] + src24[474] + src24[475] + src24[476] + src24[477] + src24[478] + src24[479] + src24[480] + src24[481] + src24[482] + src24[483] + src24[484] + src24[485])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255] + src25[256] + src25[257] + src25[258] + src25[259] + src25[260] + src25[261] + src25[262] + src25[263] + src25[264] + src25[265] + src25[266] + src25[267] + src25[268] + src25[269] + src25[270] + src25[271] + src25[272] + src25[273] + src25[274] + src25[275] + src25[276] + src25[277] + src25[278] + src25[279] + src25[280] + src25[281] + src25[282] + src25[283] + src25[284] + src25[285] + src25[286] + src25[287] + src25[288] + src25[289] + src25[290] + src25[291] + src25[292] + src25[293] + src25[294] + src25[295] + src25[296] + src25[297] + src25[298] + src25[299] + src25[300] + src25[301] + src25[302] + src25[303] + src25[304] + src25[305] + src25[306] + src25[307] + src25[308] + src25[309] + src25[310] + src25[311] + src25[312] + src25[313] + src25[314] + src25[315] + src25[316] + src25[317] + src25[318] + src25[319] + src25[320] + src25[321] + src25[322] + src25[323] + src25[324] + src25[325] + src25[326] + src25[327] + src25[328] + src25[329] + src25[330] + src25[331] + src25[332] + src25[333] + src25[334] + src25[335] + src25[336] + src25[337] + src25[338] + src25[339] + src25[340] + src25[341] + src25[342] + src25[343] + src25[344] + src25[345] + src25[346] + src25[347] + src25[348] + src25[349] + src25[350] + src25[351] + src25[352] + src25[353] + src25[354] + src25[355] + src25[356] + src25[357] + src25[358] + src25[359] + src25[360] + src25[361] + src25[362] + src25[363] + src25[364] + src25[365] + src25[366] + src25[367] + src25[368] + src25[369] + src25[370] + src25[371] + src25[372] + src25[373] + src25[374] + src25[375] + src25[376] + src25[377] + src25[378] + src25[379] + src25[380] + src25[381] + src25[382] + src25[383] + src25[384] + src25[385] + src25[386] + src25[387] + src25[388] + src25[389] + src25[390] + src25[391] + src25[392] + src25[393] + src25[394] + src25[395] + src25[396] + src25[397] + src25[398] + src25[399] + src25[400] + src25[401] + src25[402] + src25[403] + src25[404] + src25[405] + src25[406] + src25[407] + src25[408] + src25[409] + src25[410] + src25[411] + src25[412] + src25[413] + src25[414] + src25[415] + src25[416] + src25[417] + src25[418] + src25[419] + src25[420] + src25[421] + src25[422] + src25[423] + src25[424] + src25[425] + src25[426] + src25[427] + src25[428] + src25[429] + src25[430] + src25[431] + src25[432] + src25[433] + src25[434] + src25[435] + src25[436] + src25[437] + src25[438] + src25[439] + src25[440] + src25[441] + src25[442] + src25[443] + src25[444] + src25[445] + src25[446] + src25[447] + src25[448] + src25[449] + src25[450] + src25[451] + src25[452] + src25[453] + src25[454] + src25[455] + src25[456] + src25[457] + src25[458] + src25[459] + src25[460] + src25[461] + src25[462] + src25[463] + src25[464] + src25[465] + src25[466] + src25[467] + src25[468] + src25[469] + src25[470] + src25[471] + src25[472] + src25[473] + src25[474] + src25[475] + src25[476] + src25[477] + src25[478] + src25[479] + src25[480] + src25[481] + src25[482] + src25[483] + src25[484] + src25[485])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255] + src26[256] + src26[257] + src26[258] + src26[259] + src26[260] + src26[261] + src26[262] + src26[263] + src26[264] + src26[265] + src26[266] + src26[267] + src26[268] + src26[269] + src26[270] + src26[271] + src26[272] + src26[273] + src26[274] + src26[275] + src26[276] + src26[277] + src26[278] + src26[279] + src26[280] + src26[281] + src26[282] + src26[283] + src26[284] + src26[285] + src26[286] + src26[287] + src26[288] + src26[289] + src26[290] + src26[291] + src26[292] + src26[293] + src26[294] + src26[295] + src26[296] + src26[297] + src26[298] + src26[299] + src26[300] + src26[301] + src26[302] + src26[303] + src26[304] + src26[305] + src26[306] + src26[307] + src26[308] + src26[309] + src26[310] + src26[311] + src26[312] + src26[313] + src26[314] + src26[315] + src26[316] + src26[317] + src26[318] + src26[319] + src26[320] + src26[321] + src26[322] + src26[323] + src26[324] + src26[325] + src26[326] + src26[327] + src26[328] + src26[329] + src26[330] + src26[331] + src26[332] + src26[333] + src26[334] + src26[335] + src26[336] + src26[337] + src26[338] + src26[339] + src26[340] + src26[341] + src26[342] + src26[343] + src26[344] + src26[345] + src26[346] + src26[347] + src26[348] + src26[349] + src26[350] + src26[351] + src26[352] + src26[353] + src26[354] + src26[355] + src26[356] + src26[357] + src26[358] + src26[359] + src26[360] + src26[361] + src26[362] + src26[363] + src26[364] + src26[365] + src26[366] + src26[367] + src26[368] + src26[369] + src26[370] + src26[371] + src26[372] + src26[373] + src26[374] + src26[375] + src26[376] + src26[377] + src26[378] + src26[379] + src26[380] + src26[381] + src26[382] + src26[383] + src26[384] + src26[385] + src26[386] + src26[387] + src26[388] + src26[389] + src26[390] + src26[391] + src26[392] + src26[393] + src26[394] + src26[395] + src26[396] + src26[397] + src26[398] + src26[399] + src26[400] + src26[401] + src26[402] + src26[403] + src26[404] + src26[405] + src26[406] + src26[407] + src26[408] + src26[409] + src26[410] + src26[411] + src26[412] + src26[413] + src26[414] + src26[415] + src26[416] + src26[417] + src26[418] + src26[419] + src26[420] + src26[421] + src26[422] + src26[423] + src26[424] + src26[425] + src26[426] + src26[427] + src26[428] + src26[429] + src26[430] + src26[431] + src26[432] + src26[433] + src26[434] + src26[435] + src26[436] + src26[437] + src26[438] + src26[439] + src26[440] + src26[441] + src26[442] + src26[443] + src26[444] + src26[445] + src26[446] + src26[447] + src26[448] + src26[449] + src26[450] + src26[451] + src26[452] + src26[453] + src26[454] + src26[455] + src26[456] + src26[457] + src26[458] + src26[459] + src26[460] + src26[461] + src26[462] + src26[463] + src26[464] + src26[465] + src26[466] + src26[467] + src26[468] + src26[469] + src26[470] + src26[471] + src26[472] + src26[473] + src26[474] + src26[475] + src26[476] + src26[477] + src26[478] + src26[479] + src26[480] + src26[481] + src26[482] + src26[483] + src26[484] + src26[485])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255] + src27[256] + src27[257] + src27[258] + src27[259] + src27[260] + src27[261] + src27[262] + src27[263] + src27[264] + src27[265] + src27[266] + src27[267] + src27[268] + src27[269] + src27[270] + src27[271] + src27[272] + src27[273] + src27[274] + src27[275] + src27[276] + src27[277] + src27[278] + src27[279] + src27[280] + src27[281] + src27[282] + src27[283] + src27[284] + src27[285] + src27[286] + src27[287] + src27[288] + src27[289] + src27[290] + src27[291] + src27[292] + src27[293] + src27[294] + src27[295] + src27[296] + src27[297] + src27[298] + src27[299] + src27[300] + src27[301] + src27[302] + src27[303] + src27[304] + src27[305] + src27[306] + src27[307] + src27[308] + src27[309] + src27[310] + src27[311] + src27[312] + src27[313] + src27[314] + src27[315] + src27[316] + src27[317] + src27[318] + src27[319] + src27[320] + src27[321] + src27[322] + src27[323] + src27[324] + src27[325] + src27[326] + src27[327] + src27[328] + src27[329] + src27[330] + src27[331] + src27[332] + src27[333] + src27[334] + src27[335] + src27[336] + src27[337] + src27[338] + src27[339] + src27[340] + src27[341] + src27[342] + src27[343] + src27[344] + src27[345] + src27[346] + src27[347] + src27[348] + src27[349] + src27[350] + src27[351] + src27[352] + src27[353] + src27[354] + src27[355] + src27[356] + src27[357] + src27[358] + src27[359] + src27[360] + src27[361] + src27[362] + src27[363] + src27[364] + src27[365] + src27[366] + src27[367] + src27[368] + src27[369] + src27[370] + src27[371] + src27[372] + src27[373] + src27[374] + src27[375] + src27[376] + src27[377] + src27[378] + src27[379] + src27[380] + src27[381] + src27[382] + src27[383] + src27[384] + src27[385] + src27[386] + src27[387] + src27[388] + src27[389] + src27[390] + src27[391] + src27[392] + src27[393] + src27[394] + src27[395] + src27[396] + src27[397] + src27[398] + src27[399] + src27[400] + src27[401] + src27[402] + src27[403] + src27[404] + src27[405] + src27[406] + src27[407] + src27[408] + src27[409] + src27[410] + src27[411] + src27[412] + src27[413] + src27[414] + src27[415] + src27[416] + src27[417] + src27[418] + src27[419] + src27[420] + src27[421] + src27[422] + src27[423] + src27[424] + src27[425] + src27[426] + src27[427] + src27[428] + src27[429] + src27[430] + src27[431] + src27[432] + src27[433] + src27[434] + src27[435] + src27[436] + src27[437] + src27[438] + src27[439] + src27[440] + src27[441] + src27[442] + src27[443] + src27[444] + src27[445] + src27[446] + src27[447] + src27[448] + src27[449] + src27[450] + src27[451] + src27[452] + src27[453] + src27[454] + src27[455] + src27[456] + src27[457] + src27[458] + src27[459] + src27[460] + src27[461] + src27[462] + src27[463] + src27[464] + src27[465] + src27[466] + src27[467] + src27[468] + src27[469] + src27[470] + src27[471] + src27[472] + src27[473] + src27[474] + src27[475] + src27[476] + src27[477] + src27[478] + src27[479] + src27[480] + src27[481] + src27[482] + src27[483] + src27[484] + src27[485])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255] + src28[256] + src28[257] + src28[258] + src28[259] + src28[260] + src28[261] + src28[262] + src28[263] + src28[264] + src28[265] + src28[266] + src28[267] + src28[268] + src28[269] + src28[270] + src28[271] + src28[272] + src28[273] + src28[274] + src28[275] + src28[276] + src28[277] + src28[278] + src28[279] + src28[280] + src28[281] + src28[282] + src28[283] + src28[284] + src28[285] + src28[286] + src28[287] + src28[288] + src28[289] + src28[290] + src28[291] + src28[292] + src28[293] + src28[294] + src28[295] + src28[296] + src28[297] + src28[298] + src28[299] + src28[300] + src28[301] + src28[302] + src28[303] + src28[304] + src28[305] + src28[306] + src28[307] + src28[308] + src28[309] + src28[310] + src28[311] + src28[312] + src28[313] + src28[314] + src28[315] + src28[316] + src28[317] + src28[318] + src28[319] + src28[320] + src28[321] + src28[322] + src28[323] + src28[324] + src28[325] + src28[326] + src28[327] + src28[328] + src28[329] + src28[330] + src28[331] + src28[332] + src28[333] + src28[334] + src28[335] + src28[336] + src28[337] + src28[338] + src28[339] + src28[340] + src28[341] + src28[342] + src28[343] + src28[344] + src28[345] + src28[346] + src28[347] + src28[348] + src28[349] + src28[350] + src28[351] + src28[352] + src28[353] + src28[354] + src28[355] + src28[356] + src28[357] + src28[358] + src28[359] + src28[360] + src28[361] + src28[362] + src28[363] + src28[364] + src28[365] + src28[366] + src28[367] + src28[368] + src28[369] + src28[370] + src28[371] + src28[372] + src28[373] + src28[374] + src28[375] + src28[376] + src28[377] + src28[378] + src28[379] + src28[380] + src28[381] + src28[382] + src28[383] + src28[384] + src28[385] + src28[386] + src28[387] + src28[388] + src28[389] + src28[390] + src28[391] + src28[392] + src28[393] + src28[394] + src28[395] + src28[396] + src28[397] + src28[398] + src28[399] + src28[400] + src28[401] + src28[402] + src28[403] + src28[404] + src28[405] + src28[406] + src28[407] + src28[408] + src28[409] + src28[410] + src28[411] + src28[412] + src28[413] + src28[414] + src28[415] + src28[416] + src28[417] + src28[418] + src28[419] + src28[420] + src28[421] + src28[422] + src28[423] + src28[424] + src28[425] + src28[426] + src28[427] + src28[428] + src28[429] + src28[430] + src28[431] + src28[432] + src28[433] + src28[434] + src28[435] + src28[436] + src28[437] + src28[438] + src28[439] + src28[440] + src28[441] + src28[442] + src28[443] + src28[444] + src28[445] + src28[446] + src28[447] + src28[448] + src28[449] + src28[450] + src28[451] + src28[452] + src28[453] + src28[454] + src28[455] + src28[456] + src28[457] + src28[458] + src28[459] + src28[460] + src28[461] + src28[462] + src28[463] + src28[464] + src28[465] + src28[466] + src28[467] + src28[468] + src28[469] + src28[470] + src28[471] + src28[472] + src28[473] + src28[474] + src28[475] + src28[476] + src28[477] + src28[478] + src28[479] + src28[480] + src28[481] + src28[482] + src28[483] + src28[484] + src28[485])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255] + src29[256] + src29[257] + src29[258] + src29[259] + src29[260] + src29[261] + src29[262] + src29[263] + src29[264] + src29[265] + src29[266] + src29[267] + src29[268] + src29[269] + src29[270] + src29[271] + src29[272] + src29[273] + src29[274] + src29[275] + src29[276] + src29[277] + src29[278] + src29[279] + src29[280] + src29[281] + src29[282] + src29[283] + src29[284] + src29[285] + src29[286] + src29[287] + src29[288] + src29[289] + src29[290] + src29[291] + src29[292] + src29[293] + src29[294] + src29[295] + src29[296] + src29[297] + src29[298] + src29[299] + src29[300] + src29[301] + src29[302] + src29[303] + src29[304] + src29[305] + src29[306] + src29[307] + src29[308] + src29[309] + src29[310] + src29[311] + src29[312] + src29[313] + src29[314] + src29[315] + src29[316] + src29[317] + src29[318] + src29[319] + src29[320] + src29[321] + src29[322] + src29[323] + src29[324] + src29[325] + src29[326] + src29[327] + src29[328] + src29[329] + src29[330] + src29[331] + src29[332] + src29[333] + src29[334] + src29[335] + src29[336] + src29[337] + src29[338] + src29[339] + src29[340] + src29[341] + src29[342] + src29[343] + src29[344] + src29[345] + src29[346] + src29[347] + src29[348] + src29[349] + src29[350] + src29[351] + src29[352] + src29[353] + src29[354] + src29[355] + src29[356] + src29[357] + src29[358] + src29[359] + src29[360] + src29[361] + src29[362] + src29[363] + src29[364] + src29[365] + src29[366] + src29[367] + src29[368] + src29[369] + src29[370] + src29[371] + src29[372] + src29[373] + src29[374] + src29[375] + src29[376] + src29[377] + src29[378] + src29[379] + src29[380] + src29[381] + src29[382] + src29[383] + src29[384] + src29[385] + src29[386] + src29[387] + src29[388] + src29[389] + src29[390] + src29[391] + src29[392] + src29[393] + src29[394] + src29[395] + src29[396] + src29[397] + src29[398] + src29[399] + src29[400] + src29[401] + src29[402] + src29[403] + src29[404] + src29[405] + src29[406] + src29[407] + src29[408] + src29[409] + src29[410] + src29[411] + src29[412] + src29[413] + src29[414] + src29[415] + src29[416] + src29[417] + src29[418] + src29[419] + src29[420] + src29[421] + src29[422] + src29[423] + src29[424] + src29[425] + src29[426] + src29[427] + src29[428] + src29[429] + src29[430] + src29[431] + src29[432] + src29[433] + src29[434] + src29[435] + src29[436] + src29[437] + src29[438] + src29[439] + src29[440] + src29[441] + src29[442] + src29[443] + src29[444] + src29[445] + src29[446] + src29[447] + src29[448] + src29[449] + src29[450] + src29[451] + src29[452] + src29[453] + src29[454] + src29[455] + src29[456] + src29[457] + src29[458] + src29[459] + src29[460] + src29[461] + src29[462] + src29[463] + src29[464] + src29[465] + src29[466] + src29[467] + src29[468] + src29[469] + src29[470] + src29[471] + src29[472] + src29[473] + src29[474] + src29[475] + src29[476] + src29[477] + src29[478] + src29[479] + src29[480] + src29[481] + src29[482] + src29[483] + src29[484] + src29[485])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255] + src30[256] + src30[257] + src30[258] + src30[259] + src30[260] + src30[261] + src30[262] + src30[263] + src30[264] + src30[265] + src30[266] + src30[267] + src30[268] + src30[269] + src30[270] + src30[271] + src30[272] + src30[273] + src30[274] + src30[275] + src30[276] + src30[277] + src30[278] + src30[279] + src30[280] + src30[281] + src30[282] + src30[283] + src30[284] + src30[285] + src30[286] + src30[287] + src30[288] + src30[289] + src30[290] + src30[291] + src30[292] + src30[293] + src30[294] + src30[295] + src30[296] + src30[297] + src30[298] + src30[299] + src30[300] + src30[301] + src30[302] + src30[303] + src30[304] + src30[305] + src30[306] + src30[307] + src30[308] + src30[309] + src30[310] + src30[311] + src30[312] + src30[313] + src30[314] + src30[315] + src30[316] + src30[317] + src30[318] + src30[319] + src30[320] + src30[321] + src30[322] + src30[323] + src30[324] + src30[325] + src30[326] + src30[327] + src30[328] + src30[329] + src30[330] + src30[331] + src30[332] + src30[333] + src30[334] + src30[335] + src30[336] + src30[337] + src30[338] + src30[339] + src30[340] + src30[341] + src30[342] + src30[343] + src30[344] + src30[345] + src30[346] + src30[347] + src30[348] + src30[349] + src30[350] + src30[351] + src30[352] + src30[353] + src30[354] + src30[355] + src30[356] + src30[357] + src30[358] + src30[359] + src30[360] + src30[361] + src30[362] + src30[363] + src30[364] + src30[365] + src30[366] + src30[367] + src30[368] + src30[369] + src30[370] + src30[371] + src30[372] + src30[373] + src30[374] + src30[375] + src30[376] + src30[377] + src30[378] + src30[379] + src30[380] + src30[381] + src30[382] + src30[383] + src30[384] + src30[385] + src30[386] + src30[387] + src30[388] + src30[389] + src30[390] + src30[391] + src30[392] + src30[393] + src30[394] + src30[395] + src30[396] + src30[397] + src30[398] + src30[399] + src30[400] + src30[401] + src30[402] + src30[403] + src30[404] + src30[405] + src30[406] + src30[407] + src30[408] + src30[409] + src30[410] + src30[411] + src30[412] + src30[413] + src30[414] + src30[415] + src30[416] + src30[417] + src30[418] + src30[419] + src30[420] + src30[421] + src30[422] + src30[423] + src30[424] + src30[425] + src30[426] + src30[427] + src30[428] + src30[429] + src30[430] + src30[431] + src30[432] + src30[433] + src30[434] + src30[435] + src30[436] + src30[437] + src30[438] + src30[439] + src30[440] + src30[441] + src30[442] + src30[443] + src30[444] + src30[445] + src30[446] + src30[447] + src30[448] + src30[449] + src30[450] + src30[451] + src30[452] + src30[453] + src30[454] + src30[455] + src30[456] + src30[457] + src30[458] + src30[459] + src30[460] + src30[461] + src30[462] + src30[463] + src30[464] + src30[465] + src30[466] + src30[467] + src30[468] + src30[469] + src30[470] + src30[471] + src30[472] + src30[473] + src30[474] + src30[475] + src30[476] + src30[477] + src30[478] + src30[479] + src30[480] + src30[481] + src30[482] + src30[483] + src30[484] + src30[485])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255] + src31[256] + src31[257] + src31[258] + src31[259] + src31[260] + src31[261] + src31[262] + src31[263] + src31[264] + src31[265] + src31[266] + src31[267] + src31[268] + src31[269] + src31[270] + src31[271] + src31[272] + src31[273] + src31[274] + src31[275] + src31[276] + src31[277] + src31[278] + src31[279] + src31[280] + src31[281] + src31[282] + src31[283] + src31[284] + src31[285] + src31[286] + src31[287] + src31[288] + src31[289] + src31[290] + src31[291] + src31[292] + src31[293] + src31[294] + src31[295] + src31[296] + src31[297] + src31[298] + src31[299] + src31[300] + src31[301] + src31[302] + src31[303] + src31[304] + src31[305] + src31[306] + src31[307] + src31[308] + src31[309] + src31[310] + src31[311] + src31[312] + src31[313] + src31[314] + src31[315] + src31[316] + src31[317] + src31[318] + src31[319] + src31[320] + src31[321] + src31[322] + src31[323] + src31[324] + src31[325] + src31[326] + src31[327] + src31[328] + src31[329] + src31[330] + src31[331] + src31[332] + src31[333] + src31[334] + src31[335] + src31[336] + src31[337] + src31[338] + src31[339] + src31[340] + src31[341] + src31[342] + src31[343] + src31[344] + src31[345] + src31[346] + src31[347] + src31[348] + src31[349] + src31[350] + src31[351] + src31[352] + src31[353] + src31[354] + src31[355] + src31[356] + src31[357] + src31[358] + src31[359] + src31[360] + src31[361] + src31[362] + src31[363] + src31[364] + src31[365] + src31[366] + src31[367] + src31[368] + src31[369] + src31[370] + src31[371] + src31[372] + src31[373] + src31[374] + src31[375] + src31[376] + src31[377] + src31[378] + src31[379] + src31[380] + src31[381] + src31[382] + src31[383] + src31[384] + src31[385] + src31[386] + src31[387] + src31[388] + src31[389] + src31[390] + src31[391] + src31[392] + src31[393] + src31[394] + src31[395] + src31[396] + src31[397] + src31[398] + src31[399] + src31[400] + src31[401] + src31[402] + src31[403] + src31[404] + src31[405] + src31[406] + src31[407] + src31[408] + src31[409] + src31[410] + src31[411] + src31[412] + src31[413] + src31[414] + src31[415] + src31[416] + src31[417] + src31[418] + src31[419] + src31[420] + src31[421] + src31[422] + src31[423] + src31[424] + src31[425] + src31[426] + src31[427] + src31[428] + src31[429] + src31[430] + src31[431] + src31[432] + src31[433] + src31[434] + src31[435] + src31[436] + src31[437] + src31[438] + src31[439] + src31[440] + src31[441] + src31[442] + src31[443] + src31[444] + src31[445] + src31[446] + src31[447] + src31[448] + src31[449] + src31[450] + src31[451] + src31[452] + src31[453] + src31[454] + src31[455] + src31[456] + src31[457] + src31[458] + src31[459] + src31[460] + src31[461] + src31[462] + src31[463] + src31[464] + src31[465] + src31[466] + src31[467] + src31[468] + src31[469] + src31[470] + src31[471] + src31[472] + src31[473] + src31[474] + src31[475] + src31[476] + src31[477] + src31[478] + src31[479] + src31[480] + src31[481] + src31[482] + src31[483] + src31[484] + src31[485])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63] + src32[64] + src32[65] + src32[66] + src32[67] + src32[68] + src32[69] + src32[70] + src32[71] + src32[72] + src32[73] + src32[74] + src32[75] + src32[76] + src32[77] + src32[78] + src32[79] + src32[80] + src32[81] + src32[82] + src32[83] + src32[84] + src32[85] + src32[86] + src32[87] + src32[88] + src32[89] + src32[90] + src32[91] + src32[92] + src32[93] + src32[94] + src32[95] + src32[96] + src32[97] + src32[98] + src32[99] + src32[100] + src32[101] + src32[102] + src32[103] + src32[104] + src32[105] + src32[106] + src32[107] + src32[108] + src32[109] + src32[110] + src32[111] + src32[112] + src32[113] + src32[114] + src32[115] + src32[116] + src32[117] + src32[118] + src32[119] + src32[120] + src32[121] + src32[122] + src32[123] + src32[124] + src32[125] + src32[126] + src32[127] + src32[128] + src32[129] + src32[130] + src32[131] + src32[132] + src32[133] + src32[134] + src32[135] + src32[136] + src32[137] + src32[138] + src32[139] + src32[140] + src32[141] + src32[142] + src32[143] + src32[144] + src32[145] + src32[146] + src32[147] + src32[148] + src32[149] + src32[150] + src32[151] + src32[152] + src32[153] + src32[154] + src32[155] + src32[156] + src32[157] + src32[158] + src32[159] + src32[160] + src32[161] + src32[162] + src32[163] + src32[164] + src32[165] + src32[166] + src32[167] + src32[168] + src32[169] + src32[170] + src32[171] + src32[172] + src32[173] + src32[174] + src32[175] + src32[176] + src32[177] + src32[178] + src32[179] + src32[180] + src32[181] + src32[182] + src32[183] + src32[184] + src32[185] + src32[186] + src32[187] + src32[188] + src32[189] + src32[190] + src32[191] + src32[192] + src32[193] + src32[194] + src32[195] + src32[196] + src32[197] + src32[198] + src32[199] + src32[200] + src32[201] + src32[202] + src32[203] + src32[204] + src32[205] + src32[206] + src32[207] + src32[208] + src32[209] + src32[210] + src32[211] + src32[212] + src32[213] + src32[214] + src32[215] + src32[216] + src32[217] + src32[218] + src32[219] + src32[220] + src32[221] + src32[222] + src32[223] + src32[224] + src32[225] + src32[226] + src32[227] + src32[228] + src32[229] + src32[230] + src32[231] + src32[232] + src32[233] + src32[234] + src32[235] + src32[236] + src32[237] + src32[238] + src32[239] + src32[240] + src32[241] + src32[242] + src32[243] + src32[244] + src32[245] + src32[246] + src32[247] + src32[248] + src32[249] + src32[250] + src32[251] + src32[252] + src32[253] + src32[254] + src32[255] + src32[256] + src32[257] + src32[258] + src32[259] + src32[260] + src32[261] + src32[262] + src32[263] + src32[264] + src32[265] + src32[266] + src32[267] + src32[268] + src32[269] + src32[270] + src32[271] + src32[272] + src32[273] + src32[274] + src32[275] + src32[276] + src32[277] + src32[278] + src32[279] + src32[280] + src32[281] + src32[282] + src32[283] + src32[284] + src32[285] + src32[286] + src32[287] + src32[288] + src32[289] + src32[290] + src32[291] + src32[292] + src32[293] + src32[294] + src32[295] + src32[296] + src32[297] + src32[298] + src32[299] + src32[300] + src32[301] + src32[302] + src32[303] + src32[304] + src32[305] + src32[306] + src32[307] + src32[308] + src32[309] + src32[310] + src32[311] + src32[312] + src32[313] + src32[314] + src32[315] + src32[316] + src32[317] + src32[318] + src32[319] + src32[320] + src32[321] + src32[322] + src32[323] + src32[324] + src32[325] + src32[326] + src32[327] + src32[328] + src32[329] + src32[330] + src32[331] + src32[332] + src32[333] + src32[334] + src32[335] + src32[336] + src32[337] + src32[338] + src32[339] + src32[340] + src32[341] + src32[342] + src32[343] + src32[344] + src32[345] + src32[346] + src32[347] + src32[348] + src32[349] + src32[350] + src32[351] + src32[352] + src32[353] + src32[354] + src32[355] + src32[356] + src32[357] + src32[358] + src32[359] + src32[360] + src32[361] + src32[362] + src32[363] + src32[364] + src32[365] + src32[366] + src32[367] + src32[368] + src32[369] + src32[370] + src32[371] + src32[372] + src32[373] + src32[374] + src32[375] + src32[376] + src32[377] + src32[378] + src32[379] + src32[380] + src32[381] + src32[382] + src32[383] + src32[384] + src32[385] + src32[386] + src32[387] + src32[388] + src32[389] + src32[390] + src32[391] + src32[392] + src32[393] + src32[394] + src32[395] + src32[396] + src32[397] + src32[398] + src32[399] + src32[400] + src32[401] + src32[402] + src32[403] + src32[404] + src32[405] + src32[406] + src32[407] + src32[408] + src32[409] + src32[410] + src32[411] + src32[412] + src32[413] + src32[414] + src32[415] + src32[416] + src32[417] + src32[418] + src32[419] + src32[420] + src32[421] + src32[422] + src32[423] + src32[424] + src32[425] + src32[426] + src32[427] + src32[428] + src32[429] + src32[430] + src32[431] + src32[432] + src32[433] + src32[434] + src32[435] + src32[436] + src32[437] + src32[438] + src32[439] + src32[440] + src32[441] + src32[442] + src32[443] + src32[444] + src32[445] + src32[446] + src32[447] + src32[448] + src32[449] + src32[450] + src32[451] + src32[452] + src32[453] + src32[454] + src32[455] + src32[456] + src32[457] + src32[458] + src32[459] + src32[460] + src32[461] + src32[462] + src32[463] + src32[464] + src32[465] + src32[466] + src32[467] + src32[468] + src32[469] + src32[470] + src32[471] + src32[472] + src32[473] + src32[474] + src32[475] + src32[476] + src32[477] + src32[478] + src32[479] + src32[480] + src32[481] + src32[482] + src32[483] + src32[484] + src32[485])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63] + src33[64] + src33[65] + src33[66] + src33[67] + src33[68] + src33[69] + src33[70] + src33[71] + src33[72] + src33[73] + src33[74] + src33[75] + src33[76] + src33[77] + src33[78] + src33[79] + src33[80] + src33[81] + src33[82] + src33[83] + src33[84] + src33[85] + src33[86] + src33[87] + src33[88] + src33[89] + src33[90] + src33[91] + src33[92] + src33[93] + src33[94] + src33[95] + src33[96] + src33[97] + src33[98] + src33[99] + src33[100] + src33[101] + src33[102] + src33[103] + src33[104] + src33[105] + src33[106] + src33[107] + src33[108] + src33[109] + src33[110] + src33[111] + src33[112] + src33[113] + src33[114] + src33[115] + src33[116] + src33[117] + src33[118] + src33[119] + src33[120] + src33[121] + src33[122] + src33[123] + src33[124] + src33[125] + src33[126] + src33[127] + src33[128] + src33[129] + src33[130] + src33[131] + src33[132] + src33[133] + src33[134] + src33[135] + src33[136] + src33[137] + src33[138] + src33[139] + src33[140] + src33[141] + src33[142] + src33[143] + src33[144] + src33[145] + src33[146] + src33[147] + src33[148] + src33[149] + src33[150] + src33[151] + src33[152] + src33[153] + src33[154] + src33[155] + src33[156] + src33[157] + src33[158] + src33[159] + src33[160] + src33[161] + src33[162] + src33[163] + src33[164] + src33[165] + src33[166] + src33[167] + src33[168] + src33[169] + src33[170] + src33[171] + src33[172] + src33[173] + src33[174] + src33[175] + src33[176] + src33[177] + src33[178] + src33[179] + src33[180] + src33[181] + src33[182] + src33[183] + src33[184] + src33[185] + src33[186] + src33[187] + src33[188] + src33[189] + src33[190] + src33[191] + src33[192] + src33[193] + src33[194] + src33[195] + src33[196] + src33[197] + src33[198] + src33[199] + src33[200] + src33[201] + src33[202] + src33[203] + src33[204] + src33[205] + src33[206] + src33[207] + src33[208] + src33[209] + src33[210] + src33[211] + src33[212] + src33[213] + src33[214] + src33[215] + src33[216] + src33[217] + src33[218] + src33[219] + src33[220] + src33[221] + src33[222] + src33[223] + src33[224] + src33[225] + src33[226] + src33[227] + src33[228] + src33[229] + src33[230] + src33[231] + src33[232] + src33[233] + src33[234] + src33[235] + src33[236] + src33[237] + src33[238] + src33[239] + src33[240] + src33[241] + src33[242] + src33[243] + src33[244] + src33[245] + src33[246] + src33[247] + src33[248] + src33[249] + src33[250] + src33[251] + src33[252] + src33[253] + src33[254] + src33[255] + src33[256] + src33[257] + src33[258] + src33[259] + src33[260] + src33[261] + src33[262] + src33[263] + src33[264] + src33[265] + src33[266] + src33[267] + src33[268] + src33[269] + src33[270] + src33[271] + src33[272] + src33[273] + src33[274] + src33[275] + src33[276] + src33[277] + src33[278] + src33[279] + src33[280] + src33[281] + src33[282] + src33[283] + src33[284] + src33[285] + src33[286] + src33[287] + src33[288] + src33[289] + src33[290] + src33[291] + src33[292] + src33[293] + src33[294] + src33[295] + src33[296] + src33[297] + src33[298] + src33[299] + src33[300] + src33[301] + src33[302] + src33[303] + src33[304] + src33[305] + src33[306] + src33[307] + src33[308] + src33[309] + src33[310] + src33[311] + src33[312] + src33[313] + src33[314] + src33[315] + src33[316] + src33[317] + src33[318] + src33[319] + src33[320] + src33[321] + src33[322] + src33[323] + src33[324] + src33[325] + src33[326] + src33[327] + src33[328] + src33[329] + src33[330] + src33[331] + src33[332] + src33[333] + src33[334] + src33[335] + src33[336] + src33[337] + src33[338] + src33[339] + src33[340] + src33[341] + src33[342] + src33[343] + src33[344] + src33[345] + src33[346] + src33[347] + src33[348] + src33[349] + src33[350] + src33[351] + src33[352] + src33[353] + src33[354] + src33[355] + src33[356] + src33[357] + src33[358] + src33[359] + src33[360] + src33[361] + src33[362] + src33[363] + src33[364] + src33[365] + src33[366] + src33[367] + src33[368] + src33[369] + src33[370] + src33[371] + src33[372] + src33[373] + src33[374] + src33[375] + src33[376] + src33[377] + src33[378] + src33[379] + src33[380] + src33[381] + src33[382] + src33[383] + src33[384] + src33[385] + src33[386] + src33[387] + src33[388] + src33[389] + src33[390] + src33[391] + src33[392] + src33[393] + src33[394] + src33[395] + src33[396] + src33[397] + src33[398] + src33[399] + src33[400] + src33[401] + src33[402] + src33[403] + src33[404] + src33[405] + src33[406] + src33[407] + src33[408] + src33[409] + src33[410] + src33[411] + src33[412] + src33[413] + src33[414] + src33[415] + src33[416] + src33[417] + src33[418] + src33[419] + src33[420] + src33[421] + src33[422] + src33[423] + src33[424] + src33[425] + src33[426] + src33[427] + src33[428] + src33[429] + src33[430] + src33[431] + src33[432] + src33[433] + src33[434] + src33[435] + src33[436] + src33[437] + src33[438] + src33[439] + src33[440] + src33[441] + src33[442] + src33[443] + src33[444] + src33[445] + src33[446] + src33[447] + src33[448] + src33[449] + src33[450] + src33[451] + src33[452] + src33[453] + src33[454] + src33[455] + src33[456] + src33[457] + src33[458] + src33[459] + src33[460] + src33[461] + src33[462] + src33[463] + src33[464] + src33[465] + src33[466] + src33[467] + src33[468] + src33[469] + src33[470] + src33[471] + src33[472] + src33[473] + src33[474] + src33[475] + src33[476] + src33[477] + src33[478] + src33[479] + src33[480] + src33[481] + src33[482] + src33[483] + src33[484] + src33[485])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63] + src34[64] + src34[65] + src34[66] + src34[67] + src34[68] + src34[69] + src34[70] + src34[71] + src34[72] + src34[73] + src34[74] + src34[75] + src34[76] + src34[77] + src34[78] + src34[79] + src34[80] + src34[81] + src34[82] + src34[83] + src34[84] + src34[85] + src34[86] + src34[87] + src34[88] + src34[89] + src34[90] + src34[91] + src34[92] + src34[93] + src34[94] + src34[95] + src34[96] + src34[97] + src34[98] + src34[99] + src34[100] + src34[101] + src34[102] + src34[103] + src34[104] + src34[105] + src34[106] + src34[107] + src34[108] + src34[109] + src34[110] + src34[111] + src34[112] + src34[113] + src34[114] + src34[115] + src34[116] + src34[117] + src34[118] + src34[119] + src34[120] + src34[121] + src34[122] + src34[123] + src34[124] + src34[125] + src34[126] + src34[127] + src34[128] + src34[129] + src34[130] + src34[131] + src34[132] + src34[133] + src34[134] + src34[135] + src34[136] + src34[137] + src34[138] + src34[139] + src34[140] + src34[141] + src34[142] + src34[143] + src34[144] + src34[145] + src34[146] + src34[147] + src34[148] + src34[149] + src34[150] + src34[151] + src34[152] + src34[153] + src34[154] + src34[155] + src34[156] + src34[157] + src34[158] + src34[159] + src34[160] + src34[161] + src34[162] + src34[163] + src34[164] + src34[165] + src34[166] + src34[167] + src34[168] + src34[169] + src34[170] + src34[171] + src34[172] + src34[173] + src34[174] + src34[175] + src34[176] + src34[177] + src34[178] + src34[179] + src34[180] + src34[181] + src34[182] + src34[183] + src34[184] + src34[185] + src34[186] + src34[187] + src34[188] + src34[189] + src34[190] + src34[191] + src34[192] + src34[193] + src34[194] + src34[195] + src34[196] + src34[197] + src34[198] + src34[199] + src34[200] + src34[201] + src34[202] + src34[203] + src34[204] + src34[205] + src34[206] + src34[207] + src34[208] + src34[209] + src34[210] + src34[211] + src34[212] + src34[213] + src34[214] + src34[215] + src34[216] + src34[217] + src34[218] + src34[219] + src34[220] + src34[221] + src34[222] + src34[223] + src34[224] + src34[225] + src34[226] + src34[227] + src34[228] + src34[229] + src34[230] + src34[231] + src34[232] + src34[233] + src34[234] + src34[235] + src34[236] + src34[237] + src34[238] + src34[239] + src34[240] + src34[241] + src34[242] + src34[243] + src34[244] + src34[245] + src34[246] + src34[247] + src34[248] + src34[249] + src34[250] + src34[251] + src34[252] + src34[253] + src34[254] + src34[255] + src34[256] + src34[257] + src34[258] + src34[259] + src34[260] + src34[261] + src34[262] + src34[263] + src34[264] + src34[265] + src34[266] + src34[267] + src34[268] + src34[269] + src34[270] + src34[271] + src34[272] + src34[273] + src34[274] + src34[275] + src34[276] + src34[277] + src34[278] + src34[279] + src34[280] + src34[281] + src34[282] + src34[283] + src34[284] + src34[285] + src34[286] + src34[287] + src34[288] + src34[289] + src34[290] + src34[291] + src34[292] + src34[293] + src34[294] + src34[295] + src34[296] + src34[297] + src34[298] + src34[299] + src34[300] + src34[301] + src34[302] + src34[303] + src34[304] + src34[305] + src34[306] + src34[307] + src34[308] + src34[309] + src34[310] + src34[311] + src34[312] + src34[313] + src34[314] + src34[315] + src34[316] + src34[317] + src34[318] + src34[319] + src34[320] + src34[321] + src34[322] + src34[323] + src34[324] + src34[325] + src34[326] + src34[327] + src34[328] + src34[329] + src34[330] + src34[331] + src34[332] + src34[333] + src34[334] + src34[335] + src34[336] + src34[337] + src34[338] + src34[339] + src34[340] + src34[341] + src34[342] + src34[343] + src34[344] + src34[345] + src34[346] + src34[347] + src34[348] + src34[349] + src34[350] + src34[351] + src34[352] + src34[353] + src34[354] + src34[355] + src34[356] + src34[357] + src34[358] + src34[359] + src34[360] + src34[361] + src34[362] + src34[363] + src34[364] + src34[365] + src34[366] + src34[367] + src34[368] + src34[369] + src34[370] + src34[371] + src34[372] + src34[373] + src34[374] + src34[375] + src34[376] + src34[377] + src34[378] + src34[379] + src34[380] + src34[381] + src34[382] + src34[383] + src34[384] + src34[385] + src34[386] + src34[387] + src34[388] + src34[389] + src34[390] + src34[391] + src34[392] + src34[393] + src34[394] + src34[395] + src34[396] + src34[397] + src34[398] + src34[399] + src34[400] + src34[401] + src34[402] + src34[403] + src34[404] + src34[405] + src34[406] + src34[407] + src34[408] + src34[409] + src34[410] + src34[411] + src34[412] + src34[413] + src34[414] + src34[415] + src34[416] + src34[417] + src34[418] + src34[419] + src34[420] + src34[421] + src34[422] + src34[423] + src34[424] + src34[425] + src34[426] + src34[427] + src34[428] + src34[429] + src34[430] + src34[431] + src34[432] + src34[433] + src34[434] + src34[435] + src34[436] + src34[437] + src34[438] + src34[439] + src34[440] + src34[441] + src34[442] + src34[443] + src34[444] + src34[445] + src34[446] + src34[447] + src34[448] + src34[449] + src34[450] + src34[451] + src34[452] + src34[453] + src34[454] + src34[455] + src34[456] + src34[457] + src34[458] + src34[459] + src34[460] + src34[461] + src34[462] + src34[463] + src34[464] + src34[465] + src34[466] + src34[467] + src34[468] + src34[469] + src34[470] + src34[471] + src34[472] + src34[473] + src34[474] + src34[475] + src34[476] + src34[477] + src34[478] + src34[479] + src34[480] + src34[481] + src34[482] + src34[483] + src34[484] + src34[485])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63] + src35[64] + src35[65] + src35[66] + src35[67] + src35[68] + src35[69] + src35[70] + src35[71] + src35[72] + src35[73] + src35[74] + src35[75] + src35[76] + src35[77] + src35[78] + src35[79] + src35[80] + src35[81] + src35[82] + src35[83] + src35[84] + src35[85] + src35[86] + src35[87] + src35[88] + src35[89] + src35[90] + src35[91] + src35[92] + src35[93] + src35[94] + src35[95] + src35[96] + src35[97] + src35[98] + src35[99] + src35[100] + src35[101] + src35[102] + src35[103] + src35[104] + src35[105] + src35[106] + src35[107] + src35[108] + src35[109] + src35[110] + src35[111] + src35[112] + src35[113] + src35[114] + src35[115] + src35[116] + src35[117] + src35[118] + src35[119] + src35[120] + src35[121] + src35[122] + src35[123] + src35[124] + src35[125] + src35[126] + src35[127] + src35[128] + src35[129] + src35[130] + src35[131] + src35[132] + src35[133] + src35[134] + src35[135] + src35[136] + src35[137] + src35[138] + src35[139] + src35[140] + src35[141] + src35[142] + src35[143] + src35[144] + src35[145] + src35[146] + src35[147] + src35[148] + src35[149] + src35[150] + src35[151] + src35[152] + src35[153] + src35[154] + src35[155] + src35[156] + src35[157] + src35[158] + src35[159] + src35[160] + src35[161] + src35[162] + src35[163] + src35[164] + src35[165] + src35[166] + src35[167] + src35[168] + src35[169] + src35[170] + src35[171] + src35[172] + src35[173] + src35[174] + src35[175] + src35[176] + src35[177] + src35[178] + src35[179] + src35[180] + src35[181] + src35[182] + src35[183] + src35[184] + src35[185] + src35[186] + src35[187] + src35[188] + src35[189] + src35[190] + src35[191] + src35[192] + src35[193] + src35[194] + src35[195] + src35[196] + src35[197] + src35[198] + src35[199] + src35[200] + src35[201] + src35[202] + src35[203] + src35[204] + src35[205] + src35[206] + src35[207] + src35[208] + src35[209] + src35[210] + src35[211] + src35[212] + src35[213] + src35[214] + src35[215] + src35[216] + src35[217] + src35[218] + src35[219] + src35[220] + src35[221] + src35[222] + src35[223] + src35[224] + src35[225] + src35[226] + src35[227] + src35[228] + src35[229] + src35[230] + src35[231] + src35[232] + src35[233] + src35[234] + src35[235] + src35[236] + src35[237] + src35[238] + src35[239] + src35[240] + src35[241] + src35[242] + src35[243] + src35[244] + src35[245] + src35[246] + src35[247] + src35[248] + src35[249] + src35[250] + src35[251] + src35[252] + src35[253] + src35[254] + src35[255] + src35[256] + src35[257] + src35[258] + src35[259] + src35[260] + src35[261] + src35[262] + src35[263] + src35[264] + src35[265] + src35[266] + src35[267] + src35[268] + src35[269] + src35[270] + src35[271] + src35[272] + src35[273] + src35[274] + src35[275] + src35[276] + src35[277] + src35[278] + src35[279] + src35[280] + src35[281] + src35[282] + src35[283] + src35[284] + src35[285] + src35[286] + src35[287] + src35[288] + src35[289] + src35[290] + src35[291] + src35[292] + src35[293] + src35[294] + src35[295] + src35[296] + src35[297] + src35[298] + src35[299] + src35[300] + src35[301] + src35[302] + src35[303] + src35[304] + src35[305] + src35[306] + src35[307] + src35[308] + src35[309] + src35[310] + src35[311] + src35[312] + src35[313] + src35[314] + src35[315] + src35[316] + src35[317] + src35[318] + src35[319] + src35[320] + src35[321] + src35[322] + src35[323] + src35[324] + src35[325] + src35[326] + src35[327] + src35[328] + src35[329] + src35[330] + src35[331] + src35[332] + src35[333] + src35[334] + src35[335] + src35[336] + src35[337] + src35[338] + src35[339] + src35[340] + src35[341] + src35[342] + src35[343] + src35[344] + src35[345] + src35[346] + src35[347] + src35[348] + src35[349] + src35[350] + src35[351] + src35[352] + src35[353] + src35[354] + src35[355] + src35[356] + src35[357] + src35[358] + src35[359] + src35[360] + src35[361] + src35[362] + src35[363] + src35[364] + src35[365] + src35[366] + src35[367] + src35[368] + src35[369] + src35[370] + src35[371] + src35[372] + src35[373] + src35[374] + src35[375] + src35[376] + src35[377] + src35[378] + src35[379] + src35[380] + src35[381] + src35[382] + src35[383] + src35[384] + src35[385] + src35[386] + src35[387] + src35[388] + src35[389] + src35[390] + src35[391] + src35[392] + src35[393] + src35[394] + src35[395] + src35[396] + src35[397] + src35[398] + src35[399] + src35[400] + src35[401] + src35[402] + src35[403] + src35[404] + src35[405] + src35[406] + src35[407] + src35[408] + src35[409] + src35[410] + src35[411] + src35[412] + src35[413] + src35[414] + src35[415] + src35[416] + src35[417] + src35[418] + src35[419] + src35[420] + src35[421] + src35[422] + src35[423] + src35[424] + src35[425] + src35[426] + src35[427] + src35[428] + src35[429] + src35[430] + src35[431] + src35[432] + src35[433] + src35[434] + src35[435] + src35[436] + src35[437] + src35[438] + src35[439] + src35[440] + src35[441] + src35[442] + src35[443] + src35[444] + src35[445] + src35[446] + src35[447] + src35[448] + src35[449] + src35[450] + src35[451] + src35[452] + src35[453] + src35[454] + src35[455] + src35[456] + src35[457] + src35[458] + src35[459] + src35[460] + src35[461] + src35[462] + src35[463] + src35[464] + src35[465] + src35[466] + src35[467] + src35[468] + src35[469] + src35[470] + src35[471] + src35[472] + src35[473] + src35[474] + src35[475] + src35[476] + src35[477] + src35[478] + src35[479] + src35[480] + src35[481] + src35[482] + src35[483] + src35[484] + src35[485])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63] + src36[64] + src36[65] + src36[66] + src36[67] + src36[68] + src36[69] + src36[70] + src36[71] + src36[72] + src36[73] + src36[74] + src36[75] + src36[76] + src36[77] + src36[78] + src36[79] + src36[80] + src36[81] + src36[82] + src36[83] + src36[84] + src36[85] + src36[86] + src36[87] + src36[88] + src36[89] + src36[90] + src36[91] + src36[92] + src36[93] + src36[94] + src36[95] + src36[96] + src36[97] + src36[98] + src36[99] + src36[100] + src36[101] + src36[102] + src36[103] + src36[104] + src36[105] + src36[106] + src36[107] + src36[108] + src36[109] + src36[110] + src36[111] + src36[112] + src36[113] + src36[114] + src36[115] + src36[116] + src36[117] + src36[118] + src36[119] + src36[120] + src36[121] + src36[122] + src36[123] + src36[124] + src36[125] + src36[126] + src36[127] + src36[128] + src36[129] + src36[130] + src36[131] + src36[132] + src36[133] + src36[134] + src36[135] + src36[136] + src36[137] + src36[138] + src36[139] + src36[140] + src36[141] + src36[142] + src36[143] + src36[144] + src36[145] + src36[146] + src36[147] + src36[148] + src36[149] + src36[150] + src36[151] + src36[152] + src36[153] + src36[154] + src36[155] + src36[156] + src36[157] + src36[158] + src36[159] + src36[160] + src36[161] + src36[162] + src36[163] + src36[164] + src36[165] + src36[166] + src36[167] + src36[168] + src36[169] + src36[170] + src36[171] + src36[172] + src36[173] + src36[174] + src36[175] + src36[176] + src36[177] + src36[178] + src36[179] + src36[180] + src36[181] + src36[182] + src36[183] + src36[184] + src36[185] + src36[186] + src36[187] + src36[188] + src36[189] + src36[190] + src36[191] + src36[192] + src36[193] + src36[194] + src36[195] + src36[196] + src36[197] + src36[198] + src36[199] + src36[200] + src36[201] + src36[202] + src36[203] + src36[204] + src36[205] + src36[206] + src36[207] + src36[208] + src36[209] + src36[210] + src36[211] + src36[212] + src36[213] + src36[214] + src36[215] + src36[216] + src36[217] + src36[218] + src36[219] + src36[220] + src36[221] + src36[222] + src36[223] + src36[224] + src36[225] + src36[226] + src36[227] + src36[228] + src36[229] + src36[230] + src36[231] + src36[232] + src36[233] + src36[234] + src36[235] + src36[236] + src36[237] + src36[238] + src36[239] + src36[240] + src36[241] + src36[242] + src36[243] + src36[244] + src36[245] + src36[246] + src36[247] + src36[248] + src36[249] + src36[250] + src36[251] + src36[252] + src36[253] + src36[254] + src36[255] + src36[256] + src36[257] + src36[258] + src36[259] + src36[260] + src36[261] + src36[262] + src36[263] + src36[264] + src36[265] + src36[266] + src36[267] + src36[268] + src36[269] + src36[270] + src36[271] + src36[272] + src36[273] + src36[274] + src36[275] + src36[276] + src36[277] + src36[278] + src36[279] + src36[280] + src36[281] + src36[282] + src36[283] + src36[284] + src36[285] + src36[286] + src36[287] + src36[288] + src36[289] + src36[290] + src36[291] + src36[292] + src36[293] + src36[294] + src36[295] + src36[296] + src36[297] + src36[298] + src36[299] + src36[300] + src36[301] + src36[302] + src36[303] + src36[304] + src36[305] + src36[306] + src36[307] + src36[308] + src36[309] + src36[310] + src36[311] + src36[312] + src36[313] + src36[314] + src36[315] + src36[316] + src36[317] + src36[318] + src36[319] + src36[320] + src36[321] + src36[322] + src36[323] + src36[324] + src36[325] + src36[326] + src36[327] + src36[328] + src36[329] + src36[330] + src36[331] + src36[332] + src36[333] + src36[334] + src36[335] + src36[336] + src36[337] + src36[338] + src36[339] + src36[340] + src36[341] + src36[342] + src36[343] + src36[344] + src36[345] + src36[346] + src36[347] + src36[348] + src36[349] + src36[350] + src36[351] + src36[352] + src36[353] + src36[354] + src36[355] + src36[356] + src36[357] + src36[358] + src36[359] + src36[360] + src36[361] + src36[362] + src36[363] + src36[364] + src36[365] + src36[366] + src36[367] + src36[368] + src36[369] + src36[370] + src36[371] + src36[372] + src36[373] + src36[374] + src36[375] + src36[376] + src36[377] + src36[378] + src36[379] + src36[380] + src36[381] + src36[382] + src36[383] + src36[384] + src36[385] + src36[386] + src36[387] + src36[388] + src36[389] + src36[390] + src36[391] + src36[392] + src36[393] + src36[394] + src36[395] + src36[396] + src36[397] + src36[398] + src36[399] + src36[400] + src36[401] + src36[402] + src36[403] + src36[404] + src36[405] + src36[406] + src36[407] + src36[408] + src36[409] + src36[410] + src36[411] + src36[412] + src36[413] + src36[414] + src36[415] + src36[416] + src36[417] + src36[418] + src36[419] + src36[420] + src36[421] + src36[422] + src36[423] + src36[424] + src36[425] + src36[426] + src36[427] + src36[428] + src36[429] + src36[430] + src36[431] + src36[432] + src36[433] + src36[434] + src36[435] + src36[436] + src36[437] + src36[438] + src36[439] + src36[440] + src36[441] + src36[442] + src36[443] + src36[444] + src36[445] + src36[446] + src36[447] + src36[448] + src36[449] + src36[450] + src36[451] + src36[452] + src36[453] + src36[454] + src36[455] + src36[456] + src36[457] + src36[458] + src36[459] + src36[460] + src36[461] + src36[462] + src36[463] + src36[464] + src36[465] + src36[466] + src36[467] + src36[468] + src36[469] + src36[470] + src36[471] + src36[472] + src36[473] + src36[474] + src36[475] + src36[476] + src36[477] + src36[478] + src36[479] + src36[480] + src36[481] + src36[482] + src36[483] + src36[484] + src36[485])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63] + src37[64] + src37[65] + src37[66] + src37[67] + src37[68] + src37[69] + src37[70] + src37[71] + src37[72] + src37[73] + src37[74] + src37[75] + src37[76] + src37[77] + src37[78] + src37[79] + src37[80] + src37[81] + src37[82] + src37[83] + src37[84] + src37[85] + src37[86] + src37[87] + src37[88] + src37[89] + src37[90] + src37[91] + src37[92] + src37[93] + src37[94] + src37[95] + src37[96] + src37[97] + src37[98] + src37[99] + src37[100] + src37[101] + src37[102] + src37[103] + src37[104] + src37[105] + src37[106] + src37[107] + src37[108] + src37[109] + src37[110] + src37[111] + src37[112] + src37[113] + src37[114] + src37[115] + src37[116] + src37[117] + src37[118] + src37[119] + src37[120] + src37[121] + src37[122] + src37[123] + src37[124] + src37[125] + src37[126] + src37[127] + src37[128] + src37[129] + src37[130] + src37[131] + src37[132] + src37[133] + src37[134] + src37[135] + src37[136] + src37[137] + src37[138] + src37[139] + src37[140] + src37[141] + src37[142] + src37[143] + src37[144] + src37[145] + src37[146] + src37[147] + src37[148] + src37[149] + src37[150] + src37[151] + src37[152] + src37[153] + src37[154] + src37[155] + src37[156] + src37[157] + src37[158] + src37[159] + src37[160] + src37[161] + src37[162] + src37[163] + src37[164] + src37[165] + src37[166] + src37[167] + src37[168] + src37[169] + src37[170] + src37[171] + src37[172] + src37[173] + src37[174] + src37[175] + src37[176] + src37[177] + src37[178] + src37[179] + src37[180] + src37[181] + src37[182] + src37[183] + src37[184] + src37[185] + src37[186] + src37[187] + src37[188] + src37[189] + src37[190] + src37[191] + src37[192] + src37[193] + src37[194] + src37[195] + src37[196] + src37[197] + src37[198] + src37[199] + src37[200] + src37[201] + src37[202] + src37[203] + src37[204] + src37[205] + src37[206] + src37[207] + src37[208] + src37[209] + src37[210] + src37[211] + src37[212] + src37[213] + src37[214] + src37[215] + src37[216] + src37[217] + src37[218] + src37[219] + src37[220] + src37[221] + src37[222] + src37[223] + src37[224] + src37[225] + src37[226] + src37[227] + src37[228] + src37[229] + src37[230] + src37[231] + src37[232] + src37[233] + src37[234] + src37[235] + src37[236] + src37[237] + src37[238] + src37[239] + src37[240] + src37[241] + src37[242] + src37[243] + src37[244] + src37[245] + src37[246] + src37[247] + src37[248] + src37[249] + src37[250] + src37[251] + src37[252] + src37[253] + src37[254] + src37[255] + src37[256] + src37[257] + src37[258] + src37[259] + src37[260] + src37[261] + src37[262] + src37[263] + src37[264] + src37[265] + src37[266] + src37[267] + src37[268] + src37[269] + src37[270] + src37[271] + src37[272] + src37[273] + src37[274] + src37[275] + src37[276] + src37[277] + src37[278] + src37[279] + src37[280] + src37[281] + src37[282] + src37[283] + src37[284] + src37[285] + src37[286] + src37[287] + src37[288] + src37[289] + src37[290] + src37[291] + src37[292] + src37[293] + src37[294] + src37[295] + src37[296] + src37[297] + src37[298] + src37[299] + src37[300] + src37[301] + src37[302] + src37[303] + src37[304] + src37[305] + src37[306] + src37[307] + src37[308] + src37[309] + src37[310] + src37[311] + src37[312] + src37[313] + src37[314] + src37[315] + src37[316] + src37[317] + src37[318] + src37[319] + src37[320] + src37[321] + src37[322] + src37[323] + src37[324] + src37[325] + src37[326] + src37[327] + src37[328] + src37[329] + src37[330] + src37[331] + src37[332] + src37[333] + src37[334] + src37[335] + src37[336] + src37[337] + src37[338] + src37[339] + src37[340] + src37[341] + src37[342] + src37[343] + src37[344] + src37[345] + src37[346] + src37[347] + src37[348] + src37[349] + src37[350] + src37[351] + src37[352] + src37[353] + src37[354] + src37[355] + src37[356] + src37[357] + src37[358] + src37[359] + src37[360] + src37[361] + src37[362] + src37[363] + src37[364] + src37[365] + src37[366] + src37[367] + src37[368] + src37[369] + src37[370] + src37[371] + src37[372] + src37[373] + src37[374] + src37[375] + src37[376] + src37[377] + src37[378] + src37[379] + src37[380] + src37[381] + src37[382] + src37[383] + src37[384] + src37[385] + src37[386] + src37[387] + src37[388] + src37[389] + src37[390] + src37[391] + src37[392] + src37[393] + src37[394] + src37[395] + src37[396] + src37[397] + src37[398] + src37[399] + src37[400] + src37[401] + src37[402] + src37[403] + src37[404] + src37[405] + src37[406] + src37[407] + src37[408] + src37[409] + src37[410] + src37[411] + src37[412] + src37[413] + src37[414] + src37[415] + src37[416] + src37[417] + src37[418] + src37[419] + src37[420] + src37[421] + src37[422] + src37[423] + src37[424] + src37[425] + src37[426] + src37[427] + src37[428] + src37[429] + src37[430] + src37[431] + src37[432] + src37[433] + src37[434] + src37[435] + src37[436] + src37[437] + src37[438] + src37[439] + src37[440] + src37[441] + src37[442] + src37[443] + src37[444] + src37[445] + src37[446] + src37[447] + src37[448] + src37[449] + src37[450] + src37[451] + src37[452] + src37[453] + src37[454] + src37[455] + src37[456] + src37[457] + src37[458] + src37[459] + src37[460] + src37[461] + src37[462] + src37[463] + src37[464] + src37[465] + src37[466] + src37[467] + src37[468] + src37[469] + src37[470] + src37[471] + src37[472] + src37[473] + src37[474] + src37[475] + src37[476] + src37[477] + src37[478] + src37[479] + src37[480] + src37[481] + src37[482] + src37[483] + src37[484] + src37[485])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63] + src38[64] + src38[65] + src38[66] + src38[67] + src38[68] + src38[69] + src38[70] + src38[71] + src38[72] + src38[73] + src38[74] + src38[75] + src38[76] + src38[77] + src38[78] + src38[79] + src38[80] + src38[81] + src38[82] + src38[83] + src38[84] + src38[85] + src38[86] + src38[87] + src38[88] + src38[89] + src38[90] + src38[91] + src38[92] + src38[93] + src38[94] + src38[95] + src38[96] + src38[97] + src38[98] + src38[99] + src38[100] + src38[101] + src38[102] + src38[103] + src38[104] + src38[105] + src38[106] + src38[107] + src38[108] + src38[109] + src38[110] + src38[111] + src38[112] + src38[113] + src38[114] + src38[115] + src38[116] + src38[117] + src38[118] + src38[119] + src38[120] + src38[121] + src38[122] + src38[123] + src38[124] + src38[125] + src38[126] + src38[127] + src38[128] + src38[129] + src38[130] + src38[131] + src38[132] + src38[133] + src38[134] + src38[135] + src38[136] + src38[137] + src38[138] + src38[139] + src38[140] + src38[141] + src38[142] + src38[143] + src38[144] + src38[145] + src38[146] + src38[147] + src38[148] + src38[149] + src38[150] + src38[151] + src38[152] + src38[153] + src38[154] + src38[155] + src38[156] + src38[157] + src38[158] + src38[159] + src38[160] + src38[161] + src38[162] + src38[163] + src38[164] + src38[165] + src38[166] + src38[167] + src38[168] + src38[169] + src38[170] + src38[171] + src38[172] + src38[173] + src38[174] + src38[175] + src38[176] + src38[177] + src38[178] + src38[179] + src38[180] + src38[181] + src38[182] + src38[183] + src38[184] + src38[185] + src38[186] + src38[187] + src38[188] + src38[189] + src38[190] + src38[191] + src38[192] + src38[193] + src38[194] + src38[195] + src38[196] + src38[197] + src38[198] + src38[199] + src38[200] + src38[201] + src38[202] + src38[203] + src38[204] + src38[205] + src38[206] + src38[207] + src38[208] + src38[209] + src38[210] + src38[211] + src38[212] + src38[213] + src38[214] + src38[215] + src38[216] + src38[217] + src38[218] + src38[219] + src38[220] + src38[221] + src38[222] + src38[223] + src38[224] + src38[225] + src38[226] + src38[227] + src38[228] + src38[229] + src38[230] + src38[231] + src38[232] + src38[233] + src38[234] + src38[235] + src38[236] + src38[237] + src38[238] + src38[239] + src38[240] + src38[241] + src38[242] + src38[243] + src38[244] + src38[245] + src38[246] + src38[247] + src38[248] + src38[249] + src38[250] + src38[251] + src38[252] + src38[253] + src38[254] + src38[255] + src38[256] + src38[257] + src38[258] + src38[259] + src38[260] + src38[261] + src38[262] + src38[263] + src38[264] + src38[265] + src38[266] + src38[267] + src38[268] + src38[269] + src38[270] + src38[271] + src38[272] + src38[273] + src38[274] + src38[275] + src38[276] + src38[277] + src38[278] + src38[279] + src38[280] + src38[281] + src38[282] + src38[283] + src38[284] + src38[285] + src38[286] + src38[287] + src38[288] + src38[289] + src38[290] + src38[291] + src38[292] + src38[293] + src38[294] + src38[295] + src38[296] + src38[297] + src38[298] + src38[299] + src38[300] + src38[301] + src38[302] + src38[303] + src38[304] + src38[305] + src38[306] + src38[307] + src38[308] + src38[309] + src38[310] + src38[311] + src38[312] + src38[313] + src38[314] + src38[315] + src38[316] + src38[317] + src38[318] + src38[319] + src38[320] + src38[321] + src38[322] + src38[323] + src38[324] + src38[325] + src38[326] + src38[327] + src38[328] + src38[329] + src38[330] + src38[331] + src38[332] + src38[333] + src38[334] + src38[335] + src38[336] + src38[337] + src38[338] + src38[339] + src38[340] + src38[341] + src38[342] + src38[343] + src38[344] + src38[345] + src38[346] + src38[347] + src38[348] + src38[349] + src38[350] + src38[351] + src38[352] + src38[353] + src38[354] + src38[355] + src38[356] + src38[357] + src38[358] + src38[359] + src38[360] + src38[361] + src38[362] + src38[363] + src38[364] + src38[365] + src38[366] + src38[367] + src38[368] + src38[369] + src38[370] + src38[371] + src38[372] + src38[373] + src38[374] + src38[375] + src38[376] + src38[377] + src38[378] + src38[379] + src38[380] + src38[381] + src38[382] + src38[383] + src38[384] + src38[385] + src38[386] + src38[387] + src38[388] + src38[389] + src38[390] + src38[391] + src38[392] + src38[393] + src38[394] + src38[395] + src38[396] + src38[397] + src38[398] + src38[399] + src38[400] + src38[401] + src38[402] + src38[403] + src38[404] + src38[405] + src38[406] + src38[407] + src38[408] + src38[409] + src38[410] + src38[411] + src38[412] + src38[413] + src38[414] + src38[415] + src38[416] + src38[417] + src38[418] + src38[419] + src38[420] + src38[421] + src38[422] + src38[423] + src38[424] + src38[425] + src38[426] + src38[427] + src38[428] + src38[429] + src38[430] + src38[431] + src38[432] + src38[433] + src38[434] + src38[435] + src38[436] + src38[437] + src38[438] + src38[439] + src38[440] + src38[441] + src38[442] + src38[443] + src38[444] + src38[445] + src38[446] + src38[447] + src38[448] + src38[449] + src38[450] + src38[451] + src38[452] + src38[453] + src38[454] + src38[455] + src38[456] + src38[457] + src38[458] + src38[459] + src38[460] + src38[461] + src38[462] + src38[463] + src38[464] + src38[465] + src38[466] + src38[467] + src38[468] + src38[469] + src38[470] + src38[471] + src38[472] + src38[473] + src38[474] + src38[475] + src38[476] + src38[477] + src38[478] + src38[479] + src38[480] + src38[481] + src38[482] + src38[483] + src38[484] + src38[485])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63] + src39[64] + src39[65] + src39[66] + src39[67] + src39[68] + src39[69] + src39[70] + src39[71] + src39[72] + src39[73] + src39[74] + src39[75] + src39[76] + src39[77] + src39[78] + src39[79] + src39[80] + src39[81] + src39[82] + src39[83] + src39[84] + src39[85] + src39[86] + src39[87] + src39[88] + src39[89] + src39[90] + src39[91] + src39[92] + src39[93] + src39[94] + src39[95] + src39[96] + src39[97] + src39[98] + src39[99] + src39[100] + src39[101] + src39[102] + src39[103] + src39[104] + src39[105] + src39[106] + src39[107] + src39[108] + src39[109] + src39[110] + src39[111] + src39[112] + src39[113] + src39[114] + src39[115] + src39[116] + src39[117] + src39[118] + src39[119] + src39[120] + src39[121] + src39[122] + src39[123] + src39[124] + src39[125] + src39[126] + src39[127] + src39[128] + src39[129] + src39[130] + src39[131] + src39[132] + src39[133] + src39[134] + src39[135] + src39[136] + src39[137] + src39[138] + src39[139] + src39[140] + src39[141] + src39[142] + src39[143] + src39[144] + src39[145] + src39[146] + src39[147] + src39[148] + src39[149] + src39[150] + src39[151] + src39[152] + src39[153] + src39[154] + src39[155] + src39[156] + src39[157] + src39[158] + src39[159] + src39[160] + src39[161] + src39[162] + src39[163] + src39[164] + src39[165] + src39[166] + src39[167] + src39[168] + src39[169] + src39[170] + src39[171] + src39[172] + src39[173] + src39[174] + src39[175] + src39[176] + src39[177] + src39[178] + src39[179] + src39[180] + src39[181] + src39[182] + src39[183] + src39[184] + src39[185] + src39[186] + src39[187] + src39[188] + src39[189] + src39[190] + src39[191] + src39[192] + src39[193] + src39[194] + src39[195] + src39[196] + src39[197] + src39[198] + src39[199] + src39[200] + src39[201] + src39[202] + src39[203] + src39[204] + src39[205] + src39[206] + src39[207] + src39[208] + src39[209] + src39[210] + src39[211] + src39[212] + src39[213] + src39[214] + src39[215] + src39[216] + src39[217] + src39[218] + src39[219] + src39[220] + src39[221] + src39[222] + src39[223] + src39[224] + src39[225] + src39[226] + src39[227] + src39[228] + src39[229] + src39[230] + src39[231] + src39[232] + src39[233] + src39[234] + src39[235] + src39[236] + src39[237] + src39[238] + src39[239] + src39[240] + src39[241] + src39[242] + src39[243] + src39[244] + src39[245] + src39[246] + src39[247] + src39[248] + src39[249] + src39[250] + src39[251] + src39[252] + src39[253] + src39[254] + src39[255] + src39[256] + src39[257] + src39[258] + src39[259] + src39[260] + src39[261] + src39[262] + src39[263] + src39[264] + src39[265] + src39[266] + src39[267] + src39[268] + src39[269] + src39[270] + src39[271] + src39[272] + src39[273] + src39[274] + src39[275] + src39[276] + src39[277] + src39[278] + src39[279] + src39[280] + src39[281] + src39[282] + src39[283] + src39[284] + src39[285] + src39[286] + src39[287] + src39[288] + src39[289] + src39[290] + src39[291] + src39[292] + src39[293] + src39[294] + src39[295] + src39[296] + src39[297] + src39[298] + src39[299] + src39[300] + src39[301] + src39[302] + src39[303] + src39[304] + src39[305] + src39[306] + src39[307] + src39[308] + src39[309] + src39[310] + src39[311] + src39[312] + src39[313] + src39[314] + src39[315] + src39[316] + src39[317] + src39[318] + src39[319] + src39[320] + src39[321] + src39[322] + src39[323] + src39[324] + src39[325] + src39[326] + src39[327] + src39[328] + src39[329] + src39[330] + src39[331] + src39[332] + src39[333] + src39[334] + src39[335] + src39[336] + src39[337] + src39[338] + src39[339] + src39[340] + src39[341] + src39[342] + src39[343] + src39[344] + src39[345] + src39[346] + src39[347] + src39[348] + src39[349] + src39[350] + src39[351] + src39[352] + src39[353] + src39[354] + src39[355] + src39[356] + src39[357] + src39[358] + src39[359] + src39[360] + src39[361] + src39[362] + src39[363] + src39[364] + src39[365] + src39[366] + src39[367] + src39[368] + src39[369] + src39[370] + src39[371] + src39[372] + src39[373] + src39[374] + src39[375] + src39[376] + src39[377] + src39[378] + src39[379] + src39[380] + src39[381] + src39[382] + src39[383] + src39[384] + src39[385] + src39[386] + src39[387] + src39[388] + src39[389] + src39[390] + src39[391] + src39[392] + src39[393] + src39[394] + src39[395] + src39[396] + src39[397] + src39[398] + src39[399] + src39[400] + src39[401] + src39[402] + src39[403] + src39[404] + src39[405] + src39[406] + src39[407] + src39[408] + src39[409] + src39[410] + src39[411] + src39[412] + src39[413] + src39[414] + src39[415] + src39[416] + src39[417] + src39[418] + src39[419] + src39[420] + src39[421] + src39[422] + src39[423] + src39[424] + src39[425] + src39[426] + src39[427] + src39[428] + src39[429] + src39[430] + src39[431] + src39[432] + src39[433] + src39[434] + src39[435] + src39[436] + src39[437] + src39[438] + src39[439] + src39[440] + src39[441] + src39[442] + src39[443] + src39[444] + src39[445] + src39[446] + src39[447] + src39[448] + src39[449] + src39[450] + src39[451] + src39[452] + src39[453] + src39[454] + src39[455] + src39[456] + src39[457] + src39[458] + src39[459] + src39[460] + src39[461] + src39[462] + src39[463] + src39[464] + src39[465] + src39[466] + src39[467] + src39[468] + src39[469] + src39[470] + src39[471] + src39[472] + src39[473] + src39[474] + src39[475] + src39[476] + src39[477] + src39[478] + src39[479] + src39[480] + src39[481] + src39[482] + src39[483] + src39[484] + src39[485])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63] + src40[64] + src40[65] + src40[66] + src40[67] + src40[68] + src40[69] + src40[70] + src40[71] + src40[72] + src40[73] + src40[74] + src40[75] + src40[76] + src40[77] + src40[78] + src40[79] + src40[80] + src40[81] + src40[82] + src40[83] + src40[84] + src40[85] + src40[86] + src40[87] + src40[88] + src40[89] + src40[90] + src40[91] + src40[92] + src40[93] + src40[94] + src40[95] + src40[96] + src40[97] + src40[98] + src40[99] + src40[100] + src40[101] + src40[102] + src40[103] + src40[104] + src40[105] + src40[106] + src40[107] + src40[108] + src40[109] + src40[110] + src40[111] + src40[112] + src40[113] + src40[114] + src40[115] + src40[116] + src40[117] + src40[118] + src40[119] + src40[120] + src40[121] + src40[122] + src40[123] + src40[124] + src40[125] + src40[126] + src40[127] + src40[128] + src40[129] + src40[130] + src40[131] + src40[132] + src40[133] + src40[134] + src40[135] + src40[136] + src40[137] + src40[138] + src40[139] + src40[140] + src40[141] + src40[142] + src40[143] + src40[144] + src40[145] + src40[146] + src40[147] + src40[148] + src40[149] + src40[150] + src40[151] + src40[152] + src40[153] + src40[154] + src40[155] + src40[156] + src40[157] + src40[158] + src40[159] + src40[160] + src40[161] + src40[162] + src40[163] + src40[164] + src40[165] + src40[166] + src40[167] + src40[168] + src40[169] + src40[170] + src40[171] + src40[172] + src40[173] + src40[174] + src40[175] + src40[176] + src40[177] + src40[178] + src40[179] + src40[180] + src40[181] + src40[182] + src40[183] + src40[184] + src40[185] + src40[186] + src40[187] + src40[188] + src40[189] + src40[190] + src40[191] + src40[192] + src40[193] + src40[194] + src40[195] + src40[196] + src40[197] + src40[198] + src40[199] + src40[200] + src40[201] + src40[202] + src40[203] + src40[204] + src40[205] + src40[206] + src40[207] + src40[208] + src40[209] + src40[210] + src40[211] + src40[212] + src40[213] + src40[214] + src40[215] + src40[216] + src40[217] + src40[218] + src40[219] + src40[220] + src40[221] + src40[222] + src40[223] + src40[224] + src40[225] + src40[226] + src40[227] + src40[228] + src40[229] + src40[230] + src40[231] + src40[232] + src40[233] + src40[234] + src40[235] + src40[236] + src40[237] + src40[238] + src40[239] + src40[240] + src40[241] + src40[242] + src40[243] + src40[244] + src40[245] + src40[246] + src40[247] + src40[248] + src40[249] + src40[250] + src40[251] + src40[252] + src40[253] + src40[254] + src40[255] + src40[256] + src40[257] + src40[258] + src40[259] + src40[260] + src40[261] + src40[262] + src40[263] + src40[264] + src40[265] + src40[266] + src40[267] + src40[268] + src40[269] + src40[270] + src40[271] + src40[272] + src40[273] + src40[274] + src40[275] + src40[276] + src40[277] + src40[278] + src40[279] + src40[280] + src40[281] + src40[282] + src40[283] + src40[284] + src40[285] + src40[286] + src40[287] + src40[288] + src40[289] + src40[290] + src40[291] + src40[292] + src40[293] + src40[294] + src40[295] + src40[296] + src40[297] + src40[298] + src40[299] + src40[300] + src40[301] + src40[302] + src40[303] + src40[304] + src40[305] + src40[306] + src40[307] + src40[308] + src40[309] + src40[310] + src40[311] + src40[312] + src40[313] + src40[314] + src40[315] + src40[316] + src40[317] + src40[318] + src40[319] + src40[320] + src40[321] + src40[322] + src40[323] + src40[324] + src40[325] + src40[326] + src40[327] + src40[328] + src40[329] + src40[330] + src40[331] + src40[332] + src40[333] + src40[334] + src40[335] + src40[336] + src40[337] + src40[338] + src40[339] + src40[340] + src40[341] + src40[342] + src40[343] + src40[344] + src40[345] + src40[346] + src40[347] + src40[348] + src40[349] + src40[350] + src40[351] + src40[352] + src40[353] + src40[354] + src40[355] + src40[356] + src40[357] + src40[358] + src40[359] + src40[360] + src40[361] + src40[362] + src40[363] + src40[364] + src40[365] + src40[366] + src40[367] + src40[368] + src40[369] + src40[370] + src40[371] + src40[372] + src40[373] + src40[374] + src40[375] + src40[376] + src40[377] + src40[378] + src40[379] + src40[380] + src40[381] + src40[382] + src40[383] + src40[384] + src40[385] + src40[386] + src40[387] + src40[388] + src40[389] + src40[390] + src40[391] + src40[392] + src40[393] + src40[394] + src40[395] + src40[396] + src40[397] + src40[398] + src40[399] + src40[400] + src40[401] + src40[402] + src40[403] + src40[404] + src40[405] + src40[406] + src40[407] + src40[408] + src40[409] + src40[410] + src40[411] + src40[412] + src40[413] + src40[414] + src40[415] + src40[416] + src40[417] + src40[418] + src40[419] + src40[420] + src40[421] + src40[422] + src40[423] + src40[424] + src40[425] + src40[426] + src40[427] + src40[428] + src40[429] + src40[430] + src40[431] + src40[432] + src40[433] + src40[434] + src40[435] + src40[436] + src40[437] + src40[438] + src40[439] + src40[440] + src40[441] + src40[442] + src40[443] + src40[444] + src40[445] + src40[446] + src40[447] + src40[448] + src40[449] + src40[450] + src40[451] + src40[452] + src40[453] + src40[454] + src40[455] + src40[456] + src40[457] + src40[458] + src40[459] + src40[460] + src40[461] + src40[462] + src40[463] + src40[464] + src40[465] + src40[466] + src40[467] + src40[468] + src40[469] + src40[470] + src40[471] + src40[472] + src40[473] + src40[474] + src40[475] + src40[476] + src40[477] + src40[478] + src40[479] + src40[480] + src40[481] + src40[482] + src40[483] + src40[484] + src40[485])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63] + src41[64] + src41[65] + src41[66] + src41[67] + src41[68] + src41[69] + src41[70] + src41[71] + src41[72] + src41[73] + src41[74] + src41[75] + src41[76] + src41[77] + src41[78] + src41[79] + src41[80] + src41[81] + src41[82] + src41[83] + src41[84] + src41[85] + src41[86] + src41[87] + src41[88] + src41[89] + src41[90] + src41[91] + src41[92] + src41[93] + src41[94] + src41[95] + src41[96] + src41[97] + src41[98] + src41[99] + src41[100] + src41[101] + src41[102] + src41[103] + src41[104] + src41[105] + src41[106] + src41[107] + src41[108] + src41[109] + src41[110] + src41[111] + src41[112] + src41[113] + src41[114] + src41[115] + src41[116] + src41[117] + src41[118] + src41[119] + src41[120] + src41[121] + src41[122] + src41[123] + src41[124] + src41[125] + src41[126] + src41[127] + src41[128] + src41[129] + src41[130] + src41[131] + src41[132] + src41[133] + src41[134] + src41[135] + src41[136] + src41[137] + src41[138] + src41[139] + src41[140] + src41[141] + src41[142] + src41[143] + src41[144] + src41[145] + src41[146] + src41[147] + src41[148] + src41[149] + src41[150] + src41[151] + src41[152] + src41[153] + src41[154] + src41[155] + src41[156] + src41[157] + src41[158] + src41[159] + src41[160] + src41[161] + src41[162] + src41[163] + src41[164] + src41[165] + src41[166] + src41[167] + src41[168] + src41[169] + src41[170] + src41[171] + src41[172] + src41[173] + src41[174] + src41[175] + src41[176] + src41[177] + src41[178] + src41[179] + src41[180] + src41[181] + src41[182] + src41[183] + src41[184] + src41[185] + src41[186] + src41[187] + src41[188] + src41[189] + src41[190] + src41[191] + src41[192] + src41[193] + src41[194] + src41[195] + src41[196] + src41[197] + src41[198] + src41[199] + src41[200] + src41[201] + src41[202] + src41[203] + src41[204] + src41[205] + src41[206] + src41[207] + src41[208] + src41[209] + src41[210] + src41[211] + src41[212] + src41[213] + src41[214] + src41[215] + src41[216] + src41[217] + src41[218] + src41[219] + src41[220] + src41[221] + src41[222] + src41[223] + src41[224] + src41[225] + src41[226] + src41[227] + src41[228] + src41[229] + src41[230] + src41[231] + src41[232] + src41[233] + src41[234] + src41[235] + src41[236] + src41[237] + src41[238] + src41[239] + src41[240] + src41[241] + src41[242] + src41[243] + src41[244] + src41[245] + src41[246] + src41[247] + src41[248] + src41[249] + src41[250] + src41[251] + src41[252] + src41[253] + src41[254] + src41[255] + src41[256] + src41[257] + src41[258] + src41[259] + src41[260] + src41[261] + src41[262] + src41[263] + src41[264] + src41[265] + src41[266] + src41[267] + src41[268] + src41[269] + src41[270] + src41[271] + src41[272] + src41[273] + src41[274] + src41[275] + src41[276] + src41[277] + src41[278] + src41[279] + src41[280] + src41[281] + src41[282] + src41[283] + src41[284] + src41[285] + src41[286] + src41[287] + src41[288] + src41[289] + src41[290] + src41[291] + src41[292] + src41[293] + src41[294] + src41[295] + src41[296] + src41[297] + src41[298] + src41[299] + src41[300] + src41[301] + src41[302] + src41[303] + src41[304] + src41[305] + src41[306] + src41[307] + src41[308] + src41[309] + src41[310] + src41[311] + src41[312] + src41[313] + src41[314] + src41[315] + src41[316] + src41[317] + src41[318] + src41[319] + src41[320] + src41[321] + src41[322] + src41[323] + src41[324] + src41[325] + src41[326] + src41[327] + src41[328] + src41[329] + src41[330] + src41[331] + src41[332] + src41[333] + src41[334] + src41[335] + src41[336] + src41[337] + src41[338] + src41[339] + src41[340] + src41[341] + src41[342] + src41[343] + src41[344] + src41[345] + src41[346] + src41[347] + src41[348] + src41[349] + src41[350] + src41[351] + src41[352] + src41[353] + src41[354] + src41[355] + src41[356] + src41[357] + src41[358] + src41[359] + src41[360] + src41[361] + src41[362] + src41[363] + src41[364] + src41[365] + src41[366] + src41[367] + src41[368] + src41[369] + src41[370] + src41[371] + src41[372] + src41[373] + src41[374] + src41[375] + src41[376] + src41[377] + src41[378] + src41[379] + src41[380] + src41[381] + src41[382] + src41[383] + src41[384] + src41[385] + src41[386] + src41[387] + src41[388] + src41[389] + src41[390] + src41[391] + src41[392] + src41[393] + src41[394] + src41[395] + src41[396] + src41[397] + src41[398] + src41[399] + src41[400] + src41[401] + src41[402] + src41[403] + src41[404] + src41[405] + src41[406] + src41[407] + src41[408] + src41[409] + src41[410] + src41[411] + src41[412] + src41[413] + src41[414] + src41[415] + src41[416] + src41[417] + src41[418] + src41[419] + src41[420] + src41[421] + src41[422] + src41[423] + src41[424] + src41[425] + src41[426] + src41[427] + src41[428] + src41[429] + src41[430] + src41[431] + src41[432] + src41[433] + src41[434] + src41[435] + src41[436] + src41[437] + src41[438] + src41[439] + src41[440] + src41[441] + src41[442] + src41[443] + src41[444] + src41[445] + src41[446] + src41[447] + src41[448] + src41[449] + src41[450] + src41[451] + src41[452] + src41[453] + src41[454] + src41[455] + src41[456] + src41[457] + src41[458] + src41[459] + src41[460] + src41[461] + src41[462] + src41[463] + src41[464] + src41[465] + src41[466] + src41[467] + src41[468] + src41[469] + src41[470] + src41[471] + src41[472] + src41[473] + src41[474] + src41[475] + src41[476] + src41[477] + src41[478] + src41[479] + src41[480] + src41[481] + src41[482] + src41[483] + src41[484] + src41[485])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63] + src42[64] + src42[65] + src42[66] + src42[67] + src42[68] + src42[69] + src42[70] + src42[71] + src42[72] + src42[73] + src42[74] + src42[75] + src42[76] + src42[77] + src42[78] + src42[79] + src42[80] + src42[81] + src42[82] + src42[83] + src42[84] + src42[85] + src42[86] + src42[87] + src42[88] + src42[89] + src42[90] + src42[91] + src42[92] + src42[93] + src42[94] + src42[95] + src42[96] + src42[97] + src42[98] + src42[99] + src42[100] + src42[101] + src42[102] + src42[103] + src42[104] + src42[105] + src42[106] + src42[107] + src42[108] + src42[109] + src42[110] + src42[111] + src42[112] + src42[113] + src42[114] + src42[115] + src42[116] + src42[117] + src42[118] + src42[119] + src42[120] + src42[121] + src42[122] + src42[123] + src42[124] + src42[125] + src42[126] + src42[127] + src42[128] + src42[129] + src42[130] + src42[131] + src42[132] + src42[133] + src42[134] + src42[135] + src42[136] + src42[137] + src42[138] + src42[139] + src42[140] + src42[141] + src42[142] + src42[143] + src42[144] + src42[145] + src42[146] + src42[147] + src42[148] + src42[149] + src42[150] + src42[151] + src42[152] + src42[153] + src42[154] + src42[155] + src42[156] + src42[157] + src42[158] + src42[159] + src42[160] + src42[161] + src42[162] + src42[163] + src42[164] + src42[165] + src42[166] + src42[167] + src42[168] + src42[169] + src42[170] + src42[171] + src42[172] + src42[173] + src42[174] + src42[175] + src42[176] + src42[177] + src42[178] + src42[179] + src42[180] + src42[181] + src42[182] + src42[183] + src42[184] + src42[185] + src42[186] + src42[187] + src42[188] + src42[189] + src42[190] + src42[191] + src42[192] + src42[193] + src42[194] + src42[195] + src42[196] + src42[197] + src42[198] + src42[199] + src42[200] + src42[201] + src42[202] + src42[203] + src42[204] + src42[205] + src42[206] + src42[207] + src42[208] + src42[209] + src42[210] + src42[211] + src42[212] + src42[213] + src42[214] + src42[215] + src42[216] + src42[217] + src42[218] + src42[219] + src42[220] + src42[221] + src42[222] + src42[223] + src42[224] + src42[225] + src42[226] + src42[227] + src42[228] + src42[229] + src42[230] + src42[231] + src42[232] + src42[233] + src42[234] + src42[235] + src42[236] + src42[237] + src42[238] + src42[239] + src42[240] + src42[241] + src42[242] + src42[243] + src42[244] + src42[245] + src42[246] + src42[247] + src42[248] + src42[249] + src42[250] + src42[251] + src42[252] + src42[253] + src42[254] + src42[255] + src42[256] + src42[257] + src42[258] + src42[259] + src42[260] + src42[261] + src42[262] + src42[263] + src42[264] + src42[265] + src42[266] + src42[267] + src42[268] + src42[269] + src42[270] + src42[271] + src42[272] + src42[273] + src42[274] + src42[275] + src42[276] + src42[277] + src42[278] + src42[279] + src42[280] + src42[281] + src42[282] + src42[283] + src42[284] + src42[285] + src42[286] + src42[287] + src42[288] + src42[289] + src42[290] + src42[291] + src42[292] + src42[293] + src42[294] + src42[295] + src42[296] + src42[297] + src42[298] + src42[299] + src42[300] + src42[301] + src42[302] + src42[303] + src42[304] + src42[305] + src42[306] + src42[307] + src42[308] + src42[309] + src42[310] + src42[311] + src42[312] + src42[313] + src42[314] + src42[315] + src42[316] + src42[317] + src42[318] + src42[319] + src42[320] + src42[321] + src42[322] + src42[323] + src42[324] + src42[325] + src42[326] + src42[327] + src42[328] + src42[329] + src42[330] + src42[331] + src42[332] + src42[333] + src42[334] + src42[335] + src42[336] + src42[337] + src42[338] + src42[339] + src42[340] + src42[341] + src42[342] + src42[343] + src42[344] + src42[345] + src42[346] + src42[347] + src42[348] + src42[349] + src42[350] + src42[351] + src42[352] + src42[353] + src42[354] + src42[355] + src42[356] + src42[357] + src42[358] + src42[359] + src42[360] + src42[361] + src42[362] + src42[363] + src42[364] + src42[365] + src42[366] + src42[367] + src42[368] + src42[369] + src42[370] + src42[371] + src42[372] + src42[373] + src42[374] + src42[375] + src42[376] + src42[377] + src42[378] + src42[379] + src42[380] + src42[381] + src42[382] + src42[383] + src42[384] + src42[385] + src42[386] + src42[387] + src42[388] + src42[389] + src42[390] + src42[391] + src42[392] + src42[393] + src42[394] + src42[395] + src42[396] + src42[397] + src42[398] + src42[399] + src42[400] + src42[401] + src42[402] + src42[403] + src42[404] + src42[405] + src42[406] + src42[407] + src42[408] + src42[409] + src42[410] + src42[411] + src42[412] + src42[413] + src42[414] + src42[415] + src42[416] + src42[417] + src42[418] + src42[419] + src42[420] + src42[421] + src42[422] + src42[423] + src42[424] + src42[425] + src42[426] + src42[427] + src42[428] + src42[429] + src42[430] + src42[431] + src42[432] + src42[433] + src42[434] + src42[435] + src42[436] + src42[437] + src42[438] + src42[439] + src42[440] + src42[441] + src42[442] + src42[443] + src42[444] + src42[445] + src42[446] + src42[447] + src42[448] + src42[449] + src42[450] + src42[451] + src42[452] + src42[453] + src42[454] + src42[455] + src42[456] + src42[457] + src42[458] + src42[459] + src42[460] + src42[461] + src42[462] + src42[463] + src42[464] + src42[465] + src42[466] + src42[467] + src42[468] + src42[469] + src42[470] + src42[471] + src42[472] + src42[473] + src42[474] + src42[475] + src42[476] + src42[477] + src42[478] + src42[479] + src42[480] + src42[481] + src42[482] + src42[483] + src42[484] + src42[485])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63] + src43[64] + src43[65] + src43[66] + src43[67] + src43[68] + src43[69] + src43[70] + src43[71] + src43[72] + src43[73] + src43[74] + src43[75] + src43[76] + src43[77] + src43[78] + src43[79] + src43[80] + src43[81] + src43[82] + src43[83] + src43[84] + src43[85] + src43[86] + src43[87] + src43[88] + src43[89] + src43[90] + src43[91] + src43[92] + src43[93] + src43[94] + src43[95] + src43[96] + src43[97] + src43[98] + src43[99] + src43[100] + src43[101] + src43[102] + src43[103] + src43[104] + src43[105] + src43[106] + src43[107] + src43[108] + src43[109] + src43[110] + src43[111] + src43[112] + src43[113] + src43[114] + src43[115] + src43[116] + src43[117] + src43[118] + src43[119] + src43[120] + src43[121] + src43[122] + src43[123] + src43[124] + src43[125] + src43[126] + src43[127] + src43[128] + src43[129] + src43[130] + src43[131] + src43[132] + src43[133] + src43[134] + src43[135] + src43[136] + src43[137] + src43[138] + src43[139] + src43[140] + src43[141] + src43[142] + src43[143] + src43[144] + src43[145] + src43[146] + src43[147] + src43[148] + src43[149] + src43[150] + src43[151] + src43[152] + src43[153] + src43[154] + src43[155] + src43[156] + src43[157] + src43[158] + src43[159] + src43[160] + src43[161] + src43[162] + src43[163] + src43[164] + src43[165] + src43[166] + src43[167] + src43[168] + src43[169] + src43[170] + src43[171] + src43[172] + src43[173] + src43[174] + src43[175] + src43[176] + src43[177] + src43[178] + src43[179] + src43[180] + src43[181] + src43[182] + src43[183] + src43[184] + src43[185] + src43[186] + src43[187] + src43[188] + src43[189] + src43[190] + src43[191] + src43[192] + src43[193] + src43[194] + src43[195] + src43[196] + src43[197] + src43[198] + src43[199] + src43[200] + src43[201] + src43[202] + src43[203] + src43[204] + src43[205] + src43[206] + src43[207] + src43[208] + src43[209] + src43[210] + src43[211] + src43[212] + src43[213] + src43[214] + src43[215] + src43[216] + src43[217] + src43[218] + src43[219] + src43[220] + src43[221] + src43[222] + src43[223] + src43[224] + src43[225] + src43[226] + src43[227] + src43[228] + src43[229] + src43[230] + src43[231] + src43[232] + src43[233] + src43[234] + src43[235] + src43[236] + src43[237] + src43[238] + src43[239] + src43[240] + src43[241] + src43[242] + src43[243] + src43[244] + src43[245] + src43[246] + src43[247] + src43[248] + src43[249] + src43[250] + src43[251] + src43[252] + src43[253] + src43[254] + src43[255] + src43[256] + src43[257] + src43[258] + src43[259] + src43[260] + src43[261] + src43[262] + src43[263] + src43[264] + src43[265] + src43[266] + src43[267] + src43[268] + src43[269] + src43[270] + src43[271] + src43[272] + src43[273] + src43[274] + src43[275] + src43[276] + src43[277] + src43[278] + src43[279] + src43[280] + src43[281] + src43[282] + src43[283] + src43[284] + src43[285] + src43[286] + src43[287] + src43[288] + src43[289] + src43[290] + src43[291] + src43[292] + src43[293] + src43[294] + src43[295] + src43[296] + src43[297] + src43[298] + src43[299] + src43[300] + src43[301] + src43[302] + src43[303] + src43[304] + src43[305] + src43[306] + src43[307] + src43[308] + src43[309] + src43[310] + src43[311] + src43[312] + src43[313] + src43[314] + src43[315] + src43[316] + src43[317] + src43[318] + src43[319] + src43[320] + src43[321] + src43[322] + src43[323] + src43[324] + src43[325] + src43[326] + src43[327] + src43[328] + src43[329] + src43[330] + src43[331] + src43[332] + src43[333] + src43[334] + src43[335] + src43[336] + src43[337] + src43[338] + src43[339] + src43[340] + src43[341] + src43[342] + src43[343] + src43[344] + src43[345] + src43[346] + src43[347] + src43[348] + src43[349] + src43[350] + src43[351] + src43[352] + src43[353] + src43[354] + src43[355] + src43[356] + src43[357] + src43[358] + src43[359] + src43[360] + src43[361] + src43[362] + src43[363] + src43[364] + src43[365] + src43[366] + src43[367] + src43[368] + src43[369] + src43[370] + src43[371] + src43[372] + src43[373] + src43[374] + src43[375] + src43[376] + src43[377] + src43[378] + src43[379] + src43[380] + src43[381] + src43[382] + src43[383] + src43[384] + src43[385] + src43[386] + src43[387] + src43[388] + src43[389] + src43[390] + src43[391] + src43[392] + src43[393] + src43[394] + src43[395] + src43[396] + src43[397] + src43[398] + src43[399] + src43[400] + src43[401] + src43[402] + src43[403] + src43[404] + src43[405] + src43[406] + src43[407] + src43[408] + src43[409] + src43[410] + src43[411] + src43[412] + src43[413] + src43[414] + src43[415] + src43[416] + src43[417] + src43[418] + src43[419] + src43[420] + src43[421] + src43[422] + src43[423] + src43[424] + src43[425] + src43[426] + src43[427] + src43[428] + src43[429] + src43[430] + src43[431] + src43[432] + src43[433] + src43[434] + src43[435] + src43[436] + src43[437] + src43[438] + src43[439] + src43[440] + src43[441] + src43[442] + src43[443] + src43[444] + src43[445] + src43[446] + src43[447] + src43[448] + src43[449] + src43[450] + src43[451] + src43[452] + src43[453] + src43[454] + src43[455] + src43[456] + src43[457] + src43[458] + src43[459] + src43[460] + src43[461] + src43[462] + src43[463] + src43[464] + src43[465] + src43[466] + src43[467] + src43[468] + src43[469] + src43[470] + src43[471] + src43[472] + src43[473] + src43[474] + src43[475] + src43[476] + src43[477] + src43[478] + src43[479] + src43[480] + src43[481] + src43[482] + src43[483] + src43[484] + src43[485])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63] + src44[64] + src44[65] + src44[66] + src44[67] + src44[68] + src44[69] + src44[70] + src44[71] + src44[72] + src44[73] + src44[74] + src44[75] + src44[76] + src44[77] + src44[78] + src44[79] + src44[80] + src44[81] + src44[82] + src44[83] + src44[84] + src44[85] + src44[86] + src44[87] + src44[88] + src44[89] + src44[90] + src44[91] + src44[92] + src44[93] + src44[94] + src44[95] + src44[96] + src44[97] + src44[98] + src44[99] + src44[100] + src44[101] + src44[102] + src44[103] + src44[104] + src44[105] + src44[106] + src44[107] + src44[108] + src44[109] + src44[110] + src44[111] + src44[112] + src44[113] + src44[114] + src44[115] + src44[116] + src44[117] + src44[118] + src44[119] + src44[120] + src44[121] + src44[122] + src44[123] + src44[124] + src44[125] + src44[126] + src44[127] + src44[128] + src44[129] + src44[130] + src44[131] + src44[132] + src44[133] + src44[134] + src44[135] + src44[136] + src44[137] + src44[138] + src44[139] + src44[140] + src44[141] + src44[142] + src44[143] + src44[144] + src44[145] + src44[146] + src44[147] + src44[148] + src44[149] + src44[150] + src44[151] + src44[152] + src44[153] + src44[154] + src44[155] + src44[156] + src44[157] + src44[158] + src44[159] + src44[160] + src44[161] + src44[162] + src44[163] + src44[164] + src44[165] + src44[166] + src44[167] + src44[168] + src44[169] + src44[170] + src44[171] + src44[172] + src44[173] + src44[174] + src44[175] + src44[176] + src44[177] + src44[178] + src44[179] + src44[180] + src44[181] + src44[182] + src44[183] + src44[184] + src44[185] + src44[186] + src44[187] + src44[188] + src44[189] + src44[190] + src44[191] + src44[192] + src44[193] + src44[194] + src44[195] + src44[196] + src44[197] + src44[198] + src44[199] + src44[200] + src44[201] + src44[202] + src44[203] + src44[204] + src44[205] + src44[206] + src44[207] + src44[208] + src44[209] + src44[210] + src44[211] + src44[212] + src44[213] + src44[214] + src44[215] + src44[216] + src44[217] + src44[218] + src44[219] + src44[220] + src44[221] + src44[222] + src44[223] + src44[224] + src44[225] + src44[226] + src44[227] + src44[228] + src44[229] + src44[230] + src44[231] + src44[232] + src44[233] + src44[234] + src44[235] + src44[236] + src44[237] + src44[238] + src44[239] + src44[240] + src44[241] + src44[242] + src44[243] + src44[244] + src44[245] + src44[246] + src44[247] + src44[248] + src44[249] + src44[250] + src44[251] + src44[252] + src44[253] + src44[254] + src44[255] + src44[256] + src44[257] + src44[258] + src44[259] + src44[260] + src44[261] + src44[262] + src44[263] + src44[264] + src44[265] + src44[266] + src44[267] + src44[268] + src44[269] + src44[270] + src44[271] + src44[272] + src44[273] + src44[274] + src44[275] + src44[276] + src44[277] + src44[278] + src44[279] + src44[280] + src44[281] + src44[282] + src44[283] + src44[284] + src44[285] + src44[286] + src44[287] + src44[288] + src44[289] + src44[290] + src44[291] + src44[292] + src44[293] + src44[294] + src44[295] + src44[296] + src44[297] + src44[298] + src44[299] + src44[300] + src44[301] + src44[302] + src44[303] + src44[304] + src44[305] + src44[306] + src44[307] + src44[308] + src44[309] + src44[310] + src44[311] + src44[312] + src44[313] + src44[314] + src44[315] + src44[316] + src44[317] + src44[318] + src44[319] + src44[320] + src44[321] + src44[322] + src44[323] + src44[324] + src44[325] + src44[326] + src44[327] + src44[328] + src44[329] + src44[330] + src44[331] + src44[332] + src44[333] + src44[334] + src44[335] + src44[336] + src44[337] + src44[338] + src44[339] + src44[340] + src44[341] + src44[342] + src44[343] + src44[344] + src44[345] + src44[346] + src44[347] + src44[348] + src44[349] + src44[350] + src44[351] + src44[352] + src44[353] + src44[354] + src44[355] + src44[356] + src44[357] + src44[358] + src44[359] + src44[360] + src44[361] + src44[362] + src44[363] + src44[364] + src44[365] + src44[366] + src44[367] + src44[368] + src44[369] + src44[370] + src44[371] + src44[372] + src44[373] + src44[374] + src44[375] + src44[376] + src44[377] + src44[378] + src44[379] + src44[380] + src44[381] + src44[382] + src44[383] + src44[384] + src44[385] + src44[386] + src44[387] + src44[388] + src44[389] + src44[390] + src44[391] + src44[392] + src44[393] + src44[394] + src44[395] + src44[396] + src44[397] + src44[398] + src44[399] + src44[400] + src44[401] + src44[402] + src44[403] + src44[404] + src44[405] + src44[406] + src44[407] + src44[408] + src44[409] + src44[410] + src44[411] + src44[412] + src44[413] + src44[414] + src44[415] + src44[416] + src44[417] + src44[418] + src44[419] + src44[420] + src44[421] + src44[422] + src44[423] + src44[424] + src44[425] + src44[426] + src44[427] + src44[428] + src44[429] + src44[430] + src44[431] + src44[432] + src44[433] + src44[434] + src44[435] + src44[436] + src44[437] + src44[438] + src44[439] + src44[440] + src44[441] + src44[442] + src44[443] + src44[444] + src44[445] + src44[446] + src44[447] + src44[448] + src44[449] + src44[450] + src44[451] + src44[452] + src44[453] + src44[454] + src44[455] + src44[456] + src44[457] + src44[458] + src44[459] + src44[460] + src44[461] + src44[462] + src44[463] + src44[464] + src44[465] + src44[466] + src44[467] + src44[468] + src44[469] + src44[470] + src44[471] + src44[472] + src44[473] + src44[474] + src44[475] + src44[476] + src44[477] + src44[478] + src44[479] + src44[480] + src44[481] + src44[482] + src44[483] + src44[484] + src44[485])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63] + src45[64] + src45[65] + src45[66] + src45[67] + src45[68] + src45[69] + src45[70] + src45[71] + src45[72] + src45[73] + src45[74] + src45[75] + src45[76] + src45[77] + src45[78] + src45[79] + src45[80] + src45[81] + src45[82] + src45[83] + src45[84] + src45[85] + src45[86] + src45[87] + src45[88] + src45[89] + src45[90] + src45[91] + src45[92] + src45[93] + src45[94] + src45[95] + src45[96] + src45[97] + src45[98] + src45[99] + src45[100] + src45[101] + src45[102] + src45[103] + src45[104] + src45[105] + src45[106] + src45[107] + src45[108] + src45[109] + src45[110] + src45[111] + src45[112] + src45[113] + src45[114] + src45[115] + src45[116] + src45[117] + src45[118] + src45[119] + src45[120] + src45[121] + src45[122] + src45[123] + src45[124] + src45[125] + src45[126] + src45[127] + src45[128] + src45[129] + src45[130] + src45[131] + src45[132] + src45[133] + src45[134] + src45[135] + src45[136] + src45[137] + src45[138] + src45[139] + src45[140] + src45[141] + src45[142] + src45[143] + src45[144] + src45[145] + src45[146] + src45[147] + src45[148] + src45[149] + src45[150] + src45[151] + src45[152] + src45[153] + src45[154] + src45[155] + src45[156] + src45[157] + src45[158] + src45[159] + src45[160] + src45[161] + src45[162] + src45[163] + src45[164] + src45[165] + src45[166] + src45[167] + src45[168] + src45[169] + src45[170] + src45[171] + src45[172] + src45[173] + src45[174] + src45[175] + src45[176] + src45[177] + src45[178] + src45[179] + src45[180] + src45[181] + src45[182] + src45[183] + src45[184] + src45[185] + src45[186] + src45[187] + src45[188] + src45[189] + src45[190] + src45[191] + src45[192] + src45[193] + src45[194] + src45[195] + src45[196] + src45[197] + src45[198] + src45[199] + src45[200] + src45[201] + src45[202] + src45[203] + src45[204] + src45[205] + src45[206] + src45[207] + src45[208] + src45[209] + src45[210] + src45[211] + src45[212] + src45[213] + src45[214] + src45[215] + src45[216] + src45[217] + src45[218] + src45[219] + src45[220] + src45[221] + src45[222] + src45[223] + src45[224] + src45[225] + src45[226] + src45[227] + src45[228] + src45[229] + src45[230] + src45[231] + src45[232] + src45[233] + src45[234] + src45[235] + src45[236] + src45[237] + src45[238] + src45[239] + src45[240] + src45[241] + src45[242] + src45[243] + src45[244] + src45[245] + src45[246] + src45[247] + src45[248] + src45[249] + src45[250] + src45[251] + src45[252] + src45[253] + src45[254] + src45[255] + src45[256] + src45[257] + src45[258] + src45[259] + src45[260] + src45[261] + src45[262] + src45[263] + src45[264] + src45[265] + src45[266] + src45[267] + src45[268] + src45[269] + src45[270] + src45[271] + src45[272] + src45[273] + src45[274] + src45[275] + src45[276] + src45[277] + src45[278] + src45[279] + src45[280] + src45[281] + src45[282] + src45[283] + src45[284] + src45[285] + src45[286] + src45[287] + src45[288] + src45[289] + src45[290] + src45[291] + src45[292] + src45[293] + src45[294] + src45[295] + src45[296] + src45[297] + src45[298] + src45[299] + src45[300] + src45[301] + src45[302] + src45[303] + src45[304] + src45[305] + src45[306] + src45[307] + src45[308] + src45[309] + src45[310] + src45[311] + src45[312] + src45[313] + src45[314] + src45[315] + src45[316] + src45[317] + src45[318] + src45[319] + src45[320] + src45[321] + src45[322] + src45[323] + src45[324] + src45[325] + src45[326] + src45[327] + src45[328] + src45[329] + src45[330] + src45[331] + src45[332] + src45[333] + src45[334] + src45[335] + src45[336] + src45[337] + src45[338] + src45[339] + src45[340] + src45[341] + src45[342] + src45[343] + src45[344] + src45[345] + src45[346] + src45[347] + src45[348] + src45[349] + src45[350] + src45[351] + src45[352] + src45[353] + src45[354] + src45[355] + src45[356] + src45[357] + src45[358] + src45[359] + src45[360] + src45[361] + src45[362] + src45[363] + src45[364] + src45[365] + src45[366] + src45[367] + src45[368] + src45[369] + src45[370] + src45[371] + src45[372] + src45[373] + src45[374] + src45[375] + src45[376] + src45[377] + src45[378] + src45[379] + src45[380] + src45[381] + src45[382] + src45[383] + src45[384] + src45[385] + src45[386] + src45[387] + src45[388] + src45[389] + src45[390] + src45[391] + src45[392] + src45[393] + src45[394] + src45[395] + src45[396] + src45[397] + src45[398] + src45[399] + src45[400] + src45[401] + src45[402] + src45[403] + src45[404] + src45[405] + src45[406] + src45[407] + src45[408] + src45[409] + src45[410] + src45[411] + src45[412] + src45[413] + src45[414] + src45[415] + src45[416] + src45[417] + src45[418] + src45[419] + src45[420] + src45[421] + src45[422] + src45[423] + src45[424] + src45[425] + src45[426] + src45[427] + src45[428] + src45[429] + src45[430] + src45[431] + src45[432] + src45[433] + src45[434] + src45[435] + src45[436] + src45[437] + src45[438] + src45[439] + src45[440] + src45[441] + src45[442] + src45[443] + src45[444] + src45[445] + src45[446] + src45[447] + src45[448] + src45[449] + src45[450] + src45[451] + src45[452] + src45[453] + src45[454] + src45[455] + src45[456] + src45[457] + src45[458] + src45[459] + src45[460] + src45[461] + src45[462] + src45[463] + src45[464] + src45[465] + src45[466] + src45[467] + src45[468] + src45[469] + src45[470] + src45[471] + src45[472] + src45[473] + src45[474] + src45[475] + src45[476] + src45[477] + src45[478] + src45[479] + src45[480] + src45[481] + src45[482] + src45[483] + src45[484] + src45[485])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63] + src46[64] + src46[65] + src46[66] + src46[67] + src46[68] + src46[69] + src46[70] + src46[71] + src46[72] + src46[73] + src46[74] + src46[75] + src46[76] + src46[77] + src46[78] + src46[79] + src46[80] + src46[81] + src46[82] + src46[83] + src46[84] + src46[85] + src46[86] + src46[87] + src46[88] + src46[89] + src46[90] + src46[91] + src46[92] + src46[93] + src46[94] + src46[95] + src46[96] + src46[97] + src46[98] + src46[99] + src46[100] + src46[101] + src46[102] + src46[103] + src46[104] + src46[105] + src46[106] + src46[107] + src46[108] + src46[109] + src46[110] + src46[111] + src46[112] + src46[113] + src46[114] + src46[115] + src46[116] + src46[117] + src46[118] + src46[119] + src46[120] + src46[121] + src46[122] + src46[123] + src46[124] + src46[125] + src46[126] + src46[127] + src46[128] + src46[129] + src46[130] + src46[131] + src46[132] + src46[133] + src46[134] + src46[135] + src46[136] + src46[137] + src46[138] + src46[139] + src46[140] + src46[141] + src46[142] + src46[143] + src46[144] + src46[145] + src46[146] + src46[147] + src46[148] + src46[149] + src46[150] + src46[151] + src46[152] + src46[153] + src46[154] + src46[155] + src46[156] + src46[157] + src46[158] + src46[159] + src46[160] + src46[161] + src46[162] + src46[163] + src46[164] + src46[165] + src46[166] + src46[167] + src46[168] + src46[169] + src46[170] + src46[171] + src46[172] + src46[173] + src46[174] + src46[175] + src46[176] + src46[177] + src46[178] + src46[179] + src46[180] + src46[181] + src46[182] + src46[183] + src46[184] + src46[185] + src46[186] + src46[187] + src46[188] + src46[189] + src46[190] + src46[191] + src46[192] + src46[193] + src46[194] + src46[195] + src46[196] + src46[197] + src46[198] + src46[199] + src46[200] + src46[201] + src46[202] + src46[203] + src46[204] + src46[205] + src46[206] + src46[207] + src46[208] + src46[209] + src46[210] + src46[211] + src46[212] + src46[213] + src46[214] + src46[215] + src46[216] + src46[217] + src46[218] + src46[219] + src46[220] + src46[221] + src46[222] + src46[223] + src46[224] + src46[225] + src46[226] + src46[227] + src46[228] + src46[229] + src46[230] + src46[231] + src46[232] + src46[233] + src46[234] + src46[235] + src46[236] + src46[237] + src46[238] + src46[239] + src46[240] + src46[241] + src46[242] + src46[243] + src46[244] + src46[245] + src46[246] + src46[247] + src46[248] + src46[249] + src46[250] + src46[251] + src46[252] + src46[253] + src46[254] + src46[255] + src46[256] + src46[257] + src46[258] + src46[259] + src46[260] + src46[261] + src46[262] + src46[263] + src46[264] + src46[265] + src46[266] + src46[267] + src46[268] + src46[269] + src46[270] + src46[271] + src46[272] + src46[273] + src46[274] + src46[275] + src46[276] + src46[277] + src46[278] + src46[279] + src46[280] + src46[281] + src46[282] + src46[283] + src46[284] + src46[285] + src46[286] + src46[287] + src46[288] + src46[289] + src46[290] + src46[291] + src46[292] + src46[293] + src46[294] + src46[295] + src46[296] + src46[297] + src46[298] + src46[299] + src46[300] + src46[301] + src46[302] + src46[303] + src46[304] + src46[305] + src46[306] + src46[307] + src46[308] + src46[309] + src46[310] + src46[311] + src46[312] + src46[313] + src46[314] + src46[315] + src46[316] + src46[317] + src46[318] + src46[319] + src46[320] + src46[321] + src46[322] + src46[323] + src46[324] + src46[325] + src46[326] + src46[327] + src46[328] + src46[329] + src46[330] + src46[331] + src46[332] + src46[333] + src46[334] + src46[335] + src46[336] + src46[337] + src46[338] + src46[339] + src46[340] + src46[341] + src46[342] + src46[343] + src46[344] + src46[345] + src46[346] + src46[347] + src46[348] + src46[349] + src46[350] + src46[351] + src46[352] + src46[353] + src46[354] + src46[355] + src46[356] + src46[357] + src46[358] + src46[359] + src46[360] + src46[361] + src46[362] + src46[363] + src46[364] + src46[365] + src46[366] + src46[367] + src46[368] + src46[369] + src46[370] + src46[371] + src46[372] + src46[373] + src46[374] + src46[375] + src46[376] + src46[377] + src46[378] + src46[379] + src46[380] + src46[381] + src46[382] + src46[383] + src46[384] + src46[385] + src46[386] + src46[387] + src46[388] + src46[389] + src46[390] + src46[391] + src46[392] + src46[393] + src46[394] + src46[395] + src46[396] + src46[397] + src46[398] + src46[399] + src46[400] + src46[401] + src46[402] + src46[403] + src46[404] + src46[405] + src46[406] + src46[407] + src46[408] + src46[409] + src46[410] + src46[411] + src46[412] + src46[413] + src46[414] + src46[415] + src46[416] + src46[417] + src46[418] + src46[419] + src46[420] + src46[421] + src46[422] + src46[423] + src46[424] + src46[425] + src46[426] + src46[427] + src46[428] + src46[429] + src46[430] + src46[431] + src46[432] + src46[433] + src46[434] + src46[435] + src46[436] + src46[437] + src46[438] + src46[439] + src46[440] + src46[441] + src46[442] + src46[443] + src46[444] + src46[445] + src46[446] + src46[447] + src46[448] + src46[449] + src46[450] + src46[451] + src46[452] + src46[453] + src46[454] + src46[455] + src46[456] + src46[457] + src46[458] + src46[459] + src46[460] + src46[461] + src46[462] + src46[463] + src46[464] + src46[465] + src46[466] + src46[467] + src46[468] + src46[469] + src46[470] + src46[471] + src46[472] + src46[473] + src46[474] + src46[475] + src46[476] + src46[477] + src46[478] + src46[479] + src46[480] + src46[481] + src46[482] + src46[483] + src46[484] + src46[485])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63] + src47[64] + src47[65] + src47[66] + src47[67] + src47[68] + src47[69] + src47[70] + src47[71] + src47[72] + src47[73] + src47[74] + src47[75] + src47[76] + src47[77] + src47[78] + src47[79] + src47[80] + src47[81] + src47[82] + src47[83] + src47[84] + src47[85] + src47[86] + src47[87] + src47[88] + src47[89] + src47[90] + src47[91] + src47[92] + src47[93] + src47[94] + src47[95] + src47[96] + src47[97] + src47[98] + src47[99] + src47[100] + src47[101] + src47[102] + src47[103] + src47[104] + src47[105] + src47[106] + src47[107] + src47[108] + src47[109] + src47[110] + src47[111] + src47[112] + src47[113] + src47[114] + src47[115] + src47[116] + src47[117] + src47[118] + src47[119] + src47[120] + src47[121] + src47[122] + src47[123] + src47[124] + src47[125] + src47[126] + src47[127] + src47[128] + src47[129] + src47[130] + src47[131] + src47[132] + src47[133] + src47[134] + src47[135] + src47[136] + src47[137] + src47[138] + src47[139] + src47[140] + src47[141] + src47[142] + src47[143] + src47[144] + src47[145] + src47[146] + src47[147] + src47[148] + src47[149] + src47[150] + src47[151] + src47[152] + src47[153] + src47[154] + src47[155] + src47[156] + src47[157] + src47[158] + src47[159] + src47[160] + src47[161] + src47[162] + src47[163] + src47[164] + src47[165] + src47[166] + src47[167] + src47[168] + src47[169] + src47[170] + src47[171] + src47[172] + src47[173] + src47[174] + src47[175] + src47[176] + src47[177] + src47[178] + src47[179] + src47[180] + src47[181] + src47[182] + src47[183] + src47[184] + src47[185] + src47[186] + src47[187] + src47[188] + src47[189] + src47[190] + src47[191] + src47[192] + src47[193] + src47[194] + src47[195] + src47[196] + src47[197] + src47[198] + src47[199] + src47[200] + src47[201] + src47[202] + src47[203] + src47[204] + src47[205] + src47[206] + src47[207] + src47[208] + src47[209] + src47[210] + src47[211] + src47[212] + src47[213] + src47[214] + src47[215] + src47[216] + src47[217] + src47[218] + src47[219] + src47[220] + src47[221] + src47[222] + src47[223] + src47[224] + src47[225] + src47[226] + src47[227] + src47[228] + src47[229] + src47[230] + src47[231] + src47[232] + src47[233] + src47[234] + src47[235] + src47[236] + src47[237] + src47[238] + src47[239] + src47[240] + src47[241] + src47[242] + src47[243] + src47[244] + src47[245] + src47[246] + src47[247] + src47[248] + src47[249] + src47[250] + src47[251] + src47[252] + src47[253] + src47[254] + src47[255] + src47[256] + src47[257] + src47[258] + src47[259] + src47[260] + src47[261] + src47[262] + src47[263] + src47[264] + src47[265] + src47[266] + src47[267] + src47[268] + src47[269] + src47[270] + src47[271] + src47[272] + src47[273] + src47[274] + src47[275] + src47[276] + src47[277] + src47[278] + src47[279] + src47[280] + src47[281] + src47[282] + src47[283] + src47[284] + src47[285] + src47[286] + src47[287] + src47[288] + src47[289] + src47[290] + src47[291] + src47[292] + src47[293] + src47[294] + src47[295] + src47[296] + src47[297] + src47[298] + src47[299] + src47[300] + src47[301] + src47[302] + src47[303] + src47[304] + src47[305] + src47[306] + src47[307] + src47[308] + src47[309] + src47[310] + src47[311] + src47[312] + src47[313] + src47[314] + src47[315] + src47[316] + src47[317] + src47[318] + src47[319] + src47[320] + src47[321] + src47[322] + src47[323] + src47[324] + src47[325] + src47[326] + src47[327] + src47[328] + src47[329] + src47[330] + src47[331] + src47[332] + src47[333] + src47[334] + src47[335] + src47[336] + src47[337] + src47[338] + src47[339] + src47[340] + src47[341] + src47[342] + src47[343] + src47[344] + src47[345] + src47[346] + src47[347] + src47[348] + src47[349] + src47[350] + src47[351] + src47[352] + src47[353] + src47[354] + src47[355] + src47[356] + src47[357] + src47[358] + src47[359] + src47[360] + src47[361] + src47[362] + src47[363] + src47[364] + src47[365] + src47[366] + src47[367] + src47[368] + src47[369] + src47[370] + src47[371] + src47[372] + src47[373] + src47[374] + src47[375] + src47[376] + src47[377] + src47[378] + src47[379] + src47[380] + src47[381] + src47[382] + src47[383] + src47[384] + src47[385] + src47[386] + src47[387] + src47[388] + src47[389] + src47[390] + src47[391] + src47[392] + src47[393] + src47[394] + src47[395] + src47[396] + src47[397] + src47[398] + src47[399] + src47[400] + src47[401] + src47[402] + src47[403] + src47[404] + src47[405] + src47[406] + src47[407] + src47[408] + src47[409] + src47[410] + src47[411] + src47[412] + src47[413] + src47[414] + src47[415] + src47[416] + src47[417] + src47[418] + src47[419] + src47[420] + src47[421] + src47[422] + src47[423] + src47[424] + src47[425] + src47[426] + src47[427] + src47[428] + src47[429] + src47[430] + src47[431] + src47[432] + src47[433] + src47[434] + src47[435] + src47[436] + src47[437] + src47[438] + src47[439] + src47[440] + src47[441] + src47[442] + src47[443] + src47[444] + src47[445] + src47[446] + src47[447] + src47[448] + src47[449] + src47[450] + src47[451] + src47[452] + src47[453] + src47[454] + src47[455] + src47[456] + src47[457] + src47[458] + src47[459] + src47[460] + src47[461] + src47[462] + src47[463] + src47[464] + src47[465] + src47[466] + src47[467] + src47[468] + src47[469] + src47[470] + src47[471] + src47[472] + src47[473] + src47[474] + src47[475] + src47[476] + src47[477] + src47[478] + src47[479] + src47[480] + src47[481] + src47[482] + src47[483] + src47[484] + src47[485])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63] + src48[64] + src48[65] + src48[66] + src48[67] + src48[68] + src48[69] + src48[70] + src48[71] + src48[72] + src48[73] + src48[74] + src48[75] + src48[76] + src48[77] + src48[78] + src48[79] + src48[80] + src48[81] + src48[82] + src48[83] + src48[84] + src48[85] + src48[86] + src48[87] + src48[88] + src48[89] + src48[90] + src48[91] + src48[92] + src48[93] + src48[94] + src48[95] + src48[96] + src48[97] + src48[98] + src48[99] + src48[100] + src48[101] + src48[102] + src48[103] + src48[104] + src48[105] + src48[106] + src48[107] + src48[108] + src48[109] + src48[110] + src48[111] + src48[112] + src48[113] + src48[114] + src48[115] + src48[116] + src48[117] + src48[118] + src48[119] + src48[120] + src48[121] + src48[122] + src48[123] + src48[124] + src48[125] + src48[126] + src48[127] + src48[128] + src48[129] + src48[130] + src48[131] + src48[132] + src48[133] + src48[134] + src48[135] + src48[136] + src48[137] + src48[138] + src48[139] + src48[140] + src48[141] + src48[142] + src48[143] + src48[144] + src48[145] + src48[146] + src48[147] + src48[148] + src48[149] + src48[150] + src48[151] + src48[152] + src48[153] + src48[154] + src48[155] + src48[156] + src48[157] + src48[158] + src48[159] + src48[160] + src48[161] + src48[162] + src48[163] + src48[164] + src48[165] + src48[166] + src48[167] + src48[168] + src48[169] + src48[170] + src48[171] + src48[172] + src48[173] + src48[174] + src48[175] + src48[176] + src48[177] + src48[178] + src48[179] + src48[180] + src48[181] + src48[182] + src48[183] + src48[184] + src48[185] + src48[186] + src48[187] + src48[188] + src48[189] + src48[190] + src48[191] + src48[192] + src48[193] + src48[194] + src48[195] + src48[196] + src48[197] + src48[198] + src48[199] + src48[200] + src48[201] + src48[202] + src48[203] + src48[204] + src48[205] + src48[206] + src48[207] + src48[208] + src48[209] + src48[210] + src48[211] + src48[212] + src48[213] + src48[214] + src48[215] + src48[216] + src48[217] + src48[218] + src48[219] + src48[220] + src48[221] + src48[222] + src48[223] + src48[224] + src48[225] + src48[226] + src48[227] + src48[228] + src48[229] + src48[230] + src48[231] + src48[232] + src48[233] + src48[234] + src48[235] + src48[236] + src48[237] + src48[238] + src48[239] + src48[240] + src48[241] + src48[242] + src48[243] + src48[244] + src48[245] + src48[246] + src48[247] + src48[248] + src48[249] + src48[250] + src48[251] + src48[252] + src48[253] + src48[254] + src48[255] + src48[256] + src48[257] + src48[258] + src48[259] + src48[260] + src48[261] + src48[262] + src48[263] + src48[264] + src48[265] + src48[266] + src48[267] + src48[268] + src48[269] + src48[270] + src48[271] + src48[272] + src48[273] + src48[274] + src48[275] + src48[276] + src48[277] + src48[278] + src48[279] + src48[280] + src48[281] + src48[282] + src48[283] + src48[284] + src48[285] + src48[286] + src48[287] + src48[288] + src48[289] + src48[290] + src48[291] + src48[292] + src48[293] + src48[294] + src48[295] + src48[296] + src48[297] + src48[298] + src48[299] + src48[300] + src48[301] + src48[302] + src48[303] + src48[304] + src48[305] + src48[306] + src48[307] + src48[308] + src48[309] + src48[310] + src48[311] + src48[312] + src48[313] + src48[314] + src48[315] + src48[316] + src48[317] + src48[318] + src48[319] + src48[320] + src48[321] + src48[322] + src48[323] + src48[324] + src48[325] + src48[326] + src48[327] + src48[328] + src48[329] + src48[330] + src48[331] + src48[332] + src48[333] + src48[334] + src48[335] + src48[336] + src48[337] + src48[338] + src48[339] + src48[340] + src48[341] + src48[342] + src48[343] + src48[344] + src48[345] + src48[346] + src48[347] + src48[348] + src48[349] + src48[350] + src48[351] + src48[352] + src48[353] + src48[354] + src48[355] + src48[356] + src48[357] + src48[358] + src48[359] + src48[360] + src48[361] + src48[362] + src48[363] + src48[364] + src48[365] + src48[366] + src48[367] + src48[368] + src48[369] + src48[370] + src48[371] + src48[372] + src48[373] + src48[374] + src48[375] + src48[376] + src48[377] + src48[378] + src48[379] + src48[380] + src48[381] + src48[382] + src48[383] + src48[384] + src48[385] + src48[386] + src48[387] + src48[388] + src48[389] + src48[390] + src48[391] + src48[392] + src48[393] + src48[394] + src48[395] + src48[396] + src48[397] + src48[398] + src48[399] + src48[400] + src48[401] + src48[402] + src48[403] + src48[404] + src48[405] + src48[406] + src48[407] + src48[408] + src48[409] + src48[410] + src48[411] + src48[412] + src48[413] + src48[414] + src48[415] + src48[416] + src48[417] + src48[418] + src48[419] + src48[420] + src48[421] + src48[422] + src48[423] + src48[424] + src48[425] + src48[426] + src48[427] + src48[428] + src48[429] + src48[430] + src48[431] + src48[432] + src48[433] + src48[434] + src48[435] + src48[436] + src48[437] + src48[438] + src48[439] + src48[440] + src48[441] + src48[442] + src48[443] + src48[444] + src48[445] + src48[446] + src48[447] + src48[448] + src48[449] + src48[450] + src48[451] + src48[452] + src48[453] + src48[454] + src48[455] + src48[456] + src48[457] + src48[458] + src48[459] + src48[460] + src48[461] + src48[462] + src48[463] + src48[464] + src48[465] + src48[466] + src48[467] + src48[468] + src48[469] + src48[470] + src48[471] + src48[472] + src48[473] + src48[474] + src48[475] + src48[476] + src48[477] + src48[478] + src48[479] + src48[480] + src48[481] + src48[482] + src48[483] + src48[484] + src48[485])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63] + src49[64] + src49[65] + src49[66] + src49[67] + src49[68] + src49[69] + src49[70] + src49[71] + src49[72] + src49[73] + src49[74] + src49[75] + src49[76] + src49[77] + src49[78] + src49[79] + src49[80] + src49[81] + src49[82] + src49[83] + src49[84] + src49[85] + src49[86] + src49[87] + src49[88] + src49[89] + src49[90] + src49[91] + src49[92] + src49[93] + src49[94] + src49[95] + src49[96] + src49[97] + src49[98] + src49[99] + src49[100] + src49[101] + src49[102] + src49[103] + src49[104] + src49[105] + src49[106] + src49[107] + src49[108] + src49[109] + src49[110] + src49[111] + src49[112] + src49[113] + src49[114] + src49[115] + src49[116] + src49[117] + src49[118] + src49[119] + src49[120] + src49[121] + src49[122] + src49[123] + src49[124] + src49[125] + src49[126] + src49[127] + src49[128] + src49[129] + src49[130] + src49[131] + src49[132] + src49[133] + src49[134] + src49[135] + src49[136] + src49[137] + src49[138] + src49[139] + src49[140] + src49[141] + src49[142] + src49[143] + src49[144] + src49[145] + src49[146] + src49[147] + src49[148] + src49[149] + src49[150] + src49[151] + src49[152] + src49[153] + src49[154] + src49[155] + src49[156] + src49[157] + src49[158] + src49[159] + src49[160] + src49[161] + src49[162] + src49[163] + src49[164] + src49[165] + src49[166] + src49[167] + src49[168] + src49[169] + src49[170] + src49[171] + src49[172] + src49[173] + src49[174] + src49[175] + src49[176] + src49[177] + src49[178] + src49[179] + src49[180] + src49[181] + src49[182] + src49[183] + src49[184] + src49[185] + src49[186] + src49[187] + src49[188] + src49[189] + src49[190] + src49[191] + src49[192] + src49[193] + src49[194] + src49[195] + src49[196] + src49[197] + src49[198] + src49[199] + src49[200] + src49[201] + src49[202] + src49[203] + src49[204] + src49[205] + src49[206] + src49[207] + src49[208] + src49[209] + src49[210] + src49[211] + src49[212] + src49[213] + src49[214] + src49[215] + src49[216] + src49[217] + src49[218] + src49[219] + src49[220] + src49[221] + src49[222] + src49[223] + src49[224] + src49[225] + src49[226] + src49[227] + src49[228] + src49[229] + src49[230] + src49[231] + src49[232] + src49[233] + src49[234] + src49[235] + src49[236] + src49[237] + src49[238] + src49[239] + src49[240] + src49[241] + src49[242] + src49[243] + src49[244] + src49[245] + src49[246] + src49[247] + src49[248] + src49[249] + src49[250] + src49[251] + src49[252] + src49[253] + src49[254] + src49[255] + src49[256] + src49[257] + src49[258] + src49[259] + src49[260] + src49[261] + src49[262] + src49[263] + src49[264] + src49[265] + src49[266] + src49[267] + src49[268] + src49[269] + src49[270] + src49[271] + src49[272] + src49[273] + src49[274] + src49[275] + src49[276] + src49[277] + src49[278] + src49[279] + src49[280] + src49[281] + src49[282] + src49[283] + src49[284] + src49[285] + src49[286] + src49[287] + src49[288] + src49[289] + src49[290] + src49[291] + src49[292] + src49[293] + src49[294] + src49[295] + src49[296] + src49[297] + src49[298] + src49[299] + src49[300] + src49[301] + src49[302] + src49[303] + src49[304] + src49[305] + src49[306] + src49[307] + src49[308] + src49[309] + src49[310] + src49[311] + src49[312] + src49[313] + src49[314] + src49[315] + src49[316] + src49[317] + src49[318] + src49[319] + src49[320] + src49[321] + src49[322] + src49[323] + src49[324] + src49[325] + src49[326] + src49[327] + src49[328] + src49[329] + src49[330] + src49[331] + src49[332] + src49[333] + src49[334] + src49[335] + src49[336] + src49[337] + src49[338] + src49[339] + src49[340] + src49[341] + src49[342] + src49[343] + src49[344] + src49[345] + src49[346] + src49[347] + src49[348] + src49[349] + src49[350] + src49[351] + src49[352] + src49[353] + src49[354] + src49[355] + src49[356] + src49[357] + src49[358] + src49[359] + src49[360] + src49[361] + src49[362] + src49[363] + src49[364] + src49[365] + src49[366] + src49[367] + src49[368] + src49[369] + src49[370] + src49[371] + src49[372] + src49[373] + src49[374] + src49[375] + src49[376] + src49[377] + src49[378] + src49[379] + src49[380] + src49[381] + src49[382] + src49[383] + src49[384] + src49[385] + src49[386] + src49[387] + src49[388] + src49[389] + src49[390] + src49[391] + src49[392] + src49[393] + src49[394] + src49[395] + src49[396] + src49[397] + src49[398] + src49[399] + src49[400] + src49[401] + src49[402] + src49[403] + src49[404] + src49[405] + src49[406] + src49[407] + src49[408] + src49[409] + src49[410] + src49[411] + src49[412] + src49[413] + src49[414] + src49[415] + src49[416] + src49[417] + src49[418] + src49[419] + src49[420] + src49[421] + src49[422] + src49[423] + src49[424] + src49[425] + src49[426] + src49[427] + src49[428] + src49[429] + src49[430] + src49[431] + src49[432] + src49[433] + src49[434] + src49[435] + src49[436] + src49[437] + src49[438] + src49[439] + src49[440] + src49[441] + src49[442] + src49[443] + src49[444] + src49[445] + src49[446] + src49[447] + src49[448] + src49[449] + src49[450] + src49[451] + src49[452] + src49[453] + src49[454] + src49[455] + src49[456] + src49[457] + src49[458] + src49[459] + src49[460] + src49[461] + src49[462] + src49[463] + src49[464] + src49[465] + src49[466] + src49[467] + src49[468] + src49[469] + src49[470] + src49[471] + src49[472] + src49[473] + src49[474] + src49[475] + src49[476] + src49[477] + src49[478] + src49[479] + src49[480] + src49[481] + src49[482] + src49[483] + src49[484] + src49[485])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63] + src50[64] + src50[65] + src50[66] + src50[67] + src50[68] + src50[69] + src50[70] + src50[71] + src50[72] + src50[73] + src50[74] + src50[75] + src50[76] + src50[77] + src50[78] + src50[79] + src50[80] + src50[81] + src50[82] + src50[83] + src50[84] + src50[85] + src50[86] + src50[87] + src50[88] + src50[89] + src50[90] + src50[91] + src50[92] + src50[93] + src50[94] + src50[95] + src50[96] + src50[97] + src50[98] + src50[99] + src50[100] + src50[101] + src50[102] + src50[103] + src50[104] + src50[105] + src50[106] + src50[107] + src50[108] + src50[109] + src50[110] + src50[111] + src50[112] + src50[113] + src50[114] + src50[115] + src50[116] + src50[117] + src50[118] + src50[119] + src50[120] + src50[121] + src50[122] + src50[123] + src50[124] + src50[125] + src50[126] + src50[127] + src50[128] + src50[129] + src50[130] + src50[131] + src50[132] + src50[133] + src50[134] + src50[135] + src50[136] + src50[137] + src50[138] + src50[139] + src50[140] + src50[141] + src50[142] + src50[143] + src50[144] + src50[145] + src50[146] + src50[147] + src50[148] + src50[149] + src50[150] + src50[151] + src50[152] + src50[153] + src50[154] + src50[155] + src50[156] + src50[157] + src50[158] + src50[159] + src50[160] + src50[161] + src50[162] + src50[163] + src50[164] + src50[165] + src50[166] + src50[167] + src50[168] + src50[169] + src50[170] + src50[171] + src50[172] + src50[173] + src50[174] + src50[175] + src50[176] + src50[177] + src50[178] + src50[179] + src50[180] + src50[181] + src50[182] + src50[183] + src50[184] + src50[185] + src50[186] + src50[187] + src50[188] + src50[189] + src50[190] + src50[191] + src50[192] + src50[193] + src50[194] + src50[195] + src50[196] + src50[197] + src50[198] + src50[199] + src50[200] + src50[201] + src50[202] + src50[203] + src50[204] + src50[205] + src50[206] + src50[207] + src50[208] + src50[209] + src50[210] + src50[211] + src50[212] + src50[213] + src50[214] + src50[215] + src50[216] + src50[217] + src50[218] + src50[219] + src50[220] + src50[221] + src50[222] + src50[223] + src50[224] + src50[225] + src50[226] + src50[227] + src50[228] + src50[229] + src50[230] + src50[231] + src50[232] + src50[233] + src50[234] + src50[235] + src50[236] + src50[237] + src50[238] + src50[239] + src50[240] + src50[241] + src50[242] + src50[243] + src50[244] + src50[245] + src50[246] + src50[247] + src50[248] + src50[249] + src50[250] + src50[251] + src50[252] + src50[253] + src50[254] + src50[255] + src50[256] + src50[257] + src50[258] + src50[259] + src50[260] + src50[261] + src50[262] + src50[263] + src50[264] + src50[265] + src50[266] + src50[267] + src50[268] + src50[269] + src50[270] + src50[271] + src50[272] + src50[273] + src50[274] + src50[275] + src50[276] + src50[277] + src50[278] + src50[279] + src50[280] + src50[281] + src50[282] + src50[283] + src50[284] + src50[285] + src50[286] + src50[287] + src50[288] + src50[289] + src50[290] + src50[291] + src50[292] + src50[293] + src50[294] + src50[295] + src50[296] + src50[297] + src50[298] + src50[299] + src50[300] + src50[301] + src50[302] + src50[303] + src50[304] + src50[305] + src50[306] + src50[307] + src50[308] + src50[309] + src50[310] + src50[311] + src50[312] + src50[313] + src50[314] + src50[315] + src50[316] + src50[317] + src50[318] + src50[319] + src50[320] + src50[321] + src50[322] + src50[323] + src50[324] + src50[325] + src50[326] + src50[327] + src50[328] + src50[329] + src50[330] + src50[331] + src50[332] + src50[333] + src50[334] + src50[335] + src50[336] + src50[337] + src50[338] + src50[339] + src50[340] + src50[341] + src50[342] + src50[343] + src50[344] + src50[345] + src50[346] + src50[347] + src50[348] + src50[349] + src50[350] + src50[351] + src50[352] + src50[353] + src50[354] + src50[355] + src50[356] + src50[357] + src50[358] + src50[359] + src50[360] + src50[361] + src50[362] + src50[363] + src50[364] + src50[365] + src50[366] + src50[367] + src50[368] + src50[369] + src50[370] + src50[371] + src50[372] + src50[373] + src50[374] + src50[375] + src50[376] + src50[377] + src50[378] + src50[379] + src50[380] + src50[381] + src50[382] + src50[383] + src50[384] + src50[385] + src50[386] + src50[387] + src50[388] + src50[389] + src50[390] + src50[391] + src50[392] + src50[393] + src50[394] + src50[395] + src50[396] + src50[397] + src50[398] + src50[399] + src50[400] + src50[401] + src50[402] + src50[403] + src50[404] + src50[405] + src50[406] + src50[407] + src50[408] + src50[409] + src50[410] + src50[411] + src50[412] + src50[413] + src50[414] + src50[415] + src50[416] + src50[417] + src50[418] + src50[419] + src50[420] + src50[421] + src50[422] + src50[423] + src50[424] + src50[425] + src50[426] + src50[427] + src50[428] + src50[429] + src50[430] + src50[431] + src50[432] + src50[433] + src50[434] + src50[435] + src50[436] + src50[437] + src50[438] + src50[439] + src50[440] + src50[441] + src50[442] + src50[443] + src50[444] + src50[445] + src50[446] + src50[447] + src50[448] + src50[449] + src50[450] + src50[451] + src50[452] + src50[453] + src50[454] + src50[455] + src50[456] + src50[457] + src50[458] + src50[459] + src50[460] + src50[461] + src50[462] + src50[463] + src50[464] + src50[465] + src50[466] + src50[467] + src50[468] + src50[469] + src50[470] + src50[471] + src50[472] + src50[473] + src50[474] + src50[475] + src50[476] + src50[477] + src50[478] + src50[479] + src50[480] + src50[481] + src50[482] + src50[483] + src50[484] + src50[485])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63] + src51[64] + src51[65] + src51[66] + src51[67] + src51[68] + src51[69] + src51[70] + src51[71] + src51[72] + src51[73] + src51[74] + src51[75] + src51[76] + src51[77] + src51[78] + src51[79] + src51[80] + src51[81] + src51[82] + src51[83] + src51[84] + src51[85] + src51[86] + src51[87] + src51[88] + src51[89] + src51[90] + src51[91] + src51[92] + src51[93] + src51[94] + src51[95] + src51[96] + src51[97] + src51[98] + src51[99] + src51[100] + src51[101] + src51[102] + src51[103] + src51[104] + src51[105] + src51[106] + src51[107] + src51[108] + src51[109] + src51[110] + src51[111] + src51[112] + src51[113] + src51[114] + src51[115] + src51[116] + src51[117] + src51[118] + src51[119] + src51[120] + src51[121] + src51[122] + src51[123] + src51[124] + src51[125] + src51[126] + src51[127] + src51[128] + src51[129] + src51[130] + src51[131] + src51[132] + src51[133] + src51[134] + src51[135] + src51[136] + src51[137] + src51[138] + src51[139] + src51[140] + src51[141] + src51[142] + src51[143] + src51[144] + src51[145] + src51[146] + src51[147] + src51[148] + src51[149] + src51[150] + src51[151] + src51[152] + src51[153] + src51[154] + src51[155] + src51[156] + src51[157] + src51[158] + src51[159] + src51[160] + src51[161] + src51[162] + src51[163] + src51[164] + src51[165] + src51[166] + src51[167] + src51[168] + src51[169] + src51[170] + src51[171] + src51[172] + src51[173] + src51[174] + src51[175] + src51[176] + src51[177] + src51[178] + src51[179] + src51[180] + src51[181] + src51[182] + src51[183] + src51[184] + src51[185] + src51[186] + src51[187] + src51[188] + src51[189] + src51[190] + src51[191] + src51[192] + src51[193] + src51[194] + src51[195] + src51[196] + src51[197] + src51[198] + src51[199] + src51[200] + src51[201] + src51[202] + src51[203] + src51[204] + src51[205] + src51[206] + src51[207] + src51[208] + src51[209] + src51[210] + src51[211] + src51[212] + src51[213] + src51[214] + src51[215] + src51[216] + src51[217] + src51[218] + src51[219] + src51[220] + src51[221] + src51[222] + src51[223] + src51[224] + src51[225] + src51[226] + src51[227] + src51[228] + src51[229] + src51[230] + src51[231] + src51[232] + src51[233] + src51[234] + src51[235] + src51[236] + src51[237] + src51[238] + src51[239] + src51[240] + src51[241] + src51[242] + src51[243] + src51[244] + src51[245] + src51[246] + src51[247] + src51[248] + src51[249] + src51[250] + src51[251] + src51[252] + src51[253] + src51[254] + src51[255] + src51[256] + src51[257] + src51[258] + src51[259] + src51[260] + src51[261] + src51[262] + src51[263] + src51[264] + src51[265] + src51[266] + src51[267] + src51[268] + src51[269] + src51[270] + src51[271] + src51[272] + src51[273] + src51[274] + src51[275] + src51[276] + src51[277] + src51[278] + src51[279] + src51[280] + src51[281] + src51[282] + src51[283] + src51[284] + src51[285] + src51[286] + src51[287] + src51[288] + src51[289] + src51[290] + src51[291] + src51[292] + src51[293] + src51[294] + src51[295] + src51[296] + src51[297] + src51[298] + src51[299] + src51[300] + src51[301] + src51[302] + src51[303] + src51[304] + src51[305] + src51[306] + src51[307] + src51[308] + src51[309] + src51[310] + src51[311] + src51[312] + src51[313] + src51[314] + src51[315] + src51[316] + src51[317] + src51[318] + src51[319] + src51[320] + src51[321] + src51[322] + src51[323] + src51[324] + src51[325] + src51[326] + src51[327] + src51[328] + src51[329] + src51[330] + src51[331] + src51[332] + src51[333] + src51[334] + src51[335] + src51[336] + src51[337] + src51[338] + src51[339] + src51[340] + src51[341] + src51[342] + src51[343] + src51[344] + src51[345] + src51[346] + src51[347] + src51[348] + src51[349] + src51[350] + src51[351] + src51[352] + src51[353] + src51[354] + src51[355] + src51[356] + src51[357] + src51[358] + src51[359] + src51[360] + src51[361] + src51[362] + src51[363] + src51[364] + src51[365] + src51[366] + src51[367] + src51[368] + src51[369] + src51[370] + src51[371] + src51[372] + src51[373] + src51[374] + src51[375] + src51[376] + src51[377] + src51[378] + src51[379] + src51[380] + src51[381] + src51[382] + src51[383] + src51[384] + src51[385] + src51[386] + src51[387] + src51[388] + src51[389] + src51[390] + src51[391] + src51[392] + src51[393] + src51[394] + src51[395] + src51[396] + src51[397] + src51[398] + src51[399] + src51[400] + src51[401] + src51[402] + src51[403] + src51[404] + src51[405] + src51[406] + src51[407] + src51[408] + src51[409] + src51[410] + src51[411] + src51[412] + src51[413] + src51[414] + src51[415] + src51[416] + src51[417] + src51[418] + src51[419] + src51[420] + src51[421] + src51[422] + src51[423] + src51[424] + src51[425] + src51[426] + src51[427] + src51[428] + src51[429] + src51[430] + src51[431] + src51[432] + src51[433] + src51[434] + src51[435] + src51[436] + src51[437] + src51[438] + src51[439] + src51[440] + src51[441] + src51[442] + src51[443] + src51[444] + src51[445] + src51[446] + src51[447] + src51[448] + src51[449] + src51[450] + src51[451] + src51[452] + src51[453] + src51[454] + src51[455] + src51[456] + src51[457] + src51[458] + src51[459] + src51[460] + src51[461] + src51[462] + src51[463] + src51[464] + src51[465] + src51[466] + src51[467] + src51[468] + src51[469] + src51[470] + src51[471] + src51[472] + src51[473] + src51[474] + src51[475] + src51[476] + src51[477] + src51[478] + src51[479] + src51[480] + src51[481] + src51[482] + src51[483] + src51[484] + src51[485])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63] + src52[64] + src52[65] + src52[66] + src52[67] + src52[68] + src52[69] + src52[70] + src52[71] + src52[72] + src52[73] + src52[74] + src52[75] + src52[76] + src52[77] + src52[78] + src52[79] + src52[80] + src52[81] + src52[82] + src52[83] + src52[84] + src52[85] + src52[86] + src52[87] + src52[88] + src52[89] + src52[90] + src52[91] + src52[92] + src52[93] + src52[94] + src52[95] + src52[96] + src52[97] + src52[98] + src52[99] + src52[100] + src52[101] + src52[102] + src52[103] + src52[104] + src52[105] + src52[106] + src52[107] + src52[108] + src52[109] + src52[110] + src52[111] + src52[112] + src52[113] + src52[114] + src52[115] + src52[116] + src52[117] + src52[118] + src52[119] + src52[120] + src52[121] + src52[122] + src52[123] + src52[124] + src52[125] + src52[126] + src52[127] + src52[128] + src52[129] + src52[130] + src52[131] + src52[132] + src52[133] + src52[134] + src52[135] + src52[136] + src52[137] + src52[138] + src52[139] + src52[140] + src52[141] + src52[142] + src52[143] + src52[144] + src52[145] + src52[146] + src52[147] + src52[148] + src52[149] + src52[150] + src52[151] + src52[152] + src52[153] + src52[154] + src52[155] + src52[156] + src52[157] + src52[158] + src52[159] + src52[160] + src52[161] + src52[162] + src52[163] + src52[164] + src52[165] + src52[166] + src52[167] + src52[168] + src52[169] + src52[170] + src52[171] + src52[172] + src52[173] + src52[174] + src52[175] + src52[176] + src52[177] + src52[178] + src52[179] + src52[180] + src52[181] + src52[182] + src52[183] + src52[184] + src52[185] + src52[186] + src52[187] + src52[188] + src52[189] + src52[190] + src52[191] + src52[192] + src52[193] + src52[194] + src52[195] + src52[196] + src52[197] + src52[198] + src52[199] + src52[200] + src52[201] + src52[202] + src52[203] + src52[204] + src52[205] + src52[206] + src52[207] + src52[208] + src52[209] + src52[210] + src52[211] + src52[212] + src52[213] + src52[214] + src52[215] + src52[216] + src52[217] + src52[218] + src52[219] + src52[220] + src52[221] + src52[222] + src52[223] + src52[224] + src52[225] + src52[226] + src52[227] + src52[228] + src52[229] + src52[230] + src52[231] + src52[232] + src52[233] + src52[234] + src52[235] + src52[236] + src52[237] + src52[238] + src52[239] + src52[240] + src52[241] + src52[242] + src52[243] + src52[244] + src52[245] + src52[246] + src52[247] + src52[248] + src52[249] + src52[250] + src52[251] + src52[252] + src52[253] + src52[254] + src52[255] + src52[256] + src52[257] + src52[258] + src52[259] + src52[260] + src52[261] + src52[262] + src52[263] + src52[264] + src52[265] + src52[266] + src52[267] + src52[268] + src52[269] + src52[270] + src52[271] + src52[272] + src52[273] + src52[274] + src52[275] + src52[276] + src52[277] + src52[278] + src52[279] + src52[280] + src52[281] + src52[282] + src52[283] + src52[284] + src52[285] + src52[286] + src52[287] + src52[288] + src52[289] + src52[290] + src52[291] + src52[292] + src52[293] + src52[294] + src52[295] + src52[296] + src52[297] + src52[298] + src52[299] + src52[300] + src52[301] + src52[302] + src52[303] + src52[304] + src52[305] + src52[306] + src52[307] + src52[308] + src52[309] + src52[310] + src52[311] + src52[312] + src52[313] + src52[314] + src52[315] + src52[316] + src52[317] + src52[318] + src52[319] + src52[320] + src52[321] + src52[322] + src52[323] + src52[324] + src52[325] + src52[326] + src52[327] + src52[328] + src52[329] + src52[330] + src52[331] + src52[332] + src52[333] + src52[334] + src52[335] + src52[336] + src52[337] + src52[338] + src52[339] + src52[340] + src52[341] + src52[342] + src52[343] + src52[344] + src52[345] + src52[346] + src52[347] + src52[348] + src52[349] + src52[350] + src52[351] + src52[352] + src52[353] + src52[354] + src52[355] + src52[356] + src52[357] + src52[358] + src52[359] + src52[360] + src52[361] + src52[362] + src52[363] + src52[364] + src52[365] + src52[366] + src52[367] + src52[368] + src52[369] + src52[370] + src52[371] + src52[372] + src52[373] + src52[374] + src52[375] + src52[376] + src52[377] + src52[378] + src52[379] + src52[380] + src52[381] + src52[382] + src52[383] + src52[384] + src52[385] + src52[386] + src52[387] + src52[388] + src52[389] + src52[390] + src52[391] + src52[392] + src52[393] + src52[394] + src52[395] + src52[396] + src52[397] + src52[398] + src52[399] + src52[400] + src52[401] + src52[402] + src52[403] + src52[404] + src52[405] + src52[406] + src52[407] + src52[408] + src52[409] + src52[410] + src52[411] + src52[412] + src52[413] + src52[414] + src52[415] + src52[416] + src52[417] + src52[418] + src52[419] + src52[420] + src52[421] + src52[422] + src52[423] + src52[424] + src52[425] + src52[426] + src52[427] + src52[428] + src52[429] + src52[430] + src52[431] + src52[432] + src52[433] + src52[434] + src52[435] + src52[436] + src52[437] + src52[438] + src52[439] + src52[440] + src52[441] + src52[442] + src52[443] + src52[444] + src52[445] + src52[446] + src52[447] + src52[448] + src52[449] + src52[450] + src52[451] + src52[452] + src52[453] + src52[454] + src52[455] + src52[456] + src52[457] + src52[458] + src52[459] + src52[460] + src52[461] + src52[462] + src52[463] + src52[464] + src52[465] + src52[466] + src52[467] + src52[468] + src52[469] + src52[470] + src52[471] + src52[472] + src52[473] + src52[474] + src52[475] + src52[476] + src52[477] + src52[478] + src52[479] + src52[480] + src52[481] + src52[482] + src52[483] + src52[484] + src52[485])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63] + src53[64] + src53[65] + src53[66] + src53[67] + src53[68] + src53[69] + src53[70] + src53[71] + src53[72] + src53[73] + src53[74] + src53[75] + src53[76] + src53[77] + src53[78] + src53[79] + src53[80] + src53[81] + src53[82] + src53[83] + src53[84] + src53[85] + src53[86] + src53[87] + src53[88] + src53[89] + src53[90] + src53[91] + src53[92] + src53[93] + src53[94] + src53[95] + src53[96] + src53[97] + src53[98] + src53[99] + src53[100] + src53[101] + src53[102] + src53[103] + src53[104] + src53[105] + src53[106] + src53[107] + src53[108] + src53[109] + src53[110] + src53[111] + src53[112] + src53[113] + src53[114] + src53[115] + src53[116] + src53[117] + src53[118] + src53[119] + src53[120] + src53[121] + src53[122] + src53[123] + src53[124] + src53[125] + src53[126] + src53[127] + src53[128] + src53[129] + src53[130] + src53[131] + src53[132] + src53[133] + src53[134] + src53[135] + src53[136] + src53[137] + src53[138] + src53[139] + src53[140] + src53[141] + src53[142] + src53[143] + src53[144] + src53[145] + src53[146] + src53[147] + src53[148] + src53[149] + src53[150] + src53[151] + src53[152] + src53[153] + src53[154] + src53[155] + src53[156] + src53[157] + src53[158] + src53[159] + src53[160] + src53[161] + src53[162] + src53[163] + src53[164] + src53[165] + src53[166] + src53[167] + src53[168] + src53[169] + src53[170] + src53[171] + src53[172] + src53[173] + src53[174] + src53[175] + src53[176] + src53[177] + src53[178] + src53[179] + src53[180] + src53[181] + src53[182] + src53[183] + src53[184] + src53[185] + src53[186] + src53[187] + src53[188] + src53[189] + src53[190] + src53[191] + src53[192] + src53[193] + src53[194] + src53[195] + src53[196] + src53[197] + src53[198] + src53[199] + src53[200] + src53[201] + src53[202] + src53[203] + src53[204] + src53[205] + src53[206] + src53[207] + src53[208] + src53[209] + src53[210] + src53[211] + src53[212] + src53[213] + src53[214] + src53[215] + src53[216] + src53[217] + src53[218] + src53[219] + src53[220] + src53[221] + src53[222] + src53[223] + src53[224] + src53[225] + src53[226] + src53[227] + src53[228] + src53[229] + src53[230] + src53[231] + src53[232] + src53[233] + src53[234] + src53[235] + src53[236] + src53[237] + src53[238] + src53[239] + src53[240] + src53[241] + src53[242] + src53[243] + src53[244] + src53[245] + src53[246] + src53[247] + src53[248] + src53[249] + src53[250] + src53[251] + src53[252] + src53[253] + src53[254] + src53[255] + src53[256] + src53[257] + src53[258] + src53[259] + src53[260] + src53[261] + src53[262] + src53[263] + src53[264] + src53[265] + src53[266] + src53[267] + src53[268] + src53[269] + src53[270] + src53[271] + src53[272] + src53[273] + src53[274] + src53[275] + src53[276] + src53[277] + src53[278] + src53[279] + src53[280] + src53[281] + src53[282] + src53[283] + src53[284] + src53[285] + src53[286] + src53[287] + src53[288] + src53[289] + src53[290] + src53[291] + src53[292] + src53[293] + src53[294] + src53[295] + src53[296] + src53[297] + src53[298] + src53[299] + src53[300] + src53[301] + src53[302] + src53[303] + src53[304] + src53[305] + src53[306] + src53[307] + src53[308] + src53[309] + src53[310] + src53[311] + src53[312] + src53[313] + src53[314] + src53[315] + src53[316] + src53[317] + src53[318] + src53[319] + src53[320] + src53[321] + src53[322] + src53[323] + src53[324] + src53[325] + src53[326] + src53[327] + src53[328] + src53[329] + src53[330] + src53[331] + src53[332] + src53[333] + src53[334] + src53[335] + src53[336] + src53[337] + src53[338] + src53[339] + src53[340] + src53[341] + src53[342] + src53[343] + src53[344] + src53[345] + src53[346] + src53[347] + src53[348] + src53[349] + src53[350] + src53[351] + src53[352] + src53[353] + src53[354] + src53[355] + src53[356] + src53[357] + src53[358] + src53[359] + src53[360] + src53[361] + src53[362] + src53[363] + src53[364] + src53[365] + src53[366] + src53[367] + src53[368] + src53[369] + src53[370] + src53[371] + src53[372] + src53[373] + src53[374] + src53[375] + src53[376] + src53[377] + src53[378] + src53[379] + src53[380] + src53[381] + src53[382] + src53[383] + src53[384] + src53[385] + src53[386] + src53[387] + src53[388] + src53[389] + src53[390] + src53[391] + src53[392] + src53[393] + src53[394] + src53[395] + src53[396] + src53[397] + src53[398] + src53[399] + src53[400] + src53[401] + src53[402] + src53[403] + src53[404] + src53[405] + src53[406] + src53[407] + src53[408] + src53[409] + src53[410] + src53[411] + src53[412] + src53[413] + src53[414] + src53[415] + src53[416] + src53[417] + src53[418] + src53[419] + src53[420] + src53[421] + src53[422] + src53[423] + src53[424] + src53[425] + src53[426] + src53[427] + src53[428] + src53[429] + src53[430] + src53[431] + src53[432] + src53[433] + src53[434] + src53[435] + src53[436] + src53[437] + src53[438] + src53[439] + src53[440] + src53[441] + src53[442] + src53[443] + src53[444] + src53[445] + src53[446] + src53[447] + src53[448] + src53[449] + src53[450] + src53[451] + src53[452] + src53[453] + src53[454] + src53[455] + src53[456] + src53[457] + src53[458] + src53[459] + src53[460] + src53[461] + src53[462] + src53[463] + src53[464] + src53[465] + src53[466] + src53[467] + src53[468] + src53[469] + src53[470] + src53[471] + src53[472] + src53[473] + src53[474] + src53[475] + src53[476] + src53[477] + src53[478] + src53[479] + src53[480] + src53[481] + src53[482] + src53[483] + src53[484] + src53[485])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63] + src54[64] + src54[65] + src54[66] + src54[67] + src54[68] + src54[69] + src54[70] + src54[71] + src54[72] + src54[73] + src54[74] + src54[75] + src54[76] + src54[77] + src54[78] + src54[79] + src54[80] + src54[81] + src54[82] + src54[83] + src54[84] + src54[85] + src54[86] + src54[87] + src54[88] + src54[89] + src54[90] + src54[91] + src54[92] + src54[93] + src54[94] + src54[95] + src54[96] + src54[97] + src54[98] + src54[99] + src54[100] + src54[101] + src54[102] + src54[103] + src54[104] + src54[105] + src54[106] + src54[107] + src54[108] + src54[109] + src54[110] + src54[111] + src54[112] + src54[113] + src54[114] + src54[115] + src54[116] + src54[117] + src54[118] + src54[119] + src54[120] + src54[121] + src54[122] + src54[123] + src54[124] + src54[125] + src54[126] + src54[127] + src54[128] + src54[129] + src54[130] + src54[131] + src54[132] + src54[133] + src54[134] + src54[135] + src54[136] + src54[137] + src54[138] + src54[139] + src54[140] + src54[141] + src54[142] + src54[143] + src54[144] + src54[145] + src54[146] + src54[147] + src54[148] + src54[149] + src54[150] + src54[151] + src54[152] + src54[153] + src54[154] + src54[155] + src54[156] + src54[157] + src54[158] + src54[159] + src54[160] + src54[161] + src54[162] + src54[163] + src54[164] + src54[165] + src54[166] + src54[167] + src54[168] + src54[169] + src54[170] + src54[171] + src54[172] + src54[173] + src54[174] + src54[175] + src54[176] + src54[177] + src54[178] + src54[179] + src54[180] + src54[181] + src54[182] + src54[183] + src54[184] + src54[185] + src54[186] + src54[187] + src54[188] + src54[189] + src54[190] + src54[191] + src54[192] + src54[193] + src54[194] + src54[195] + src54[196] + src54[197] + src54[198] + src54[199] + src54[200] + src54[201] + src54[202] + src54[203] + src54[204] + src54[205] + src54[206] + src54[207] + src54[208] + src54[209] + src54[210] + src54[211] + src54[212] + src54[213] + src54[214] + src54[215] + src54[216] + src54[217] + src54[218] + src54[219] + src54[220] + src54[221] + src54[222] + src54[223] + src54[224] + src54[225] + src54[226] + src54[227] + src54[228] + src54[229] + src54[230] + src54[231] + src54[232] + src54[233] + src54[234] + src54[235] + src54[236] + src54[237] + src54[238] + src54[239] + src54[240] + src54[241] + src54[242] + src54[243] + src54[244] + src54[245] + src54[246] + src54[247] + src54[248] + src54[249] + src54[250] + src54[251] + src54[252] + src54[253] + src54[254] + src54[255] + src54[256] + src54[257] + src54[258] + src54[259] + src54[260] + src54[261] + src54[262] + src54[263] + src54[264] + src54[265] + src54[266] + src54[267] + src54[268] + src54[269] + src54[270] + src54[271] + src54[272] + src54[273] + src54[274] + src54[275] + src54[276] + src54[277] + src54[278] + src54[279] + src54[280] + src54[281] + src54[282] + src54[283] + src54[284] + src54[285] + src54[286] + src54[287] + src54[288] + src54[289] + src54[290] + src54[291] + src54[292] + src54[293] + src54[294] + src54[295] + src54[296] + src54[297] + src54[298] + src54[299] + src54[300] + src54[301] + src54[302] + src54[303] + src54[304] + src54[305] + src54[306] + src54[307] + src54[308] + src54[309] + src54[310] + src54[311] + src54[312] + src54[313] + src54[314] + src54[315] + src54[316] + src54[317] + src54[318] + src54[319] + src54[320] + src54[321] + src54[322] + src54[323] + src54[324] + src54[325] + src54[326] + src54[327] + src54[328] + src54[329] + src54[330] + src54[331] + src54[332] + src54[333] + src54[334] + src54[335] + src54[336] + src54[337] + src54[338] + src54[339] + src54[340] + src54[341] + src54[342] + src54[343] + src54[344] + src54[345] + src54[346] + src54[347] + src54[348] + src54[349] + src54[350] + src54[351] + src54[352] + src54[353] + src54[354] + src54[355] + src54[356] + src54[357] + src54[358] + src54[359] + src54[360] + src54[361] + src54[362] + src54[363] + src54[364] + src54[365] + src54[366] + src54[367] + src54[368] + src54[369] + src54[370] + src54[371] + src54[372] + src54[373] + src54[374] + src54[375] + src54[376] + src54[377] + src54[378] + src54[379] + src54[380] + src54[381] + src54[382] + src54[383] + src54[384] + src54[385] + src54[386] + src54[387] + src54[388] + src54[389] + src54[390] + src54[391] + src54[392] + src54[393] + src54[394] + src54[395] + src54[396] + src54[397] + src54[398] + src54[399] + src54[400] + src54[401] + src54[402] + src54[403] + src54[404] + src54[405] + src54[406] + src54[407] + src54[408] + src54[409] + src54[410] + src54[411] + src54[412] + src54[413] + src54[414] + src54[415] + src54[416] + src54[417] + src54[418] + src54[419] + src54[420] + src54[421] + src54[422] + src54[423] + src54[424] + src54[425] + src54[426] + src54[427] + src54[428] + src54[429] + src54[430] + src54[431] + src54[432] + src54[433] + src54[434] + src54[435] + src54[436] + src54[437] + src54[438] + src54[439] + src54[440] + src54[441] + src54[442] + src54[443] + src54[444] + src54[445] + src54[446] + src54[447] + src54[448] + src54[449] + src54[450] + src54[451] + src54[452] + src54[453] + src54[454] + src54[455] + src54[456] + src54[457] + src54[458] + src54[459] + src54[460] + src54[461] + src54[462] + src54[463] + src54[464] + src54[465] + src54[466] + src54[467] + src54[468] + src54[469] + src54[470] + src54[471] + src54[472] + src54[473] + src54[474] + src54[475] + src54[476] + src54[477] + src54[478] + src54[479] + src54[480] + src54[481] + src54[482] + src54[483] + src54[484] + src54[485])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63] + src55[64] + src55[65] + src55[66] + src55[67] + src55[68] + src55[69] + src55[70] + src55[71] + src55[72] + src55[73] + src55[74] + src55[75] + src55[76] + src55[77] + src55[78] + src55[79] + src55[80] + src55[81] + src55[82] + src55[83] + src55[84] + src55[85] + src55[86] + src55[87] + src55[88] + src55[89] + src55[90] + src55[91] + src55[92] + src55[93] + src55[94] + src55[95] + src55[96] + src55[97] + src55[98] + src55[99] + src55[100] + src55[101] + src55[102] + src55[103] + src55[104] + src55[105] + src55[106] + src55[107] + src55[108] + src55[109] + src55[110] + src55[111] + src55[112] + src55[113] + src55[114] + src55[115] + src55[116] + src55[117] + src55[118] + src55[119] + src55[120] + src55[121] + src55[122] + src55[123] + src55[124] + src55[125] + src55[126] + src55[127] + src55[128] + src55[129] + src55[130] + src55[131] + src55[132] + src55[133] + src55[134] + src55[135] + src55[136] + src55[137] + src55[138] + src55[139] + src55[140] + src55[141] + src55[142] + src55[143] + src55[144] + src55[145] + src55[146] + src55[147] + src55[148] + src55[149] + src55[150] + src55[151] + src55[152] + src55[153] + src55[154] + src55[155] + src55[156] + src55[157] + src55[158] + src55[159] + src55[160] + src55[161] + src55[162] + src55[163] + src55[164] + src55[165] + src55[166] + src55[167] + src55[168] + src55[169] + src55[170] + src55[171] + src55[172] + src55[173] + src55[174] + src55[175] + src55[176] + src55[177] + src55[178] + src55[179] + src55[180] + src55[181] + src55[182] + src55[183] + src55[184] + src55[185] + src55[186] + src55[187] + src55[188] + src55[189] + src55[190] + src55[191] + src55[192] + src55[193] + src55[194] + src55[195] + src55[196] + src55[197] + src55[198] + src55[199] + src55[200] + src55[201] + src55[202] + src55[203] + src55[204] + src55[205] + src55[206] + src55[207] + src55[208] + src55[209] + src55[210] + src55[211] + src55[212] + src55[213] + src55[214] + src55[215] + src55[216] + src55[217] + src55[218] + src55[219] + src55[220] + src55[221] + src55[222] + src55[223] + src55[224] + src55[225] + src55[226] + src55[227] + src55[228] + src55[229] + src55[230] + src55[231] + src55[232] + src55[233] + src55[234] + src55[235] + src55[236] + src55[237] + src55[238] + src55[239] + src55[240] + src55[241] + src55[242] + src55[243] + src55[244] + src55[245] + src55[246] + src55[247] + src55[248] + src55[249] + src55[250] + src55[251] + src55[252] + src55[253] + src55[254] + src55[255] + src55[256] + src55[257] + src55[258] + src55[259] + src55[260] + src55[261] + src55[262] + src55[263] + src55[264] + src55[265] + src55[266] + src55[267] + src55[268] + src55[269] + src55[270] + src55[271] + src55[272] + src55[273] + src55[274] + src55[275] + src55[276] + src55[277] + src55[278] + src55[279] + src55[280] + src55[281] + src55[282] + src55[283] + src55[284] + src55[285] + src55[286] + src55[287] + src55[288] + src55[289] + src55[290] + src55[291] + src55[292] + src55[293] + src55[294] + src55[295] + src55[296] + src55[297] + src55[298] + src55[299] + src55[300] + src55[301] + src55[302] + src55[303] + src55[304] + src55[305] + src55[306] + src55[307] + src55[308] + src55[309] + src55[310] + src55[311] + src55[312] + src55[313] + src55[314] + src55[315] + src55[316] + src55[317] + src55[318] + src55[319] + src55[320] + src55[321] + src55[322] + src55[323] + src55[324] + src55[325] + src55[326] + src55[327] + src55[328] + src55[329] + src55[330] + src55[331] + src55[332] + src55[333] + src55[334] + src55[335] + src55[336] + src55[337] + src55[338] + src55[339] + src55[340] + src55[341] + src55[342] + src55[343] + src55[344] + src55[345] + src55[346] + src55[347] + src55[348] + src55[349] + src55[350] + src55[351] + src55[352] + src55[353] + src55[354] + src55[355] + src55[356] + src55[357] + src55[358] + src55[359] + src55[360] + src55[361] + src55[362] + src55[363] + src55[364] + src55[365] + src55[366] + src55[367] + src55[368] + src55[369] + src55[370] + src55[371] + src55[372] + src55[373] + src55[374] + src55[375] + src55[376] + src55[377] + src55[378] + src55[379] + src55[380] + src55[381] + src55[382] + src55[383] + src55[384] + src55[385] + src55[386] + src55[387] + src55[388] + src55[389] + src55[390] + src55[391] + src55[392] + src55[393] + src55[394] + src55[395] + src55[396] + src55[397] + src55[398] + src55[399] + src55[400] + src55[401] + src55[402] + src55[403] + src55[404] + src55[405] + src55[406] + src55[407] + src55[408] + src55[409] + src55[410] + src55[411] + src55[412] + src55[413] + src55[414] + src55[415] + src55[416] + src55[417] + src55[418] + src55[419] + src55[420] + src55[421] + src55[422] + src55[423] + src55[424] + src55[425] + src55[426] + src55[427] + src55[428] + src55[429] + src55[430] + src55[431] + src55[432] + src55[433] + src55[434] + src55[435] + src55[436] + src55[437] + src55[438] + src55[439] + src55[440] + src55[441] + src55[442] + src55[443] + src55[444] + src55[445] + src55[446] + src55[447] + src55[448] + src55[449] + src55[450] + src55[451] + src55[452] + src55[453] + src55[454] + src55[455] + src55[456] + src55[457] + src55[458] + src55[459] + src55[460] + src55[461] + src55[462] + src55[463] + src55[464] + src55[465] + src55[466] + src55[467] + src55[468] + src55[469] + src55[470] + src55[471] + src55[472] + src55[473] + src55[474] + src55[475] + src55[476] + src55[477] + src55[478] + src55[479] + src55[480] + src55[481] + src55[482] + src55[483] + src55[484] + src55[485])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63] + src56[64] + src56[65] + src56[66] + src56[67] + src56[68] + src56[69] + src56[70] + src56[71] + src56[72] + src56[73] + src56[74] + src56[75] + src56[76] + src56[77] + src56[78] + src56[79] + src56[80] + src56[81] + src56[82] + src56[83] + src56[84] + src56[85] + src56[86] + src56[87] + src56[88] + src56[89] + src56[90] + src56[91] + src56[92] + src56[93] + src56[94] + src56[95] + src56[96] + src56[97] + src56[98] + src56[99] + src56[100] + src56[101] + src56[102] + src56[103] + src56[104] + src56[105] + src56[106] + src56[107] + src56[108] + src56[109] + src56[110] + src56[111] + src56[112] + src56[113] + src56[114] + src56[115] + src56[116] + src56[117] + src56[118] + src56[119] + src56[120] + src56[121] + src56[122] + src56[123] + src56[124] + src56[125] + src56[126] + src56[127] + src56[128] + src56[129] + src56[130] + src56[131] + src56[132] + src56[133] + src56[134] + src56[135] + src56[136] + src56[137] + src56[138] + src56[139] + src56[140] + src56[141] + src56[142] + src56[143] + src56[144] + src56[145] + src56[146] + src56[147] + src56[148] + src56[149] + src56[150] + src56[151] + src56[152] + src56[153] + src56[154] + src56[155] + src56[156] + src56[157] + src56[158] + src56[159] + src56[160] + src56[161] + src56[162] + src56[163] + src56[164] + src56[165] + src56[166] + src56[167] + src56[168] + src56[169] + src56[170] + src56[171] + src56[172] + src56[173] + src56[174] + src56[175] + src56[176] + src56[177] + src56[178] + src56[179] + src56[180] + src56[181] + src56[182] + src56[183] + src56[184] + src56[185] + src56[186] + src56[187] + src56[188] + src56[189] + src56[190] + src56[191] + src56[192] + src56[193] + src56[194] + src56[195] + src56[196] + src56[197] + src56[198] + src56[199] + src56[200] + src56[201] + src56[202] + src56[203] + src56[204] + src56[205] + src56[206] + src56[207] + src56[208] + src56[209] + src56[210] + src56[211] + src56[212] + src56[213] + src56[214] + src56[215] + src56[216] + src56[217] + src56[218] + src56[219] + src56[220] + src56[221] + src56[222] + src56[223] + src56[224] + src56[225] + src56[226] + src56[227] + src56[228] + src56[229] + src56[230] + src56[231] + src56[232] + src56[233] + src56[234] + src56[235] + src56[236] + src56[237] + src56[238] + src56[239] + src56[240] + src56[241] + src56[242] + src56[243] + src56[244] + src56[245] + src56[246] + src56[247] + src56[248] + src56[249] + src56[250] + src56[251] + src56[252] + src56[253] + src56[254] + src56[255] + src56[256] + src56[257] + src56[258] + src56[259] + src56[260] + src56[261] + src56[262] + src56[263] + src56[264] + src56[265] + src56[266] + src56[267] + src56[268] + src56[269] + src56[270] + src56[271] + src56[272] + src56[273] + src56[274] + src56[275] + src56[276] + src56[277] + src56[278] + src56[279] + src56[280] + src56[281] + src56[282] + src56[283] + src56[284] + src56[285] + src56[286] + src56[287] + src56[288] + src56[289] + src56[290] + src56[291] + src56[292] + src56[293] + src56[294] + src56[295] + src56[296] + src56[297] + src56[298] + src56[299] + src56[300] + src56[301] + src56[302] + src56[303] + src56[304] + src56[305] + src56[306] + src56[307] + src56[308] + src56[309] + src56[310] + src56[311] + src56[312] + src56[313] + src56[314] + src56[315] + src56[316] + src56[317] + src56[318] + src56[319] + src56[320] + src56[321] + src56[322] + src56[323] + src56[324] + src56[325] + src56[326] + src56[327] + src56[328] + src56[329] + src56[330] + src56[331] + src56[332] + src56[333] + src56[334] + src56[335] + src56[336] + src56[337] + src56[338] + src56[339] + src56[340] + src56[341] + src56[342] + src56[343] + src56[344] + src56[345] + src56[346] + src56[347] + src56[348] + src56[349] + src56[350] + src56[351] + src56[352] + src56[353] + src56[354] + src56[355] + src56[356] + src56[357] + src56[358] + src56[359] + src56[360] + src56[361] + src56[362] + src56[363] + src56[364] + src56[365] + src56[366] + src56[367] + src56[368] + src56[369] + src56[370] + src56[371] + src56[372] + src56[373] + src56[374] + src56[375] + src56[376] + src56[377] + src56[378] + src56[379] + src56[380] + src56[381] + src56[382] + src56[383] + src56[384] + src56[385] + src56[386] + src56[387] + src56[388] + src56[389] + src56[390] + src56[391] + src56[392] + src56[393] + src56[394] + src56[395] + src56[396] + src56[397] + src56[398] + src56[399] + src56[400] + src56[401] + src56[402] + src56[403] + src56[404] + src56[405] + src56[406] + src56[407] + src56[408] + src56[409] + src56[410] + src56[411] + src56[412] + src56[413] + src56[414] + src56[415] + src56[416] + src56[417] + src56[418] + src56[419] + src56[420] + src56[421] + src56[422] + src56[423] + src56[424] + src56[425] + src56[426] + src56[427] + src56[428] + src56[429] + src56[430] + src56[431] + src56[432] + src56[433] + src56[434] + src56[435] + src56[436] + src56[437] + src56[438] + src56[439] + src56[440] + src56[441] + src56[442] + src56[443] + src56[444] + src56[445] + src56[446] + src56[447] + src56[448] + src56[449] + src56[450] + src56[451] + src56[452] + src56[453] + src56[454] + src56[455] + src56[456] + src56[457] + src56[458] + src56[459] + src56[460] + src56[461] + src56[462] + src56[463] + src56[464] + src56[465] + src56[466] + src56[467] + src56[468] + src56[469] + src56[470] + src56[471] + src56[472] + src56[473] + src56[474] + src56[475] + src56[476] + src56[477] + src56[478] + src56[479] + src56[480] + src56[481] + src56[482] + src56[483] + src56[484] + src56[485])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63] + src57[64] + src57[65] + src57[66] + src57[67] + src57[68] + src57[69] + src57[70] + src57[71] + src57[72] + src57[73] + src57[74] + src57[75] + src57[76] + src57[77] + src57[78] + src57[79] + src57[80] + src57[81] + src57[82] + src57[83] + src57[84] + src57[85] + src57[86] + src57[87] + src57[88] + src57[89] + src57[90] + src57[91] + src57[92] + src57[93] + src57[94] + src57[95] + src57[96] + src57[97] + src57[98] + src57[99] + src57[100] + src57[101] + src57[102] + src57[103] + src57[104] + src57[105] + src57[106] + src57[107] + src57[108] + src57[109] + src57[110] + src57[111] + src57[112] + src57[113] + src57[114] + src57[115] + src57[116] + src57[117] + src57[118] + src57[119] + src57[120] + src57[121] + src57[122] + src57[123] + src57[124] + src57[125] + src57[126] + src57[127] + src57[128] + src57[129] + src57[130] + src57[131] + src57[132] + src57[133] + src57[134] + src57[135] + src57[136] + src57[137] + src57[138] + src57[139] + src57[140] + src57[141] + src57[142] + src57[143] + src57[144] + src57[145] + src57[146] + src57[147] + src57[148] + src57[149] + src57[150] + src57[151] + src57[152] + src57[153] + src57[154] + src57[155] + src57[156] + src57[157] + src57[158] + src57[159] + src57[160] + src57[161] + src57[162] + src57[163] + src57[164] + src57[165] + src57[166] + src57[167] + src57[168] + src57[169] + src57[170] + src57[171] + src57[172] + src57[173] + src57[174] + src57[175] + src57[176] + src57[177] + src57[178] + src57[179] + src57[180] + src57[181] + src57[182] + src57[183] + src57[184] + src57[185] + src57[186] + src57[187] + src57[188] + src57[189] + src57[190] + src57[191] + src57[192] + src57[193] + src57[194] + src57[195] + src57[196] + src57[197] + src57[198] + src57[199] + src57[200] + src57[201] + src57[202] + src57[203] + src57[204] + src57[205] + src57[206] + src57[207] + src57[208] + src57[209] + src57[210] + src57[211] + src57[212] + src57[213] + src57[214] + src57[215] + src57[216] + src57[217] + src57[218] + src57[219] + src57[220] + src57[221] + src57[222] + src57[223] + src57[224] + src57[225] + src57[226] + src57[227] + src57[228] + src57[229] + src57[230] + src57[231] + src57[232] + src57[233] + src57[234] + src57[235] + src57[236] + src57[237] + src57[238] + src57[239] + src57[240] + src57[241] + src57[242] + src57[243] + src57[244] + src57[245] + src57[246] + src57[247] + src57[248] + src57[249] + src57[250] + src57[251] + src57[252] + src57[253] + src57[254] + src57[255] + src57[256] + src57[257] + src57[258] + src57[259] + src57[260] + src57[261] + src57[262] + src57[263] + src57[264] + src57[265] + src57[266] + src57[267] + src57[268] + src57[269] + src57[270] + src57[271] + src57[272] + src57[273] + src57[274] + src57[275] + src57[276] + src57[277] + src57[278] + src57[279] + src57[280] + src57[281] + src57[282] + src57[283] + src57[284] + src57[285] + src57[286] + src57[287] + src57[288] + src57[289] + src57[290] + src57[291] + src57[292] + src57[293] + src57[294] + src57[295] + src57[296] + src57[297] + src57[298] + src57[299] + src57[300] + src57[301] + src57[302] + src57[303] + src57[304] + src57[305] + src57[306] + src57[307] + src57[308] + src57[309] + src57[310] + src57[311] + src57[312] + src57[313] + src57[314] + src57[315] + src57[316] + src57[317] + src57[318] + src57[319] + src57[320] + src57[321] + src57[322] + src57[323] + src57[324] + src57[325] + src57[326] + src57[327] + src57[328] + src57[329] + src57[330] + src57[331] + src57[332] + src57[333] + src57[334] + src57[335] + src57[336] + src57[337] + src57[338] + src57[339] + src57[340] + src57[341] + src57[342] + src57[343] + src57[344] + src57[345] + src57[346] + src57[347] + src57[348] + src57[349] + src57[350] + src57[351] + src57[352] + src57[353] + src57[354] + src57[355] + src57[356] + src57[357] + src57[358] + src57[359] + src57[360] + src57[361] + src57[362] + src57[363] + src57[364] + src57[365] + src57[366] + src57[367] + src57[368] + src57[369] + src57[370] + src57[371] + src57[372] + src57[373] + src57[374] + src57[375] + src57[376] + src57[377] + src57[378] + src57[379] + src57[380] + src57[381] + src57[382] + src57[383] + src57[384] + src57[385] + src57[386] + src57[387] + src57[388] + src57[389] + src57[390] + src57[391] + src57[392] + src57[393] + src57[394] + src57[395] + src57[396] + src57[397] + src57[398] + src57[399] + src57[400] + src57[401] + src57[402] + src57[403] + src57[404] + src57[405] + src57[406] + src57[407] + src57[408] + src57[409] + src57[410] + src57[411] + src57[412] + src57[413] + src57[414] + src57[415] + src57[416] + src57[417] + src57[418] + src57[419] + src57[420] + src57[421] + src57[422] + src57[423] + src57[424] + src57[425] + src57[426] + src57[427] + src57[428] + src57[429] + src57[430] + src57[431] + src57[432] + src57[433] + src57[434] + src57[435] + src57[436] + src57[437] + src57[438] + src57[439] + src57[440] + src57[441] + src57[442] + src57[443] + src57[444] + src57[445] + src57[446] + src57[447] + src57[448] + src57[449] + src57[450] + src57[451] + src57[452] + src57[453] + src57[454] + src57[455] + src57[456] + src57[457] + src57[458] + src57[459] + src57[460] + src57[461] + src57[462] + src57[463] + src57[464] + src57[465] + src57[466] + src57[467] + src57[468] + src57[469] + src57[470] + src57[471] + src57[472] + src57[473] + src57[474] + src57[475] + src57[476] + src57[477] + src57[478] + src57[479] + src57[480] + src57[481] + src57[482] + src57[483] + src57[484] + src57[485])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63] + src58[64] + src58[65] + src58[66] + src58[67] + src58[68] + src58[69] + src58[70] + src58[71] + src58[72] + src58[73] + src58[74] + src58[75] + src58[76] + src58[77] + src58[78] + src58[79] + src58[80] + src58[81] + src58[82] + src58[83] + src58[84] + src58[85] + src58[86] + src58[87] + src58[88] + src58[89] + src58[90] + src58[91] + src58[92] + src58[93] + src58[94] + src58[95] + src58[96] + src58[97] + src58[98] + src58[99] + src58[100] + src58[101] + src58[102] + src58[103] + src58[104] + src58[105] + src58[106] + src58[107] + src58[108] + src58[109] + src58[110] + src58[111] + src58[112] + src58[113] + src58[114] + src58[115] + src58[116] + src58[117] + src58[118] + src58[119] + src58[120] + src58[121] + src58[122] + src58[123] + src58[124] + src58[125] + src58[126] + src58[127] + src58[128] + src58[129] + src58[130] + src58[131] + src58[132] + src58[133] + src58[134] + src58[135] + src58[136] + src58[137] + src58[138] + src58[139] + src58[140] + src58[141] + src58[142] + src58[143] + src58[144] + src58[145] + src58[146] + src58[147] + src58[148] + src58[149] + src58[150] + src58[151] + src58[152] + src58[153] + src58[154] + src58[155] + src58[156] + src58[157] + src58[158] + src58[159] + src58[160] + src58[161] + src58[162] + src58[163] + src58[164] + src58[165] + src58[166] + src58[167] + src58[168] + src58[169] + src58[170] + src58[171] + src58[172] + src58[173] + src58[174] + src58[175] + src58[176] + src58[177] + src58[178] + src58[179] + src58[180] + src58[181] + src58[182] + src58[183] + src58[184] + src58[185] + src58[186] + src58[187] + src58[188] + src58[189] + src58[190] + src58[191] + src58[192] + src58[193] + src58[194] + src58[195] + src58[196] + src58[197] + src58[198] + src58[199] + src58[200] + src58[201] + src58[202] + src58[203] + src58[204] + src58[205] + src58[206] + src58[207] + src58[208] + src58[209] + src58[210] + src58[211] + src58[212] + src58[213] + src58[214] + src58[215] + src58[216] + src58[217] + src58[218] + src58[219] + src58[220] + src58[221] + src58[222] + src58[223] + src58[224] + src58[225] + src58[226] + src58[227] + src58[228] + src58[229] + src58[230] + src58[231] + src58[232] + src58[233] + src58[234] + src58[235] + src58[236] + src58[237] + src58[238] + src58[239] + src58[240] + src58[241] + src58[242] + src58[243] + src58[244] + src58[245] + src58[246] + src58[247] + src58[248] + src58[249] + src58[250] + src58[251] + src58[252] + src58[253] + src58[254] + src58[255] + src58[256] + src58[257] + src58[258] + src58[259] + src58[260] + src58[261] + src58[262] + src58[263] + src58[264] + src58[265] + src58[266] + src58[267] + src58[268] + src58[269] + src58[270] + src58[271] + src58[272] + src58[273] + src58[274] + src58[275] + src58[276] + src58[277] + src58[278] + src58[279] + src58[280] + src58[281] + src58[282] + src58[283] + src58[284] + src58[285] + src58[286] + src58[287] + src58[288] + src58[289] + src58[290] + src58[291] + src58[292] + src58[293] + src58[294] + src58[295] + src58[296] + src58[297] + src58[298] + src58[299] + src58[300] + src58[301] + src58[302] + src58[303] + src58[304] + src58[305] + src58[306] + src58[307] + src58[308] + src58[309] + src58[310] + src58[311] + src58[312] + src58[313] + src58[314] + src58[315] + src58[316] + src58[317] + src58[318] + src58[319] + src58[320] + src58[321] + src58[322] + src58[323] + src58[324] + src58[325] + src58[326] + src58[327] + src58[328] + src58[329] + src58[330] + src58[331] + src58[332] + src58[333] + src58[334] + src58[335] + src58[336] + src58[337] + src58[338] + src58[339] + src58[340] + src58[341] + src58[342] + src58[343] + src58[344] + src58[345] + src58[346] + src58[347] + src58[348] + src58[349] + src58[350] + src58[351] + src58[352] + src58[353] + src58[354] + src58[355] + src58[356] + src58[357] + src58[358] + src58[359] + src58[360] + src58[361] + src58[362] + src58[363] + src58[364] + src58[365] + src58[366] + src58[367] + src58[368] + src58[369] + src58[370] + src58[371] + src58[372] + src58[373] + src58[374] + src58[375] + src58[376] + src58[377] + src58[378] + src58[379] + src58[380] + src58[381] + src58[382] + src58[383] + src58[384] + src58[385] + src58[386] + src58[387] + src58[388] + src58[389] + src58[390] + src58[391] + src58[392] + src58[393] + src58[394] + src58[395] + src58[396] + src58[397] + src58[398] + src58[399] + src58[400] + src58[401] + src58[402] + src58[403] + src58[404] + src58[405] + src58[406] + src58[407] + src58[408] + src58[409] + src58[410] + src58[411] + src58[412] + src58[413] + src58[414] + src58[415] + src58[416] + src58[417] + src58[418] + src58[419] + src58[420] + src58[421] + src58[422] + src58[423] + src58[424] + src58[425] + src58[426] + src58[427] + src58[428] + src58[429] + src58[430] + src58[431] + src58[432] + src58[433] + src58[434] + src58[435] + src58[436] + src58[437] + src58[438] + src58[439] + src58[440] + src58[441] + src58[442] + src58[443] + src58[444] + src58[445] + src58[446] + src58[447] + src58[448] + src58[449] + src58[450] + src58[451] + src58[452] + src58[453] + src58[454] + src58[455] + src58[456] + src58[457] + src58[458] + src58[459] + src58[460] + src58[461] + src58[462] + src58[463] + src58[464] + src58[465] + src58[466] + src58[467] + src58[468] + src58[469] + src58[470] + src58[471] + src58[472] + src58[473] + src58[474] + src58[475] + src58[476] + src58[477] + src58[478] + src58[479] + src58[480] + src58[481] + src58[482] + src58[483] + src58[484] + src58[485])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63] + src59[64] + src59[65] + src59[66] + src59[67] + src59[68] + src59[69] + src59[70] + src59[71] + src59[72] + src59[73] + src59[74] + src59[75] + src59[76] + src59[77] + src59[78] + src59[79] + src59[80] + src59[81] + src59[82] + src59[83] + src59[84] + src59[85] + src59[86] + src59[87] + src59[88] + src59[89] + src59[90] + src59[91] + src59[92] + src59[93] + src59[94] + src59[95] + src59[96] + src59[97] + src59[98] + src59[99] + src59[100] + src59[101] + src59[102] + src59[103] + src59[104] + src59[105] + src59[106] + src59[107] + src59[108] + src59[109] + src59[110] + src59[111] + src59[112] + src59[113] + src59[114] + src59[115] + src59[116] + src59[117] + src59[118] + src59[119] + src59[120] + src59[121] + src59[122] + src59[123] + src59[124] + src59[125] + src59[126] + src59[127] + src59[128] + src59[129] + src59[130] + src59[131] + src59[132] + src59[133] + src59[134] + src59[135] + src59[136] + src59[137] + src59[138] + src59[139] + src59[140] + src59[141] + src59[142] + src59[143] + src59[144] + src59[145] + src59[146] + src59[147] + src59[148] + src59[149] + src59[150] + src59[151] + src59[152] + src59[153] + src59[154] + src59[155] + src59[156] + src59[157] + src59[158] + src59[159] + src59[160] + src59[161] + src59[162] + src59[163] + src59[164] + src59[165] + src59[166] + src59[167] + src59[168] + src59[169] + src59[170] + src59[171] + src59[172] + src59[173] + src59[174] + src59[175] + src59[176] + src59[177] + src59[178] + src59[179] + src59[180] + src59[181] + src59[182] + src59[183] + src59[184] + src59[185] + src59[186] + src59[187] + src59[188] + src59[189] + src59[190] + src59[191] + src59[192] + src59[193] + src59[194] + src59[195] + src59[196] + src59[197] + src59[198] + src59[199] + src59[200] + src59[201] + src59[202] + src59[203] + src59[204] + src59[205] + src59[206] + src59[207] + src59[208] + src59[209] + src59[210] + src59[211] + src59[212] + src59[213] + src59[214] + src59[215] + src59[216] + src59[217] + src59[218] + src59[219] + src59[220] + src59[221] + src59[222] + src59[223] + src59[224] + src59[225] + src59[226] + src59[227] + src59[228] + src59[229] + src59[230] + src59[231] + src59[232] + src59[233] + src59[234] + src59[235] + src59[236] + src59[237] + src59[238] + src59[239] + src59[240] + src59[241] + src59[242] + src59[243] + src59[244] + src59[245] + src59[246] + src59[247] + src59[248] + src59[249] + src59[250] + src59[251] + src59[252] + src59[253] + src59[254] + src59[255] + src59[256] + src59[257] + src59[258] + src59[259] + src59[260] + src59[261] + src59[262] + src59[263] + src59[264] + src59[265] + src59[266] + src59[267] + src59[268] + src59[269] + src59[270] + src59[271] + src59[272] + src59[273] + src59[274] + src59[275] + src59[276] + src59[277] + src59[278] + src59[279] + src59[280] + src59[281] + src59[282] + src59[283] + src59[284] + src59[285] + src59[286] + src59[287] + src59[288] + src59[289] + src59[290] + src59[291] + src59[292] + src59[293] + src59[294] + src59[295] + src59[296] + src59[297] + src59[298] + src59[299] + src59[300] + src59[301] + src59[302] + src59[303] + src59[304] + src59[305] + src59[306] + src59[307] + src59[308] + src59[309] + src59[310] + src59[311] + src59[312] + src59[313] + src59[314] + src59[315] + src59[316] + src59[317] + src59[318] + src59[319] + src59[320] + src59[321] + src59[322] + src59[323] + src59[324] + src59[325] + src59[326] + src59[327] + src59[328] + src59[329] + src59[330] + src59[331] + src59[332] + src59[333] + src59[334] + src59[335] + src59[336] + src59[337] + src59[338] + src59[339] + src59[340] + src59[341] + src59[342] + src59[343] + src59[344] + src59[345] + src59[346] + src59[347] + src59[348] + src59[349] + src59[350] + src59[351] + src59[352] + src59[353] + src59[354] + src59[355] + src59[356] + src59[357] + src59[358] + src59[359] + src59[360] + src59[361] + src59[362] + src59[363] + src59[364] + src59[365] + src59[366] + src59[367] + src59[368] + src59[369] + src59[370] + src59[371] + src59[372] + src59[373] + src59[374] + src59[375] + src59[376] + src59[377] + src59[378] + src59[379] + src59[380] + src59[381] + src59[382] + src59[383] + src59[384] + src59[385] + src59[386] + src59[387] + src59[388] + src59[389] + src59[390] + src59[391] + src59[392] + src59[393] + src59[394] + src59[395] + src59[396] + src59[397] + src59[398] + src59[399] + src59[400] + src59[401] + src59[402] + src59[403] + src59[404] + src59[405] + src59[406] + src59[407] + src59[408] + src59[409] + src59[410] + src59[411] + src59[412] + src59[413] + src59[414] + src59[415] + src59[416] + src59[417] + src59[418] + src59[419] + src59[420] + src59[421] + src59[422] + src59[423] + src59[424] + src59[425] + src59[426] + src59[427] + src59[428] + src59[429] + src59[430] + src59[431] + src59[432] + src59[433] + src59[434] + src59[435] + src59[436] + src59[437] + src59[438] + src59[439] + src59[440] + src59[441] + src59[442] + src59[443] + src59[444] + src59[445] + src59[446] + src59[447] + src59[448] + src59[449] + src59[450] + src59[451] + src59[452] + src59[453] + src59[454] + src59[455] + src59[456] + src59[457] + src59[458] + src59[459] + src59[460] + src59[461] + src59[462] + src59[463] + src59[464] + src59[465] + src59[466] + src59[467] + src59[468] + src59[469] + src59[470] + src59[471] + src59[472] + src59[473] + src59[474] + src59[475] + src59[476] + src59[477] + src59[478] + src59[479] + src59[480] + src59[481] + src59[482] + src59[483] + src59[484] + src59[485])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63] + src60[64] + src60[65] + src60[66] + src60[67] + src60[68] + src60[69] + src60[70] + src60[71] + src60[72] + src60[73] + src60[74] + src60[75] + src60[76] + src60[77] + src60[78] + src60[79] + src60[80] + src60[81] + src60[82] + src60[83] + src60[84] + src60[85] + src60[86] + src60[87] + src60[88] + src60[89] + src60[90] + src60[91] + src60[92] + src60[93] + src60[94] + src60[95] + src60[96] + src60[97] + src60[98] + src60[99] + src60[100] + src60[101] + src60[102] + src60[103] + src60[104] + src60[105] + src60[106] + src60[107] + src60[108] + src60[109] + src60[110] + src60[111] + src60[112] + src60[113] + src60[114] + src60[115] + src60[116] + src60[117] + src60[118] + src60[119] + src60[120] + src60[121] + src60[122] + src60[123] + src60[124] + src60[125] + src60[126] + src60[127] + src60[128] + src60[129] + src60[130] + src60[131] + src60[132] + src60[133] + src60[134] + src60[135] + src60[136] + src60[137] + src60[138] + src60[139] + src60[140] + src60[141] + src60[142] + src60[143] + src60[144] + src60[145] + src60[146] + src60[147] + src60[148] + src60[149] + src60[150] + src60[151] + src60[152] + src60[153] + src60[154] + src60[155] + src60[156] + src60[157] + src60[158] + src60[159] + src60[160] + src60[161] + src60[162] + src60[163] + src60[164] + src60[165] + src60[166] + src60[167] + src60[168] + src60[169] + src60[170] + src60[171] + src60[172] + src60[173] + src60[174] + src60[175] + src60[176] + src60[177] + src60[178] + src60[179] + src60[180] + src60[181] + src60[182] + src60[183] + src60[184] + src60[185] + src60[186] + src60[187] + src60[188] + src60[189] + src60[190] + src60[191] + src60[192] + src60[193] + src60[194] + src60[195] + src60[196] + src60[197] + src60[198] + src60[199] + src60[200] + src60[201] + src60[202] + src60[203] + src60[204] + src60[205] + src60[206] + src60[207] + src60[208] + src60[209] + src60[210] + src60[211] + src60[212] + src60[213] + src60[214] + src60[215] + src60[216] + src60[217] + src60[218] + src60[219] + src60[220] + src60[221] + src60[222] + src60[223] + src60[224] + src60[225] + src60[226] + src60[227] + src60[228] + src60[229] + src60[230] + src60[231] + src60[232] + src60[233] + src60[234] + src60[235] + src60[236] + src60[237] + src60[238] + src60[239] + src60[240] + src60[241] + src60[242] + src60[243] + src60[244] + src60[245] + src60[246] + src60[247] + src60[248] + src60[249] + src60[250] + src60[251] + src60[252] + src60[253] + src60[254] + src60[255] + src60[256] + src60[257] + src60[258] + src60[259] + src60[260] + src60[261] + src60[262] + src60[263] + src60[264] + src60[265] + src60[266] + src60[267] + src60[268] + src60[269] + src60[270] + src60[271] + src60[272] + src60[273] + src60[274] + src60[275] + src60[276] + src60[277] + src60[278] + src60[279] + src60[280] + src60[281] + src60[282] + src60[283] + src60[284] + src60[285] + src60[286] + src60[287] + src60[288] + src60[289] + src60[290] + src60[291] + src60[292] + src60[293] + src60[294] + src60[295] + src60[296] + src60[297] + src60[298] + src60[299] + src60[300] + src60[301] + src60[302] + src60[303] + src60[304] + src60[305] + src60[306] + src60[307] + src60[308] + src60[309] + src60[310] + src60[311] + src60[312] + src60[313] + src60[314] + src60[315] + src60[316] + src60[317] + src60[318] + src60[319] + src60[320] + src60[321] + src60[322] + src60[323] + src60[324] + src60[325] + src60[326] + src60[327] + src60[328] + src60[329] + src60[330] + src60[331] + src60[332] + src60[333] + src60[334] + src60[335] + src60[336] + src60[337] + src60[338] + src60[339] + src60[340] + src60[341] + src60[342] + src60[343] + src60[344] + src60[345] + src60[346] + src60[347] + src60[348] + src60[349] + src60[350] + src60[351] + src60[352] + src60[353] + src60[354] + src60[355] + src60[356] + src60[357] + src60[358] + src60[359] + src60[360] + src60[361] + src60[362] + src60[363] + src60[364] + src60[365] + src60[366] + src60[367] + src60[368] + src60[369] + src60[370] + src60[371] + src60[372] + src60[373] + src60[374] + src60[375] + src60[376] + src60[377] + src60[378] + src60[379] + src60[380] + src60[381] + src60[382] + src60[383] + src60[384] + src60[385] + src60[386] + src60[387] + src60[388] + src60[389] + src60[390] + src60[391] + src60[392] + src60[393] + src60[394] + src60[395] + src60[396] + src60[397] + src60[398] + src60[399] + src60[400] + src60[401] + src60[402] + src60[403] + src60[404] + src60[405] + src60[406] + src60[407] + src60[408] + src60[409] + src60[410] + src60[411] + src60[412] + src60[413] + src60[414] + src60[415] + src60[416] + src60[417] + src60[418] + src60[419] + src60[420] + src60[421] + src60[422] + src60[423] + src60[424] + src60[425] + src60[426] + src60[427] + src60[428] + src60[429] + src60[430] + src60[431] + src60[432] + src60[433] + src60[434] + src60[435] + src60[436] + src60[437] + src60[438] + src60[439] + src60[440] + src60[441] + src60[442] + src60[443] + src60[444] + src60[445] + src60[446] + src60[447] + src60[448] + src60[449] + src60[450] + src60[451] + src60[452] + src60[453] + src60[454] + src60[455] + src60[456] + src60[457] + src60[458] + src60[459] + src60[460] + src60[461] + src60[462] + src60[463] + src60[464] + src60[465] + src60[466] + src60[467] + src60[468] + src60[469] + src60[470] + src60[471] + src60[472] + src60[473] + src60[474] + src60[475] + src60[476] + src60[477] + src60[478] + src60[479] + src60[480] + src60[481] + src60[482] + src60[483] + src60[484] + src60[485])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63] + src61[64] + src61[65] + src61[66] + src61[67] + src61[68] + src61[69] + src61[70] + src61[71] + src61[72] + src61[73] + src61[74] + src61[75] + src61[76] + src61[77] + src61[78] + src61[79] + src61[80] + src61[81] + src61[82] + src61[83] + src61[84] + src61[85] + src61[86] + src61[87] + src61[88] + src61[89] + src61[90] + src61[91] + src61[92] + src61[93] + src61[94] + src61[95] + src61[96] + src61[97] + src61[98] + src61[99] + src61[100] + src61[101] + src61[102] + src61[103] + src61[104] + src61[105] + src61[106] + src61[107] + src61[108] + src61[109] + src61[110] + src61[111] + src61[112] + src61[113] + src61[114] + src61[115] + src61[116] + src61[117] + src61[118] + src61[119] + src61[120] + src61[121] + src61[122] + src61[123] + src61[124] + src61[125] + src61[126] + src61[127] + src61[128] + src61[129] + src61[130] + src61[131] + src61[132] + src61[133] + src61[134] + src61[135] + src61[136] + src61[137] + src61[138] + src61[139] + src61[140] + src61[141] + src61[142] + src61[143] + src61[144] + src61[145] + src61[146] + src61[147] + src61[148] + src61[149] + src61[150] + src61[151] + src61[152] + src61[153] + src61[154] + src61[155] + src61[156] + src61[157] + src61[158] + src61[159] + src61[160] + src61[161] + src61[162] + src61[163] + src61[164] + src61[165] + src61[166] + src61[167] + src61[168] + src61[169] + src61[170] + src61[171] + src61[172] + src61[173] + src61[174] + src61[175] + src61[176] + src61[177] + src61[178] + src61[179] + src61[180] + src61[181] + src61[182] + src61[183] + src61[184] + src61[185] + src61[186] + src61[187] + src61[188] + src61[189] + src61[190] + src61[191] + src61[192] + src61[193] + src61[194] + src61[195] + src61[196] + src61[197] + src61[198] + src61[199] + src61[200] + src61[201] + src61[202] + src61[203] + src61[204] + src61[205] + src61[206] + src61[207] + src61[208] + src61[209] + src61[210] + src61[211] + src61[212] + src61[213] + src61[214] + src61[215] + src61[216] + src61[217] + src61[218] + src61[219] + src61[220] + src61[221] + src61[222] + src61[223] + src61[224] + src61[225] + src61[226] + src61[227] + src61[228] + src61[229] + src61[230] + src61[231] + src61[232] + src61[233] + src61[234] + src61[235] + src61[236] + src61[237] + src61[238] + src61[239] + src61[240] + src61[241] + src61[242] + src61[243] + src61[244] + src61[245] + src61[246] + src61[247] + src61[248] + src61[249] + src61[250] + src61[251] + src61[252] + src61[253] + src61[254] + src61[255] + src61[256] + src61[257] + src61[258] + src61[259] + src61[260] + src61[261] + src61[262] + src61[263] + src61[264] + src61[265] + src61[266] + src61[267] + src61[268] + src61[269] + src61[270] + src61[271] + src61[272] + src61[273] + src61[274] + src61[275] + src61[276] + src61[277] + src61[278] + src61[279] + src61[280] + src61[281] + src61[282] + src61[283] + src61[284] + src61[285] + src61[286] + src61[287] + src61[288] + src61[289] + src61[290] + src61[291] + src61[292] + src61[293] + src61[294] + src61[295] + src61[296] + src61[297] + src61[298] + src61[299] + src61[300] + src61[301] + src61[302] + src61[303] + src61[304] + src61[305] + src61[306] + src61[307] + src61[308] + src61[309] + src61[310] + src61[311] + src61[312] + src61[313] + src61[314] + src61[315] + src61[316] + src61[317] + src61[318] + src61[319] + src61[320] + src61[321] + src61[322] + src61[323] + src61[324] + src61[325] + src61[326] + src61[327] + src61[328] + src61[329] + src61[330] + src61[331] + src61[332] + src61[333] + src61[334] + src61[335] + src61[336] + src61[337] + src61[338] + src61[339] + src61[340] + src61[341] + src61[342] + src61[343] + src61[344] + src61[345] + src61[346] + src61[347] + src61[348] + src61[349] + src61[350] + src61[351] + src61[352] + src61[353] + src61[354] + src61[355] + src61[356] + src61[357] + src61[358] + src61[359] + src61[360] + src61[361] + src61[362] + src61[363] + src61[364] + src61[365] + src61[366] + src61[367] + src61[368] + src61[369] + src61[370] + src61[371] + src61[372] + src61[373] + src61[374] + src61[375] + src61[376] + src61[377] + src61[378] + src61[379] + src61[380] + src61[381] + src61[382] + src61[383] + src61[384] + src61[385] + src61[386] + src61[387] + src61[388] + src61[389] + src61[390] + src61[391] + src61[392] + src61[393] + src61[394] + src61[395] + src61[396] + src61[397] + src61[398] + src61[399] + src61[400] + src61[401] + src61[402] + src61[403] + src61[404] + src61[405] + src61[406] + src61[407] + src61[408] + src61[409] + src61[410] + src61[411] + src61[412] + src61[413] + src61[414] + src61[415] + src61[416] + src61[417] + src61[418] + src61[419] + src61[420] + src61[421] + src61[422] + src61[423] + src61[424] + src61[425] + src61[426] + src61[427] + src61[428] + src61[429] + src61[430] + src61[431] + src61[432] + src61[433] + src61[434] + src61[435] + src61[436] + src61[437] + src61[438] + src61[439] + src61[440] + src61[441] + src61[442] + src61[443] + src61[444] + src61[445] + src61[446] + src61[447] + src61[448] + src61[449] + src61[450] + src61[451] + src61[452] + src61[453] + src61[454] + src61[455] + src61[456] + src61[457] + src61[458] + src61[459] + src61[460] + src61[461] + src61[462] + src61[463] + src61[464] + src61[465] + src61[466] + src61[467] + src61[468] + src61[469] + src61[470] + src61[471] + src61[472] + src61[473] + src61[474] + src61[475] + src61[476] + src61[477] + src61[478] + src61[479] + src61[480] + src61[481] + src61[482] + src61[483] + src61[484] + src61[485])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63] + src62[64] + src62[65] + src62[66] + src62[67] + src62[68] + src62[69] + src62[70] + src62[71] + src62[72] + src62[73] + src62[74] + src62[75] + src62[76] + src62[77] + src62[78] + src62[79] + src62[80] + src62[81] + src62[82] + src62[83] + src62[84] + src62[85] + src62[86] + src62[87] + src62[88] + src62[89] + src62[90] + src62[91] + src62[92] + src62[93] + src62[94] + src62[95] + src62[96] + src62[97] + src62[98] + src62[99] + src62[100] + src62[101] + src62[102] + src62[103] + src62[104] + src62[105] + src62[106] + src62[107] + src62[108] + src62[109] + src62[110] + src62[111] + src62[112] + src62[113] + src62[114] + src62[115] + src62[116] + src62[117] + src62[118] + src62[119] + src62[120] + src62[121] + src62[122] + src62[123] + src62[124] + src62[125] + src62[126] + src62[127] + src62[128] + src62[129] + src62[130] + src62[131] + src62[132] + src62[133] + src62[134] + src62[135] + src62[136] + src62[137] + src62[138] + src62[139] + src62[140] + src62[141] + src62[142] + src62[143] + src62[144] + src62[145] + src62[146] + src62[147] + src62[148] + src62[149] + src62[150] + src62[151] + src62[152] + src62[153] + src62[154] + src62[155] + src62[156] + src62[157] + src62[158] + src62[159] + src62[160] + src62[161] + src62[162] + src62[163] + src62[164] + src62[165] + src62[166] + src62[167] + src62[168] + src62[169] + src62[170] + src62[171] + src62[172] + src62[173] + src62[174] + src62[175] + src62[176] + src62[177] + src62[178] + src62[179] + src62[180] + src62[181] + src62[182] + src62[183] + src62[184] + src62[185] + src62[186] + src62[187] + src62[188] + src62[189] + src62[190] + src62[191] + src62[192] + src62[193] + src62[194] + src62[195] + src62[196] + src62[197] + src62[198] + src62[199] + src62[200] + src62[201] + src62[202] + src62[203] + src62[204] + src62[205] + src62[206] + src62[207] + src62[208] + src62[209] + src62[210] + src62[211] + src62[212] + src62[213] + src62[214] + src62[215] + src62[216] + src62[217] + src62[218] + src62[219] + src62[220] + src62[221] + src62[222] + src62[223] + src62[224] + src62[225] + src62[226] + src62[227] + src62[228] + src62[229] + src62[230] + src62[231] + src62[232] + src62[233] + src62[234] + src62[235] + src62[236] + src62[237] + src62[238] + src62[239] + src62[240] + src62[241] + src62[242] + src62[243] + src62[244] + src62[245] + src62[246] + src62[247] + src62[248] + src62[249] + src62[250] + src62[251] + src62[252] + src62[253] + src62[254] + src62[255] + src62[256] + src62[257] + src62[258] + src62[259] + src62[260] + src62[261] + src62[262] + src62[263] + src62[264] + src62[265] + src62[266] + src62[267] + src62[268] + src62[269] + src62[270] + src62[271] + src62[272] + src62[273] + src62[274] + src62[275] + src62[276] + src62[277] + src62[278] + src62[279] + src62[280] + src62[281] + src62[282] + src62[283] + src62[284] + src62[285] + src62[286] + src62[287] + src62[288] + src62[289] + src62[290] + src62[291] + src62[292] + src62[293] + src62[294] + src62[295] + src62[296] + src62[297] + src62[298] + src62[299] + src62[300] + src62[301] + src62[302] + src62[303] + src62[304] + src62[305] + src62[306] + src62[307] + src62[308] + src62[309] + src62[310] + src62[311] + src62[312] + src62[313] + src62[314] + src62[315] + src62[316] + src62[317] + src62[318] + src62[319] + src62[320] + src62[321] + src62[322] + src62[323] + src62[324] + src62[325] + src62[326] + src62[327] + src62[328] + src62[329] + src62[330] + src62[331] + src62[332] + src62[333] + src62[334] + src62[335] + src62[336] + src62[337] + src62[338] + src62[339] + src62[340] + src62[341] + src62[342] + src62[343] + src62[344] + src62[345] + src62[346] + src62[347] + src62[348] + src62[349] + src62[350] + src62[351] + src62[352] + src62[353] + src62[354] + src62[355] + src62[356] + src62[357] + src62[358] + src62[359] + src62[360] + src62[361] + src62[362] + src62[363] + src62[364] + src62[365] + src62[366] + src62[367] + src62[368] + src62[369] + src62[370] + src62[371] + src62[372] + src62[373] + src62[374] + src62[375] + src62[376] + src62[377] + src62[378] + src62[379] + src62[380] + src62[381] + src62[382] + src62[383] + src62[384] + src62[385] + src62[386] + src62[387] + src62[388] + src62[389] + src62[390] + src62[391] + src62[392] + src62[393] + src62[394] + src62[395] + src62[396] + src62[397] + src62[398] + src62[399] + src62[400] + src62[401] + src62[402] + src62[403] + src62[404] + src62[405] + src62[406] + src62[407] + src62[408] + src62[409] + src62[410] + src62[411] + src62[412] + src62[413] + src62[414] + src62[415] + src62[416] + src62[417] + src62[418] + src62[419] + src62[420] + src62[421] + src62[422] + src62[423] + src62[424] + src62[425] + src62[426] + src62[427] + src62[428] + src62[429] + src62[430] + src62[431] + src62[432] + src62[433] + src62[434] + src62[435] + src62[436] + src62[437] + src62[438] + src62[439] + src62[440] + src62[441] + src62[442] + src62[443] + src62[444] + src62[445] + src62[446] + src62[447] + src62[448] + src62[449] + src62[450] + src62[451] + src62[452] + src62[453] + src62[454] + src62[455] + src62[456] + src62[457] + src62[458] + src62[459] + src62[460] + src62[461] + src62[462] + src62[463] + src62[464] + src62[465] + src62[466] + src62[467] + src62[468] + src62[469] + src62[470] + src62[471] + src62[472] + src62[473] + src62[474] + src62[475] + src62[476] + src62[477] + src62[478] + src62[479] + src62[480] + src62[481] + src62[482] + src62[483] + src62[484] + src62[485])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63] + src63[64] + src63[65] + src63[66] + src63[67] + src63[68] + src63[69] + src63[70] + src63[71] + src63[72] + src63[73] + src63[74] + src63[75] + src63[76] + src63[77] + src63[78] + src63[79] + src63[80] + src63[81] + src63[82] + src63[83] + src63[84] + src63[85] + src63[86] + src63[87] + src63[88] + src63[89] + src63[90] + src63[91] + src63[92] + src63[93] + src63[94] + src63[95] + src63[96] + src63[97] + src63[98] + src63[99] + src63[100] + src63[101] + src63[102] + src63[103] + src63[104] + src63[105] + src63[106] + src63[107] + src63[108] + src63[109] + src63[110] + src63[111] + src63[112] + src63[113] + src63[114] + src63[115] + src63[116] + src63[117] + src63[118] + src63[119] + src63[120] + src63[121] + src63[122] + src63[123] + src63[124] + src63[125] + src63[126] + src63[127] + src63[128] + src63[129] + src63[130] + src63[131] + src63[132] + src63[133] + src63[134] + src63[135] + src63[136] + src63[137] + src63[138] + src63[139] + src63[140] + src63[141] + src63[142] + src63[143] + src63[144] + src63[145] + src63[146] + src63[147] + src63[148] + src63[149] + src63[150] + src63[151] + src63[152] + src63[153] + src63[154] + src63[155] + src63[156] + src63[157] + src63[158] + src63[159] + src63[160] + src63[161] + src63[162] + src63[163] + src63[164] + src63[165] + src63[166] + src63[167] + src63[168] + src63[169] + src63[170] + src63[171] + src63[172] + src63[173] + src63[174] + src63[175] + src63[176] + src63[177] + src63[178] + src63[179] + src63[180] + src63[181] + src63[182] + src63[183] + src63[184] + src63[185] + src63[186] + src63[187] + src63[188] + src63[189] + src63[190] + src63[191] + src63[192] + src63[193] + src63[194] + src63[195] + src63[196] + src63[197] + src63[198] + src63[199] + src63[200] + src63[201] + src63[202] + src63[203] + src63[204] + src63[205] + src63[206] + src63[207] + src63[208] + src63[209] + src63[210] + src63[211] + src63[212] + src63[213] + src63[214] + src63[215] + src63[216] + src63[217] + src63[218] + src63[219] + src63[220] + src63[221] + src63[222] + src63[223] + src63[224] + src63[225] + src63[226] + src63[227] + src63[228] + src63[229] + src63[230] + src63[231] + src63[232] + src63[233] + src63[234] + src63[235] + src63[236] + src63[237] + src63[238] + src63[239] + src63[240] + src63[241] + src63[242] + src63[243] + src63[244] + src63[245] + src63[246] + src63[247] + src63[248] + src63[249] + src63[250] + src63[251] + src63[252] + src63[253] + src63[254] + src63[255] + src63[256] + src63[257] + src63[258] + src63[259] + src63[260] + src63[261] + src63[262] + src63[263] + src63[264] + src63[265] + src63[266] + src63[267] + src63[268] + src63[269] + src63[270] + src63[271] + src63[272] + src63[273] + src63[274] + src63[275] + src63[276] + src63[277] + src63[278] + src63[279] + src63[280] + src63[281] + src63[282] + src63[283] + src63[284] + src63[285] + src63[286] + src63[287] + src63[288] + src63[289] + src63[290] + src63[291] + src63[292] + src63[293] + src63[294] + src63[295] + src63[296] + src63[297] + src63[298] + src63[299] + src63[300] + src63[301] + src63[302] + src63[303] + src63[304] + src63[305] + src63[306] + src63[307] + src63[308] + src63[309] + src63[310] + src63[311] + src63[312] + src63[313] + src63[314] + src63[315] + src63[316] + src63[317] + src63[318] + src63[319] + src63[320] + src63[321] + src63[322] + src63[323] + src63[324] + src63[325] + src63[326] + src63[327] + src63[328] + src63[329] + src63[330] + src63[331] + src63[332] + src63[333] + src63[334] + src63[335] + src63[336] + src63[337] + src63[338] + src63[339] + src63[340] + src63[341] + src63[342] + src63[343] + src63[344] + src63[345] + src63[346] + src63[347] + src63[348] + src63[349] + src63[350] + src63[351] + src63[352] + src63[353] + src63[354] + src63[355] + src63[356] + src63[357] + src63[358] + src63[359] + src63[360] + src63[361] + src63[362] + src63[363] + src63[364] + src63[365] + src63[366] + src63[367] + src63[368] + src63[369] + src63[370] + src63[371] + src63[372] + src63[373] + src63[374] + src63[375] + src63[376] + src63[377] + src63[378] + src63[379] + src63[380] + src63[381] + src63[382] + src63[383] + src63[384] + src63[385] + src63[386] + src63[387] + src63[388] + src63[389] + src63[390] + src63[391] + src63[392] + src63[393] + src63[394] + src63[395] + src63[396] + src63[397] + src63[398] + src63[399] + src63[400] + src63[401] + src63[402] + src63[403] + src63[404] + src63[405] + src63[406] + src63[407] + src63[408] + src63[409] + src63[410] + src63[411] + src63[412] + src63[413] + src63[414] + src63[415] + src63[416] + src63[417] + src63[418] + src63[419] + src63[420] + src63[421] + src63[422] + src63[423] + src63[424] + src63[425] + src63[426] + src63[427] + src63[428] + src63[429] + src63[430] + src63[431] + src63[432] + src63[433] + src63[434] + src63[435] + src63[436] + src63[437] + src63[438] + src63[439] + src63[440] + src63[441] + src63[442] + src63[443] + src63[444] + src63[445] + src63[446] + src63[447] + src63[448] + src63[449] + src63[450] + src63[451] + src63[452] + src63[453] + src63[454] + src63[455] + src63[456] + src63[457] + src63[458] + src63[459] + src63[460] + src63[461] + src63[462] + src63[463] + src63[464] + src63[465] + src63[466] + src63[467] + src63[468] + src63[469] + src63[470] + src63[471] + src63[472] + src63[473] + src63[474] + src63[475] + src63[476] + src63[477] + src63[478] + src63[479] + src63[480] + src63[481] + src63[482] + src63[483] + src63[484] + src63[485])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69) + ((dst70[0])<<70) + ((dst71[0])<<71) + ((dst72[0])<<72);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h7f2b80ba386822b37c7039f05f0ac3cfba3c03405803ec087b019329ddca2abb89f1d553274eece4c733ef0f01d338c6b34cefeaf03131160fdcf32af33f951961a3a184bbf4607c96079895fcab768f69db9dcb51573c165db2c8f22aab45a2311bb2305d63a9994fef4b12a01956405d0c64618e00f5852517370d0b86437cbee0437e83644e5d8e0c56b7e9773d2d3b08fa7811899e4d771bdca4d88d98f8a5b600ef21a62bd9134445d71827d00a11bdac30909b95bed272e88f1f3af0c1b154d5b6dac1c1c4a30aa536e2d7edb0cd89e5f203ed1e38772b8be0dc785103664d273c19e69fdaf3ffafd7c797aa944ff036975805cb202de9fe778c08f9f08baf2d4ee9a5fd513495dc945546b11b264199083b0a0deb958b2a9cebba8a38f62bc341cbca76519e206039ebeb14bcef02ec01ccd8a28369fc69bccd43870f6b039e47332c64461b09fb0854c7d67b2af6b527da36f75dff65edcd2e75692bc2d80bf94a18bd28278dd4d3d52d13d761daccad4fb9a20e602279f33a7c71b8998d1eeb19ddd7b01cf31a06381e15e8058e57c66aaf141f2c894149939a37ffb5fa9f3ffd4b9960e265be94d2c6e3fd6e7429a70a4ea67f628fbab8d2656d387b37f93495bb1497c6dc845b376917a3eb256b76befdded2454b1bf05b57787360cb897f4d0de941c24ad7fe9b7587a5d0251b387ea815d4631bfdf80e69fd8c9f47a1ad0cc5ddf96955103df7e017728c81bf4e8e54b6d07f9a69bd64f91b53da18eae0b81813efa2eb3b2c7fa72e0fe7d0c55b1b0bd13d6fb5f37a92fbdfed7808c4cb5d9573ad2cdfcf3ae5d8c1a59781b810326c756a8a893e2f1e065ceaf346d41774762c56856dd9f7159c9f6c6b79178c305f4dd0a62ec20c9eaf7fb20fdaf4a24f960a5bb8539d0030d7e645d53a1c694b01de72c118eb3d44830481b6136c2ff4cb128d5e669bf2234edef16546e12e0e7c8904aeffa35f9d03a14f790a7521dcd309109f1853c8bb8abd070a57ab63339681ac49fdff0404d3341b418032e8abced7ee0f94bec6332cf6d849fa81c1a6aea987be1dce480e2f9d2cf391d56af0a333ef8396106216a54ef0ecf105c6c956457d97561f64400f7a34a920678b5c87c4076d9ee808a2784ae03c1bd4a101ee10e7348126bbef9f51b843f8ee6dfc2ac95e0741cf1892bc0c87bda904e48eeee5423e805e450685a62be0dd45943abc92ea1b23c900b9e4f9c5eaf3e5df6c0964e8c25ca6c11f97726e78451a8290574ea72f5b09d8e26261686ef663a5af8ce94ed477d11f04ccca9f94b1966f8b29ec8134f856b8a52994d3c87763972655a13e1a33b2656be7da362cc6fe9c0eb1384af855953d92a9eff401b07f229c26455e33be0100796098d0c787ada16e4b8df3988e2c9b2bf5412f0fc8db595593c0cb1cf29f24c0c1b7ceb5e59a78b1ccdc013d07539662e25e811acb3b0b6b1b18563c7bcbca07a17139033f93f85c3f80411ef5c049e0faf678b02d4d5b229ae7c1c3cd0fc0b1d8e51fd44a1807c1e797c7b1aca6a789f89430dc4cf08fb63298ecdff47ce53f0855ee44bb30633ba7980bac516fa90b51ccdee96feb2aac95ce5e8ab13aa2dc58b8674a51df57d4c7ae4c6962eb7751181cf4cf024fce1ed411e8fbbbcb4544f5e9141d3ff57d2471f8310e872f9f3773296052b2c6af99ea0d5cb5236ba4cb28cdb76be42321babd8bed57dd02a67ef6b66249f8f99e5ce7e8be0ce816fb12e9225ab3c072a418a4777f4311dc0531b03a1f8791c2d124a573c68c48da7bd4443850e423d715cd0f4c8222e79d2c1abf1188a1d3cd418a23986e3ef87a19e4017087b6ea368ba296e1fcb75f520db540ea131754adfd3b2b552de346fd8c38123e532223964cb091dcf4d422c76cdc017711c8d9366ceceaa206d66f4b6994d955e38528c8118c51ed73ade23b87caa705c17f753079707bd4fca4ed80b678779c4d9b7f0f0bca9720490ca6cc6fd31aa7462622ef8f597dd8cede03fee524e1886d3be82761d28959655744cc21576d1fc2498ce17c0994c2a85a88aca3245568affd9c380b431e1ed5d92528123e0b5f9821ef4d57c204f15a9e383eecc8c895bf41fd48695ed5328ab2b623d44ba40587dca5066b719a719c39048a6c5207119aa7bb694c2aa13979fe85b5f7ce039055eed48a5ed6105a17d49abdd9fadbde06ffb14751fe5647952f63e07b035b78c72cdc2df81e5fc8ecf0c8c38b0cd05912ae695c498dce781bbaa0be9edfa7665de348d0460a08013ac462d4b3c6420936524c3ebb91348b56c33ffbaa10aee1f0c96d466dfa14cdadfd51d69712aa405cc5a1f5e35a4402ea39374eb78d3852c036b5f130a5b1571945c746d63243385ed23e4f82e0d1f948f5668a51fcf3e1a37fba380cd81cce494f5beddc560204d589303755cf38e7464129727136c6bafe81395db0db44794021c1e24fb958e1769f8e72f83a24fc8eb7634ab1fc23ce14771bcc92c64d7c15b891cc438726a757e18b242f96232f348425e702b5c1c49984d244945b69fb469f2b20ad414044a52003f1f036dcce35df67d67bd931e8bc0685711561a0e000a9084038f5d52c37b84c5343961444d129f857ea2a113d63c0c05c900bfca5296f2027213b2132b07277dfa593a3940fac7f81d42262cffd43756202d1dfac329e528d4d5b7fb25f47fa5fcec0ecb7eb8ac5342f6a64d3d536433f58f8a1f721fdd447d2c6a1682f6eb4d4f2f50dae332f6fdf23c835116a924414fad708a617f00490c23b4058319ac5358c67b40c97bd37cbad0b1b5d3c774448f8d459120e780f4da86a16c1ecbca369b6292fedd2292ba5a8c9ae98a625af16ef8970a231ea5eb7af2e60a593dc9932e959861a35f468f02bdc4b0fd9c25ebef4a048a3e200eba97a9a62e6f80e1a30eb25e1e202e24d9a3f7f85f8159c60066570f3f8b509efd2495708a5834a3f1ddc8210159bb95f3c6db2166b9cfc324e963e2e8b2412fe2ee44d2c9205a2a608d90162c48c91b191384c83467a48e74e503babb98f836e6ccf5947c48f2610a9e0aa1e76eb369a5d27b2a9516ce1c53e64e84b53e0afddb824e791af6d5aabf866b28af5cb46f294e162ef3f9220bd47725a1153074453713c7ed6f94543e334120196e6cfed79cf78414033799f0e139f42b3be807f6dce03151211fe4676ba03cf53bffbb178012274766010dec5a3ac8b126b9f48b6b3443d2520c78550612b5abfc6d2da7464b538a8636ce33c95c24ba8a5e937353e71e8f5928b0ed11c0d66d131c44594e5ad1264e094cc5fa72e9ed4a37ab638dc8caa63e49e0095a614e43b55f838d96aa9cc51a19ef579d9fd386ab3756b84379758a19b7516de286570e778b50d9ed56f8ad5ed4ba42b5b453dceebee7dea3960c4aa575449a750ba2c3437dcb2f6d68b73efed01adcd62f31e3059c3a362c0b35d5c741d3833a5473247bf832922ea2bf84f1a67da43837643624de65ff09b78f3c73170994fdd22cb0d3b416044f38e14072ac7deaa6e3c010225851959225a1eb220c0c59b619d5cf493ed50fcb49a53f38203891de029e8e2745df79ac29b1526522d6b2632d648856fa710d7a5336a01caf9fef0b7a94b8b998e895e1937e9e97132addbeeb13d0834dd7b4aeb7de4e30880520db5980fbda51a5bff05783daa2115c6c22ecab75a621fe4191e4e9b6ea61e0dc76a52cab7d5e6c35e49894e1a7f9c4af1146f83aefe3a9b02a7b3640f8a7c1e3b379434c6d36b6e9aa3207380aaba7281f6635400f4282538cf6708bcc0c5d786c07c5d14ded58122c5084489d1e9854062f44f954f50ff83c29fa8d80711f9fafd3b7038b06fec8f568a735fe26b552d51a63d6c0b90e06afad8e588d9001a621cbdfc039127b9d49cb6fd7378b26052f6c680d58908d0fe4feaac78c2e70e22d9c01f47abd398436a8d8ad22085b335c317e300f5dba422ec0d422158fd0be9bd73cfe1377c1b88ca9e4a2f5361bd2fceef274c7eff811fee2c32c44617495bb73e62101e71dda2331f813937820f3a982a456ee57107f4956dd3ff4b29a5e960e2922d10efeb8bc377b8f5a5ab562413bd4370221b9b909347cab7bce5c9e66e29b105a1c48d6f35d1885585c52962421e1cafed19c701904450315fcbef0f5abc92b1ec26167543bdb8daa0ee1d406d0f0a18d79ad1e054923e01b44207678f9e84987f1092fe161fcfe2e081e7976068c0d9c0c4d98ef92f8fadc18eb2e4ec162f6aa4e2f4f79386ced607d9802f4f668a863c04407a074274cfb619f90aeff670e3d0b31985c4f028722fa9b0d48ffd95b0fcc0dd96a614492e9fb16f675804fb2d9c3dc2d1e902250a3d80b0cdc632f5b945c2ce762d501030dd1fc3efb022095de07a932c284630c1c7212e658ab2eaf6e3a04664df87dbb6d5d09a9bc5b81b94d800eae7c43cb7fee48b19d907850932946c06552a313f26f1687943ac413dc843711c9e9255f7e81bd52c6316f959564bb86e4dde1cad6b59fa2bb6c63c32658bcb1c44d296e72c077e83d999212c2d7f0eeb5dae64ce6954086ad8b0f8317034a6124e023a4aa4413bb9a4f1ce8caf2fdcd96996b5113420a4f85487de5404c8881c0906fd901c392d33a84671858496a24db43896b86149fc9fcf4e6babc547d757cb06a82097208e9469984e7587c6d30a9e761bcb99513bd3c3f134c6ccf7644ee8926f902706f67a7d76aebd3402c2be501fa3c2819949181181d8daf5e569cd05d4413a63aeed214c04f6274344f44c54bd3bfd736c1466a2b6122e62c419337852c21c418c65a0f32e434b28dc052095c462311845d62ce9db4d8587b31bd6f5d48a89068fc62eb4e7a00948e1aee35287a9d587e29fb4aae7e779136c54c898a9a032bd78779db03782213f5434a5f1606a7b844d3610fa4b13e0d3ac36a85968d66a5d4c1e4bf64e1b7e47ee2dcda1b7479309b5ad2bd5da6bec5f574c1d9285a48ec27003f7f4b12564d9736787bb86f78b7e7cbd4862d33e0fb9fdee1a36541e8eabce675f0282fd8228c8b06cacd273da871dd94daa6d0448f429addeda75b8fb2ba94b11f417a203075961e6bbee58bec3c8d68c8e315830647e2c72c7bb22361def16bf381ff28d0dee6feb72e82b9deb3527855f38a580872f11d907e1583c32e6016973ea7df59cfc1a88a422268af1c72bc00e89e97cd48bd38ebe5932ad009743fa574f25211eb6293a11890dead645686205d46f41224071fcb1a8c57ac8022fe68bbb4e2fa33f323c4e18dd221200d395f59bea8849e918b7a856eb1e9b7b9105e422d166bf02618a81dbc9fe5f037d9aadc76dd778c551015a20709132447cafe444e2a02085ba027ac6da3feb2959872856d044e546c4691363a6736f0e8012270591306afc0b5a157c1768d6db74080ac5c72e22d4a0d69aa7f4dfab4dc73e81a24739077e9b7750d3c585fe0baa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3210c223ee4abea4b7975b7cb5a5f0e8e39f85218c588bb10a94ada36ad5fc295da513461568af5ff277e4477048bda7d6b95e5f2c289bf68f0afa9cdd45a1249ca8fe99a5e732e37f865d834ebd430c9f3043e4f3fc6becec4211b0fa335fbd03f9039634e0c4f58f46d2a8ca7e29b1f2ecff84a6a145f92e8f850953eb7786ca1d50e7d68e103ff2df092f4dc146c50a038efc510be48d791f87e6c8a36168a79d9e4feb1abe19529b8f5b090808404977b7c388d56bf1eaa7a5104a6d10a650e30ad47a8305d2aacb21fa5036306b74986685f770207402849d8527218d85c3efa8b08decf29ab39ac8932551a57357b2a67d2af92cf6ce92b8a1a797ed316f063f4980398e16e136ece5e62f9798f5723c3b969474dfbd3658709137e2c7606be425a9b4c7e1ab54c02a11f3a1157bec0774cefe7035b0d1a06ed9733bb5952891e3e4ef85b774baff27226aeb23ff4b5c174e220ddfaf08362e0dca5a8d17565221d3e1093b85934a57eac074a5427797d26d91fcfd6cd03af9a640145c543e46150301769b5054c0476cbee2c72a0fe75c288e21a74a80f4a865d95123b7cd58a95c33866c73900f63fcb8f6b3d288a1080a38e16f0538c1259db51c4aefa95ce7c4b3a53f3001c106f1a81d449ac114623ee85ac2a55dee043f0072889e16f5a5a5ce6e1de26df4b1dcbec9b230cc6727822891c1d00259212f013a3396be87d7294b740c27dbbf79682ccf03fcef521f341d090c8fee5381fdfc142f7951e2885719b69e0b26928a1263f0db244163ce561611631732166d7c7cba3f20a87e99b70abf40de4019ed5a8c5dcf03ce5d98d103ccf8c1a0826f556ac81d55a0d003138a84564c92f762fb0d5f69d1ef488f3b7906e9c17fcab5426c42fff1e7a1b00896d47cab3155a88a324682f762a06b9e28f8c9906f294ab8266b2d12639173f769ebea89b4cdbb695ad4f53ef61707ff4f3e82c310fa6b5808ec04d6565d12d384b124b0c1b0fb9c5233c089442cdf9496279455d8e206f68b2f15a8f6dbb6c1d643169c831578f35b730ad8a57518ade799aa3220162318d90717312e536b179b303377746757db92e687acfb5ea91c5675b6472b620514f9dd2c5366158d0a3cab17238eb08c74396b299d11b6a033edabf9955fc30ba0b335ed389852863fb2e8dde6852fa17a1853ca9e603955a63252b97e758c42cb0bc0584c51a6c7163b87d542e3341da1c277d571ae746b9196ba56199aef3ad87c1dd3e7edfdb078ba48a429247b2c465e1d9c61ca714cbd181824466166ebace2333128b2f7b4c1481947241afca3e6a8ea84451343646090a48d52080271e1e2d65f865ff68bfacacfe453f37551b717cbd7a12e492322ad5f4afabf0cab778493b952209eb04ebf5f3c3f989e80cddf9835dbdf051aa47d2395b04d0f2109c5488de820f36791f104ae1cad03b125df7076d14f3084d3ced725ab704a1c7f7b11e802feaacec332fe0b5bf35a5f8167ad176b74d7c6eb97334a381d7b127255a695fcfbaa6ade78fffc50f7a4a32cf043eb8082ac0e6b3ea7ec813ea34a1cc5bab1fe52f68191e1e78daebaf14da88628080ea8e446d2edab13a4a569c927cfc336ee831241c4d98d3b93a9d9bcd742538ad8c95b8ad87c23f413760d67556e838fb3ed56d246c4565218f7df81d57b9e23aae3c8e26ac8748eb3dcd78b9f072cd65787661730bd285f9d440acb9b0c9612ab6fd3a8293f205141563ba961a29fb1ccce1e1726af648a6b0674c8533d31e7a3d5177a0d8bd6d0ae48e2e9c6b8800e5ba72030ef7350847a3ccba8753c80f8969cd68f80727086c2bd1a69b7579196b608afd72822fba81c4d31b783ceb6510a42088ee7f7fcee8f68a09c6eaa70ad13daa05d8fc5236e59f42badcc84646d9526f7b3de792677e536bf7ce1c6f500b1e571af393d4f47491e0318860ec653f3f60ccd028ca642f68042f2ad667443d6a1d25ba9c44fd664823f8df10d61acdbb4e543241fb8ecf744cd0640ea6e0612c508fcaa0ceba4a0f090737e779ce36ab97368a529777d8cfb7762cb36d79036603ded2a12e827285e84e2a7cbfd9ec3d834a87f4644e62058a7224e6d89247dc89cd37643d84e6699aa13fc004cdb96da5c00c9ff12790165350ce9543514cc52f23b690be381c2aaa891d7eae22285741b36f9bc7b1c1f8b8bd2bdeb9ed588332a4e31726c4d8cfd5e3f5e9218c6703ecd45dbda2969bf60f31fb1869be49cf47fcbe863c336ae97cd91ad69489a1bb2eafa908100b6b9cae010b39e04fb577998af16d7db8d1deb568d71c2ce82b71fe843deb261b1858471af65485001200f087b1af7800719dff64e3bd8e2576b419afb3e3f007e0195be6f2867feea5b524a58d107c29e41c40fa02744f44f365d66bc14686363bd290ad4f00b24354a69d26bedf8506e083e2046a591d791d271f900403cbccea6448508899b719e7671cf7190ca0d06287d36df65dc2a88b9fe3627cea1c60a42bd2b3dc6309333a8dac7ecd15946411278caafa4dc94310260a83b84fe7c2197f881b6906ed7d79ac9665c1dd6bd5af6e0f86f540fec629eee509b860681c3c040de2a3c6aadf494901a35b9caacf2b165727bf989b3792c49fc1d89c8c7572f6bf83b331e6a3624d94b78c68f70aec344d24e09587c469238ebe0d4893fd6debf5ce5e30663e7bfb401f2dd774237bcb9e6d8c2bd96a1e33cdfd30d41f7be2c25d57036eafa9be04bb194a86f9fb2ed25c8f413e06b8369978a7c3d16c99080dc49caba9396c6328d974fda475c9ae7d20c5ca28cc4f9067407b002cb7a28448bdfb3e6c59f626f87cfa419d5cc37d0bef47c3b5554d098a966e27c8c102ffca41614b60cfa7036ea983fa4997b42de1d9d62a114a93358e69ca4adb35d40f36229c9453983cf2c68c23bd0ca979a13e260d0e3936ec65004b28451d3eb88626458b2ac2fce35b9344868830101ed0af5a6a7f719d50f2ed26ad76d50842c18d36dc27208093b51765d195e05577dfa236cc959a53a475f76a8449c19a2f66a4a4cd362ec8be0c296159d92369ad2f4509e017f3496f4acc784dbe15b5008e65d31ed94e857d77a3f1ddb8da5502e5735cb4466597be7133305aa50541d0ccfbdccda6ded9facdf0f75d64f97962845161c917155857b1b064b61afce5a18d28a8832a501126b14087798f943a8c06b0a3e79e1b996ed98971b5abefd551cb153b53d70de34d8083188e6da240f2a3d784e50aba8e76f6d7fe0f77068a8d9fd294ae822a990f96258f7d9ded555353ca06e4f441937a3db8c92541b7ab34d5abe8295c5d5e0d46861e5448cb9d284c2f6f2e0ab5b5460cb6be8a245a1c44aa5258c8d09ce0c622616607f07a5b92f675e4c48018537f4c9838c54334fce7793bec83f7d443c8a6a815f2871e9fb858e5aefdc3241ba259ea3d49a28fd11905d55245a8209a2d8ba237d1ff5aac51bea1b23b81a5fba9fd0164a9c055c9db857dc7310267647571339d45f9390dc12844ce565b2e64fb5baa95c46f0c8c007e0f5c45ca3cf0770f7b00f34418f48965fa73be4a6b1f0001baa692a4d4b28d0e9e26e5accca6d70d5f032980a67498ce1a6dea65959b2b69a2337de8beb3e8ff9526e689f735d8867a8aeb940c594d763ed13d070762f09b7395db2dcd513445bba3ba38944f512e73cb059d869d0071c31ff7463af567fd5f43a014a0cdece199139301261f0474a6b22804dec06cc10cc699cab1e8ffb18fe4c0cfdd3a8500e8745e7281b7e63c74b476a57419206c910fc91946d0adc082af163970ec9e0c73c26934866274f5030f19759b5db450ab8fbb27bcabc5aa49b7ce6a5092c4111b996791dca50d65b065213194747d7c31b569455ef099c84f7c788a68a929f84d62dd8718193f7441fbfb826bf43a8b77d63e69ada9b07818e389b03401997c6dc8251984056611ccaf74d732e7cf684f97035941c962cd06aa1fc0c05c8093aae9347f1aa01d2e624751124c575b2225b6c4a17c3603dd8dab7a50296848f33b0d5a8ee8d8f78ed1aa1b34e55d205eeeed4f4e24b6038bffd2d5d970ca2934b8c9e01298c5601300a23ed577c4be46a2ed43d4cadc7711269a31dd84c2469a21456ea9bfa877c24558e55636bca046630af20ecf9e7787c44a44dd95be1e085da6ad940048be1bf5a9b6acf9bcee2d1b37cf2223e6a12f80a2b729839d69025eb1ed5f176b3e1243cc17dab2b27901fcd74df6fe1465a6045298e119edc4f4760cff557dd2ba096e84995dfbcb814f6dfe6897ece60a6ddfd2e4a418493768e5346ac26291734335a9afc7fc1dcf659c1864158b42a96266a6629fec9ea1389900d80a9c294829f93d761a5288258cf5ae128c086e64b615b92e794748ace6013573b8d8a2640b654a463f51fb9fb854dcbae3a3a4eb6755451c5e1b9c1fd562126d32c7f370d2a431d7758965ca434644950f11bd938d3b4a4a34d0675c275df74819c4b918f1bce8655b48ae78b1e8463de36c2d2946e2ca799079578e7fc779a8ef423e1687d9272386f96126f7d5f50e173d86ab388d80f73aa7b83bc9c71dd2c031d664408cf934e4adb6053f7f6082f2f6969124705850d0aea7b890c1aac1215c85574f8018866f6db931ba05bd577fde77fdf56aea94df2e00db28a95b6275354e2ed7e7a634572744b8d9e49b5b942623bf2c51cd9e46f910532ede7fdcd5c13335caf199c4143a052f500ff18424c54de784e249d5bc719cc503af1bcc7733944478b0d77913ef9cfdaea58ca0390fc80c83c9a683e9e67e521495f73eb76450ef147c81c985baede25d9533f6f0a3a4a01005dbf6786b49958fe08bd1aa62e1e8566cecc80f598df65278932178ca8359931956fa9226b049bce26a9070c2ea0481e241ae12a31af29246ae298d7bbcc6b16c13e08e2cbaf1145407e579c9e1864096624d635e99d92b37a79bcb3ce5a8d44ddf605f3501c15b707dd568537a1d8074066edcd6e3625ab66b32ddc66246a69f7fd7ad1be1053c2a0e46a8667ba17d17400d0a639bd86d0b17aa04d223f338750911875544c5a04a7ca1d17b850ddfaeae2d31340a71d26832c1a06e6fa06ab75f494de38928673339f1ebf9d6dc9474aec735b3b7abbbb19604365ae3d8b9bd4367284ac049d533509b4c1b180698444e24fb62c210bc65db5baa39c46aee764b06a986b43b8c5ba856738f383425a480fb4954ba217df2d228558f50528d0aca89f3196dae46cbc4b0c00c80826a04856f0cf34fe2c85022e92cd17ba6c60f210ba466fbc41df10232f3ca4f3fa68d8424165779aafb55b4f4d08de232f02846dbca017f995291d66c0a134ab9726f64922ad2d0e22beb38c91c4c76522dae73ab527340f5a528e8a84f64d240bed0c1a3d0bbe21187e86738bebefb859f6e76bcd0f8d603356106f82f6590a3cbeb224420aaa2d5275b5ba8d93392d63;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h60ec1c5c7f46213005c3cddaab5483bcede0caa609822d4c6340b950b74c80ca2f4303e8e621c9f8e2bf033144fa828792a77dc3e67bb4e2b03bc360b90779230521cc9a6e4786a83fc480e7867eff01c12f15ede2394f83676e39ab331cd079d0a52d58efd75cb006252c24936620158661f5d167d082465bc2a62437c43b947b0e654d2bb84ab2d3097db648b68d1566a9f3f6bdd191c5982c8bde5b6df9662b6750bff3feb986a20dc10629f933713a7f273de81d8ab3509a26d511e8e6926b95c3c4f73da49e1ca51806fd40cf037cab9a9ad29649b3dd77299f9325286abf2a2c996a3573ff079ecb14595e920f1bf1014bafa3f2bdea3ef320dff24bea8f64c47aaba505f2fc823c1533a29aa73c5618d1de03aed21ee420e490e65ac85991c94eca953274c732d9a33e01bd9369d6368a9d38e7dbbb9e58d18d0c91e87ee181b79bb087dac8a0bf8ffd2bf134a087421290b3bb04cbea42db65ae453869858e18cefd1b32b62f2b318f6310c2d0cfc7740c9a89c6187af89985e531c4e9b120ab97897260a732fcb59d978709954fc793d34abc820f33000c7748b29536004b923be7c10d9af633f9c55354c01ba9aebce45e2f857d6dcc9bc8d4ce6f4dd46d1158f059a84ed585d9e0acd7076e8453323eecb9be802c8fbcf312630d06f9821ae1bfc21ea8a19e6668ddd32287308492c0646e954a6b65450a513b4f7701078f5691bf08936fed5f3531a1e3c97acf7363a80d2264e8399b71be68b2b0ee17fd4a4b2a453b6a33e303983aea0d489f260ca1e272f1f6bdcc3d21cbee5e034ed1610bb7c909a2c60fa79aed1e08a87845a6b418a06ca08c0123bfa8fa01d522b1e1e1555ec77aacc77be5e83eeb2f8d76cd987a3cf72c903f40333e5da8e5599eeed7e6150bee794cab1a742edc3d3fa23adcbddde077a3d5864d558e73f791509aa7efefd6e5ebabdbc17da90048a1c1562dab4189f62a522c546c7f143ca71cf153d7f109c9ae848838a7e307fbff8f74a3c3e9b905bdd8a32f57dfa4438e3541166790dd7a8f9a41ad461523fd7721e00c6a39a36f9a5019f5ae3ad205c7ba42aa347b83a601aaabd03c5944e9a2cf610315f0d8d77c10763980a79eb4c36a1c1365e697fd61f9dd317cb7bbf78f15ce50094f8fc0eb73174620989547268207197bbfdab2f194e11e46159abb3bc8a304b6582aa98e593aba169814a727c21437193c7fa8a2f097368f736a7b4f0e72f75d5d5ce2bf47a9cf9b7e07521a1d3efa97d6207d84f4a35a3a9fb2deac1a34d5fc3816a3ac54f890c0ab69fa0660958be65b90ebda4b09c8ba5ea4dd03c15f9345d0be7a89c8e54251ab979131482a15f33e783bf2f30763112e89e0a85ccd0508a6aef6875293c6ecc53b0866b63029ac433f1f4408a93b92937d4e45697be7b3d96c8d61e0a16ddb426c53acb9b2ac12a6ef0c3127e835b707e7dfeee365dc8c04db0dd4c4789483dd087c3c3663fa27decd40453c7e9100c4cb1800ca79570b151c5199ca919bab92f746866b1d80af3a8be339b628e783c25bdb7a199f3ab523c901d580115467b810779f4f3a26a92c2db672b7a426d76dc418c3785be743e87fe1d278a394e57024a429c5fb67916dc15b355f0b18ac61189f9a8571430df493fc5f0d352d786976897c5967b949e482baf8d5d2c3e5f74806ab49e60a7cd742497ad0b8a1b0113b6766aed3cedc9184f35668aa10469f065d47919cfa524186cdc7eebfc87d5eb4a575d943a1d157f23487ce512b69c13ccd614a0cd6a52e41a3dc8866052eb8cbb23d1667f22c21c562f4211453cf773159bdce0fc122ad6e2f7abb66a573a961c909b2579a1a87d4bdb77b6f310ebfe5e013f25c954765604caa3ca431e5f4fdc11d26618e3d0a345a631ed0bae93f3d15535b598ccba65e11666f033707f17c4e693e2193c45031bc3c2cdea882c047dc74f82cae5ad1bcab9281b59de21a1ea7f6468f4dcc4bd081dce9fa4f276f9b644551ea94fcb23ba5e4c3c87bef6a33d4baad1d5bf6eee7d008f295072e1201d409e44d7621a51671ea25905d397af7e188f200fef9b2f231461bbdb9c4334180c5c6d23b35a1f2d91d5dab3900fe6e187ce79d2d726875fc0f0476cc730adee875f8c0b16aab556011916db96059c5793211af63d08d7e6aed6793e1847e9f2469eca0a33ce297ad8164c02dbb2c5695d02c25186ee9060754e2aff4762ba5d00c5a647823642c2354279135f60a96566ddb61b3c8ac016bdb821f42639fd5c7d702e205a4f5c36f68d5569947e469f45c6ab521e901e32c07989add109e1158c4f9b4368c5e361b3e3d6c2eb49b2b1a5695d8eba87014d441809741d64bc92f007b2bda2d54710901b0fded9ec36c10a77558ed5ef9747f8a97f20c42c366cdc43dc55619f887ff7938a7b60da97d4e9da290a041f1c53053d82124c685d69dae9ae8935de1029026d42e2d4dc919d5b615d28e6bbe7515ffb99bb5e441e0c8c36afa854d5dba68f9d6d156c6c0f468968fd7fbbaa8e48eddafdf27972552ecf0ee46828495f17bcc11b9d62ef555d86375f88c675a0d5373afed162c5c0ca60d7e89fd559654f17291588a86ef2bf3b7e5bb1d07339072d68a6cfb07ce2201d71de19c08397b35352c553bdc4abc1784d0a4405d884d4ef7b69a6288c52a805e12aebf797ac87557673717f0a51dde144885dd9fcbb2a10c63f405b13927e5a9bfae91832570505274f0ce3856963f8fbf4127e179640204ca9d761b8d55e8695c911345a671724efc5273e5c7fb2d8a7e30851b6d8db89080eef0f6b11a6a804be448f21ca17227d0650885a189696e05137ed07a0ff0d8d5e8b38de9f29d00feccf41f6a5875899a7007bdfad6e1c279c5173fea6edb8c7e99fd8d488c162cf4efd41dee34e122337c28ec907fdce3f15f719e6715110c1d19fac85276b51ce938745974f179d1b43605004f4db917ae3f581bc35ec50dee06f85bb1e67500e588fca98f55bd45b9eefe9bc6a41129f058e7e221458eb9a9da2dc38583aaf8b0dfb181e35a6aa1d309f7e6685dc13c27583c206e120df077537f3585a2dee1a8970598e4b88f22ac1801ae3d329e39657f50811651476960f685603fb2a02a22b272dccc201bccab60213f476b82ca9dada9c46fe6b1fccb0a9e8aec2e1db72ffac44e3e3c9d8d3a7cc897e9dbc146e31887d4e2ddd8f0d1fa03c3741bd56aa8fa03fa8d809f5517344ad003bff53a40a47633ff9d9de3040a6183c05bd6727e66dae93915d3e625cc10ad67fcca35fa12b7da09ede2273713c012a6f0ad1a132194eafccd6dbc4e9086d1169296470cf87523091cee358c77ac8ab75789000467ddee0e6780fe8c75ab497c25b67e7eaac2c1e957ada2314fba85d419a4002daddd34451af600632f59934c6fe61572d47eb57b8791a60c57ebf6fec181b408735f870b45c2e936f7dbbe05937c28a0425b691180d354af7b3a8e756e95c320e6dbacc44a0c3d36308169ee855915ce597d2d835c99649ec624feaa5b35213b666ae5e8f012f255f6802e9bfebb0823bb66578d6efa1b60f23a4e2d15d5e6d52888768819c76a4f38d1947c9296939ff437256e03477620634232e7c7faf60cc3f4ea9cc1248cb8b5e6a532d16fd637f1fe57f7a33c5f504a2c0caadbacf554d855722607c31a60774370d887c747e0bdda77ea793b3ca261e93421a4f0d39e49ca258b3ddb6d55245de289a79ed59f0a11ba0ecba52c4bf8af2087b85f5199064e7e5348254345ddba4cda8e10116a4539c8ca784422b6bce0591006a78da038419f5fac795bff45ef5894ef4705c9c4a5ec6c06324a3c723ec9d88de3e90a48bf260a63ec71c58ab8b0a674c943400a0236a2caa2b340706358464fe9cba82c0c362ceb249e4f50db827e387c07bf45bc12890c5162b6f6dd9a3b2c6adb4c66a57580b775dd239a83d2889effd95ef42e77299c2ed44d8e7049232e755c2dc8e9cb062551d77490d86640248317dbf4035dc348fb17cae668a8f4af0b3b77f21ff0337eac17b10b8503284c9bc593e0c3f0f9cf9a8acc8b62904b18b0c69e9e717ccd2deba1ce61453c019865966485d2abfd7e02e8649ead27e4c60a980a8888856344e8048df4cae9cb1563cbde89c9ff3367bd6761550bc20f05fecabdef2b9cdfc49107a2c2d897ab5a7a31f0e56b42b37f312f222db87ca9db318b0afbdfcd790604d237950e112598bb94665560197e33fc80f56bae8359c62e85b8024c58b28356f0635a95051d0b5c225bc60b0c92bae0d7405d50ef75ee94c30576cbb6d9c0629e69ddfe3874b4fa70e53cccae31cad60801bdbc545025f7aeb6cf45bdc5bca92177834d223a71362204453a676141c29d7fce27209dfca5599185fdce2e2bbb1bb6a2892fe0d09071bc17d5411c01dd173853d8faf1e834b4cbf89e46fa031d5ba9483e2a6b7f70cc1fc04390417682474cff2d2b715b7418c648b2abe122fea0493af5da0500cda20d8abac12b068eba76cd73d8bbeaedd996c6bb2d1de2631805696130c1b7e7390dc11a1068613ff15787a9cb765ce4e26afd1b445676353669642fdbd92a9e46e4542c79c9732cd175ac84c6bb8b70634d89f64432061c35c56ea32d276f626e138bbcd0b923677533db9b953fdfe40e3f195c65710864d4a3840d20bc87cec0e9c7af0911fea9ce7cd13ca28672ed5b5aaab614626d2124dcd7d7367b065726c64aaa0e75098a0b079358884e4e7855675f9af035a34682d3cb1be58c28944b5f3f1785eb8486843efcdd966dcc01371ce9afda6146937dcdc0adc6361851f6c8d861bd282d40d6c0a241e7e62e397c5540c9adf79e0a99ca7288541abf4e411e29d990b1aba9ac569aa6806871370e2944ff5250bb0345f0200d2dd0274ef836964e0da7f9ecc5261cd91382383e8a2233cc1c1ed2db4112000c6629f659ca81ecdb9e7d9632aaca5d5423a43b87d0f565868c0fb4987c5188985e554791f67ac0ac95b65a252e1a724549be26f258c430ab8d8fae2c493e8ecafd5d02893526e6f0ba2fdf1aab3b666c9290f85652e3ebe9de2365cecbe85a6e5c34ee9c97cdfa0c9c18d0e3f76cdf09f25afc7daa3e10732942e30255fbd63d79b8afe4c960f98b09553e48c75868a19f4b7f4966174e005d8039d20d03f8b65190b506c5dd7c7c70a9d13b078626c681aed411c43d2c84240e438f7a2fe412257573cec755c38c4ab94ce223233b5a5aba432cf0dd44d4f4bf4dff853238dccc59bdc67dbb7ae52f327066288e6e2967528b777045289ffea4e28df6397a5980c5fb2f054fbf15e4ef35560b9e4c20014266242bb7508919c637e7f109af658af74f0d080658aef2a245ac0bc42c06510a8be39b820137f30a00796bb22f43c6ea2240190184fa1fb1c3a1e5e316888e3bec1ad1b923416601b9e6d7dda7b004cc9886ece001e2c1f79221febdd4e43c97;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h9e3f0db35408c7aca1c6d887faf520c22b4365a14a2d8ef1f478c03634b116e89b4c84bb9f841b95c0ab7b8f0661a4ec643ff96b0a29c61338bb73fa75b05af1bffd036d2f6e9c5704b5e038871ec9287fff12f63839a311ae066fa52816da5bf310afb2d7e327cd8105e8fa6347f18a596c9f435c194c422a0cced09a0a7410bd97324ed3ce3e28b3ca728a75cd65ba5f55839ba226990ce2a55c2674dfbe9e249bd6bdbcefd6c55f8c894aeaa048e563905297723be12b3cb488cf8fa525e671da7dd72def6e43e896e1bacf1ae3f645c3eeb1642f722f620336aa9d3d8c4059d13f6d4b5bdf4b9818220d601499f9f2c446ce110c3ceba7cbad01bfdc0a997d235e65f37271cefe48f01adb5fe9f17301dda5c4161d633bb94ba7a975157d0e044e6f8fcd1b8632f2969da47b61468152bb67c5d1e71d7ee179013c747278547ddb7da02c8d0d26c7f32895d4248166a0be26492a29816c841c25cb8dc9c689cc4eee0a13185fc5c16df0ecf0b7c4be034a59068403d00149f9bc24caeb8a6522c31994bc842c82ce07c5d8ba04c666db6fa0f026eb72c0725f583ed389c911b8738b068106017c415382b410db0f20ef8320980ef411f7b2ab9991418a005ba4474c43313ebfd6cd0d8d96ef8a40444c81fe45ddcde6a4a7eb978444f58509d349d781b94debfdaf07a8a1c9f11ef739b4c1696d6fe387695567cfa8af11c2e718adeec403da572abf18b1d34cefa7266f7cea7f8f159ea34e90970c2d21749559221ab556e1a86ec4bb6a4d6625f707ccf05eae6d24a67bf5a36ec39d89852ac30bff8cbec681b83563df52b457f744a2f9cb5f2adf90f40b39143642478540751de042db6acfafbfc9cefb4332d0ce6aa0d24097ebab789071839cc68995f3180870b8e0e4ec41cc7e59b0a59a9ff47a97fc06e5f28d5b3bcdecd8d4b1ffa5f8c38443eddc7e8b82872d78adc871ef84ee4d47c8d9c5a7517c2d2f39a0eb758e0814b0c0f8be6607dfbf5bb9520ec2755a7f5ec7ca7c0c2cb667873e73a7dd505cc301430a8e08c0bc46a2d370211b4331ab57f8d962802383fec0c5b8bb9116354de48fa76b6ebd05caaa79b1b439eab41b84dbcbecf1835f7dd619df9ef04f5bb695aec6ead831463ce27246c286c259e21540affd156399a6d113f1f509e464f2f037329175dcb113a273d0b45bfb25f93a9b57c4f476e0ab4974a32e0edb1bc6c100548a2c1f0e42e216dd39bc52fb7fe142c8eb816fb79f47b5cd4bb394a8471ecd8b496200095993ace752327c1869b891b3dc4e7f2e7983cbb93714f62f30bc0c14d3db95bc2f999556fa3f8429173c125748d846acc83adffa2f7d35d8c5d98cb223fafcddf2ae1e066f55a30e4ccc4a779ad864c7ef2332b02f92b7fa7a9bbb90f00db3d20d991fcf562cca00e26ef6604ba3fe994e51572fb93d54878c8b99a31dddca7d7650a67d4c05b0f08ede1f7ee62ed006befab6ad9654b39b1c17839e75d2d089936e7e1bbc36adde651c290525f09f95708b925039bfe9e955cd32e737f14b98b9603ad2ed7d6ab9cf909b9fe719675dadcce7fee3b9e09ff37dd3938d25ab2905e0a62932eeca7fb150f0d8c0fcb3925018b7391eb888fa7f78ebcafd754e725f2ea4cbc53e2caf01f7a181dbd2c84b37b0370dbd09354f330e0adaae42fa825d8a55b111dbe08a4fe0070b9d842a664bcfad52bbb09131bf66770cd074ef4d52506d09889b0c9b70dfb2e66b7f157a6f29dbc5b638b77d4b34153befde8ed72f1a2c8c4d713930d39645bd73f0f92f3458842520b27f6220e93b953f07c721812d59556ac455871202c901adc302cab9926b5c537e53b85bf98295a2f9cd36e4ef6907ff535c0362c68e78457ed23ea9e728b37dccbd1cc4173742208142af463a2f559fccca8b1250ff783e93d4b028ed621778643d372a2b77724a8e3a05e16deb5f466049861d045f51fd806755c75286ae7aaa7c64922cba2cac52c4b859d67a49da69a74c8b7da7f8ebcd24f8dc47592187222083d9b3cf922597ac13c46fb7000a3beef5d50d76cd28fe3a77061e5477e3675e0e8eb34d2589a996bea93ccd4e84d9bd095705af10c98596a45964f9d1b4a9cf1ac74d8ac3158bb7a6f0beb0ba8b8f9911b66311dfe960924c89174a1487ff783a6a7c48e0e2984f3852affd384ef8d1c88f825653a9e6cc47a84145a0dea59820fd956a87c217a14a3ea913543be44c1097e7cffe83e80293ebcfe9c16d85d274034aa849672e0af15d244e7cbc896c0c4109b87b54d2667e0c902ecf28a68e04fea2ecd4099e9e46f864cef472b8b52bd1a3bb55039e7cea30b3c4fccfeb1a3e42ad4057ea9106ae657cf057ab91b28e5ddb3ea00ab79ad101012098f6c768b618cafc0c728942e217c9cb459d5b725d6019bb03c9c53ff3d0633e07bd677974b473156c0ab4cf16e56a691944f6ce9884c959e6fb6fc17276ed15a406b520e5c9c0627f43b12e2c6ab86d676ef0f1d3705999edc39b98b1951ab09db5818180314d69983662b95b6c9606419b3d81e98fe65fe347599051f3ac13731f1b22d21788aebfbe32594af195515d2956901f28044818b0be12db969dceb5e72c712e834768c0361ccf344339d889b6123eda9d980991f43f75922fac0ed13aea2dee42310ae112005b881a864a383af1de162b63af66aebbfc66e16979830ae50d12bafbc814cd13a3477e54b9417b5304f1528f7f349f60cfe22e715259ca16fa0ad489fbbf3fbc68c28e162deef9a1d4c8dc0403fab701c6a7bff6ed9388b976e034d78e49acfdcb2cb30622efe2acffee5ee95e538b76484ce6b6bb75e8a8b0e2736e3a82a6fa6103c8127de3a4f80154f2070410c8f07039867991c4a33b61de49941363a2f393cdb55b5bd925f15af829363ca0ab10020bce5c56a3230d8599a6828c218c7739255543ec9a0f3f2a72d09581b00d90e488376598e1eb7cf1c3fce825c8f221fe16e446e59f7da3a2b3264a75d06e95f5ee77d2679bc8efb1121aee4df94f1d74c2f3e111d354ea937e0b8d2a71286f04f8847a850885e8b2bad8923e9bf6ac639766841737b2c9dca5c43aad42a44a53e75c26048748836a2b074f4be658f2d8dce5b581684079d9d7535137f1924bff2b6945661fbeb76bd7f8707bcbdbea7bb2339aa50bdc50bb23687f2b7781f6845714a4e87bde068da847ba901b578ba86ad43669a449542aef7701cd7bdb3425452a604a40c2a465e72ff26cfa77c1198491697f5512d341c497001c99548e84e00168dd850b01bfbc9934b982ce0b9e3d6dae9ed00fde375ac47783a35d462aa52d2d10d380b3d0b3b594bbb0a6b8c50d7bb5d88428c81cd7f6bbe8ddc11cefb32e1740a09b93e1c4adcb80313f498e719e49685ad76eb8a7948731a412a149345c4afa4919531d36afa7078c45842bde07bf1711fc53c0397dd97e954cc18b246616b5c1e59ba53a3fefe2fbdcf1b74c860082b19e17b28b77b61dab066b5c5ff1f6e50148232f46dde2581af14621e79d1a0b27ef8e9de642ca7a9bad1c1651116cadf617fe9043893a5309f1a2068050cf9f185769f0f139be676c1f0fe982d786998df3418b5924c390bdd87d0a128bd31204c9551848b3357ee5a2fad7b83de439fbb108761228e0378ee7eb9ba3a1e16200c6f9c38362ca3d0eff5ca1c19c791ba8ecfdc166f087c9418bb2794965296ac55b2191d0c26e60bb832c1d5bb3a7764a05d85732fdfcf384f335e4b371735459c763e59b9bd89e0197ccc53e70155e5494dd65bc91df528c86a814fc9f2df070b761db71a49ccbe82c23d4edc05cddaaeb69b467d21acd9c0d9b97cb99c1eddb97c7b2009cf0dfddec266aad523f10c17941769adf2cea11ca962181baed11a1fc6a0af48c22bdb8674d75b5fa7dd8e807d201d382e5650868b2889409f7db58af55f98f1d53aaa48268dcf6ff81d9283f8ca885f300e575b45669a750d113295e399cc7c58f489859ed8a79376dc26ab42f747cbe59550c025a43e8715ced85e106a22ac7082541dcdcbb8cc72cc672f8e7636fdf7d1238b2f10a11c2c10fd659bea6408d0fcc248ecee5697d5231cc31bbc5bf964f492d5c8924c351e6e6e370ad84d637522c89884abbbf7c6988d28afcaca5f1b36bca111c4d8f33be8443bbe618b7f8570098acc75a7f369654f4fb0cfcc54c99828f3dab6cf5d3c2813a319223bc638954d2f18cfbf0944205423ece5def92490b7804ce5d2a793dfe706d397adf3ee16e3e51866e79b5cac86e3f3bcfbee79dfa8664b689e6d3f77565d2d4d4088f7cf6b4f642c96d2a69c0182aefa887b7faa2579be920652ca08a687dffe23c78489f1735faae6af53f1ce05651a49e04ff41f47bc306f42b04de60c0df7d41eec9ba1691d786a12b5dcb08a064e5746f4a8662116f2fd670e7e18a341ce6d65bf93c19d2a1b91f2ddc6cd14822ee4a0acd7dc79cfeefe16cd8d551637f54d72e145a8eb98afdcc484de1cdb2eae06d4b805b2137940e7d55eaeb63eca0ca6c00d941bfd5d2321eee3b211c1f488267372da4f07e8d4b2e3fc2119535c383d426edff22b8e72a2b5b25dc40e10781251b20dac1611a5693816037bf61dcd11ddb0f5b4bbc557ed5634cb54f23ff4c26c151e89d75a784943520dc8b2599a45e88587a6deb539c125ddb14803d2f07020154b03d181b4f3ba20074c411529cf2e9d03cf2fe1f4ee93b51a95508994c0717ff3c3cc1e1e53c3777a670f23d7e1d542195131dc39ada5017bb64021e6f61e847a69092ec638ebb0d11f946b83d1920ac2eeedc5d58100efa0f264281a570a0c747b3784d9e9d64a8ca404a41946686b790bcd730526711bf19d1ed113e7bf041d1a82c32de5c801ffbcf014aa47871a20d730a5d6f40b9ad4772af58d8e821f774a6152d3b9a6abd0f2a506bbf9d7406e18cb01a8c4aa191004e84277178c168e5674dae64cd2bcf0e9204e7d8866534fe439eafa3d96f9efa104e3e46ca84e55b2fbb7ca587f359fc8952fcac868cc09816f8854aff72dfaff1a348397c45b80674bc2e4320658db62f649f245ffd2306db90726d443fdf30d0f96a9809e1ec2995e5292bf4dcd77b29e72b73d44c478f7c8cebaa91723206093d9f104c8f032c43feb740307232440f201d395a9eb318ea5e4146395b662066ddcec0232d2e8242046fc25276cf471341a57684b2448a544bbfd8854fd2b46d43ca92ea7a41718efc77b181535de56353f3063aedf0a386db5849eadd4bf1db5d2755136c76e14205764321c7456c06bb04c2ca2e9fc05231ac2a76d3edd7565da9281a7caaa75f596ff98e576294a170c6b737139f83e2e7720754708ffbc68dda890f57f5f8b949c34d6a1b9910ed934c79a8e7b60486caa01c96e050963eceed17545616ca5bb47d60e78986fb01eb2d7157c88fdec4205aba7ea21866bffe8fc418196d5f5c89411a70becd9e3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hb565d6f23e061def550417b48a4e3b77bb06bbe46e7b4ab083e109bc15fd869f2e9a39372eb804d4bbef316d0e9923404f95c75896b2d230c07120e628d47211490842a67e1256cb3fbc820c71b0890cdf222f603dac818f838ba78c71cbf67622af328f739da4c454e42bd5abb6d634779e5462962f8cf9d5645a245f49d0f046b7bc08c7a1dc04e7137654c5e3c128e624001eec63245d8def06736cb5f82cb9e538086aff3f60e9da190a4efaf2f53f152881877714e815a47f19ad376969360353c772dfe5a4c7ae7a5d0f883dc806c031bc6243ae3ec88a576032c39b732fb34a6fa3ba0be4b73f8a3f5177094ab4dea12cdef3e76b274645592bef88eb1221d269c4eccf4306ec143ae4157578affb0fcfdd492a3d1296372bff4fdd27fdece852e3b0549f07e71155e48c90be9d07f08e5f8e0e292624519661a14f8e481ebf071d9e2d6f83c4857964af4ca2f9261be32821ec9a6c973e969622df52c02801065aa5a4871aabd188b008cdaed3481116a223991978e2494dd89a749f33e68ab5c57c514d0a52aa6b0c2ff1560113f00dabbfe3acf7009bc38b61b5eab76cc94bc7fffe08b8291d0fc7e4ec91102b39e7838667ed4795ba40ea654c0c97f8e48d87910871918d4251f3b93f2bb7a6e1561107da66d2fdd9facead7c659b4941c19dd91eb2f97512ecf794393f17d2de9f06c5e40d92e09668adebdd2015a445af0eb36c88acbe024d589f2735fbf27727f6c722512da765511c94cb52c9491dd21cd69be685e695abe34537447f1c7d7827762ea3f5f0f5d0e37c5660c7dfffc6a341f42a946ce575999b459190c61752cac1c52759a0abcc30076ced82c95d21d3195017bbe630de12142023dd6a7dec63522e1d218a74d1ac6986a48ad105f9092135e7e800b1d09240573956c2ae7ceb6bd48509879ffa5149b57d34f0379fb7ade628b48644b1927a580761ac0d81b8c8b77a5df7080936987f3e136c631c22beb1960d1d507684f741acc4f1a34a5dabc923f272be173af6e60404c6efd6cb9ef7b3e235e352ef0eeef8c0d414443ce127962693a08eb9a0cc46ef646decdf35c336a4ac13e1b4811c40ab1173d886d793473b5be221c2f3984f7d8a969656472f2832da439171a1e9da3ee090c787886ee525241d611a0b8047dcf9113917fd0956ec371cc0df4f2d8baabce9e37e4342b682429231d81ee96df97eef12018a85677d85bfae1ed8b6a59fb0be7b0c5838fee776ce1b87cfffb9cf18085b6bc05f0ee45942b3ca5945a123153d85a5f6bb90af0a501e71779f836dc2d02428b95684ca161729c7c47c71cd1bb86c66b7636b79358da73a1016e5d0f311470c152be69c9f408deca3fe023c1a7b3a44087c01847587f5b1072abe69015861e6f4c15c65f5d2359e92717767a2a0b782ce3350dc455ce6e92edc44d39e18eb750408859a7e2a9ee59da23f7ac67e2a116644a77911baa6431eeec7daa667625b65f325b6490e9d4f26ebc545e7df3036e26867ee0fe160c797689654e4ebd40e22b538958d82baf9376dcfaea906309493bf35d3e7dc4caeea3f7910dcad6176fd144305e75d10fc54ed668ba5071f941b4ee392d8d50dea96255b96886511759864b00b84eeea8eaec9b3d939d51249a7cccaf2da6e124848cf0d85bd8c53bfce1c8ff46e254f3e77a2a30bda6a625562b8fd2ffd69511051d9f9fa9d93d508ff95f874ccc64e568f430cf0accac682bcce602c9cef2c72e542001ce3aed9c43751e9851b9836e77f3ca439538883ce8b8711a98b4209960b4e57c7baeae509c6b0826994a06673140e0298502c52722738875ca79b2395d31b10305af663b9119d598b2f0911f76d2892557a528830eb8a7cac58815dc7536f793fdd3b0fe0bec1120a1a21911d037b86f46656b3aab8e91b4d0125e7e93866bbbabf0d4966334d78f0e8b036c4a14da78fda04966f301d26534060d99bf3b0ce1f65184f663d25ad26e23c1425cd56b96136756cc6d62ce0a6b0008cde8be83e8d9b55dfee642419ac3541a0370548e52336b789a500f6645e14469243521282deb7e6c621fe02177538597711306536c7451b33b2595bd7a1d07a146226be3c27614e6f48a39fc1ccdf7f2a7f61ae59423b54a0f5b472295397d9d313364d4c0f3a3a0209dc75eed38f3fee99ed61d6d195661c3efbc3fb27d37a32976a5d77de26afb92ed97ebfaa78170a0db498e31096ffeb6d44322ed9860095c5ea59aa7abfd757f782b246936e28ea0b125304c032605e4e769e65cf6624713001046ee9890ba0e3b1067f8434d3be80e1ebf3bca5d64107a2abecb444b6834cd9700e59cdfc33818ebb58c8e379f77c419f6b90dee128fa30fc1eb60c92619b2f770664ebe936d5e3325d3302142adff26d528f6c7d4622b856b9060f67644cd2b6315d50857c61c4f9b11e490e553a29b4c91527a8d1faae11cd369a6a1f4a85b6bc2771f79e4608a807effc44907db0b645a7463a07aaee3835311171c22ba92ccffcaddf9579f528084117090131017a6f18d418bcbc54bad68fb5a6f888fa3249310487e69a7f0b3cca4d6c37b37916aaacb072f7446fbbba4f84c12928018512b512a18b9f3beed7b4bbfb4c3b2d4ff4c7614c23099f535e3eb1f6b8deaae321cc4fded8264ee329c56de1b0cf29f959f82469680f9a15c30c620e04b40a96450c249863bd1b3c2cd5eaad68aaa1000a6c8e400d64ad489f3d83b42b08146840cfcb73a4eb74ee179316e9c920a13b1af561fafdbef1eaf6e0127fe71fa18b0744920a8c536668728afe44faaf87862a03315a15b628f43aa41add22af83467d2adab7c4e73911f8b2f68963b2824e6c514f3025aa375f1a63a738963fafc2da1bb155d12e1a90934db2472c20cfe9e9541b4528c9b59b1088b0fe30e4fec16de5f79f6eaba40748bf805ada38a856095f884b28c8954af09d11435e22061f50ec77d4500de624a49ddf32b1ffa3bc861506df0e3928e5c3f6ae27d121e969611893b23cccf9df99571087d7eec2aef7248a36a4a048d660c0db4efd1d576bce0df66967b9f83aa7be7aa3b0bc193e1fc8d942d07b0e9288e65a72cdc1fe729eed0bf9680d5cd6f7e82081c3e52b2837872c863ff019d7783eac0f1364abe0f2018b1b3c68aea5c522c038ac62719210f1529339817eb9e44e5ae98cfee27b7e6cfc136f3f42bdd824a452294c0d8f78d023023799ea26eeec0e85ea29817caa653d5aad31f65cac08a449478f207219cb8e24bb5f40f58e7ad8ab16fad437b4ef531a16c286b05bb50494fec6ddee9a0182390bcaefbe951673fd9532e3ee1b9ea487b875ec62018197108f221e5ca48b123b222d4393017a75aacfb4faf234e0129287ac82535270dc1b9abd84891a9a8c854015883d773c01ca1275dddf72a4c389e9e01f39581c2cfed5b3ed0e045deeab6d98f311da77683dfb2518781b39beeafec36c08e84b5a4a74b007770dea90c476d70589c6ff66d473b431ac3410ab03655bf92ece46f4edcd8ecf16d7118a2985877d43101eff03a6a05847b5c41369a49a84bc01fbc233fb8af4001614f6a061e2d3b2149e2bf10439ea8cf579b6978b11fe462d36e6e2a92c2b8736828ff8a878a3892504000b98f83bf7722f95120e4b19a0cbdd0a508cd01be11283de33997c6cd3e8e20a6e56f44b4a7a90beae536ef06fe10af219d8c154cfe9ad275f46cff2210732f78620aac86c5bb3b40ad23551c0803261b05a84f26ed3ca8c1e815d194e4779cdac89961b1c1f2625a99bba0ecdde2eb2de81fb495fdebcd18b56bc844cdc07473c85da6882691d66f220a4dd201d448003ea0e51455e0b40218a30d63c890c9b2782284169f1a259514c3885bae41cf1009d71fea7b16c5ba8b013e2f79d418426b37b8479cf5bb51f30f614ad057a313b6b19be302b991ff7b6b8480ab102110233a17a971366b1c1e74fc525ed6215f981e3833ed506126ce31a865f0f4cdb5d713208976cf1542c2600a0d60a17c5557fc5423cf3adeb07dcad7f62531bd42e1330984da2b2dfcb0cfb983517f6b6128265ae4f222b0f3d3d8e2813b6f842cc523b18d7674c8ba2e16233b10a82de6df1a467cc8aa3715c27bffd71dc344f47040853487e81c77c1c7a7a35834eb1787b80942923cb9588e6533d56ad98c963b66b7bd674d952ab1cce93df017eedce8fd5ca76410e7fdd4a230a8435fee62946d52d60c1b09aa9ad25c1b18c4cab72dc3825e106b4a34508fcea64cb23defc50141f135c76852a1da2496eec2ef43438d497fee482c03e08cc5d769fe51d8dd9ef75ae4b5e868003b8268844ca83219d9e97de884b21520953babd7477a35698fe47b5340bba38106dc139a5ee801b93718dca9f1e54981e5be22a2dfacc23c6c8ff706d561e0c2b2ec5f609a91fa28a4976160d3c7008c2ad8f6847c80e53e73c65e4433d6d85d3ba0ac45cdf93292d5bb6d618f9094cb028f9f99a7114c817cffdbf630e1059c0b14fd8c1ec2d0f6added1b4bcd088447160806a1e87d67998d3641947b0e5e3af59085d21abbd16eff751b5c07b00d23138af141efc06a2112f68132cef6b0758d158bf56d4d8457685b392689813e8f38430b3590e8be9a75bfe15a19d58daf982357fa93cdd359531a1a326a2b0bd4f9e93d2b07d31d71f3a544e04da28398ab4b7316e0a9c1fba32154799a4500d88494176d0592a37dbb5bdd8c781f6020ffc0f961f2f0d7853ee2a1cf53e9f0561532d6b8ac1ccc89b87407f8975d032a908af9fd3ebbc9eab1dfb68b3eba773a34605a67cbd891118cb0827fc186cb83532b83d0a4d95fa64a9b41c5faa35b3bd579902afbd121f27398946e0ab0b09c115119e09ba90785c683434f5524bfca6897b3137a76c12703a4c09ef37280cf07f031b49889b92e0dfb7c5dbb5936c450f79f140b2067f2b483e96fd6e9217d48729876ff9eec40a21d84287846b7c099f6eeac10cb09b8dbb28a1eb8b4b39f7b85136bedc32f2f7b295a959b06292f5bfb12ef04f44d5166849dedd768671bb4455b515c6dfad6e9215ad41693cb71cc98d2b26c72833505446ff7a01ef913ba29e46506cbed2bc740c0ccc38ffac19cfa58e3a55604298994eaa42e9dc3442c93905a3aef0121e16767d7ae3709feea58459c2b8698390c81721e29fa67935206d4834e8da1eb03ab5cf21736689caea052cfda646e5d8a0466385eba043fcdf8a2966d21b070f63a8371867ba4238171fa96abb1193918d3beea7b8ba1b460f094381728422be235a4151f23939a7ec054d45049a0e4f115ba61cfbf26c5b74c0943f2c017093029dd57186dead25f4f6d94532d34140fcfdd62e3451b91188a44f8a8a11358d599437a542e54a937df64aece65bce8039a6f1d9f8cdbc2ecf5e6e465ebcc431770330484eeb4636eaa5ae73dbc7104798d78d84d8e9df5bc0daeb27d5df99b9c5f4dd1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h2e06b2d63cbe42ce314192a1afc6013833ac06c50413dffe0602d5d8ca776d57a63f4c8dd1dae6e4b4d1a1352d1c3aee70c2c189e287a4509015c78117f6cfdd18a0310efc1536e1e3e85f4c233c345aa3e7a997eeb0cf8ccebc4d13665621bd26565cf7343dbf76ca2eaa9e5cbfe127e65790325fd24e4397936ab2b24ae877e0074ed833a4c6403dcdd135b2b2722ac0edae9d55fe4486e600cc975c53ad3fbca5660761ba56f22be0016c35b8cffa6c51c013d23f0a4dc5501e553068fc48f0a9a2bade6422cf3a3ed2b38f147988bd7383ccb07a73ea825847f7c4650d924a8b57fbfb947e43cf044be152336e100e2e09fe904049fd5fc3e60647665c869a457da8ea61c6c7c0c7a2e1df7094764333ae4fc31c47295147b77c09c8bac9f03b8d137473821b5a184a06fe143410cc37e34e4414f7f31e3022a2d5d3d9d756d667d77742efd383479b45c0066b74a2405974d9094e1a3056821fa0ffe056b8edbdd551011c844ba018735205212d19ec0afa354831eb039026e5111f7f43fa00f52c5d9b3d15effa41a53219cd2e4e26eed885622241b0b75ba55528b0d07f598002af4dcdb9d94ad4f7b7e50d2047aca1bf1ecadeadc7051f16c798cf871e65187f27a1033695e7137b8b7e8b97cbd3fe330dbe83f013db8c35908931e5ba6c21ce405ae72520a0ca7a38f8cc25a3be4e9e1735208c7931249b1dee9b291e8a65295b5c2eb3bccd0220f33e162fc54f354f77292a802ae30ea1f589ce8ebc8e56bbdcc264dd7a469aac406f98df8a00fd1eb20e88ca7534047a9f2c91fa424db526a483c4690bf858d8a08d0d4916525e162076acfede1acd2f09287054228ec8f759649aba2443d6e1ea15a5e716a6979f80493a99f15f41bf07108a00694fa9f77b696be24939775b110e83a835d73f1de53070224f3580c5c7d5814f6996f516747fc38ff6c82dc2984793990a6bdaaebbf4279874a6beea3e7544bd23d6808381c3690e13f791ed99b8c17c297e9ab299ae3daf31f8e1bc17154ac1d6176eae863a1925e83701e7b761c4ea64460d9ec0cc6602dfc388645cb0f7343bf8497d6ee6863d2240049b14bd142355cbf8723f3e9875fe41ef9bdca4ca606d5292beaf7cd236e85f19a4f4b521e02ac8a93af23ade050d5013d4baaa459815d19e85ad711a5cd1cc0d6032d364433775a5112619d56c9fc589f7d0d2541a150c101f15413d829480ba716dc1e84cad68301d867878f3ac597b388af79f3358a124a579a5c7660562acc91ff2c05ebc157d6c3232d02b82051dfb7b5e724f17b77e1ee50e781577e05ec11fbd6f87c3a50ab7cd074b6e1ab9fe923fbc6d1b97c88a7db966b37bd601333339d07cf8caf9f8b46a8d1a4dd79827dea766952bf90e48ff48f934a2d371146880e294407cf9f31e3afea27a7f962ff446b4f4de2cc3e42414ae1b522e1b87f40c22a224aafb3efce8263c9602b6bff20bc9980bc1e43be7c0734da4fe0496f94aa15b414bb83b2605785974cdbe46098a9ee6aa07665607ae0589e26a943861dabecd2b6249fa1841262108750d90e63bb7820ffe5ddfb72df79c5e4ac6f448f470de987abfa38b932885c8c41006aa64064615fad5a01eac3929b6a45250b956c65f97bbdbaf115e8c1f4923cee6021a981c3d39b3a695b7c333fa8722f457a79d7d03bc33c89164048a701c6ae8a7b823daa1bb44d2c64381a0e5eca62a3b5b2ccab3f0fb76c78b4b9004056cd82b0427d8fbb8596e37b1eb99eff95fca4d63af67d25ec486397a45cbf1b275681d464b4d0e9aca07ebb589a017fe165b6d68d57025dfa1a3b737c3b393f8be1cbc9674b1f037bd7120a6f2f245fa857dfeef95c7be6870840216fd9c2f35344df85f886a8c0aade3e99a1e4b92daf436fe0ffcbd0a2214ce90ead48ee8dbfdffabbab6836927ccca0ccf21b88765e36ee839631b652c3a2af1fff0b4bdf93674037efd18a2c1cc7187c8b69a2051fd093465b4c202533c5bcbf030816b513180c7bdabf87429fd8370b8dbecfabce942314e3cc5ca4c2617913ff3be957961fc7bfa7db7c847f2af9cb4753b5909b05b8fe1567244b8a5967cc5cd76d111a040c07e596e838a265e281807259951225c756132128fff48ada0a62508b5e7fafef57f59a1d423517e37d6997745e64eb938754fc17920641d3b2845c65ac5ba7d6e72b58c73aed85a7f280183e4fa6780d6e75abf0a6c02f4ecdd851d643d6fc977c04a5e9a9905291afae292f836acde0bd5399f75249801e90a914fbdbb5f04efcb8e87a3b346dedcfc057c36e6e6f34bbb7832224a2fa97bfc223952721231b406969352b25c22f718d23aa6bdeb518c63c04e8d1c8ddafe8f58e8f56308ab215e275937e7dd06439dc75533fd2ccd6214597fe71c1c77f435d1048f91c562ed80e0c0f58104c3b2e352635cf566573aa6846792d28ff00129cb26cc4e61eedbb6ef1250509dcbf4f6c80a2bbc368d0bccca9b0fecbb82a0272e1c2c11c9e4e641bac6d37bc44bdad56f77282578b73970f71563745e338c985ea2833bf8acfda2357e879b8cee1fd7b849d36e4126d58597570b144e31250e478749801ae72010200ad4cd586d9394b70063bdde18a39f9cb49f6d0d332689ae8a12220b636b225cb816ab40e785d1765c682f7107a1bb603f48a56b1280f0c1c3738cbc835f3a4d3fc6cc36523597dead4e783bab7af66fd8a985608c6bfa756d971579be8444c4503cb4dda6fda39cb77bcccf5a632c081b5d4f0c6161f2c56f6ae9e0bc8d1d6aaf2c09561bf39afd5781fa896c389270592fc0366ba710771931c531d21ca51ffc497a5b83f2722ee15ca03df6789c7ba97b30ca1f4aebf78f81033e5f107127d17eb4be1565e116011b6e3a77eafd44171a79335af103772000c21d042aa5e7b6a638b6b4b69c21e6a86fcd7e992c1ca626f5edc7c0ad25ef2fb28199bbd0ccb9c87b524935bb8c485608f76ac137f310eccae6a8093fb1450772f00013cbc6d78b6f37b7a74fcb9e5f1a8da082252caf1c0806e8672cf2451a952f8d28cc0f287ab64cc6872f4a4a5a9ff9a121399d39c31a4ac8ebe233f531d60fb34053619b2096739450c12c12c592302999c2cf02def382fa999d80f1373ea204cfc364c30cee21f7c491f87cbd2094328a997d36378b60b714eacdf57f6ac0ff1dbdb4077fa6aeefa22ebbf122550ca221af1e1b465a4deac73aad2f0be273d472e8ca76e68a516d4e330be1b8eb0d26b6c39629b64cf9377c8346db12ac8c86aec9c4f20af6329e6a6a1092488206dce29bb9787bcd1c9430bd2d2e76cf6a030c5f600c3f37c06c72689285d8cddc8f0f9c05e8ec82eb861cf9782a23de586e511f31ce2cd665c827fceac1e67d4c377433b2666bd79a68f29f4f714c6a35ecfcc9ab035fa0dca79e75cf1a28156475464c10943527bc6a4f42874dc7f0c17784b83d0a91794283136c265ddb36269416064c775cfb1c3688ac435c9707fde7e3fbabd192560ea293a4539cab41400cb75a750ae2c916924453a457e6c1a87a0ddee9247d47346b466420b8c6662cf8b2c655860f7417626b04673d46096988fd290d4885a297457917f2934c69170d8dde2ad4336b618761b59abda7b9e5e4d362e0a31ee3e73e589323fe7ba52c5feb0492488c5c723ac8f0f435639c97c699678fc78822d2bdf09c1bcf35ce02ca217375ac70d5e662b76ade43fa126cf1bc43da5278fe87c21a067e1c62859cdf90579421f125dec34ffead47ee4aab250753fdadc40f7334e5b0d90fcc8fcc07300a4d5364453bbe67417db2dba345ee355ee86092d4614c1ca10bb80628e7c1cf8c8468e3e1feff617c3cd001131e9fa2e1d88148fd1c7cb622d90643b2f66d8a3a983d04077e4fe29eeffef5b357b50fa1f59a8fef5933707e1a92776a95faf50542a20540d727e463b999b8435fda341e28222c59aafe0c394a5ed640a2f631ccbd718234bbe7cf1b6309f56c01f37413338e622e301286d1f6939872ccd66a42d2298e0ba7ba3a6b533c3c83ed94b1e060a073101d50de313bbc3edbf14b8a3e7f86f43f2f41f54798db175208fb9a24d1a6391d4a87bac68e7648a439e2c53103ac347395d6cdd064719d0bffdc3a6b91cb43abe1f86e940e992f2acdb1982628480d7ee4f97971e893e309c1764c37b532af8ad947affb323feac34df1f8191dcf8c8cf1b8c437a6914efbfba5ccaceadbe10a13efd606fb51d7bee5b8eee63cfe984f1dae4d0c12bc3c87a01c35c9cd3448f5bb0197b6b97415dbfe80b05d72f3ceb1c3d2b04e14fe63641f1422a34357192c04b9394dd9cbec84df432174a45b07cb44a3c7ddab34086fa6cc2e0e1ce6ba74cc31119c659383cab5086cd2da5cdeea588ac79681b32401859eac573a40d23264d6ade18730dd88b7de7ae7b7ce81882270c73693b3ee7fa073021e66ffc78f96391d2d7a8e35983061c5ef2beeb2650f4cad9d4e3bd4e604eb13a285c6a96936a8aec8410b024795a1b1c718531d513d8e5c32a8435301069a3f74bfa2135602ab257bf9b68d88e1a8bde74e2e3091e045da0e8664be96fdf2e24999a808af1a7274709ed9e5c1851ebf7a40807ebdf97562ab16c4446704678008e97f8d43df18c33930125d967040bf94770105e03042fcf0ffc13c59efa64b180a0c1420cb4176ed96393f297191b57054f2480b63deb94a625934d762fa1a4b9eea36fbb96456aca8ef5582ebccf93eef6e4f7a9927398eb0de977a2513c9cb5e167140640c22da3f8696405799445d96fc2226519931ef5f19cb3fb2f5568a882019dab4bc6d5c8bf961977531c0f9cbb6656463dd5e0f0bcb261ed08d7581b949127821b7077d7588c96276cbd663538550a9a6e98d57d70bfcacc141afaa13afcfee324381f21093f80c0340035d1a3fbfe349daa90e4ab9d1233b48d314ad50f534a3213d1072a1ffe4439d6e80f44122d6949d9deb415bc418e1c86ac9ef276bb6134a220531d78b633cfd654cebaa46fc50340c8769127974e92395c027eec04b9ba8f5a049dcd16e5efabe587f9a049ff8bd2616c3f4470533d6f4a60f571a56f1c60ad315f1dc1fd0c7d064350938f521475902bf8e5c22ef7dc9fca0d1fb60677681f5ed9c88bf0cd9548e87444396d5b057be8dc39351a9f99b46f1a11f205e93e7eb8260930d97bb9b59cca0bf70e9059be77640debb3dc7655d8d56ec932e40203f05a220dc7be5317c6a200f1807e06aa261bb31aab2868b363ad0f0c30cfca4bac001dbf45bc9230257647787362da4152607d864f76e3a7b664a237eca91aa7bfb9d54d213be220ca5747464ba2df1115ffe7e389544548df21c38f443e582d30316d01f07d1b9f7c2ade707f072447aca5c5ef2acf22936cfc5e73801a6336c0eec0e7224f2b8f8e761370a73d52714b0ba9c8081d47f288b96def5852bc5827fdfec83c380d7cebd216b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h4e4475348053ec4e1c80fc6bbd132e189e67968a62ac02257457ccacfdbea988638a3824f0f4eb1f32f59bf9888c38806ec5e5fa5e124f342fed87cb9cb0c2a6ef15efdf3bc1a9f993785010578db6cb8846176de30cf0e50c90d9a3cfada920fa972eebb4cf815610c41169ac9ff4529a3fd165cad6dba420584926e8cb85809d229c0c53be3811aa974c1b201e4a92af17d99c4580d690c86eb666c00d12eba4e3f3eb75daa07c46130782997eab32d7be5b7a1af7a99fd9ceba9b3792f76a29c4740619587564f0b834975a25cfbcea267ca78285535dec4b1284481c61293352273dad7e48101ad42eab8424f59c959247235b7239b72fc18ff980ed9a9382b59d0bf24ba332a53700e0cffe38c5669dfa17db589c9936c73f34867f98aac08912e186c57970056ea152f2641a0ef228313292a1ed3143b3182f9c79a694bca9af389b02ae2ba20abbf085623d547d26f936df42b8df203233614fc34defa9753a5ccb3558fe612ca4ca17522560141a57a8a02fdb6f99d9ebbd0e10f98c6655f3ae4051e088c8690bfa9a6104c4859848b81bd342dc371db67d01cd36d5503c82d54eff77f478c2ac08cdc32c68b75313942e666db73780cfb020431c3273c53a5f33c35e8d1545591b76e4bd069ba1c1567f115ce72194616dc99a83d169759c1d5f95c55fcd252da329b1ad1beac0a5709f179ab918175a9f0c42354cfaa0f808012b0bdb87f1369f35b02d8661a56ed3ef3798dd056ddda2a553be6ca4aa75dd7fb974360de9ff2c26d135b267e54e5e066cd21c76b8ef3a6a15f2434c4307845a4f2fdcbfa21287591c1ad929c7c1639d0cac91e0c539f9b352d801f6bc2494d4a5ba8fd878b0da896dca24bd5192768f365123edc804e5608861dea27c1ab8839a899d20c6d7d09200adb1c59c44ab7fd4961eeaff9aafba58b185fe2004c588721f91bb216e6d619942a008a73746cb7b3a8cf6efd7d85ee4ad97e279b3163c309451c12e48fe5765c6fbaa662ab1d42475bcb1514e12bc9293120c1c29f6739f63a0df42073d1a55dee106e3fcd3f925b98c01070da9a056dcb4745cb257f0902dd57dfdfa007deda90b3f930d53d7a0b53ed08a31eeb780ef8a12fac4c11f0ab7798536c672a8f31365f44464de35e9e86408dfc55f9c2cf91aeef330fd92d141b7e88ea535a28ab7e65313868fe2132273b77c48aa9fc8535fe8140d5f4dcfde0ffa29a9612bc7f1d083f48ad6cff0ac94d32896acdb6452c68657473b7958f1cdc2d2320897b312703a11e82d3fd8465eb5f11686dc202d8ab2f769e14a7bffdf63482b956d175877edf2669f8bb8681d03bcd662e052271fe6818cec547063b52419c75d47e2a8a79e74cda5dc317ccdd52c9edc2c7874ba818fbe61d7988f7fc2c13cc79ee42d49685e67af28890ea7f8021a70d941172dfc6398439586671ba081726fd9b459acd50c06e1eb3252d489e063ffa8634a605828ce1aebfe60c060906467025811ca24e6f11bf27576a536e97e7d0aa51f5ec758a726a88cdf907344c508ec7e8bcb7dad3d3f0d76f76186000e0931551b23d9998e5968a4faa40f633a38a8f7b7f40f3631aadf50c8828858db1e152c2fdbe3d3ad4d0face9da91af0d01493aa7afc2cbd7490d5d54b1716d34bdc1f30a5180d41c8a799a5251a36f3167dd92d98e205d927885ac6a5cc83ab4754873806cfb16b08735b04283f3894584891a08b59c62f64570a24444614b99aedb10e1450c234c8e24a593d044edc2dd3019adb940ab2e20743f3338fdcbf52a64d52960cc27fab5f6298728d53073e73591c7b8c32896088181b85efcc25df0eeed1c482ce8ee6b5d4836283e175790eb978091e97293dbcef0295d810388482a2d78cf319d1f57372fe2cac35cce7f4fa908da9298e4fe9bcbc941a6ac031e96b3dd79b4d14a01f491df1a605c884ce8d0afaf33f5273b5568b859bc249b8cf06b65c45d6c61718f59c1b24e7375cd7d3228facbeef17baa66b4b7988075c5d251a8b349adf0addce196f175374e5dfa2df039e7712a54846bd8d47fd1817306a01438bd56be22a958f50b678ef8bcd17b8872b3fbe75e87b08e86e55b51da7e26bd52b62bb07bd2c8fa37090be3019634178a1f6569da82115288f55373abfc7f6bffefb7ed86834a54262027a449215585ea7fb7e6e55ef580b3b9a10fa714aa6c2f9a8d642a8c9b16ed81a0a18017204247fe070c6e47fdc3332a3e196a4b46f03385660af137b6a6f5977a71cd723fa624cdf125b79071b07d47bb7ded0c2eed566ee87b77a8967a8f3aa92a529d2b67e111666cc22e3675624f1655a513eafd5fa785a6c16d51696418cb94a994eceac694c57309a19b84d7ea17fb5156f4171b12782f642130805942ffbd7f58f084f2715df74b524d5ac60c5c5f4e487b3c95c97d1a5a8e6ef1fec3c773b02f03c18617ab175d3d267d08a8c4ec2cfcd0befe9a3de3cc50db134639ac08c38c9d8216a474867b5875f4ee9879079781aa90a7fcafd6bc3ac0445771cd82747c38a80f67711e74f7917dc333a4c14f8ff65cd0cf5c701cd2565a14dd9f1c37e3ed64f8b1af2ebc226f21bc8e779804508c84e01b8967f748f31ab70fbf580e2f582350e61e6e469ffd5a0946c997aa81d520e2eabe47de9e3f5fdcf221bb7e4ab8e32991a18b06bd74016775b0f062af444a32cfc01bb7301b8106523e7b17a0dd22dc1727caa45ea1cb0f70a2a45b1721dc4b4232e8d1ad2e53e6df56ab45892cfedb8c015c7c2221341b73a4828ac0663b3e9e2fed9acdd756a0a286d8681b69386ee401153aa1bb36df3c2cdd9a8a82c090bd0c8871eacdd0f89e45a4dcd3194fa6c16a910b49b14ba70c936cb83e5fb2d841d9ea71b05aa864477ab1f6f9694327247ef4d74773458b7486fa4f983522d0354557072cab6a8ab1894264309d62256b4b3d4f621ad0928acc94ff2070d104b80fe919eed4fb7edf6a704542aed0e47a365574c9a3fe7815ae91cc0e6abe109f78e3dcc0f59cc35a4ae3bdd66120110d37839eedd4e07887334f62854852b2e91ff11e0084a0017073c663c51b88a8b69349488263dc1cfa0d7a9f5d4a86761aa072134a4d92be7777a133ae4fdf7352cc7d8a47adad89f387228bd0205b6343e37fea3c9345a9c20ba40f7ac3ddf60dd7a2f26f4bffb93ece73c264c5598b9e2142d26e61dee67f47d1f9046ef4979059f59041c20f14f5d856ad967a14e2d52436498e60428a97aaacea1be718299549c15bafafcf55e2f4fc894c0d92e5ae3cf449243b39a563bea70a4de8882ed5d584986c6d78b283b475d04c2b05b21c237c05dfde5335c272a8e6fb0d6df09da156465000770c5411d3f919338467a4669f643cc065325d59e991e588a61771537b0e0706a4111c1ce3d6e5649d1b2d664488896ca6a1244682385ff6c4732e14d1e1d7001c7ebc4459b8a1ffadc4c6b1872d531ad7386d0bd94b56dbe5af7f903af162272953a36a40a944720a6e79d15b81df433116e6018ddfa5980c57d6b05889ac60aae8d3c9df3350ed40c01a6a310bc85dba799b8cf7acb0f8cd2c3c5f2cef6c609439d64550a1300a1788a8496263c038c591a97b633388870c82fc52b35c37c9b4ddce26c5e294e8aac7a018b1afcf0649fa503c00169b6b9875cd60e5cc4cb25f39386dbc603df9a774117c6266c94c8d9ef4ae298ed239b1ccc704ee805a27e80df317c9014b5eed5bac97ea667321fda7afa21faf82e3c7eee16c99ff3d3a26796ef9ed8284f39ffb77f8dd32e379c0d4e7236c3185aadb5bbfebfbfd61f6725844072d8ea26f64dbf67bd4dd15e6807b18a727812249a92fafd6ef42e1b2dc1cf370bacadd6b874634ae261cadd97f729ebddb045e51bd2fe30de523e47b15e8e07a139ef7186f8704d84df80cfbef421081adf8a3efdfeafde4ebcf4d1eb59ea19d31bf44c7257279921f8920e8e7943517c6241bb5fc832df8e0fe46a8a1109cc545424740ab3ecb1340a55082e0de9a1f1bde4d87ce842e9bc505af482c812bf750bba86a08d43e4f9a3cd8bfaf1226ed7390b53218972f3cd3af0debf67b7af593c8199b9629a4437a8842891810a35235663af89637078cf1df4aba998d2ee6373f0915806abb27ab0289065f212dcf15e64759a7923e41362e22be4fd037b0a6341f947b53cc1ada6ca79044a4ff78eabb350d9b7f2a52ad2b5550f13af7fe14e51617f528d41b342492b3ff3601ce6d6d4555ddee26d13b0b236cc2bba636eace68dfff3c0757c2e7f3bbcc4c92a160aa0408366cb474587c137816cd165d6c37de5dde66cc97bd7a0212c61c744fa424223e929c88d8adf1857415d48c43f92f677c77269796a43d4f5c51d59e59ea17617f095a62e7503232c67977feb04f46733bfbfea4d87a51520f8dcf138acc8c3a431d90c6f1c5f951536463ea7a7ce90f2638ccecbc45eba525e49bf73b6f1a1c0ba118f81483f1e09b224279221821f72efc0c8dc5aa5deb9b33cffb49e19088926c5cfb0365a24c15fdcef039c7132aa7e78fbc4dbbb86959e7c0b57462e7e2ef98b539771d0502d42705ffa7aa0fe3ccc0084d62d54bf33506427d7733069fa9d5db25dd77ae674a38f22a231c4eae94bf466c2c8fc4809918f2e4cd90a167bdd4f53a146ca0d40df50a2a34033e6a94783958672a624e00793d64b7110dc6a174b982ee4cc082be6524189f00bf19d9c1217bffa359da27a72b1d611a085759a188d0e3c1547731cdceeac8b510e841b2cf72061c75c858ac20da51f8e0b028fc1120daff711b7334b85febc54d7d0d95ee14df489a195e52167b7fc408fa4ee7416e40ae5c2c7ed6001967061fc54ea355c2a01a78e9757407d407eb1d11edfaa4b0dd9244edc03feb80c18215bfdaf17d16b45d433886833a91c3118cd349b4f62003f097955307b4372af18159fe9e8d4962f8e41449e0c2057b1cbbc70c271302768285785525d39f4336814e5c9a9703afeaffc6d50387aa84eccc3106085830dec676417a2e7afc3ddf739de454632270d19d82e7c66968541f9fc9e8b1a1f1ea90e7372a27dcafbbb8197e8f429cb78076d96cfd13fbbcce790b4d3c468dfc86e48345d9f210cef19ecc594507586fcb2e135f0054baee41f61c1a3881d19c648c79b8699d04198966a6d34ea8a941dc6da2fd505717fd194f19cc6f2567368fbcf92bd8379634e9cd651da812f110ed7d85cd332ba009aa4dd183a6aa476aff4863caed09acc97dbe10694a25cdc6cd4c75dc1b2ec308c10d12cddc422233cccf3c5b15d9268a73dc490dedd2ccbed8ba3970fea072d58a8bf1eda2b62599f7fef64214df4cc55efd7e38297ffa747d2d8a90347cf019ac374412fd6167289092c27191d8efd442d2910148b12c92f63bb16afc6c398d3a2ccc20f9eb7b8fae3c2ab3d6dbf1e5502d2fdef32bce1b4bbab12aa7af560e25bf09b3f7c09a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5ed64c2122baa2fad217ece090a9193d2492685024de4a2f45bc611dcc4f1c11b992b75fa251a44938e515395730c9dcce1cae294ba6347bf4801c52c7753c0edf0b8f9601396c320cc28f2ba131d7e54fcee893239c7751ca183de879f5d3984cd82cb38cf28a8b6b0ca413f670e344cbbec2d60dc5c789e59e6d8d1e717da4743fd3fab7b60e6905314b1864cbc363f4f8aa7e3943b1f02519ab7fc22241d300efb72ad4ee354e73cd940400bf0b43243d6991e49ed508344974d820e9a52363dfb5707c9aea2783d5f9b4fa272e04e9f9eff436a6156a40ac9cc444628ddb6f5405f32605c4d7efbe0eae11527259155a3d8fab10d31167e6052423059861d654223aa66c2e348130ad43ca9cbfaac56567fafaa3730697e76bf196c5a0a100db63ef2fae0b99e3c5105085ed05bce6cab0fce62791adf022cc316f9ec9ece236746dae818b458ff9610f0369caa2d35bdeb9261cf9e36e6e41b064e1c376487eafbb9490fd8b32916ccf74a804f4a354a388a6458b35a3af54f0f170b5ade21ee2c1237790735967ff657dbe2f8ad080dd82497a3680de7938a601f871c3eb29de6ea649095c67cf3f90e1c7c9d0c39c5b4f30ba9925bbb665e8a2bd2617d41b5a522d1d175ec7c4e72367e5a6c29065074a1cc8b95286f263b3b404275036d399b8355e176686193e291b80070f6d42ab9bb509f207fe6d304724ac2daa5f82ffd06a4f2a4ab7f28f5a0e6c136b4d37eba7a5cfeff9effdfdb50e36deb6d6ffc841697703cc0b511114008a1c3abe4522992c998aa9b7817e9b7acc44b620f66bbd647961960ff062fbb74d9ea3b86561d079468abaf61df28853680299556ff8f92800dd92ad3b9dc581a1ae0638a495285092914b8ff2c6c7fe9c497b90f1fbfb15567828f7aae0146446745422c25bf5751300ad868c769623ec1a3bb3599a159a48a53947ba43f19c4cb9d18756e3f942348e6efa69a647842938270a1eefea1703f89aafcd2c5b07b03de68e17f73b771e69344d274461efe4500031953955d2b223fd3bf28e016e9891a190bcb92a61205fb07643785c29872ef45f5ed0af3bf58147826ce0f174c3e6011766b0c8dc29733a2d96fe113cfa4a770193bd3632a3439d9e77d6d0d3bc8fdff641784b0fb5145637fa61eb419b1b70d6aaeed3440cdc80d05cb0adcf5fb6ec9b85e1abfe3fc4bf3712a0e45b171acbb0b582b5d033dcc425b860c2661f180608254b3c1e656607b075a1b6575ef0693785e8a943bfca38128a9fe886b6938ffefd15fc07905343b535148a35adac747deb0c6f53c8419f98b08d83290dac26d5fdfaf82d861018a151170f9a98bd69a2b8005e4bb317c517d87b15a1b2ea1bc6bde8637b43ce36e0d5b2ac84e4a155e55912c360eb871e289564b3e5fef725cf7ea7c4d7fb87b0c529dab26aa2c0e98b1b445f77d0954cbc14f7e15825824ee40f2ac24916d520780033945308376e6d2e4cd904d467b0bfd8851e2765f3abe7dbafde44ac64f3611019dce48b8b3ebb776ed3e1be35b2d383c0cdd7005da6622565b37b162508eb5b67b7f86813efda2ff5e6b7ac5714bea0e345ff0a7e5138e0db555a347c96163aad4dfd88216fdacd837636eafaa49552ad43af1f6f1f7104255a786ea6da7eab0da2b5c46cd0dad8e3f8cd13203fc054a191dbc5a902b40c9a7c65167d7900e565327121cf4a06636accd0a63cbd7030f589f38ea3ed27bcba356ee00b9b323c230cbbd4776c33ce0580015943d05be93c2d65a67cb5dd7d32fc6af91ab5de07d6d31ead964ef3d437aca3e908919a0cdaf0981f3ae78db9a2431f9e1262f86381183a6250a9373bbd4b28b34807a69cac090777c7b953b3dcd4d4cfa7aa5dffef1b0e50c093543466e7683796cd87965ee012b7698cd00e9c4d8f8465b0b636d68e5a730342ca2899e1c7169d7a3b21a59ff105b8d4c5882fe93d67ae231db9ac6817b75ec21b286fcf1471b681ab167a2df70e419656a2de6a75f75ec9de599d21e2e8d71fbef82f8fcde0e7ef0c87a3fe3e0884dffb9695b16e2cefa6e9c575643c861a935aad6fac22cbfa0104ba8688f96dd842f41bc17323f84e636b8492acdb585a7358f574dfd22481fd922ffb851fa7738c399b6e61d892c1f1a1528804008ac00fbea54756d06c0f4d12387deca789b147593dfc6d2d5e9ce5a22d05ff1512d214b933aead28847373051941b072521c2d204ebb5d8cdc77b12202c6c0834ce44d23f8a0329e3b93379e4cb4ce4a0f539f96959c6cf7e015c97a438ce5eb29b0bcf16db0fdc15f7ccda88a8248747e67ba2ba6dda54242923b8a6dae5bd16f7bda78d1a3a43afb908beec4cdf5ab4f08d2165cc80c62ed612edf594b23592d0ded353cbec4473964f21227a272b1c804cb7797b4a82719cef3b4b4386ce40c47ce3b7ac69c401a3c5c481c625e4d8761247cfb8844741aacdbcb5975eb196f95eda151bb4733c37daa3a6ec1ef5c2d8e57c91ee1dc2b78f652f66342334dfad85c43e0269db7cf42aee2ae9f60ad5adc1f33bb7742fb952750e8fb0ab1cf244d1290653e41e01a6d76fd5dee3138bb3f90738d5030a1e85527f4acd720acc603803dea09c2776acb86a80f0f6ccd5af713b3df0a52519a89df53de03fab6f15fa5e52ba23042ce6a07fb117347fff2ad1f4cb97e3ae391205a98b1ba3611d1217e8545679510e688770f1bcbcf417d5a475ecbc7af7ee854622736ad5edaf9e81ce32e78b477b57be39f8e99f0981287f96ccd56c23426a9f3887d78bcfd37038fd89ceda7fe9baceebd0c04a964a1df9712abdd52186b3067faca14c9ccb6b7d0f25024a1dd472b7120be1b5f1326da306923ef58b61309902370bff07d7fb9e75161945fd6449c88935021cf467e7773e6f00a833a2cd18920f8fe97d45becd27566287cfdcf06e034f8f316b6ee8b8e788c4025fdab6bd2ac3b93158009f975d9c19dc9deed1e9225ea5b8cd437a9bcde4725895e0909e3aa0a537ae2a78963622b5bedd6b5f4c5241192f341ae6ebc916a7eaab202f2b9d63801290b89ac81a69925d88cd943f726f8488f05075cabc205caf25344917214e293c5b3aa7c9b39c84fc669eabc377b6186ebfdfa2294007881bd38b4e0966c82b02147dd79059632544ddf67152784ffd9575d2fd2e1c3d826eaee6ede271129cbbc57f39662cfccdba6a4b8551c3744a903db9d4aa55fb35f7631f6f0a1471ec31c21c4211d1f43ab6c6668dc93f1c204196071323ad4ec3be36eae7d74295d11da3d196d5c13f7e4f515b6bd82ae7a672dec39f75d14da0224f37e1b47056aa49ffeb346f6aa7eecf139744ef98f77c8cfa73fbe0bad58335e3469be5be50b7812e2eb96616ba6c397cc2fc87168ff05bdc24206761583fbd8df854251338bc934e78ad21baee2aeb6385200497d697ef45a3201e65ab1d372686fc5123b096b93c89ef1867180e49121bcc093b1bc71a666f57ef9d83c06be1b56a59cd4b522f0f7a35c05d40da6ace3fa8ce80d8bb9d1660611444f4159d9c1a582448690626cb3f36b534a06ceb443bd8a8f869a4f236f3b951ff12a420fbcdcbc819e9d92d429905da35b7dcdbf726dbff3355bb4a4a8dfb7bd594c1d944d0e1ac4e3638d3e47a3a9d7d530e69539b48d51d7d67f34c0b37f4ee9eafc2a3f8be5460ba79fd08f2624ad7665df00dbcb9d1180338e86177ee714820ea1f48e2471e2e690ded12882736791e3d1c2329e3e6ba0f9aec5749859b05a67ef5a75ff05427a949ccde49cb0f6f7e1960f124c2a19e0e04b61ff2a57a6074d1c0e7cc28003466df8d410688a706ff3f318744ef9265b6c02d5398093c84afe9a9f8bebb6fd742c1f6508f334c1d0f4f9d407c6a0ec334cd04bd154185137f7dc3dec2e72ed5676acb5a7b0982a451a954f283e8ab462ab30a09a8adabb4cd9e557d1428f19c672cc0172983269ce53cd7832707b38ce5183e3256d9c3654b017116fe201a2ec5aa0374d0ab8a18224f18238f0aefc846358002eee864a2e2842e2903f8ffc01690a4db4f261e24e0e2385baac8dca2a8817faccd42c002eee9b9f2a420337137f7ff9346beb088ed700d8977bb6ab76e04fb3b2d035786fa9b7282e30a615f3fae605616f8ea28036f8b08113024280ae90daa0944c3f76addfaec3ed5d9b103944839bc77d510eb6b058c4be7e96298f36b1947c71456f905477a62af31b676b7b9a0f8dca292165656f8039f0abf2d98b380b64e7c6b0a59a5f7901016872060749ef58f51196730197c553978e8f520c4ff96fd63cbc555605ca1eda046dcce0a7b8bf3c1d2afa19d6939d92416e6ed4e161063699909f41b4bc8c20d5e9b4026528f419a018641ba14baba9c4458c779e6ae7e7739dfc0f4c4ff5462790b5e24247b6fda8604dedad1503ba4a6db1499c8565b8732ebe5a2db111f099591fe33812ca7155ea5b594f301418b6a39e0be36362a7bc1695a169cc900b6d3ddb6b17ef30f13d265df0a2b1a26adb35fac9939ac330b271573d7e4da2960c8ba8d5df84f5cc85be4255387ac52b8f4f2c5d455010521fa428d648873accae1fe090c821db3b8430354add551a7e2a1596a9fe387160f34e81c75752135c14b9995b0258ca35f70e41b7604cf4074ca2a5854b141f023870f0b95c2c0e409d41174e4935776725c8859d41379de73a2fa8ee74df7b05b4753e6e881f5ea6b1680a8564a9a3e6f3e84ffca685d52bb49982f034ed8acfdea5679e3de6470efc29607f33c22e95080db7ba9bfea141d751f05bb4baaa1f9a8534cb320af8e851e3bb420fab5e440032d485c983a77f8c1d58f58a58e689c7b00c568168954baab4ec936871d6978d1453a99eafbbb75ad364873e6a791c34586b7a31bdcb66a9dfd6a4380bd2618a4285c4400897a5e7edcedf72c008a033f8b03eaa4ff86e13d0993ba596687d98efa6ab223142713b0f46b2f8b48c37f6fd3b2bfb75c373570a3061e19dd3202b5de5528234ea031edec127127e10c3c2144901236ef08d8e635dd9ba317930bdb1ef25b0b5669aea9358396de1c5887e74a0a2d888f861bc89485ed96d46b0799f623015168badd1090fd43db469f8221dc7cb496fb2c2d9c2a214844aeb1de86af1337f28df560ec2c8c643eca6c284dc05ccc98dc10c559026318927821416004100f9feb78dd52373cc1fe132ecdd5accebaa13f1ddabe260a8e298bacbf74069ce90adb047b77e9843d8839157d780d6c63ce75eec93bb32a30336e442f134744d70a94a4a1c92051ee5edc9acf27e04f6eaa898591387eb505257608bbed3d59844c6f0121cd277b9266f8c824810cf7ec3748ee6b9a041a61479cecc3f107c689df01718bdb6b97577e504d14700879e10507f3baa4717ef8989130e45ae83c699e76d35a902cf161dcecab412a6f57534c3d98f94c7435bc8540471c17c48154b2193cfe0f6dbb8b85d99783a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h747854a756a84d050a87625ce929d1b34938440f4836457bf6c279eead9c2bc0ba429fae29ea8fece21185abf23dd04c8dde8ae2f58a055c2387366c7c835a54926ef1540ea45f081901bdcf205d4299670a0814dc8f0d2947467272eeec412653ac15b719b9c34c4d262d31d032af64d04e1e14134a78cc71ed89509ab02ddf7ca6dde4485302af5001d108872f80c23f43e2cbde685fa7df43b97d9b3b9d55448961afbf96fbbc644c09712cdf6f1cfeff251bc42a13911588c8b45d2182875a49a5fd16683ac20051b0982598c3c9d75e808916c7fee608d1b5baa4c180047870f2a4e0f2e50392c003440f7e0adde1750d28e57af344b7eda1fd476cee4c51f9ce5c325f6d4c931d69e6cb75904b49b358f2745c7512014b4e31ae1d987772732a0c9cafe7985f5a2761c761ebf8d18b50d1245c50ced85f2cd5b2e1e1bb084cff302a84820093b7576e6d87bfc3bf7f12a0f3ccb070d4dd9f39ba8dfac8340bb046d14b6142fdb61691b7e9cdc768ff7eee4e9c8e87d4f401d70d0ab060462213a0baa1fa2a727b45914e8d5da685c216156e31fec25556b86be05e7ba63fa6576326476f24cfcc0499546cc9abcae59756e3336bbe2897d357acc8fa4c200d163f3eaedd13fdddd8096ed09d39490afec7dc70f700c2340d1efa8f1709b9fef77af2bc10ff9e5d8d2dc1cb6f5bb8f8f0ee6b81eb19adf3ea476cc51a86a1f4dee9aada7880baef076418e9b42caffa7b3717041f1d9909dbc9e37e43ff81540ea3ce850307407eb43ef642a63a364e4ce1997477e42888cfc3c25ea0aa837d957543bcf87530c8ba35214c8e7df3d094f8e52ca2f39cdd7e6477204b2c155d407fa9c66b8085ae5e5114e3e77034bbec1c97d43536653c948277095c5a58184840ca74a0b4cdc2c050ffe526f003368d7261b6d7bfb6724e1f23845498e5d16d8af89273d0a714c39b9ba718f535072ba4571b680307e8cb2c84eba44db75855922c15fd160e8fa823ee1e4072bac663d271a212d372279de24c96de24ad107ad3b12d90d9b1d05b73a1a30cc36587e2cb51889b8a2a51f6caff78f3214367ffbee72517de16a71b56e99642346106ee665a810ea282b39c61c5b25a96b17529f7ecf1cff361ce07f7544f3af00fd81f566c912e89ddb98edffa46ad48f2eeff2d0e94916514e7b63a172fa27504a779422b42f53e3882ea40378e3647ca50ee6858ac01ab020d2a17f7682f71c81adfd058f1983922257bf08a7db764a91ab6f3b1fcc5a66bf9c0def626994066304ce03afe2ed968449e3681356cd07dfaedf31b0b87cb1907af3c8d15446909380e12a10cb8983b01774877abe86d5572e259b61c5d99515160d2e1126c46c62b4abcdbaa13f9d1d6f2835c78353418a8cba8ffbe4576b18c475ed6477a806bf45139387a1afec44e4d0a5cff85a3c7292ed1033b4535541b263637e9166c574fa9186d91aed16a343ec3850347beef5bb542a2dd6367687963ab0985c287c775e57f0c94047add5aa795a66e9753937b7c8df615778e1f1e68b9a8822e3484995244a04328e0583b4b923d831e97cb2f7f0620668c86b5b77ec161c5680de8dfce9752440933b4fe9345f3e951bfd0dc4689e8d85a74b28812d95193219aae51d4fbe747414dbc7bfe7a0bee18f2d274cc37f0714faf85170d3fd1fc7cde16a9a844a6cb62847e7e01d3e0f882edd57e851b7f399426b51ffbfc2c26d3f42624b6dbfb300702b2a5bcfbcaa2657a636a7b073f4042378ad5440c5d426d4e3767e29df54953fc2b1bc0ee08698a4e62c0f5c9d580304d622b048cf43032b75b95154cc8bfa474c8c8036cb21d0f3559743117d2faa805cd997e3a69a970623f11a035cdaf79a2d3c7bb8977914c44f7d9902a27e5d57a3cb1923cc12dedb3eddd35b4c961125faaad36c6c38f65c66e4ce4d59a9500f41873231c4b45c8f7e36e88f2ecaaf2903c2a37fcfe39e6341e3fd8c60c1987221ae778a5a10b444e9d84e033fa08acac9a50688c4ddf884c3f587d2af44b4b6f9fc224c3918864786eb2066d4af12d13f2524e288c34d59ef27dea451d81c946cb080ebf860c53ae51b9cbc37afd2f7a4718dcf7365c65b69c7d4b801f8970e250a4a420432da3a16b1c89d8a8968395a8591950b60fa1152d0c2a12f86a674d248d9d9291a78d943e50a2cdfe5d216d7f136c7f2e84215e7dd7e6f4b1615a24fdfb3392193091f0f101c0205013b5f00d657c50e128e0f54e700b6d13c3bd1f787bd0a8a86f082cdd3a5c07bdf4849a48380ce11add97fda9a8a1c9b3d87d858909a76d032dd0ca7778e52cc0ffbb114e569d4a5fb4be9a982cdb23ac22fdb97c41e6dcb9d1f2a24e904c35389d454447e499a52671da47f13972ffbfbf1656dd3a4d1ac5237109ed62b16ca8f40ac22ed39897deae55540ecf33b6d33463f2c1fd1c382290ff8e065b4b723e47da7ff07bcf34572506c6ca6cab3caec41f3b4a032d8bea9f7d2934a41cbdab7ed7c2c0da942eeeb200cd0500a4300257befa2a1c62a30fc9705bf50fd69af9edee52c65b13e53dc60f170167e615aa183b21261fa85a9418531b406e3472c081506380381e633df317c6d6a5255c519e5ac85eda6b98de2d22ee67e4851b7b305d87373181bbc2ccdb714010bdcd18febe194169fa00ca2d614d48f8e3f629659c976d6183fa909358b8ad6d082dcdc48f2e438ddc72ec71a0bc408ec9abd6c82d66b66d78c9b1d6b5261d65addc7fae57768dc3d6da593c652d82e8f1c4a6fa67f42fd256d7b9b4338790ee27fc54417e3f602671abf5c2be0f1744c0ac0f86bb7091be3a4522f31a86b762706fd9f5f7ee7ffeae871a8eef8e72c98df4f29d891356ed5f8c4b6a3cfac6e8dfefd15c443cf864f99acbb52977cf04270e595f88538e498b83797850c23083e89e3b5b7dbccdb6401def91d3345631b29b89c3d011a679bdfa26ee582c6d5ac32680875c57f456fd49ed2a8379fe2dfe0164bf59cdaea2d9d15469d6949389758b1a3336a71da9d9e0ae63985d90bc3a82a15b8d7d8f6b0675670565df2840e5cef4279fb4f34e9c00c180c049f99d8a42d31a36f36f5dea46e0a76fe01aa63fe7326e40a9518fe79b2bb770a52c8908a43b58cfe537e2be74b8f201ebed63cabe6431dde89e70ec6a638f0ad2d1556495797322072cf40ff3cb142c1d7730f2cef37354f06be62c38dc0bea4d5e5812245e2294bd35b95a86de93abc8aa07e1b8f416cfa1c3bb19599a772e668b1fb26c4d135765cac3624dd48f90c56a62ee2810814aca3a0cda7d9f8db91e0d32fe36183e715b0f0797a81882b8a1962fa801f93ead66171dc98463129c92034c2c876721af4717708e5ce46b7c523d9628371476fde507457bc7a5505be816f31227fe510fa73a22924e12215351d5fa41c25fc73b6d6085d8f381c7cfd6cef265d4738b97bafe0f3fdb9d973aebcc944f157d34707b02858aa190cbbf034c3cd68969d9391e859b604dae898142cca66b2ee2cbc11662477ebf4316fd7decd468d03905576e05beebc850f9aa1a8c1c9980e7b9f115eff3da6a64ecb39e2c2b2efd8757cce020c6995460355297bf5f106b5aa8d0814c4f73e3ae88b4db5f37705cc6495af56c27fb5a464e44882c3a97d12ac4c7814eba4f5f85dd4b41e3911c7c195a14e54943c2c56ea6118d34aa465869dcc20d90068e9cd0f621e4419ff435954235b94d6cde146500f185f3084634ab38bd3534c46ff2325b2c4ef939604cea540f3c3528aa3b9f7db2a8a9b8881a5aae6dc129d1979370037c52c81ca620a429bd3b7a7610be4a8888b812e44c8718dd4388e5de4c94152885ab998a9439bfa8d4f027220103ee5a5fbc40599d7e501c467dbbc95805ba289c257fdf15a9b6b7e59f2bb8dc68be5d01675653753d6e82ed23fdd0bc3e55a3c929c6f9fb05fb64559e5757f93781feb1c3aa115571b892733f6e97e1d76846e64b28678ea57ad3b8e71b64d2ef587ea1397cde580db50f9275d504f06b41c9c87804043832b55a0d5959776815ebe2325fbd1449817d2ab2f1d6d77310d3284ee5c19bb4ef1b0f075b70e10bf1f88bbab4385abf0c3a70d65bd6bd392c0ff443f17608294c1c207dea8c5fb2d800414719f86d7d6c27461db1fb5c8804cc3be0cf555231614d40e6d48e15f3c2a7a48caffd6dfe284839b71d7bdfe95aadd84fa28bffac0da20e393cd3bee0b95054dab7500e3d59b8c84b42b1aebd640efe05c95088e4e317d7e098a89a49816bd02f2c80989969ed5186480db4a0d34ca67ef814228bddccd067ba98993e278865ae96f84b806f702dd10e8f762e624f62591000454ddee5b9d5dbeb56fd9dbf30e2da74bb5273a33b0f5be2dcf339cf4c489ba635bb3b671049e3f1265c082722beadd83c38efa7e24b5fc83936f87ba6737ae824852eb6ec7d45293eba65db66914ec207c328a6e7777f67a369d1b2658a2d9be2dc11794d223275f0cb7fecfc7c5878457e248cd3a3e9e326e8fd15187707b20d3eb31ce3bf8929c7d33e188ef41c89becaafb3101e04fe6c78e14dbaef5565df5f652abf57627463a7ece92b0fba8d0842cfa42c1ab20efe09b643d6a30dcc51cee05c1d6d6e40f9fa716dd1983035dc8b00c5ceb4858d1d9ac7d9f17250a813eac67586296e81baa6415623a7e32a28f9505fe8b320925b7e2c83749694a4f42c2e5b835db5f7377c80f16a1badd254283c4b88d7e37e7422e8d6d7ab5af4529afecde3bbd554ced69eca389724a0114f96ccf4ae2fa4b19e58a0b688395d9ed2a1724ad481ca96cbb71b66fc6b13bf2e2f9a538ee8cbca41f13327a416c7fa78b109c8cf3cf77f078dbb78e98c4f6e51b16dcd5e7bf1c77d1af6688f61528cbc85649357973773edbd9e0f5b8a2c5dcc342d35832ae9cba695c34165f27e48e2be90f08522c22c05105d8c4606f7bdf688ea61eec2e10c654a0c0ad0b3535b79a50c828986a3c15e5894a92cc698d2dafa0f5b743b778c04fbfa28870972bc8d9f4f0b0c9b95cbe12750c8e9f8e60236febaebeae54bd17f9bc6b8ab9f722306157a17ad1a0a45488fe880f07232d67e86a69a9e853baeb1fc3e2b3a0bbc4cd8ee276667e87d6988579305b59ad900d6dbb1a6f4848a7f72419c4654653ecf1576857f6f43cabb7ace6f94411196d52c7c4a8456847e388417b3772d2fa7d62e6a576b883c9a45bb1db1cdac0f89cdb725d16ea2fa4d9fa5fd37f22c447780efaebf919616890b687329f8d15de011b7021ab87099b361c128b38b505699f4378e963f86b67c1b2e9a72847680efe0327ab6f4a25a8ea1f5fc4687baf36bd7d5dfe7c3c83b569c9c205bc0aef42388ec8ba1eeb837e33068d7ad326a921277d9c305476d7ac76634e730551acf0a00ba94e82bb39ce5b1b9813ffbd7db33771356650830413bf229b52362c5ca8fcf6426c5f0af051444b79e32a9f6b2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha2931fcd21ee3b93c73efa9cdabda00ea96dc35601a8578ea6d7b4710f002354b599b22c0dc57cd83a5736687b39bb83b99b77b6dd22bdf0014275bc8bb4f7b3906afb325b3e394c3545857c05ebf60e1864273bd3f32530341c4f441ff11b0f9308cee75002591d000c790c362f98816b4a9428f528ea0289065010a5f8782d19258cb7c182af712f3909810515002370cfb815908644c8562532888fb06df8e3d280ede8df6874cc754757c1c9e1a3c608830f458091a5ba3de5c86ac8bbdef12b2d34099fab3e6a71c4f7781ca9e19c828f72d30f61db3ead064eb87caf9923f26d6140fe32f2c1ed10bc354b5fc942b195bb6f121c55870b31517f8ce8a26a734d05b0999271f8a558e9485c49954bedeb462b3cac1de8807402fe14ff5d58ce3d7a78691552c8f691451403292c3382f6b39ff0c6f87a4782e8a793df7c91d405a2e475ca7a55aee953b9c7e48233fc63f9dee432226db3227e815847ea43710e0ef7582c40bed68e4481a00c37872d71b96afd5df802d64ab15cb060433abebb3749a946ff7100bfc28641fb8d8b855ddc9ca9502ed3d95381961bccb90d112ae149ce0f55ce96e34e30922f5160aa27993061823bdbd27afb513c5ac29f7acb054ff42b1fd481c6012fbe05b8721d1b308b9bdf80e4f010457a09f538036890fb56e99d95342a2ec69b364bea60f9571164df00ca44584c28e7386dc4a3269cf0b9e1a03fdb06ec6c3b46301c7b578e1a7cd27dd067d238a8c9e75d6f429fc92ea6830393c34e189d2fca4309b804d690089d6c17cdd65e8e13a8c72398956a6c5d6bd2b8e7eb0223deaea60334b309117182f279cc5f70388be8e05f554eb93fd6352eb21c4471babc080f12ead360964cd8e4d91b3d09bd43b2a6786793bf26ea178faba44c2ccca58f3aaa48b91a7a7cd2b553312ac8d8cd4e90b472e71c75312934fdc9e21d978cff03d9314f3003569b9f2e2159fe89dc1d69e6e62f7d9af87f33899b81b75610586ff5e11d1d0483a9470bdf71623ab5c759f2fea94a0976ffc5ee0f855acc3c48b15aaab9bfff7543abcd25f9d07586f95e02f4e3c248882fbbbb002809016cfba62f801317d0ec06965f02f4e16f35692f05c538d205f8a97da464ef86c500faeef88b2c81e410859d75899424326fd7171e150a1dec015f8e29979b5b5adb314ac9b2f32af0d0ba379aabd73e87e878813d6360940c3120378a55ae91607fc27778d22c3a10121cd0f2c215b64da2f9db8f265dd253b191bbbcc080e1be71bf1af939598d62453febcb31193915d2dbf64ee5648b7a123b609bcf6d61ba03a8ccfc5d481005abaa553ffa650622ce7d6fc4e8c47df52dcd11834df0f9db2a684ba640c7a7a86c8928963d30974ee42b4b32437c3baa926c74fec2173ee8fad9b95f7888d86b77482ce5c971e236d3e4335803dc538e16e26b487191adee68d49d8fc67c92c036363015544cb1737ce6aff973ad1c5fee3f63b217f316aa4236705f2d656321248b2b33fe527216484acf9559f55fbcff50d88036a4b549bbedfbca0e455a22a3e045f5f099c07b29efc5a6bad5537c881a08a4b28255d3691e51268696eb02fe1d33baff80c034a33c914dc26f47f0d6bd632e67e45146150612d0b39e8f127173d2e53ddf3f3aacdfe87f9cd8df953e48723232f0c31ca89ef53fca75632b11678ea28cef5d67948f505f7258d07d7f75d7aaadb086557427da168234d0ea95cdc95a9a4343c12c8fd983f38b733c151da6fd086aac770990fc5a548870397526c077a0681082811196820d4ddfa44ca4aad55626aa455ced1a84ecb651d1c2f78fc7c0e66a1e231670addbc9662fa8708213365b0caea9fa187c9054e58b795773ffdf5c48cd4ac926162a0d7fcf99f2abdef6e7a9b458320883cef8fbfe51132071c95a75a3011bed154374a48927a7c1dacc17682fc98c5bb14bb39f94a4cb54a4012d7ed1390652de995206d7b973e17b947a1bd387fd18460f2a762b12a1ebf90bee0e9ba1290f065fbbe2bcb21a97edf19ce998dccd84f32807cc09ebf55e03b8a1dc8d850e01d609f25a7d13cb24154cc4be5bbda9a002ebc7b82f1f6ad1b9bc18609f67f9f1ab15535d9aa739813f997671bc4c0d9b08afd0974b356e8edb29e1da663ce4300fdb9425365b182a37d8a3f0ac743db592f928bd1534c80b8157961553170f1f2caa8ab61dc44c308940b1c6e50c18437abd12bf93f3d19cc472e08fcf497fd4cc96dfd2d55e40946813d2c32c75f6a15ca207359ac6b9bad0b48a1567bb5e479bfb5c0ecf14bdac9f57bbcb6dd786eb99cb66b95b8eb93184472d4fffc3e782915eb220bedc95e14523c9c11f92ffc2a80dfd9ca7f626a3acbe7c657bb2cb0e1ef97be4b2f7b901535d601ea69a5e1cd276253b58cc44474637922fc34d2b678ccdf7635d95217d75a97a3716a53ad56ccb529491c37c04e7b8f9bb0ed25eb77f3dc216678f98ac2b2502306d5f1b6a14932b614494ca302f76019127baa00907b5957fc1c6c0b995f554eb454394439e73bb7ec453b4187da9000cc8cd041dd61f39cbfffa79aae587bbc42b1d99378d1b64188078a31b5737f24ea7066d60cfa27dea39819ae5942b43baab34075d68671acfa5bb2f2438f84abd0a98ef24e1b4c785c5a009a2003f9217edbf4fd4958259ed4c698b7d5b76787a40e8f19b1ced8f9477955ed53b532aec8c4a2ff4483c9a3947c61c740f5a2c1911cb1d4c9588e976d7bdd9eedcfcbfd79eda8522fca01121f7a45c26d071753c5f3bd4152ff3aff2b614e3325614bf8e1ac16d8fcd19645d0c23cbfaac6f67a5afc5d8f74e16d961ca8d0e1a795e1bf2e627dc4c90c15453f76344eb01e6909b7f57e23b96695c6ac901d7787aa0a7a6197607194e174cf4b9a25bf12782cf31d66ae8ba1662fd9494ca954886353d79602dae749ac7dbad3d75943d03cc754afa5bb5a7c967e839c6806d01628779ef2f738e17ead7437a0db6e61e3208811f38d30d7e9c8bed3fde922c61ded6b133002bda1685c0de8a030f5ca5d19079287c9d898ea65836260b4a3a9262ef7f36dd32b5078f0a7d3016df3b80ac7239b01d12fdef0aaf69beb89717cb4afaddd26616a370e105cab4593eddd78a918314db89ffda5b10611eb6ec42621f323daeac108d4fa739f6a84444417fcea1b446459c737ff05852f5b04e0f8387f0c4fa51fbad87a3df9b4d53273755633522229259641c6d2a8e3a530ab5d8fc4925b44be0e3fffa5c789a5abcdc9562ed029b71d253e2c18e751a64f6d18aa5596d489f6ca2b34b7febc014ab06a3eb04323e39abdcce66aca7b6cec8e8529a6e6407055f46ece65a3dd6a01171dfbc756a465edf9b5fd06045cd77455d338d4aa2a35148551033471ed962bb7ba2d8d903bcea9f0d554bafffaa365bdf92e39ddb8e16bb995bbe3e57c09b2413507ef8df2b306c7f4e10a975ac8334b1f771a73374b5bbb57e88d63ded5fc4061e50a7990e0e93015f2d66a4c3839c5774a810ccd2c457cc3398662f910573cedd429f7ab3345f2ee9f2f32437b4aeb28dfcdb189c39c8063296c962b3b3d826f0b09c7021ee685136bd8bed08cf03756e6e5d80bb8cced08f8012e2484bf515589b6475c5b31e7d7714f7e218434c63d87bf21fb5541a93cf9323dad2068f4c3b91a13fb07ce601001bbc617e16201f473b8a6209066a14d1c8ad1d51ee640cdffa2c27909e7a07e49674dad2c184d135102b168270990991c433bb9ee6e27cf338e073e096f8577d8b548b1e7783e64726b363e3bd4687b6acd54435f32b6bec47054d81b95fe0b2008b08fb84386dcefcf17dad40f0fe5494243371eb2ecdf605effbbe02fbe6b668f6efc7ecfbb6f40c451feeca78737964b5ab039b74b2f8a991d04205bab2749c9581090e9527165c05c8d592ae26fd45765d4edb1999c7690931f71da2784e9cc592376451a1c659067ffcdbcac1eb7d19f9306623519505be428e21feaf16735faf946302fdd1327816740aca5d4fff1b3181ac66890652b418fcd29aa29674b361da989ce6e6c9235132a09215983cae783dadd8ecb3d8af3378c27fb36830e78a5b811890deb52e56584b1014812b4f270e17047ac8d69a0070933cf1bb15ff2b7c8ea9d6d74e262d5b5d2e6d3e53992be53da891a2b0ba1ddf268eccc0467985a4dc176f807c274d743b64ae8e4be1343030a36cf67b4b7684d22ef390bc9302129f44d1e1df7bec52a1a9fc256a14c598dcdc03b0ef45bc6eae78af602bf6143de0367224fc9ab90812c4b2e2b6f56ae0b91595e4cf9f6ed91caea90c6961a7cd029d39463a3fe9029880ed906ad9a26b543fa3025499394c47da209d461c58ab8409af43bc99edcce6014adafbaa16b96f14b861a92db598dfced6f40b799a83058da32e22b6acf0558a555ff0d4c880036e22fa8ba5238a079abe174eb5f07e2ef8ed7a04cb9f44c56f64ce4c5345661686630b446c439062b8348dff0cdb483fce2cce9a90b62161f2ab4ca7cc62e5ea2e08c23dc49965a770a1109eebf0cedbe1ba2de17300c7aa1ea39348ffda54fb99f5b0b89822f838954d970f21ec6cab79171a19121cf97e5df8458e7c6b216d185157cafdb2492e2d74d0d352f20502fefbc16dc0b2ab7c93d7e2a616f5e7558960f48c31880ca52209491bdce4dc4f488e07aa21316b26864f8a5aed954eb1d05138ebb95c4358ca22b19773c9cbf8b72c7e757b2d7d95719f1d1ce6976586a8d53dfc42fefb7c47ea58167f330628b794feea3d505568c05d48d08a4f1d6b9eed4deb429f84ce1610ab86a935f5c6d831e1a2aeda9fbe785b3203e3bed21a86e071b862fe836daaa94fe3b779a7f840df801ea4158d4deb10f0d0887a378d0b222649f2925947800250f412b104537ffffec5d11624b9c3ed74bb4f598c90368b2c3c303b90c0eb2a88ad4820b22af9cab765c1a100a967ac4963bc5e0cfd95e747fef5627cba42d850e5c11259d854da3d148771136f7d005a8526d6fa3eaa1e375f45ec0e1f60304430be7ab50ec8777e7264e60cb70fb137fa0d5583a49fb94ea167f31695e46ce247b88cbca2a80f1c4576c417572e518b06b0d395615265402f5d50ca30300728dba3590c8135d6467a6e318577d430ea3feab94e99e92da784e894d479edab67ce39892735e7184759616d2e2442b34388e5ed2ff5c7774d05bf4151caee0c35d51d80c127c75cdda00a38561235e822198cdaaabc1719265c6a92d9af8b7eac85556fcf54e5a2c23faa08f5a814d9c709d4beb4cdca625163865af50d47828cd8c0c4b4497064a745797217963dbca7ee73f7335fd69bf4f6281f1a75fae0e511e7602390c98d0169d17e082dc7cf9b15ee48d51ba2c8f598467f3f910bcfd4f1e9e676cefc58faa366aedb6456fcfff4a9f0f74d932ffa2923bb8e1a7c1d7e2c0dbc87709c54a89cf5a3da6b00e746a1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h56c4ab0afdcb1c0a149a875deaa8350c359379b4cce399df02679390e52e36f28562036243c1eb0981eb1039318c5235c90ecece7e3cf363c2f923f5b784a322da7e3d84308f0659541f156ac22efafe8cd44807374ef249951507f36c89223628c442c68974ab94770e8e14114b2a9f65d09d3d9742063d4c8982cddb5f289e3345694d3fb7161795a94ef5b442ff0bcd95ebb7b71a303f0b8a074815c4523c6fb067e0bd60151b13334e2600c12b0eba732e6822746643e7985a33be6db5f92f02301528ae9d19e712f35aa53270b848bb22cb467e1366647c9c09f1302cda0647109282b600665f68ac3b4572272a90d3a05594357c06544ae15423bb48fa9bdbe7ec33386d596dea74755b7e8c11f603e50329b460ce4369c7a0ca288d5d7522ec59c6604ed56f5ce104813fa967293951b639d081c2627b823040bca777351da5fdabe24c555473e72480c56930e68550a46188621d24e3011b2fc4318ac5ba10e493331f2cfc7643b115379ae47c0fd12f90f7cb842b6646b264054032478884effd7f75d9ab644799e4a3e75f7df319cc0727288963aed40c460335406041a517d3bbb469e2416b4ed1dfcc346d3231a1c73638a8add4d2c40dc2b77d313cda47273000aac2ab2b42b0e724f0040783a78e36664b0d502b56a60dee95b3abeef24beccc0cc0a91d526cba8d7d605a2e8e015653a42a74ffb2c41b272afaf0ec7a5104098af131b290619d60ad45cdce967d6a4c20776965ba0bb47e79214dadb703639e57bea106af1ad55c39adb93fa51382db82a38b1a332075641712d5641135f5dec2b92d70b7f1227e348f16e012f9564f3cbd7797bcb6ab85ec62f0d300e414137e353e0396e4d4b34d61081bdc075efb90e906a9f0b1b1a58d0209f9fca6397a7759f88b4938ca257a5aa6b26fba03b24860b643b5ac32a3414a2c431e069dc2c3c083de047ab1b9a11a6e413b8ee45a93f33bd55106fdf58023c0f25caa2082da8dcc2dc56e7dae287c955f67569559150c2e0cbbd1e8b11115cb6a9150c5c0be5656fed5efeb7469efb88bf1e052ba0b2b1f4458944122efa49209af81d052e6ff2edf8a805d97f0dfaccbdc944e4b8d0a5803a3ebcf4d9506c5c208bc2972b2140bced9b81b60daa6807f27511ce5142544abedcd6849bf45c9853e497ae5e92f4b4378d088434980d648366093a9b034dbbd7c2feab2f511d616e456afaa3c9a41f3c2ba34fda4cbd6769d8b6d51a97d3b33480aefcf241cd1c6fbe921c828145461cebbda51f228f0a7a3c9d5dff8a7c2e915ef5fa6be46103b4282c8b4b20038d5381e4019ca60c2f81ddb6dd2273e9628033c2bb333376f27a7cc44054f13373bb3e0a46231eb0e17ecf679d22e319c656c4aeff970cd50e5ec46f122edbe65791c61a0122ad37ba2ce36c7d80acfa8a18337c838083d319191060dbbd5f03a67689f58f1f1b7965fab7ab7c5acc3d2685fedf48518f1d49cb288d610f10f0c22c7928163900b5e655d5d0abfb0f55d70af2b76439b43e7da7a1fd52d4f5cec8e49b9eba1dc6a71b380053080b07f1ee3af1e4a329d2286c16f290917d5b0302946edee5a06a9c659da9364a7adc5579c3c8a1ee60bbbf6e7fd59a459ec56559be0ef010bd066e755792d8e4d522bd286b8261895dbb13b67ebd0258791ac64aa915f704416d258e0d1adf5b3776edf33a08ea909a1816545425a99049cae52d23f9d719a1fbb16ca5316f85a6d5c59b4275ced838ba3cc7506465f635882e24865658e8a03201af3dbf03bb68846dff481b29acd73209d10118cc9ed3fd77a9949d3424a19aeb14b78a7fe5d68640abae55f49bfdbae7d7947776407ba01e6fc510eb561ee66a31ee934a4182d8341fce9684bb0506a445b4fd3c51db7e59bea6c8781478bdd4711bc70ddabf34aa687e010cdbd1d8b5c2bb0eb04b58700976a66e9bcf14e0ebdff34aea86897acbd68aa0e2c67d18cfc2a374bc4c7284339da6bfbd3684645b655fe3b97ed5d617820ee39f40192ac29d08dde8129846b131454ed7e539388af0e87b52eb2ddd5c12c87e47a35d604c6e0d2a2f8807c1244fa40a4634a488e3229f9187968cdf3f8e93723944adc3d15e80a04a1c159f2c9fe894784fe6659f29d24cd4ce46d366a6cde2891a872252688f71c7518946b98e8c961b0864f3d9b2ca7e14d862d77fcaef54324b439656405068d4378bef43e8c9852d25a0f8c31462b5986931df0ca2e9d08c7eccceb2dc6811b306ba8738b99f6911432050e10cbca0db79ee15797e63f37e8515f23e5c18719a1539bd809f188f6942cfd3c5e492a6bdd1b2614e0d2feff903e1434b28808e8b6e88adc79aef96e7311a704a47572a01016f5c8e00c91050183663052afb6ce6e13c7a81aabdd238e92325d32206aba2e09ad770ce8b0d7e50752820a1073dd7308de2c4647f241aeee7bfb52a553a0ddd99186f15ff67a7cea4b8b1ff6aa98b3859adbd1c537c12fab0e7a619b5e413f91ee97c261ed5916cb6a594f90b557b66c5905e2624069f2f0dd1fa02c9aa3d80c4c3e7d87d7ae8a8b6f52f43f8a6e8e01af40ae14361af17ee36d98dc84533b4eaf1797af683c8342ca9e6f4e0cbb05eb981abeefae88518f9928c0008de23b56ec72d0cf789a65d8539082e00ff76044fecd262ccd36785da3a47e802086dee151fbed41a95f98a9ab424e6fbf65e684d47642126e3dacc4e5fd63a57530ffbef9b8b838447d6e976af59190b434c2e1f303acd1d9ffa1ad1e09a54e6ea5d969f20a513deb2797d66c5df24dd8fb05fd8c6fb127362aca15057aecd42916b977453e6f6891b72663d0ff42b2800b60398a80ab6ea346197ddafd6287d0cfa5b57de3f73ece74d75977e5a79d74a0572de29434067768e05e079b3af19d48d27b708e4d3b8c0aa300ce455cb870d26da138ad8454628e9621aba3413f01b48f617d06730e79c75e4476cd6a672eb8ea9beca88fc060fbc44e3692c3f5ee6d8c604ae523d69d500ad0ca73351d0dcec98692ea2158ad026acb71aa26f9e68ed5eeab267f666a63046eca621633a83d7a9a0966a626aeac5fed7188074e53b83fc7d8add8f4775d051fa5c3c705abe270ebe8ac16194658921678a209067401b107c11896f85acad1cf4b8165f98d19294a594372da74ef97175e072517ebc5a93d9a91e079e530d8320f67b764157b7e3383f7934b696a82caea95b9bd4287155806828ea0f4a55a8be6c1c4777544278b12fb2ac0abcd8aa237fcc72d99418abf519d4a8dcead888fe8580449e065da20229fef903350be4150a6fa36f4485ca222693dd87639bd17ac80480b1147a47b1d193993022395c539a914774e044c1e8ce2b739863d3f03a2dfc8415310660a0ae728c310989153798838c995719f1ef7d05c8a85376786586598236da184ebc241af675cc331533179525675ad349652c9783635e42ad83273e1fa2dc8ec991117d82ae98ba24ed89cba3bbdaac4436292262e33fff38782aea15566fab813c35fb4297837d28495d490f775ce86b4b37144c15c8a97597611e18042088790dec05433f50d0a32ab51f309dd72dec71cd8db6c4c24814b35de01cb39cc65b5a3ccbc6cc00d1c18a6df1e47833afd2de38d7cedfc16afd2d2857124fd00cae46bc0f3e9f51d935702c9641b2a37430030b2b76e61e6720678572272218343dbec0331a52de0c3a5ccb4b76d5191d220a86fdf5d7667e9349156f4e72fb55ff1e6a40e260ee8bf78582acf9b8810a31e6446b5649ef535a62a35945b39e9e1adafd221e7b0cf5fb1102e332e63ab3b1a4dd048c72b4d3c89326ef0dd7c2ab86a84dad59b0a3a16e65faffee3faa2d87fa22bae143a707c97184b089b6c81412b3fbef9e328c87c61a39d2c674763ae33ae3f72a8e35f0b09f527e836fd8609dea2b6d8b75a76c28dd75ac7ea6abd85ae49fcbdb25bcef702ddeed0e7500bfd32293109e8a34265da7241a2d5fd3714101d2da96fb49d17a8100dcf3a090cb1c5f992d9a91a1e654278d12fd055cb4d549e396c26006df50cf5a6494c25acf64b935c667c39439d741424d86687fb667043d6976c75efbdc5e62127c5c5eb770efba0f179dba2da61fb57dddc13e6e1ebd7ba44631eb9d9adb076044916ee22284289c799717fe8e0ea0c40bbd3c03a5d142336e0745ff2bc8e899e0e3e11117a5cf409442f03ee67fe2d88c711804293fc922af78b0b137a2c159f8c45979ffcbdaf33b2aa62dad130258c420bd1b4b864fc2edb031d98d625c09c94f3a8eb5699f9012024efa3eb7c966c5918d425922f7cbd6199896cd5b38d815a7517e1adb51fd67a0d92acae649a664b47032b02f9e69f774e25b599081e9885f347c0a22d8d41cda9f21fb71752abf9cac5bf119eca3c0f13acda3c0d8fcf9811be31c38c8d7f515a30a15d5718ba7792dde845174926bbfd0211774a58af992c13368a7de47693cb6abf9194629772e4707a0dfbb5526402a7d1182cea5ce22e32e910ce3b5c6b8c869b187b81fbe1e2d9cc41f538e589e8deb392482192fc927ca7db8aa960a86091184f8be01a8d7038bc6dcd269e4e057a1598f60cc724314ece7dc093357c516e4915a3e2219a714e90b8f79013f0ff572dac082648462fdd44f4b8a6d1756bc715b28e63985ab1482512f4d5cd386c89b2ae55c2d3bb46a7415349e395e8b46a24133473f0ae8fa03b9464af9d156ccc5493aea36c8df88b9d9b9367e907927253ed9b7ed6078e83eb5a0cb4fd53f0c48f6eec5901b6e58bc84330966783010ba24a4cd609027780b29fedc8f37055205eb4a4a5550f826826b4b407093bedb63535824ddfe2202b89b41c7285ed4378b960ccd2194dd2d6f3ec97cee9f01251f0b1a549485e6c5b749f06dd6914c45cc51b3bffa602a781168c1121fef25fd42abc31cd06167c9498faaebf345bc57f0b05f6bb85f68568ab696a051d48dd68b876c300b8bc0dfe493f4211b16a50e91aef249ea7fabd308a4f22e61e02988f86b3759ac3901c126528727e010fab4ff8ea04eb4fd2021d47c963efd2213ed75b7a5db21bfecdefb78f996bb06f618759f8f2403dc131b125f1f534efea35a3da2e2404c9c5720d7fc863d7846b1ec7a79016d6d8b588505c08e78176fb439bde193ade6498a6e1170388381792b9f7d4852228d6e8b47f363572e68c2afd45c8d32c4bc2939e3dbf75ed68a6b12b8e5ad02e98f5c07460bf9faaab117efb53a16dc699fb6aca55e4a85bf1caa34b74a04886b193cf24369905203af08504c58c9bdc28f5626b02ea01f9793f71eb8536aefe6e84e70c5b8edc639dbecfecc708d1a26bbed0f4bf16dde35e160a831a294010b56e5571911fd2cc9bb8450405cb4e0e0c30293e8f684a9dbe1c0453c4a569719d035a9b9f6f62aef047daee00c9820822c9a44bbd01ceebe57b851893713f0761605c0df5049ac0f366d835a7a35d2c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hceb7418d41348e056c8b48eea39f445545bd62e60cbc1d9cf80180954f901e812805a5b24e2485c680c6744dcd123567adca3d165ba411b4ce56310373291c5a32189622b261c251a185c2c74a0eb408ef99f6c6291834a175f71a0609434bafa427d83fa18b99b327b821481d5150245454aaa04986191e105987716adbff1a8c36a70aad885b7668ba6c8d86de2ea684c297ffac90fa40e64f3a8a34b4126a49365f0776bfdc7e2c3f6edef2df9acd7f39af49132607b15a52d1c8e683a881977b956e96ec534d11376f632e437e1365111a50e1e6f1e4ca7b178512888ee2addc0b2b93f694171680111b870308124fcf8560d8d43fbab63d04ab3e2b26d9f1226841a1d495a428609fdb2972e809f33daa3f42651526e1423608e94ba19350086df8fa27b30d7a58129a5d67db8e55f1d5923b9811cd30aeb2794b396ebe1d7a96b2492641af10cdbda4ec1a51050da0e920d7c1721e64ac733fef0ee3151c760f7509760d6324dad7393c31d69e98f26315d0c61fbb6de048b787de64bab2bfa3cf84307c820298271b0b68fdef47c8616b32e7a7c5166552350424a97e2f18c1349cad529107e8d253da18a423fd0463ff3dd8a38bd03fc4ba363d03b7f41ac5057233297e5813056ed9eda7e6729494ad0f90dbed44f5b10c0ecb06e47b410f6efe4ee8dc071ce9f21baf1421e2d6ebfc514bc08168044ea169804e2329bba6cbfdf78c53c99e7142e6f825a4b775c31a8f3435608994a639f306bc789bde048d6c7a46b88868e2c6c8e7ebaf3b15efefe3e906fcd98c001b616bfd131b1cc714446d1e06a8d0a4225d994a4d76d722a2a72edecfd1ad0d36c7cfcd3a6b352f2ccf209de9ed0ee20323c328f3ce89e53d19b997bb5463fab2ee466ec458c3ef5fbf8d8657fb6716b6dda8710cd1d2aaab40e864b3b0506532327e6420c1ec9661b0731a72f9cf6989944c8aeaa8c8a0fb4ec7442d318b8938a13db94de610b2e4ef8e1b8e60138acc2f4bf56c6ebb0fb4d9c93c327f4d9780deb303dc1e20a3ef6c70782c9f2fb47e0be7f15a44c3ca41d57ac0aa5f039635e947f3144a81d542e3b0322e647a3dfd52979c2183c970378436b0a45fbe7e63bd86cdeaf0ffb4457c3c50f1e70511a09531f30bb224d6da147c5280d161bf88cfc361e0798e5aad25364b22eb2e0dff19428ba0b8ece6d402eb1fe248e20ca0db54bca910196c78ff30739ae9d39ef611786c0b7e1a3dc73e0b7ee872dc2316e9cdf82ae0885296e7ce13b1899b1d99ee098feb75b0ae2849f966f616c7dc0322fd7a86f2a537c28c6e3c5af1523bf77c3ef1df89b945486e6e62c0cf8d78776d676d1435c4b0689ee190b6bca03c951b50c80058c6ab4be8349e994c06c32e0f8c1d037d8c1ccae33b427c14c2d23ea74aa835da32a7a04d400afa606d3113d2c5974d8096a3d371b38a2971b4fe189ecd7732fc596125e3b5ada8019f48278ec3809a4ae829afb2b552b49ea77da5a27994ee6dd242a3ca07782bac2bd03b01e038d7e427bc598e7955468adb56e9242b4f9a638e8c5c52ba5f3a719f6779673fefc7458f90fd6b419dc1e648ae8af3f47d362bd831619ecaaeb9908def1ec072fbf580bf682a9ccd514c8e15fe2d6e5cadcd185df78a86b21c6407de8018a96313bef40aef200ba04e77fff74b2544c138467abf58cfa85853b170e24bba3e22a8a0f16edc4f7613f8e9d08b8df4759d9feb47d7fd5cfb6e534ab8a153a9f09292dc58e8ef862b7bec6c42056b9fb6a5aefb4d106e3a7cc0e9c200548d2b76edfea87b913b413eea5863f67b082b4cf1423ffb6d58daca73ffb241ca30220b42537b9089a3880c98496187551e5dc7fefe98732474868e31aa95a10eba851f81f95f0b9574e67ce5ddfcedaeff09c3bd1ea32c51ba8c616007c0b39d5a79c4370edfa358890aecf17a1cd957cd3763c36a96035f40b91573dae4cb2e7011cc7f4fb55dbe212e6bae5887d86708c4c7dac514279830498ee06e9173b9a1d7c7e38da96e555582d2a65d5735bc96c6d42eda12f5b1e6e0f5ecad505490bf505492b5036eaafc62b30fda59ceca1be2b5df16295846d6c7640455d740c3f072430c39413b5b7e3a2a8555535ceaa4363ccea39777d481b57966060d0120fa4cee96c1c7a61cedc5319aec26691619e5a59f42f91a69832a35d6cdd588847d80a65726c2021622223b23b58d28eca4687f6a4b26581c37be8cdbc78cb239bfe5276e6443196196655c5cb5dc51a465e02fc214885f38a4cb8a42b2524205010f3efcc46744487df06c0afcf98cc62a71972105c41c78020782d411d9074dbd61c7850923dd65b0c4a606d3a09d8bcfaa241fceaf612dca9d32ed883075d9ddfc99f43922f51aa5fcc94f731d4078c9a6f26695b89a375f0ce32ec829d3b5e9fcdbc9868eb89c44397abe2a45962e69db14c8274873c5bd1d3c0daa2926780964d051a0f32347910c6e956d284c04cb568c994bd4548c71cc4075ddd6bf162a3e2d4c3df0c985a6f94dbed213f70edc8f82e130f25a9e0f6095afbd391f15e6af75b772306d9264eccc5a23aad478ea457acff1b73da328d7e51a92199af596afd08da23e8c83f96a267948939b0bddd67f4bbd5869342755c3bd823fb77c6b17bd72bacc25fa78958629ced58aca739357fb9c43b52a1b4f64624d8322cf99ced4b070d67c40b70d5381b6a1ef14363bd262786fa757a1105701aa0a8937a1c484e0ee66c40eb234d6eadb6a2249eb891482fea88ed592c9193ccc55e166672d1d064acea130a9456a19ce864399178902e57721adce967ac6bf6b2ebd4af7a54ab2d816fbaa5e1f7f766a8fba1de872ce4d079e7e7d1e0b203d40b059e3ea7865d0c2dd587155ba419ff7e8381b889d7ed62db9aedd7d4a554def77f70536d0ae7d238c38c819affb770ef783c38eb841c82b5ba32a5c909414e65995d8b0f00c67142d488fb98e54973f10de59fe73dae7f953e8314b0126ae76991bd53babc2780b155d4b3969e22dc18c797bd51c57f81191ec2bd3c58db89f9d3a505b911cc989a82665c30802acd312621bad03be7e5501ed56a50509e1b0c02360e2250f2ff69817252244f576179c7c7ea35b39410b9ad6797e31b6dc329e1060f37b9325b794ab9fd86b738a6f91dccc92efed815528d9752c7dd726c27a8599dfa71164c3ad627a6c5cb8db377b2dbebab1f7b0c78accc322d9052e8f8757f51c1532e660fafae7d34baf023a87ff895bbd62988653ab8906dd3c956ad9e66001c95013846f7546cead565b607b141518e8fa70d86a2aa88cb6223f39692e3babe16d9d398e48fb00fdf6ee23cb3d84e3b2f2abb75d0cbfadcfa0f67974ab21df92752eb40f03d040e1ccdeeace6eb4268bff115303a08bf1f6b732eca46a592bcdead937c133cc7e8aa2af0561cebb39b1fa20df8cea5f971a479acaaff82bd26110c33e9c113d9e099fd892185122e3b70165bf0bc304539bf9602d7103a883b00fe546ea4987236aea80342852d57e34ac27fbfb256afa6b2758f96db8c6f93ce2f459fad8305e4c32f6f5722f4fc0aeccf65a6f62e12cb1de17c4b5ee79d7d74833a9ff439c848195c3e886f6647050bfcc2b60b8f57db21fc7d6f184200e78937a947c5e294c634d7b1a55e250bc6450eae52996ed3d2878c2167431465a62d7467dce6554e61bd26d11576f1644e6a78663aaa0410d739d67becbb44b0f9748f1ca48062e501501caa584ec724a0b7a484550ef1b1f965927f541f97ced317462b24b00390d9cc374cba9bf8748c8b825dc31a4003a87c94b7c465f6f16789d05947c9881c95beed1b0d48aa38c7625d7aa92dac83fa60add0493f7c7af07515f03707c4acf0b125bdf8012c11ad7976c0a65f3a0e9c17446db9fef261f6972de352e65c60daabf1d8c0300dbe71d1d376953441754faf553533956733cd04c79364cc1eee6f645f6d8e3f9c7f0e71ac75cc22225262df7e986b6bb9cc2645bf93a0b9efc833fbc8807598792203df2054af53634ba52adf552c31e261e798dbc1f3bc4544d8ab725ebef4b362e14b0813f570f1debf9afc718b59ece10df77ff64c6e096724e46a214c839eeed3c020ca61314322962c17347afb39e8140b9722a50bd782e189607adf79ff009e9bf6d9a6fef7099f7be0e1fb2bd4de33b7b2801fb0be78dbbb1264ad2900294a179a522afd58962c77f5cfa4fabe065c488f732211f0f134026a41d3060869af5b689799d347b6579f9434714b18369d2d8902cf1b32a698d64cacb5d46dc14f212d20f2f642e0305bf454c15302c6cab42cc8fba146ab29ff5f978fe444d8240f0c56389df54b316d5aad334972998d2da67c513a548ac902a819888b1151bca4b61513161dca0d8ad4fbd949c34fbe74cce24c2435b2bcd913add42b1da5c791247af811211e1cbeef25fe85fca1139a86f2dd7c6bf2e12f6491b12be6ba72cf9b921ccab7ee70f7c5a41b5e9cdf065830a73e1758630a25e5b7a10524e99e0d82e281ddb745918c5b6463d3f6926a9d86eb65f0a1f04c6901b38b4ffc030d2012ff4ac45357f0d2bdd4e4c45c338f8f0851527349cce9da20300d1e565c056dc3032b9293de87a61d08bf0080ec7656f3be16bb65bd9fa1e85b5a7a64a6d3e3144330f4fd30ae56f323caba839359db6f850578da2847d96591baa512f04deca95e1a66f6a74c307a92352f5d951b2db4cbfcbdfc45f83bb1756441711170a79bad5aaa28c72d5ea6d9e21fc36e8a6b81b42e94000760a36816b7b37ee247c5b9737d7ed314ede1dc2fc7fed3d030a73c85cbe11a48f95444ed3793b8071e56d60213d228cbc9279c3715106f6a11c8d6f6cef670e7cfc9330ec05fa4536a90a16b9d06e474a6fa72a272a0018de84f5bf39c682f48ad34391064f7de3c75f6c03602dd9a366060715ded6557228cac7ca4de3f5cc80f2dfb0b7923f4ec2510aafc9f0d5306ba8c3cfed5293841583b459b5ad3605724b1d92565b01b8a5f4d5e045c8dcad836d607794ed5186ab601d1e4945e4ffff9dd3e2b344ceb28ff0224b568b3c67db49106d33110ab81a54a6c43205864a4e8b967db950c472629995c8bc1d825cff5feff5b38a5c84ff4423d916f7ad12e8c1fc88f8bb4cfec13bbb7f57c3b844abbb4054510d8e1ba6da86dc1b33c74362492c44878b55a0ff9bf547ac6bffe191ecf24cf47cc7f9c677b1788923a6116144230f650bab10e4731ffee829aaf364fbd8e8de25d11f26a1a130e3f9c078d565ba44ab584f2d6c6578c319f8670be1961a76b8125e4d4bacf3b35a082fe5916a150ae1caa10da5bfd96021efb91fd880c1b834cd6dc3abaef1663b8ad49ede764ab272ee971c55cf5e96901373acfac1abb9d805fe486a5417019d455756a68d6f474e601062cf906d429f8823ade74c379de252deac40a0d6795bf9701f9707683f38c1bbf530f20e3d91c6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hfff6246b3e8f00f269609381c4d48925a46bc777bce370a95487e6f5be8663069c500f697ad9a0000e7eeec8ef9744cef601b4f5b2b6cf205e9c67387d8b7e15edf595b4551a2ccab138b91fe55ded78d99cdf90941a663e95972ec4ec207269171484b620fb7267fae78c47232abda20a352a9a4c570df1d0799670513e0a36c873b40fcaaa04372653f0c29188d769b5f4ec5c708527a4cc9f2ba41b860baea99925134819d6eb176d068eecda667d5ebac46a5f0a4d4fff703db930c43e5f01ff2750162d3173d76de939dcd09724d918560522a5aa4af5a0bae49cee6658ed5bb7d150e8480e07af1368244ba0ea99e09d8b1eb8ceb65367cd1a2952ce485205a83d7ec35275c67b49baec17fec7ab268c7aaa8612cc17337169e273e8d57cf01236f80b17a537d2369c1a610ad37fd2a2020d5e6aa843be454c93dffe33ddd4f84054e52d31c90f85739b82b7ece16803f576f167538a2c8d312bf6961abbee34f671bcf753337c21a97c3616b2910785005cf17c6a63598017ebde8366945a1e1b027286e24094c3158f1cf97a91264496f0bb0f2aa9034b77322c1f77933387d633572e390e84a9ec6096f1e2507e2ce65cdd931bddd27e3a2960d5ed618b227019b146ba2c85d1a667d956bb69a56fc5914493c5564b226117c568fcc0749e7a52837f087873a2cc165e61fbafc7206e4ccb01b0696d7c7382f73f57304e780e4f91fce034868f2e5ecc75a6fc402ab0ced170dea2b4df1fc381e42e1066eecaf89947940d4dffe66003d73ff92a8ca0285810ca3da2ea17ce86397035b536fe2939bee54bd34c752d807585985ce09dca3733a40a68d128454e93a0dbcd7ba326cdbe5667f43bafd922538cc8adce67ed948cc359a758b04792f742b80c842ea07cc8a9213034ed3939fc1b276d401d01d8cdfe8c343bfcb22af905d77c469824a798e97e78465673c296c0f2c29d68ccd9c4c2efd334a240f553cd2834c5336bc3520704cac1ecc6605082e174167efaf62d430e81bd29c8103ec3e29b5840858c3c003dc3b971c9eac6de660bbfa5eac7efa5eea6ac7261b9552dbd1c4713e2007e225be02e8703fd7c3ce547ef693dda3c9e72ceaf88909996c2470ecc8a2f6fb32b752cf47381d58ebb6bf203076ca3e3aca3391747843f0e3f0c843d70ecd15fbc09e1810c5a74e3c7328942ae5a0cca454bd222333165176489d63609635e8e99455bfcb8e163ae998abca272d9ea924b80754c3da8d63d8f09b503c36b7e9c37148c566725c966ae4d601d57ec0df8d8465f7b4186bd29237361994041d80c9b7bb261b4436158d8caa281651c6d63a6e20863d4f5c21fd4c2cc5bb9b7bd4cef7985e7f9442b196c68a61a06b2c6410ec4215c38cc87587ed1acdb618992589e46a14a6f0a56cfd6360538aab9c421d0ba03e78802300c027b64d66e94f311b986a36790eb389643cb508fe39303b35642fd30d1c3ffd888242f5f882143699725219cf853983302f84abb9d2b3d3a7eba159f3339eade612e96ba51f37c88b823f34155115872294d907d500e14f751c8173e4b19ad95dae4b13559ff70513438d9cc212d452d88f9fa3fee4b008ae56203ae2ed0c80995a4a08fafc32a865ad5fc85ebee058a624f8bbef79da34639e808e6f88e869ed61a527cfe575b699f658b96fc78e1064e9779b902d4b246967ebaec01be9832a3c19fdbf029c4537558651e38c8986676dc27ab337f4ac5b288f85f3645f34cb30578784ee31279a303ff47e7cf80b33cc97075e4cfed576eb6874d33974866a3b3c31c95fc9d76304e0d4b0f75930c9b62a0a31f9102aae370458d4f13a5a08519761e6f2bfa26b01e51a0384265af8d64de8255834efbe146aed74b7ae7ef6f72b7362e5aebef80e78979bfc9a147e44f605b306cfb6d488101b5df26bebe0b852448ab72d7d2707c3577fef2b91a022db4eb92ce07f156a87b613e2a531aab026d232096e90aaff4a21ddf586b2140a029becefc0dfd8518abdddc933c887357d824010454a5d277888da3f2e5a55214c9cacef6392156103eab0e14178a7afaa4232c6c73f4c09d6d7cbc71f4c7c7a65b7de8899cf8e9eddbb30de20318c981d323323769524f4b5bb4f119850ad3fe3c95b6b4f9900fa6d515b42e5954ad9181b4aa7984932fd6cf834d5448e8f32e62979426f71b9681a7f27e97917294b2b2fc0f199fde2c82f59d92775fc03d9748edc31486c42450eac871b865f2efd3daea773fe05a977af1db05d940faa764ce297f2a462adbd080539106a050d2125f8bb38fb164ead6e669391f517ca1c4d8aa4a53f00a47c0e6789ef7080aa96319618e9a2c0fa82949f936dbfcfc74350c674321e133580ce951e369c9256219a4b8ca26b5bea3941a7cba2ea4f1a6326b049905cd1916914254c11747ecc8d0a416df3719e1469c6dee4b2e7426c50d1ae4ef3d818d49d20a553e0717e402caad1108d0f209616a07306769fb912b4e63cd31e3b37a3150f04dd8e0924001135c63bf745928ae2c155d59f2437ac5d0dca35d9974685b0dcffebd4813e19f522cf7a7c412ca1c2e2cae4ce7df1fcfb6883ba3f6726fe399fdc3e75c6edeead5e57a94a097a8af3feaf2c8e3ebfc711cbef098e6e6adfe9d45ab29df2340d8c9cb0a70b37538edfe26558ff6163c46fb4470bcecd1952bea6d53531d4079fce57f424a1d81c9e6ca0b2fe7c4773c09acf50ba55a036784b287dbe85ea1a54011013de8178daf44f9ff22f8282c31d8b5acbe0d50fcd8ba7f9609606668aff33161c504ee27b9baaa4539fb3effe70e3e76b55ddd18abbc4fece635c8b61c7a8e94919867f8a3f72fb2c33122eff1cec7cbf27efe2163471cb56a32cad38bce401ca46201645946b5d6bdb4d1bb995863f3e11c0e94886eee0ad6fd175aff15ab3b21ebf96e98a1159cf9d2f434f0aacf41811e7e3df2ec0ead16552941d536ac556904b443bc67337984d4464f07ec91195547e6b9df2b8666f7706649391093ce67216ad780b1451b2a2ed73a262b70bbed2c8549dd1d28f8d4e96f8fd23766d13975fe1cb477f97d592be8ea60b833a4e98698504dbddd7b79ada6c545c4872e9906a69a1752aaa191ffe67ac6797068011426f74475d7de1b465397ba5cfda6a5ce0e3456b5197cf94b5fb092139134922f803b69ea9868ef6a1d94b1f846283218036c1d11073a2f5fea659d4c7affae16f58990df484b3d744b9505886c9a4ea52c7b9d7a547e459546acb52c6c4dd9b270212ba477282743ecd5a49248ab95ef8cfd0d06f81b819bca070a71e8dcbf933087fdfced557ef542cf14184b69d18eabf30c4366b042ec1d6f5b203342f0769ef9b4014e949368e30b2970dc45da55a3fe34cd9bd4816108f7da0a78d021077554b9a1c444012ea4035644821e74030829f3f2c13acb80a4f185124f9a81cc9bd3e3310a2eedbeb788f49fc9b90e5d71394dd2813f1fe6e30df93904ec820ac837837a9c148b60a0e3e9bfeb9062588288b6a6f7e23967e3199404c1c90de1491775373586119fd59e0c9d8ccba1d76a29e35e7ed6aece807726bf4d2701c6e0cc000d3993543b7cb01a61683d29dbf43445c2b947c7ee496bbf0a884b48766e0341a4a700ae0d14d0ad5406aaedcf5afdb701ad81d032b7151ee4bca1508eb2cf6a655c4d0582085fae38464ccf552c23751afbdc1aaf62d37b0b8c72fb91637fc9c56f363220d9a2764ae053bb428ac0a5f98ed0e0dc678926ce239527962fc80664b47bfa831e5ef537ec364695bc804dcd2b526b7bffee498d4df8bf413176dd074fc8068801030e7d86603a51590da10fbb9642c89ab21917712dbbe7628b7696a734485c3fdacec9285678a6e970f9371b620c29b7e7b9622c9d6f3ae42ba340b836c222b36a7e22054f90a503d243d114831a6903d05101b22823c8797224122552ae8dfafe8ae7baf354594dbe99cf0076bb876212b444459c6d1852c5900bcc3a9ce37a5d7ab43bedd7f3fdf0cf3b58690e538918b5b421a60d8eca6c2024a8fc12972fe0ac9d5deb46fb124dcfa67a60eadf2566d02c731f1bb8c07a536d67284279b3b61ef1fbcaa4fd423a09f1abc6d73e9bfd1f20d398212a35531d3dea7c8e5cbd1e2afaabec0006a8ae61da30e36b9cbd7ba34e9f97e988d8ac95d5bcfadec24fa22aec144aa3afb5e93167df6221c1f19fc8b5e14780b13f634730bda5abc19c7f0103ab4019d1b86dc51ab67d3dd844c57b09a359b7ff9df71305c02fd187567acbeec97c77d01aa24c614654eb6841ce7a59c970e5eead877e34bf94bf89ebd830369e75b7376805999e723a08a158aefbbe72b190e09662fdc5fb1ea76f67651b0e444d91b8fe8de265466ee31180fcf6c27df55ab6c885a60f3d0194e32c770f96ef0678b5cda4e4fcf65e3f133049e0ec3ba9fcaf495929220a9e73e74718060ed45ed7b5452169d21fda5081a7839aaf5be6b59257fa188cba76889dec9316a58ee4e9cfb19e1e5c8ebd666b95f761dca559cae2b778b652606e7b146c163f23ef84cf4db259c7634148884719ac0f619bd5264d9f6da2aa6647c65e662f0735677ee29bb43b93a3bf1269f09371de8c21c0baf56bd5c00dac9cc684f2323000ad5c5aa2122f3f3151e573c70fee63adea5dfcf2d8dd19251291a86417dbc9762ab0ce7c08bbba06671cb199e224478d56a70a63731a9df2852a19fc1334f08cf25fad4aa877c7fa26f33677ac9641c6511628e412e34c9be1c459bd5066e0ef26b1cbbb0ea67b2dc70f07e7d7d35edc54574469d022be8735c99c65c5bab53da8bcd7f75ed18de977a6bd4b3d43a03b9dd742c674337235e1f0764349fb4c7c4ec10d5fb0cbcf9f9f9735589b1710a84b35e325f42fac990e29bbaacb7ac55f585a6cb9266e59b9c03a118af408a98d62f522c62ca9eda4001f2bc2dcf19f7a8484909aa18f1d8968d90e2c27cf2edfa12f4e37263d551da435306c3f32856c162fc1c93a8d6edaac5bcb46ed66be9584b2d8e5b2232910e2782cee7f526cdf9d657a85a5a633dc1b0e5333c769318e81d8c4250339afc17522c3901ac9ecb256a44c72f9f9dbceae551d8bba2db5de14bb7e3c6d7bf5bdc1bc6b31edb61d0f4e019e73e13e95705ba154c3c9132c7a4b50b6bd9a0bb1915fc1356768753c069de3b9763380b09b8480b2b11d7e3a2b6f70538af62943294919b3585bc90522b0bd9eb79d6a3980bb7112ae86a5e0d9a2acca5deb809feba266c6560064a472f4f3bcf654dfb099319d58e3465006de7e9ba49c3df2d82a33dec57cb0e09af6b1ec6f19f30afb09452fc440d62a3b1d1b720081ef85ce340135e6a950bd8a852d4429d17bcac929900045d87e782f28f5b7cc544339ef7e8920fdcc59c0539b1641a0b2e1f8120c5e5cf5fd5f0d1a29ae1503df6dfcb9c639898d89184529fe0678954636d4ae3a9abaffbb14757839;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3f533916ee4676b96fdeb23776a317f033956536bcff1264c81ac1f54bfad0c430a09de3a7df25c4f4e157a5182b6754bc60b85200545b5bb31482033f7e5559d386aef8b6d59849d6ac9ea18432f0d80a4468a1c3d50de5eac95d248b7273403c996fafbc8a01d4ea65eff35a0c368a11dcebe922322d7b0ab248f76ba33d274bdcc7916ac41954d9d43c14b1ce282cf6beb372afd48315588f16b7a6219e40537f29155adfc1aa751e9a32c732647ae0bf4e4984d6b49d88d1f0e9d87e3e33df98feba788b6c40317edf81a0bd593b38c08928849c72e09ba68ae6a4646a1b05669e2000962da3fb644e51da52c00c5865911e7e99ee4c977850a175968292bd91e26e610be730baa4acd5a02b87fb1ef9043a48ebabfd30324a2aa9dbcef5ea309a10118ce7652571496277bbd31519607777aa27834d756dafb4792cb980cb14ea0edbf6cf1cc867556d1b43f2efdfb8b634390e2c1ea275e0bcb3fe113275993981b08ad05fc48d8f934e102aa467497dcf3336d5f00ae42ecbd5d5faa357fc810f713e208e310cd7e032925394f301fe937bb6472fe6af9e3f5d931129bdb6d6867d7ab30ed5df79a2afabd8cf37f4cca20788aad011d5a23eb2594a23a7051de92076db7e5d5df9668804f7127c0b7b06587423ee643e5eac8253bfb13e3653a639c1c520305f38a36e535dd4d063836dd226b86f5993195d67b095f851452ba1f640dd6b75432d7e7bb0e16d36c9e3adc206525b102c7fa2f2134257972b56d7c91781818fff895eb6ddc776088aa19829c89dc658cc3ec7d4fd48ef3e688de3d95db4a13e7ebda85aeffe2d451df9d78de81fb75289cad3fd19bd31eb69fff1e9e48e8796f6ea558d7c5873fddc20f0b3a700f717b23378923a493c40c58d441c7a8076550647948cdd2d7aa0ad10bf334ed0132e0b651d3969588490ddd4140bb30aaafc6b4601641e155e2a885bf83c7ed7a79d8f6c5eb02750e19d903e60a4149ca8b7e26532d68a2e1169bd3a21894784b3492080b79188a62261e7096f06203f2d402705d8525c55f705d1115215505c81db10fe7403fc66e32629ca4d47469bd003de0ede5c0bd624a03f2c75d220588d8a9693dfccd7c6e0277a76b439c9ea47a8d545a80d2b474206a718fc39c7addec0916c6c656cd6f087d7ce79fa392d6c6249c409fe5f97c8338a3d0769183ec281540c652edabaddac42c37ed5f296104814fe741ca766d77f77ab85bf1826113ff0053e95ae7dea6ba3fec2ae563603945db2614bfe7369546e8c2eb18a029d44b68c0bf01929910e5bb711c6fe09da21ba52ec459f26df9c2783afc2a3f88a62d7fd00729b0f57e411f7225841af941fd503aed25479aee0f22a85416b90cd51387e0e512fab6a41b8afcd78c11715dbe837805939f27849f6ba96d1c461e79e590bf77f34c66276816d6865ba8b2a415190b8a206888b4bcab3597566d2450125ab4c99d9f3722d34c490e822f08d24264a8e913c562314284bd58bff49d1fd4639f495482f205f4c26d763f455c154d40213e422096752bb869a6fe6a35eda7004a610965dc85800d01bc8d97e27637cd4f831722148c141c77ec046dde6125ab218d3e06004e75e9a07aff9014cae28d75a6f95e32f9856ec43d17a9c98c0eb1b51f7add387cc736fe5612a392a57f9816082c3bc7b7d90de8cc19a9663b2e8996e400664688bd5927484dce20a947271bbda7be51363213be4910868d303f5c7d4331139662814436edc764340ecb05c05ab41ef110b65e913b477dd5baab6311355516be03cc52b891d448d50440b2b42de065abc70ac5110c29a1873fa98d7cbad76f01bdb148d3c414cd5d1d91163263003d6c470554374c8ced1bc0051ee6ac7c3ad7355e535257bf834ce7af6406dd90ceafa601965fbe0037db7a4979f17441923f07737b8737a8c77c235e1b24758ee2c3717e7b38ed2d18030b42b75623f526ba8e92e8de72ae76904ec669402d0fd82ec8d151cddfb0fc0a8768061562c6fddfbec928cd7138f2aa3e83ed53f2dac1a47cc2b1adfc0cc0331b0ad4ecb9586674435bbf44cb1be56d2319b001f1500478b60ccd5ff93cc1b7b2d4ab080dcc9625d2fa65fa06103511c8955ea529ee13ba7c288fa10850909e5e714b064dca5171a20e16563c320c2add22570e5964600a6e5156d500765c8bc2ad7f08881188c1e9ff5f9aafaf81e260ec7771c0e36b3e23161c1164ec09fd180b9fae91db169e9de8fa85b13fc1d8bbf18972f85413aa5a60e81c7f2d89075cb1c53284076c229eb7e94f6601641b4fd83b8b78f2ed9e073adc1d3c9500df63ba2652580745d542325b060853fd8d9e6716d857a89df748ee59ef02656e5974a34d73f7e1f9117700b47a6a7e341ed537b085bab9b6e3f2bc145139ea7bc7d7a481250871b8dd8e540777005fe05c1efe126fc7b286ce6f464237585ce678b67eab3930524b9892126c0f4d5dd2611868016afaa58368b56f1bbf5693a4b627994e56f1a1783dd7b6266c4340f10672076db06f789a46e5a436526cf4432bfa286ec2a72cd8e64ccb83b2245828eb55f048a8e083d736aa8333b4f3990e06b8fbfc0f3ff5e32fa5551bfc756b259d2b21848e8a46e2f76872b9014300c51733d132fb4e7cd2cb6ee301d7767a09e58056dab9b5f6c2a61e37d9be6ffad72b4ba16a0f774de0d6359181e9a6394a87bf9c8bf0773abfb14f78cf5f912769b364ab4df6a6b546b750e5c8baebef41cd9523ec20485893f5e712fb918de0ba52d9ca1e5b23401385200a22dae1dc70644b4495d399d9a593d1b10667cf9870c43a9e0e78fbc9e722bf3b1c59e13e0f56c9ff5fc955e2ada6a98fcc348789ffa638e4e7f890e778dd6c51272ca21af99909ded4573bce40668e3598b8101e8d2f5011826dd6ab0e81addc5ea0eae7900630223cb5b66882327ffa71cd5a3b8288a845a4227a6e64143f983b596e6fb0fac85de5b2d84040e18b7b4f610368b585121f5cca738eb1a4878e7fd553cdc50b03045cf66556af9c2b99f1ace1535371bc237a7f4dfb71c392f042b2cee5a2881f1db11a717b1c945117670ad1552c07315140dee439d36bb63d9ecdf81f8078abe9f9d39ff3366aeba6af2314e38e147a7ee7675faf5c39eebcd1b4b5f2f70e63085c1d5d34a59c974ef5e6a9999e5ecd60f3a8b474d4e994cdb3ddc627346cfaf8f764e847c327f1771b01f373900dd5f088706c5f079758c64e25e03809934f011c2d558d00525b80b9f822d1291182e102206ff8d4941e9b95bb7562ddb8ae2d495fadba2c219cfa73c3e684ffda293681521d30b7ae3b8f89d38424166e4ca54dd31da00b5b7bb49fe81d9cedcf6a6697f0b33fe10ff69a36174d60f51e93e1252407f37ee257dfd36f6bfce0af31fe78c01a297a317147dff784bfd912b178d1cdf392cbb9ad940d346097fe280d654d40e6903141f2a469047a2859e6999026c9c6d40f5aaf7cf31dd6208c2267220a4f45cb98a140e8932195194c289d8c601debf9bf47d0f05c8f8768b180f20dd8147a489964571015cebcfcc2e1ff8735c4bbd9a7e827dc35da0eaac56ae74def98d3244e3c6e1bbb76506624f23fc92bb9ec7f469cc2aae5f5fa1f6c61bd86675d5e88b08dda431bc369eb8bdc4a9f25aacafc395005b1b642a09df29c8be43c257e3dcbaae47331fd19b4a36ba4ffd17ca6512f7774d9f078f8a3c443f50f537a3ca676c4767ede87f1169076d038d5657dacade1bff1dde1e478f4f21a4b97ea8a08769c6d5f4c4c27b3b52ae5973d913c29e9f5e6f71e8e58ad1f80968e5a5739695a87f52446a53896880b7bb12bc690b85de178f67debeec6dae13f0293ad6da8bfe3145de5bbe9675a9faa09bbb9312d137648a1bd27b8ba1cd772e4f11ba87a7e9d5bf06801d8b3d5538f6586049bd3d04d035d39ded99f7744b6c36f6c6286b3d04e294a72c99d9732e2eb91c10607b086faf06cf2c6bd8791d46cc447b3693ed694b580eb82e05077e2462d6a5725b6356a243d21be6b786ca5ecb6e1f0709bbd9d01a2d7350f8e340e8ed8f006799d9df004c1c766fb4cdc158ca1bedf763b3144daf44883cfe689822c98a17b1664f60242216c736768d78c8eea3f1f3149f75e8b5fd11b93898d038310a5d0b225dad870bc858721283816efd2298a656465a05fa58304b0d22a308a816fba7ef06e9e32e04de2cdc523f50e5ba34ceb382ea048a3f767cba21367b44882c04b20bd281b1233e3669ac5ba27e0bcb12ae71c9dab9938c2a027954c021814a3f40b4fdfcd0701808286f98f6d79475b5347dbbd728913ffeaf1f54d85ad09ea2f44b50261b3b9d9f8da0386a7f9ded5d0195a9ce57e41e41f276706e7df704bdd6e09cc24c731923b1f00e6ab7f00239d25fe32f13543ef130d83ffe21a7683ec48d3af31349784fc76feca249fc679c9aef3f550af4c0f5cace9537b25942d0c8100de6019492c72a5c587b5c74c6106270fa384b3fd3c89d73b483108c7c61a9869e4a0b2b07f323e0d5da674d253a7f6164e4f7e707d2ebf04fdb504a8ee1e009276b87a098a28b0b7c961da31ffb37c8fc2ac94fb0aaef456c63dde24dd91fc912d7f27bbe8a82186d37798f7e07872615436395f594ea673a223f300856c3b42631b5dcf2d07b1460a3d5a6aba85cd2c5feb0ae31977a918a178f501da59d9a2dd82234e8b583625e70a17061dd244f3de175e0049842e6b9b5c08b8b581717971b0aaed5415ffe890458ef31efd501aaebf9a5adad8c7c40b2ae9c82a1e3beafd335693887ea579d1590afc7412c1a9cffa84fa620ad68b06e5512dd425d48818514d527ca824925130b936e4a21491eb33d0568836c390cf474ad0ae1c1ac9bd7df112f2105232090b70d7d5bd2e8d5bd55636d834e19184f6e875365ff530102459397415152aa5e111f233b4312bc9522cb75543f8b135f7be6571c544f9116e02af220d4ba65b34020ce64fbdbfcfa9b509861579284e7fec981f549a0da53a231b8aae1d68b1d19496664765ca3195bbeccf96517c3e5bd5a5fdfa4f28ab56eff70d07f19c2b717294e0b9a6e10027930d37bc3ce2543f19b72e6dc2afc6251bde7a00e9768e199c69d1312735405763005b06aab25248f6400bffcbe3fae86f9d3bc36bca0c6a641d7de69e071921678bcb0c9ff47d94933a63f282c7c763356f86865df1464c1d545e80cfea11067968ac445002ba82db4b6aeee1f0772773ae62afaf270b2aaf313dd1b0fa0026512e38dc0728e265777f6024cf9bcac79a1c929443203b1c46bbb1cae259b06818dc3fc05224ef752647908c0377f3d682db1721998b44abe191f6446a4b5ae77d35daea94f7da1660b5fb4632b1d84227575dd6ff6fd9b5e7739c58868ec5769450b5cc577042d979d8663bd0d929dab4b42e7ce6ba314d6008316fdb2822bfd11bb3fcd432a4716efc79ee2c2d6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hd617d446dc4825fb956860a9a460e6a7f0167c872e34930a4ca7d4e99e0036faae0aaed5c0755863d58f63838bad0b0c10a9136c0d9f2eb3cbe050038efd5f6bbced4341493367dc3bc9d9bce92f478b132e040d092db1f882962b072f4d1c48e3dffd6effaa09449d7663a71c2edb32d23069a1d619d803625ffd113b8b5daeeb8c8b09a64fc140990484478d1c4ce39fd236b37095b2c3462ba9a83919fd9f16b1d7d7ce3785df27dc0887bbeeab1c77d96edf0e778926ffb7617aea7ddda2afff420f3fe134ac487be849cac21fffbc40e29557b5d5fe29349dc1f26bb945c5a214d592af361ce680f733829ffc79aee3bc1cf4978704bfba259033b4bc6a0e792c7c2b8d51f5b646bd27e1e08c855a4cc5a9ba29ce3c4fd5e3933505593091366137e4cd5d0e4ac0960d1df9ff39c567cdd21b1348d5921d5e5c62e9c7789265f2a3e8d6b3e9cec34f8cd32d8f31e51f4c170f2fcc31b86477a2f14c0c5becc88bdbbdd63239263f6eaec1a605b10c235d99710c7758ed6f0196d101ef5674ab6c97c8090731051fcc1df3a7cafa6a5135e1847dbb9c4e77befd7fc6246d087a4dfc70663b187a5122bb3ba1a0e38a939f6473805d3f30a4562b9a93b990aaf04234f3735f008989e5ca63ba368be07c3916b166f166ea2aeca512f433e7d62cffb54d0e608c7ad50be03671f889963a42f299aec2a01f95aad357953408e6fd7864789a6e889e0f926347d0202fc17e20bb4588f6a583f0643e3c74c77afa0cd50481ae26c6d321ec31513589b5af13cecd7cd7251b37aeff08e6722c2d10b32f8739d0d097335b87bd0b24e040ce4c2d338ed275c3ca5762d3fe7eb9ba40b6a93ab7b036a51c4c0252441f0e8030031910efa659bb7cf055dbdea18855a6eac1bab235281e841b20d889d14ffea4888d638ccbce220094901fb61fe894b778f288a957b27b0d78f7068bd011f285602caa2b4adb01c143716381b11b222ddc7c0bce887d5f7f6dc72a391cc79cb1c5e72f3174666e88b785554c977e52cb29829792468b7bb34916b94492a06c65a914b0cae00896330c7d61a14985b9a8041799fc434cd51833c5f8dff9313e942e453b86e7800e85677691eb14f562ae49d2cc7728e2e323e0f81c742c376692d0102d9942a165394c75880b78507e61c6cb122b3822f9fb468b43ff74f61d8b899c78eadc8e4e9cc2dec8f92ede4be6bffdad1e2980520ddbbad9017ce96c920f231ed88a53995a96c3aa867d9c867a17519e03e87138c49724a736b999dda7ecea9f0053d04fd2fec1f85065c9450beea86a58a91d231e1b2695002d27f522de21648c2373f31f2f7e1c0f0b55dc8178804e3d8a86981da47042e611fadf17a706cbf0d16994a10a2737a5565127a527e8811e17adb4af42bf3a1b03e33679792273442ef8980dc19dc40b548bc6af0d39beb074b20e086491b74c2137b1d3426c5076ca2afce443f2ee6fac5f2e4dc5e92fc4835040e21ee5475ab32b96d38d72d1f89c9c22f106818e6c9bd7a9c905b4d69da3f1d34ab1abaa38085f96cc25dff6149b2104037356b54053e8001474f34efadb54e25ef1a6f5d5de245acc6712d0392b064527ddde96a21e3b6968edc4ea3a20354d2b5ce287bcfd0a74d2841e428c27dd3e4b8851532ff872b369c51a47f1090945c5d38dc60454e421655e5993b78219a77f0995aeae430beccdf03f170ea44a46509bbf663e2fa3157cde4d881421188c4dfa5b9ee8602b37bde177b5283bdec279d49dfabff1e5735675fad82d4a13d69e9e6f3cbab90e832cfcb0430f49966254abe87ae420dedfe9b7fff2d045027ee7ad57229a34e337f268454d7e6dcfd5e88f92ab994beacec8a9df3b955ad62ddb3aa96aad2376c34e8d3b67b4bf771f3d205dcfa19c6aa42e425112f2d95ba9e924942543e69c59568cc8aa415950dd9ac9b0e394751c9b3679f01551dc173d6bb4f64a66407cedd9f24f6bac27833f58cba6411e5bbd34366d38bb2c0117a0c6323dce4073547817645e020a53da59a6415fd553e08df0509ac2f46f7e304fcb5dfd80097140ee9f5089c846667a0604470d1fbd96376afc7bb4d98154ce618480873baabd70bdd159acd5132610260bccc070307a78f3045dd9fbf3fafcc79af0cc9994fc0c681cad14948b41ed3bed2e8510c1fcf620fc781986208feadb6ed2cb897fe8e7cb8d2a81feb8b6d77c41a79c22cb5b9169708a6e251079a393d84351a7f9851220da8fcb70d1d5bfd339a16fadde0aa560d7cb2e674d370ddeb9085fc1a3a4cf4bf69affd3043e854a35d19ba764084352f503e6ef7c7ae49a491a8ed652e9d5b3afff362854093797b4fc9ddbca7148dc9cc6a67cb3961d2bc2d323e0df5ae85d0a468b2821dd2173baf8fad0cef29608bb52a11e9027940b7735b5a20f0356d7a4cb3bc56243bd2c5afb640d959c72e0ff3e39d55d19d820f2c4006945060a6f19b328789a2197887e7bd31a32260a21414d69b0b68e8d4545e72aeb710570770926eba1cc49cad1498431f059c4d22fa891b0067761668a9f91c32126f604796906886dcd7b4f258bf20c7712c0495d394ed165bc6cd62382f46e2a3d9ddb9d7c6bd5f668488093fb1e8595bf9e2e90d05c559acac371d9c1c5ce43213f95a2f00d4136cea6abb5348efd308ead544f64eba7ae5fa3d46d8ff36e3d7732580c67ab6e4b3c1678a285b5cf05354cdaea6de32d69003c70eeabc1fdbca4ac0e1512799cf6a51f8f280df34c9250745f584b8ba8057f292a2094b27c29d65741c9a8f7c0f9c6dbc00edb963670b5f3776112e0c82f94f1882fcbd776080b672df96a5eb8afb34111f1d2162bf16162f67932d578a12aff785af5c129adb6eb6a55e82c57608164719bc98206e38b67606754a22d1f3acdafc76b8e7d8d3d1dce4842effbae67d7abb325cf1c4d90626b22b44e892ce6badd54b129a60175900f52607d9321152292b273ad4d41ad81fdc697a39fc871fc75b298a2313945553fc29c2fee47eff88ce2f1ab22c9cfdc2130430bfcc1af81217d19a1a7f57fc8b4df09b9a0044a50b5fdeb4e672fba69129423746d140fc5bc4b06b5f77b378ff8eeb255651440185bcbefffc08c8bb9ce7d2b1be6945f90f7e70453c5450dbd0cab65ee3b97b88925cc3cde77539b0e0af93742871abac27316f108a7def98a18ec8ba37b641c7024b8529ae87b119a3e12a69298301f8b5fe9459a05375fe1e2d82e3ee905b6e56afff6f1365576189538276fe58819e0836bcd6db6ddf6bc2db6f4979951e5222d2f7bdd2503b323c71d73932106fd868748f899db09d94b86631eb5f5b7a7208fd3f00ed94fa5f3472cd26d97a7cd7b0648e07afa99317251d07140bfaad5fc236023077828768ce25c0ea7f24bc0f235b9158e3eb55fcadef3b3ca2eeceef837e13420a9a4d4caceb40b73fad831613564ea9345c23f1d595cfe10a3d15c08fc1330227af7e68770a607556a96a2290672eda0ba0317685eba69c5b0ea712f9f1b17108834bcfdce837a9668892872b91c713df68ed3e358aac4ca9be97e9288921b1496241508df73f09be72f28923eb4029b0fca5ffa8b2e42e92c4c5d3ff893ad0d9c3aba806f49890d5e2799b1764acfcfc4901606ae5f033416cb5649a6c12ce5e4b12734f8a22a410d601b0183f92b7a0a88b93ab47a1ef9b4996372195f5662643f9ffa0efa200f7a6032e49f2e7711bb64d6b12aaf21458891dc61807389ec7a2be3e3e5b4aabc1a76c4d26afe981221721479764458b4f1e96705542ba7a79eb6c9652be99c01681254f7360c0af59a825cccee922eae17d6de0f223a4ded5c979f5606d3da900f44ba6d157f04f58080e5d405a6c1e2a213d976eadec44ef498227ccc6263b9596f1b8a0eb2ca5fa09083bb2a7200ce30c10b1cfa2016e929ff659fd3088f88dd97aa027c69bd65274e2cb45e6555c340b6fff8448e23d1f4c0fe540cea904bb97ce829d3e4a8342d10b050bad8065c0f96a54ef798492148dd190c433b686359570cf5a4c7208565be1b4d40071de62d3254b2315575ac95cc6a358492c9fcc745f51eed9ab72478f2228a174dda9fb206db03f86879c856ad2438618b1ae44f0e88937353c9e19a9fdf26a8de8c0c0bbf5503672e7be197eacb1a638766862b4c07e38c31f4d5f4a2f5cf62827d1c20dc2c88bc9d4b9893032883ec315846963bcfd75ae6e144e27e89064ea0fb035c4ee67d2b1f1f9b0646ddf97decb5162eefc53ae143aefa16e96c76f582771025292703069325f9e4b2c5982682d1592eb3dd9d7d1e7c43747daf8d8fb898f5cfe720e41987f24e27b7235350a350a41a53b19def260a7229d000d361c062acddf2f3d2ad17614e320499089d4d551dfc8e443b1397030ca10e2fd68ccad874f90bc4acb6f5704637ed0294c8c4ecc6047997ba1c384b2cd8faefeeab29da574b46a1d2de5f1e45fce07f8f0c17c8590984031ae77ecdee8d6d8a87739d2b79ab9cefb3d52892a26f8ae3ea99022eff19b252eeebc102ad57e31b4838db13894efa3c1e844bfdcfdf5161a0b1dd45c627831088114c7b17ccc881f2774dbc6742886375c628e0e7e0830f03473715db3c79bd4c1a4a3b147057177c568a8b56a013817b208104966432596f3cd5a315c141c43e0d536b03aa74aa06a05a60a4edf21779632521be994c587bed76f713611ec29a59564dceca7be3da7430e7237e3f2d8193e1b000cbd0c9face28c28ffb84ccd6a22c4aaba7ba00c0b428b3c31bb105980cc68385101fcc710eddbc7858f0bee0665203cdb4dc3675bb65b7153e3a34c67574c81e0954cb8802a39da4e3d5e85acda9c1f4c177b06f8dd59a4f057d10a82eae3de7ff3952fb6220a9bf0956abd1ed266f71ea9fe73d7d97c9cb592bb348698dc613d2eaab9dd32eddea5a8c83ba02db77df4b93d5201d52911d76435b0f1bdc5d7181b63ea64a5445416d1c08fbab0facd7f57043dde940a9839eef1851fcc17c0f0f6e128a0aff0f46d353878b299e44b6f08b081052820bca1e2b4e44aabbb076ef4e05acbec671810a546cbfe62d8318ed15d16e76bf28bf153d2ee647738f2ad82afa7ed0d38d8deab8675254813b77ca959acff5ec1e46f2f40695d07f472634029aa87ae08e71484a6eeae8c6f68816447a16889d17647c3b738ee4f20af744d1dede60537ee0fb590ae7c807c6ee0096f598a26e0ea1af36cdf4dcf57fe56366e6998a64ee555a05986d21e35439e1846c64858ce19e02f9acb92b0ac182f4c5f662dd4815999a3be00c7675babde79f8b8a3d94af2051297b35120ab0ba8fad4fb583da134a110ec05e7a1ff47e098dc210399eb0332fa6c4e0ab2e960b1e8aa4c9bd19febb8f80dfca36f40540210f61fb881051022ca7c1408f9350001e2c3b0f9d4967f514c8a2f1fbad5c140eff42d5274f3dde15db8ddfe542018f6bdedc596ed2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h27f0f4fbb67eb6130e6d718716d9327429943680433c5eff8bfb38d1e9cb30a2d49e94c1f5934db1f2b6312010004bba9bafd408ba342d9ac4f106c7da74a43dfc045871f0877c15e1e691164296b8903ff9fc96152b68c09f4987380b4abed7b4b4a27cf9aa17e1ea7c9d761d23d1615776d910f94ec42aa1cf8da698c0bba7a5bad5bcbe97b8f6332dedecb79e832812e83de1b6015a0361fb7c2212ab7284dbf9f89c59827e371175fc1c85fb3a11e0cdb1c04cb9b2295fe8287a470ddc7a669ab94e9a5424b7c627dbbcd4b2122cd90002ff6e93536efa932ca879477d111b8254648db0ea7ca59b12089e5c6cd22965342faed1bad5bfc2701048de32149833a3a72e5e76c8088ebcf06ea2614e8007e9401b9ee01ab1aded2a93d4f8d20a2ecf585e3e9291dd9ee564bfa74f678308ac2434ec3e33ba2cf0b7b3729c74201ac734931a2de23577f5b69d4b455c0ae84afb212fdec5aca8027605ed65018ae60094dc67f675c6cd008b0150937d1b919bc0805483aec583c02f1b9d1642e11be43896f4b6e5c339d38427e308ae1b9fd4c0bc0674653b9cf8921cc4b8931d6a1ea3aebef8afe6d3c963d0a3f342ae9077fe326a5e81a488bc3d1ed629af833f3cfddb33351ebc728f52742b4ceb538865e2b648309856e4014dabf8373667759494ef06a4f7b3cd194e2929820e40b0f18551e7de0f54366d82c3262465f0c80f4f9a5356f82bfa3e28e7c321775b342b84c7679668935383451ba5f97075f84ee0f60a593a9bc5d354f803316682302269deaaaa46f059e5d851bac2d944fd566ee75900c7ffcbaf8018c7b7ec9b997a74767fa22ee80a9373793d29c7025b293d8f75294a8484822e2e1130096946449f642da7fb1eb393be747d16fe313b943352574d43ece2b216c35ea0d448fa58ee2f83d32e35de91204abc5b6a6e62d7c8ad8f9c1beaee68beb968bed9fd1482f5d25e58da03c427636a9a8527ddd3c6a9c3bdd8ca33a00f110fd086c879e3c3130c6985f9a28232d2cfae7ff0109d0250b32a8446d29f78a1f49595eff998af82ae6b4a3b5f6fbaf1000bce92b0d08ddfb42c4b35b28bedf83a60e7e932bb6c3f78f245e1645ea924093d43c2bb02302b1dd66015af948a53a0cc9b8c46099fe6f8a6875d090e310756d94912a7905150b564ab2b0d9bb1a6cd31468aa9f96edbb1a16d41c0263281a824f7fd3ccc31396681acd4e97c30f6b12235b4b7cbd82238f4de72aaaa1f890f5c2641c09e3e5f06be65edf97b510bcbcc02473792f7c4c7bfe5176868a6671625faa74a8268894c8787b3c65f726cf4f800a1d14bfe2f21c2d7b1743c3007bdcaa40ce2f0197cc179822421bb669113565322f13d1cf1c4f0e2594e280ac7f90c3c39e85144cbe39f0f6337306511b858fd894a727dd29f0cb588745184e5693904a200d30842ee14d2c422733f6b3c3dba0d2971a937803944329f7f7f02996d765b8e002922246601ba266d65029cbb61aee6ae46093c0ec7ba74b1275d4bba49123a230f25e23a63f99f2aa3fd09eeab4b1d96a919ec597d475f236a0b67f17d300535e56f7610bda97b5a15d4830f9f090516073ab61aba70925ad64a40d76f2f059613d7e430e587359ce69f8bb4ea53a76ec81fb054dcd4e6a01007ec5190e1947e92149e54f5b2c6c481aa823961cdabd36542f1c5c25675ff017bbf19ab7fcfc8e6b27f1342a8a581a054482fe16eb9e9c573031d1dbdf984cbecbd76f94412910094fdd49b9c9bc1ae11254da9d9903baa1219927b225535b6785dca0e816f39be3d5ec582ac264d06361645cd65edddfd100a5598a2e0736e2387b1eafd6fe818a14c15df27088ffceac8b0cd6aa496f23f6b09cb1ff1f43fe56838429df11487b5d97356a8d7e70829d921c420f62ee84c96a6677abc9beff7e6d64a54f3eb50267fc3b814b5e128546ec769d515beedfdf8f2ab75ca3d9caf580341f31d5ba7794682dd4970d86feb32500a674d23bddc658f07d468d8711f19195899d0701c9d17d28c5a9a667e332ff7951553be35d389e7478f0b8f9f5e92c35c98432c9224ec575d5955a5222105571998a51c447732ba4d4198bf8544fc0886d05e736ae15c04dfa7434bc1c27ee5de98fe981dc4facfdb3ee4445aff7ed84dd1eee57ef18339678fa23d533d222b546b7a8b978dd86f87582f668ca1baebc2fe8bab304e65ea03312ef440cdee1552085ae3a28e1440938566e0cad237b58a2a804792b78ab161b08b1221bdd6607edce4f66453b90dd266c3d183735f1787a8b1e77002b8fae37ff68af6e09f3b92330c83acd84ad900214f34b4f2f8b87a8fe57faca089a924a4f985e9facd8429d1506930ee9a2da9306d2ecfa0aa3091f0bf5ad3d0326a18bca38bdfce4850a51de0b10768c9ba4ba4f2629ffb0c96192734fdd405d399ad4b627437595ef0e9bce69baafe7aad8d0c40de7f28228a0fb972713d1b821413676f2adf65d9987e378f0707c5e58f469d2769c48c7927cb5e608e2c204bdda9a73c17f575608b24b5c0474daf381cd6df2d6340d129ed701b2263e34c6750d9a4244729b5a901f0cada5dc5f473d26990ab9806dca23be060a96862bc362b11864bd6367c6dcb2d9d69b767c00576a669318baa6ee55341747ac32ae48bc35ab9f740665c9462cf175fbef292cdb09780795b868254d59e3f1b7d15d6e268be82eb7b21c6138187e6a2151cabb4d5287c9599454263806acebb8f32aa844ed7fe0bbbbcd4485cb801830681f6a92dcb76eeaf5b1ef4e56e4918710dde5bc86c88ce6366ae4bb46d41b8d5d73313d06492fec12d7d9bdc436532595d762bdfcaf91b6f2b96ce23fb34b64c9715aa3740d1c38a98d8e1f8cf058d0b67a639713c7de3d4f97d88b141ed8dbb30283d97703ea79ca2244944fb8f7ef5f1fe3a15ed6e49e9d49550fec2bdde771a59ac4a141ed92e307e35a4afc3ef37fd4b2e34c008b83579dda1b57a881a5102d77157bf35814688c30c46e409c17bfcf9cd3386eeedd1341d570ddab9f7759f7cef17df206453d9636702d054700cdf30dbc9c88b52d2db90e6b4244e44eff2d8638ba0c04534d4f4e1d67c67204d79331ae8653dfe148166c3d94e9943f168e91aa1df0a8badaa40f721d1e5b720cea99c3018f01da3e81c81ed8764af37ec438eb91f327feee45a35bce20b67ce0b0aa8ae316c292a8f591ce0b854e1f68a41f4459090e0aedc5fdb834be4a365ec4f84e62f388790b26a13040f9e64edffcd73acbabe899ebc5ebc67c72485cb6bf8e9bfb364bc7cd87f4f887d5adcf0a6e8fe7bbd179d8f5a615da5cea1a629125f96af12ab24697ab3492effcafc6297b47954cdb73c8d82f7d2a534c8bde774d2e35be87862b346e00c2c608b43bd9a159a58b0500065a3f3f47e8c3e1a931b8fdd45a1833929bc846b0e0f08a99c33f4530d16124832a01eaceba3cda3f7341205cd86bf181425e8dddeac22ef43efe1ba10b420a8e08a28db58fd22cf533b9ff926f092594a593f5d0ab8466594e857a4210df394417fd438e2acd9176abb9918a5ea3087ad351d7f66f562b67a3b30816249c82dc24bdd67067bcf484a5906d3e5a9fe25b6708e3989fe4600c39489ce40145f204a1a30c8652217e534f5c71961ac8e965b01b4a1a84e3b07620d54dae23f11d25700d4d05e77b73b133d2603b3915be9f5c4d85d037d640f513b042367c9b5f2a959d7c9d7c130e09c66cd8b2dd8a9c3ea6847227127822cec837cd2128e6ad8502f08bc13872682ef2207748925ea0be0f4ffa5607a3f1575b48d42b7d56e26fff8a911d6f77b50d7616aea2bfb3b284603b1798f972972fa2b0bd69cbbe3ffbc904a6eca1019a7ab0b5ddc55da22682f160bb63b3bf5466523e74df057312c08ebfbf1dcd64482d71de5f7752607e32d28ccbebce41178d6f9b68fc816c0da6dbe31028cab8c945b484c4cc6aa81ddee78ef5d7573ed9a7339e0807d0a751714a4e0ff85192e9a1bab753c538e7ab7f655c5a696109953c250e11b0dff746ff4257c9b01e646862f5367e2835049755f399683b94310d6423eee11e0a357421879d1a8b8bfc2395e0463b26d071d2e1e13f1876f02db07a4daad63eafb3fea2cd79e174783e48dff1ed4db45eaebab865b134c6c77d97b642ff4cd3f45eee362e991cf9d643c2de32723535fa53f480c3e4a01ea555cfb23506918b86ff181181fa45e1af61bf04e1a71554aa0906648544f489f2499a57b07bf4fa8f4154bd68c803eae8454a7db41ed5d7087e958200b2cb41a911d48daaf30637be5da2e36d060ff0c187a5bf97c2e896f98e0d105c03eee07b101be056298c759c2eab295791438f4363a4acd51cb3467618fe4686adc25b4393fe1ed778a40c765977fc54f446c290a32cd35ebbf12a69d73a9eaff8c2757d4fde51fc712063115354a1026eead47396a699656f99b493ff2bd2ba28b4be0951638e9d86d548056bd1f59c6a700cb6c0036dacfb26e633ca12a1f3fe24c49e88c295127e547c06f859ec1f0026873f78976a1005380efef0af221317158857dab2143ba6dcdfd84368265fa9c8b078f77ae23078e7b88e2a1fdb6ded8ae2c9642a45c5e33487aa8a6c16e1f0a0370d28ae929c9117c01d779d110cd7d239e21b9308886bebe8313f37c7a99deb8d593dc93134702a169ea8782a52f08fef802c266791150bdbd44a8df35bd681de553dcefea0a09eba760547c3a7f493a7a0c9138cd8eab228e84d790361a53de9439faf019946c9f274152965509fc3bff4efef990683cc09841bd1b8f3376eda5592f8db7fe9c5f1702e8841023cfcf22256f40d39dfbbba92ff165285636cebcb6f1d00bf8acc3a28b6df3a2c70dd9d21d483fc370922001a91be57d1ba08333d9ed4328afaa3b72442c662f278f329ce7bd88e1623dbb5d1b97462789728a522767e6d96868d062ebe546e8fa644e637093057b632639f0010f24208cee4a99e34fa20688ba7262c4c3aadcd7ddc2a0bb0c84863fc4b66c268dcff8e4eb98ca5bb178c8c8c37b010762dfa33912619b653b24c417d2d9e66771d91bc7d6df06f47c91763a8a2cb49310dc0ee8e3ff0abed9cc96e493f53ca62792c6a8866cfc0a585c68a2128ac128771a9c795d7b4a14e6c3e3ec6e927bf016661ad9b28b4b8bd31406fa55366ce3a6389f91d89587e759a9a319b884438f1252855b7379c8532b1ded7db721cc0cdba6e78e4428ca8391b2a6b5810747499c9a4fe4738a37fe19944a6103e1d8e07e2437d2e40f3a045fa389a5082fe0f96007009c7d209c0b144fd96798be7b431143cda07a51c7e11abb936bca24a9b9c88f2c3a2fe5e19082687fc1f06bf6bf2bb9c2a82b517faaa3c37eed2649ac0a22f9365111ff686d8563544f3214172c0f6cb5222db8967863f3deb622588e509d603864f98fa0579bc172c3ec01f57827276056eb40caca8c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h46e73e60d49a83373de26158455e12ac7c6ffd2fe826ac02a187893942f049aee3419a6e5691a71f7baeb9d291127de0996e56e0e5f252974fdc623324ed4bed94de268da6bbad75e4233ffd21e8db9abadda0921005bdffe1dc5b957a42736c720afc367418c5811545a3ddd924e8f3657af38b1f038bdcb242bd09042063965fcd1f2c2f12d273a0851aee5425bcb6013633768dbbc761a9ed80218f6abbf809293d6f3af830702747a60cf6534ec64090fa532c91f3668e7896e9bde73ab10e873fffcba73d0c9cac2cc3aa26f1018b97b8d72f96cb473caa54a4158dbf69cbcdcb714fdc83faadb11c01506d6eedba10c7456aa8398551c3c1f769d27a823a6e7d1ce9df158e10df312063bfb35f282d4fa64e962ae13b564057cf86d9619f7a9dfb729f0d8bb1b0102a81e2024c796547db27a90329d836a59ff139c03bffeebce033f9b0071ce6603431f9c3477d9873d8bb757314d08a3b297055daba723b70691958152c3532f2e03d6399b382078c2a81eb8078c13962774508461c92e0572934ef8d6057d8f4881b4259313b2922edc6179a673aff987ce5483a25e558d30bdcb757fa227b79d2cb17ce79a4f989e02d3dd7d9099277efdffd6fedc6c278f0ee6d9327c36f6527b0ee27b06ef8d16d91570bf68449a930795b912d7977a0fc9451d6b29dafa0130fa988fac5fb4233c47ab6c098689ca5a0141409c6b81adbf5248e407993ba2cb082853a15c7107e05e69c4e6f004e29c890b7848228376e6eb68c6121c0c25d865cff579ccdc75a6feded87a2272e423a463d6d2a8b1e3596ea29722f99d97f66c56a4b09513952132a68b0e60fdacb34e5249e5097b60acce2faa98be96ee2fcea7824f699a81f9aa487466ef4ea33c93c189a46e894a3482c3be3f5672b1a1d4d7d95a9c76d07f932f3158450a2b73c215c3d9b48056540f094b6f3996cf3d1bd984e7bb0990ef729975dd3b9c4d2ef6c08c937cfe9bba769c34c6db7bf38e36ce9e63a7253c97b6f845980890bc712d30998030ba4c2300c3fc58f3549c898d4a6c7edc974066c1fc785af2df3ed755a5f090099f8e9ea5b69751b5857c7102d9f005642daf98bbbb67d77bc1a9f6c9638b172672c442f5b10183695c87043abf5ef608d129b69854eb23989399b807b99c388f839cec9b763debb92157f6d06ff4f1958e174d8e990db503f49931fda161ee7bc70108a443baf4b0faad20fba72c7e8c8dc4e63ba4c663104c85554ebdf45889d528b3c5ab8507d1266457b23cb11009af1ca957384a59630345df9cba1278381803c8407a7b21591d295949b428b0d8b45034cae68adc5417ee11be1ed4ec37cf3677e2af490cac74a1b794b433b0da960a28ae4fac93f6fc7b24095747d80ae091b51841def8c62a1b9b8565a2ad3206c9c991729b63faeb1dc408ccf53ace0c2d16b71269afcce9d0cccd86f60b18de31d09e882b35fe3a150b45b3ee5461849b00d0f5ac6c14627deeac507a7f576a05a7b943e9e6296b916adc9b338c8e65af9e555134f7fe40715a9be4e7f1045e913c3f3c68d4e5f398973adf592c39392fde58369ff5e39779df15cdb86910cea7299ae1583523ad3b03cd1a2d64a01f618b2a9ef1ff2ee7abd5332e559d2a947588946dc56941592581989fef9ae66e15ec12d763c26ad15ea7df1d465a8a942f22a15d61f1088c1404e9d1e4ece9adfb5f31316340ff2559806b03a465691e8797227349863c0f94254084b280d24847cd0cdd92b29a55d20e165963828a6c42d2535ee7f035777b21f20876eba52c553104daf9e706a2afd69b54df1f017afc4e8d840750313c70798b212a8d9104f60662f27e914b910ddf72dc01293d8d28929881e954fa2158ed10a8e0a8d6289558f9d94c6910b214ea8e9bc02316d3d25ec3c15d66c70b756b916555c2faa302e45a959d34100882caac0f01e0a00f0bb18692786294f2be93467baba9334256a5a5273d214d052a3aac02c53f2c4727529398dbf5c89c110119d036b2e53a7007d7a6b7ccc7ccc9d8dd7794edd1ddacbdf2067a3492dde8435361c5f23bd36a62beb64633da1219b4f1f5e0bbbe2fc031dfdee0859500832bb092ea2258edab70b28c0a4f71c1c47367ce468db70d1659a790d6ff67d655d462171630aadd2ef8cee1d3f44ab26dc06d6974b68d450af9a54fdc1ad3fdca76ea16cb5574b43a1ea43c00f53b5180d083f46e79bf078f45660ff250a161a98b127fec54c00d0982bce04cef50f0e0a1b018ff05eb3860dcee334e5a86c75ef1a0b4e6930edc14cf3fa5d61d84e5b950b60bed05b607ac74474746b9b9a10f96e12d8229c8cf7ababa3c506b882650bc7043bd7d6f53111fcfdff8228f227b1c8b59e2b585fa3c68d28bebc48ad0ef4ebe41676afb35f3b9acf32759f62dc16f0db09c36e68152dd344906decc246269c580e434061508a2b9c7f00461b949c00f9cb910a143db8ed8adaa137a788e81fbbf5731f83a1d3a62f6d44b9558903d5ffef24d3c9db520de89e7d5f2385707fea93339fc05b6559a81398894619755d208dd95867053c5acb727b0853f394625acb29101de8259193047ee9e5eb08922654f28d20ffcae8ae2e9da0aa30c1a862ab0df425d00b05a2cabf28307019caff1ad3f3891e71169c7b7f2531219dda2b0b92bd9da4584f2d479cf14cbd07d2b71645dcb78e7c2bbdca15aa1a7057385b850b3caa29f40a1bcfacd766b1b9f2dcdfa91365d00b3da7d299ad07138991bee96a03e2894d7ce6c4170fbf5b7d9c3b7bd8803a33b89a837ad89babdc61e1e8657826eaedd8f7ae96369e6468e9f66ff1b7a9af0b5a41a8ef129386c09a62be5bebae4540fb3d4f23e63193c9435a7577af3286cbb035dccdea49034cd6116a64935fac99c50433d84f1199b895d8904e4db23224018891298c74d68a0cb05d320e1fefda0c272961990e03051532cb073157c2efcb4bda88e6a721017142e6ab16976421978cc0f66e5de069d44dd5aabfac124038fb8e987f86b047328a0ebe44224c9ca20654cd3abe016fa1dafe280b1ddcc485d0ba3cc3c162878e05eeca9be7fe6185691cec8238246aa6db926f24eea0088c3a500794d9384b32898b6fd73257636b0cb586c16e0603f5ba51f7aa7b57cab8d82c576631afdb5b9e4cb7b70868e32817b94203b5ebef2ebdfd9b2f3ce0c2711eca2f520e3af064cc1bb1d6bc494968666a48acf92cddbcae565da6fd15b99a6f4bf06234544339248061c031468276eaa6bf4563dfe0459b7519876afdf96ffd88156a2be9a0dc983c1854911c1b38c6732faf0d0fe87ae296c75d770a2cf9c23393fb58e0aa30da22f0ffc21727467bf244f26f608051311e3649fb7c7da3ad3406c3c7a9b0c6ca2f3fa2ea86eed2c13c66e935ea70b8d085817bf3561c2fe3662af20a01084bd0c5a86f7e75b277451e9b9573a6711667232135ccd85af589b92a3755a7639fe34c778968fac19f0d9597bc3a8d2e4163a9ec6ba86fbf73d65c90b791d22a20f3bc272d691f47fac2ea146c20a215fda47330bbed4f08e7d99bb499d1728976fe74e3942c48eb269ab3c991e03834f643bcfe49bdc372d7e44b8518a4657499309a424e5919fd5b442bcec1885e463f0b9443e0cfe361df7facd506c74f9ada5def3e22e485e059947a4632770dbd819905e5c18ae6462b460e141de64a94bca501c34268afdb59d82b8a35b6911b7f08add65e11a10a7bddf18a30beec88eb2be934129c1ae71125d3deae89421899f03cc612bcc0eaedafb0aa4c983634b3012d4ece5e438af57f9298c6e7e514cba9b4c5cb010fe7a96f5d704f7fc7ace045443a964962cda4fdd2211078abc058dfbb21ca053632da9623a3297bdc4eac786f56777803fa0671767c36c304ffd1546acf62c6fb51c4d8272fb12104f77fbcdd0f7333b4725e6e790bdbba27eb2a62ea7b4bc090926c783dfba5a0987eb18bb7b4579bbf6b96e49a0d1348f3d3f061187c59d04097ff5af7de92b8e206335901a44950f2c2b6f23e1c75c078caed3912cfdfd0ee898e80cdaf49ae165ad259a4042f48fa16a1950155023251c20ef159f0ccc997b735b7abbe8ff3b2704bbd03eb7fd614c332c2511f4184b6811161f8bd9d6b53ebd121b13c35352e605b7214d683018ba83e0a4f982488609f36612338c4b5c954daed1ef59caef3d46906c4017e6af28cdcb04a89f36066d42f3571a7e21979b4c4abe854884f3ec51ef3369b4a438850250dad68ee320db9d43774cd637ad1c927e0642d07cedbff3a291913b0d496775cbafaac9b5f14a6dbb011262007d70e123fb692b09eb50786796569869633f0d0d48b36fc4120a306082d2ea88bbb35ad03d8a6a54c76f4247aa0c59e38ecc66d8988546569e8833c1759228a4a65c56e32e10596c71862085395fca1624a67d5cbfd9b944f0b9e7b425405aa69a44e7e36cfd0622c9838cc0974c20038ec5725a35b55d45e08ccb5f953ff368cb105516872379e3ad95a249ab8b7d20790df0ec8b8dc5b71447784afda13e6e650df265a14fb6312750047c9b1f9c8ed9b4a61f7749accb7472c2aba979217a6712f909847adc82dd9e47a5bb758200afa02bb049cd5b9147bd39b8d1049614d3854fd0b3733eb87ff347a5844a10abcdafbfe824bc799f34e9d56bba06a23ef9bdb362844ee6853ada5513e1d3c0f54109d2e29c1a9cecfc410b1ea7d2e5bf227cb12a7dc69d9b3f2189082d8fb797fdb41a6881a03a18042d21f15bc7fb6c0e7f41ed435dc79ef739f265f98381c6c05a6b9a029b9294d949fcf1be3602d2433aebcb948c9162ed5be0da3205e7d2dce26e9a1bb7ef2273b36f5f2e090e2930630f1cb90ce8c09695730c40b6559e0decde240534c76c137c34caab549eed30463b0fa9961cb41df11a170f532d77a67d15c1ddeb36cd3f91e3d4af144c6d8fa9b0e864e6e382488e85d839618a4eb276aec6e03f6237356f1a37a7ce46b823cd3fcffd587360ad049bcd74be7f1c1077dc8c8c182276e649f1ba52a80cea6d0ae57c89286d46b634f0b4fcd18bc420a9d11a3b9e0a3ece7402eadb730d78f6c25312d4d530ce75beda8fa45e316c6e9a14862ed57ee5bd5809c57a4afd97027ffad363ff205a3a7b3b730ec000dab834d75291a613e38c873f7eeda2b98c932e6de14c99c05091a72cc559d6bc2d44a59d1a3158732ff1c2567e4174def2884ed5dad7b172a35a6c5e5f15e27f8d3e61ba31d96a3b8d300f5a87946dbb518fe5dec29e1dfb436bd91ae36067ff23a01e4927fb06a79ac1756779a2da6d6f7c5a91fbdaf8d2f7137aab91c3c711ec9c5202dfc11e182ed0850331ac27e13d85b6e3dc570e9711918870f3411f1956bf1014948b6573b4062b2e85657ab55f37c03f925438e81a0fb8b74922b04d645894642ac98eb61efdb5991500376a9548168b5e19bf0537593d5444ea513b9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3c319c8590edaf1eb04b18d932c80ba8b0b20a283de75f5e476677522ff8d698f296d09f538f4a98cf61574308eb61140c5d1b05254419f75748a89d3f999c51064adfe984b399b65b46e15e59c762f7bff6015e3c5c3d9ba6bc27a12157b3aeaeb3ae91866c6f70c4dc5026f8262d9dcb80dd6553d506f52af4e123777fc352caf0c8624d2bb8deb03a85c444f0f4d032118ba2f3f3a2a787f1d24003f2bb88d9a1b29b186f9d5fca186926eda216415205b7f5c493a089bb4855aa41c6a769fdbf077d63ec45ad45d5d5a709e4bc27fdb43965b670a84d20a7d16a8677591cfcf333fab656ce87c6a36a9581eb8594f6d5cc3d72844de23f1a870d424aa0eee8df26e2598237ee6482561c6858e5504458ba0cbd4d811ead146ac70ad38b8e406127247b195d3ed71317de9a4e565f24a81f3fd7ba71d5065d4f37d176a9c4850456725938ac962f752ef523add282f8f731662f9dbfb97262aaa6a36d99e3b30b4251c210c19f93105e972031ca2e303846b3129813059973c4c347a3bd0af07a0782c8c26403dc5f52dfe040d6ddac3246cfcdd45a4ff32bbc7dd8b159530cb261c77fac9aaa87124c5cc4d0082d6d4021b415cba1ce84de7b59876c82d31e9723aa162df70e0188d212f59ba0fa3fcbac8206103172527a9f751d64b771341e8d127fd52f836b913a869224b67414561a628300c418d012e5a4787d20686e2345995e0ad11a1e50dcc1e474e5a4d0a59eb6f837bcc494a43c6260136c69907e6f3de6863b9520bf7adad23f4c4be173c4ee577f4473da6583b883aed72c3dc700dfda41c863d940f6d8c43a7f3317efe84163db310db9e798cf7544cba181f45a915f8fc30b6849cec0b15017f57ce6257c320813d627a9bd1b0cdd1c0f22d47c0170a48955dd6ea6b98ad25ec6c71df0068568ce6e39801bfbbf81d846cbe936178527607aba02704f3f419530b3ec643766d64ca5168395d7f1a73244f16ac6e8f1dbfbd50ace8dbc75de3f8f7b72f75068f8ad49b9a7a84d3f40510913519cfa7559978031a387ae879c5207f738f8b50f6413c38612f4d088ee539944438f57df8706148de1d83d349d4dd69e41adbec87adbdaede7f217982c426efd476aca7d40bccae882d5febfdb0fbbba3cd9332de0d743701c3033d4d39928a5d0b8b3a8a764e322326cec12ac8a77cd6b0c040836538ef3da394d10f28bdae43f367c574f57e9243df773473ec63f5920420d4a69d84bdf60f99bcc7e47eacf77b98eefd873f25ebc883277fe5aece86512ee2e83665db1c481e5dc5a165a338cc7f976be530a4e755214218063196ea9620726dfff6acdbcafd8882c5647b0ae70e518bd36af8d2b749f783a452f35e817e981cd359af454d92a8214e4396116dc172f59943af5a37d9c8b03010df3439388233dca9f870ac93b0c3fa76b3420f1d0f28bf87fe08ba88e7341de7a863cf3c21520faeb8291adf511aa3dbad748500c95cc69b7bb7a8b4b2435bebc6548db70ac23859919b0fb047e5a0109e76c5303e66837b1996e197b22b55fa86d8b0adcf00ee5becb45eb2edae5a93a6181a3c06c660b3e519428ab5ef9644a9aa9432fa0c841476e5add4c8339cf01ca546168a1b596b016bf665e2ddc392ff87ee82d8c9a00c9a62675643629f246ca3ae8cf74dbbd141ae6379cd293e46b5098ec3a0f99b0978b6bf72c3cdb3f8dbbd65952b8b7268d364355b586a8f23673fd40987d5d47cf6bac30f33098f3bf1d421d63105e26dcd0f8bf80db1b4650f2339fcec327e7a17d7e693da23f348bbaa684a04bc3132ec94f3d7965b11b689cea9c670ee2d85ba9c52f5db425aee393cc1e8ef1c423caf44c55e299f5b883bbb60c368c2dc6fe173aa0f3aaa9dbe04cc1324304783d23077b183dde17eaff5e3e221c308a4f81376b4c8bcb60dd26d1bec37799439a6464ca6eccd24bbb058a1e63934ac1b73f0973f50b50fec7bb87a71732914807e771c773394cc4a058decfd6e089ef2674164a30c2203140991be8572b92ac85a06227594d73544702900d114b9eb520f9ef7512600deaf2df250548f415f60609aa77656a654e17198d3a47572f9b39417d2b782908a3b7eb4bfd49967ee498c5d78bf7f94e153b23d41cd16c47818d19cc507c6239f6190ac5b38ae880aa7b3181193ac98dd3b9857dc76f437ac47138ae3f8c65fee05a706c6df0a4de11d65178c6031eb14e334678c52cbd1f8e5e2d278ee1405a24e79de21ea6f8e226ce3eb57c980ddf25a345981965cc46be141e34f234ffef7f5522419571fc1ead6fce19e1c99a14fd4bb8b45a7a2d40073bcad4b471b3ff386d7d84fd37fb1e7aa88dceaf3747e7821eb0537ba504933df1fc14ad756f677fb352d6b22e0c792148ac099f7a4a88042c8a9bd1c70ddaaa5cb4ca43c79cd810251af6922cd10413fbe82b48d724a05e6d6f1416c55aa10f37aed6cf35063857da1133495680328a8828286978e6023bb0c8a2c4fe2d07688c65c5643f0dd34b2a5a0e5e562b7774ee520feff352cc4278f9b79f0b4e7f86c23894e5ebe601b35aa652762adea0a80edfc5b4b5bbf426ce6759df3fbf165aa0eb057961b331ac27033d2f9db4bbc6bf2e34b123ab87d4e7df00c4ce9c7e417bfcad483096b902c5588f3eef8b3e89e1b3e6fb1d8208e5a4cd6fdc16f7e223e45ebc9b1244f523213513036949d7e1337b386aeb4f24bfdf3924f7a3427f3be778a39870033ff15c156b5a2d29773f77eb36dbf23ef9b8ec0e18b2b9932485968f54c7d2f0634b0e7f69870cd1a096846f0f91b5dfd7b0ffd83b03b0b4b7fa4420f29bb584d72d5b8234f3808e8870dcc9362e9daf3b84b5aae6d3af710f05483d2ce52b421bcf6da2b6f39b61bf6132777043017dddc5387e395b45eaea6ab3108998f99fae82e6c6f01eb66d46ad6bacd903ba1b89a59ce334d6889a92e9a4518db31dfe1e7cc4398e48c731cfa329037f7fe9769c8772ccac8298467a504014b3bca21f6b17ef7de3559b1f8e65fc2af321ea8273029b93d588b499448d993ca3b4c6fd21e8a86bcc9dad1199e178486089d65cc56db543a7f0056a2535e3a0e9b55d4d42e8c53140dfdbdcbe1b1873159fc2e0a2581540405527c42b05240b5ac8218adcda2696c64927b8ab16ee18f0fbf0a595306f803678225fdf075f622b804e91eb51c9b61084314c6e54fd16ef2b857e9cd74875f2108704325dc414b0bf02484cc271166d174d233448f052eb4ada36e07b9209d66ac2033599aa8894fb82ac55508d68b2d786c2204906e4ccb78608efdc01541752932347c1cee452e66804ef86423f42c896647b99cfa05ceb5611220a02d84865bcafa19e6a7055acfd555f63fdc7d4009e3891d42815fb166ae2f0eab67f937143d65f62adea7998bb34e5153b5692b4487e793ec7f2a38005ef8208f67001c63fc0491d3e578d130ad9d4bfaa406b7b315db2d336aa911ef00de6a9eac308e077fb6f954dafff25e2064b2242ef12c4f28702928049cd67ec45536f31d9c15bbfad4cde69eafb660f1461abd5ecb72ab0e7ccd836289ba0a3488c7fc2b0077b921d17d636f94e23f9cdfdfb6f4b23fca6fe17c2c0ae48fb0acdb66b62a46bff2d43656ebb8cf8f020310b05bfa0460a82f78e63a41a86025d49ae49be4324646f3bfa08a385cddb6d27cc423379a58283d2b0ec69e9a1d9a39e11a6e8177c87e92b9d5321254d844f22ecfd7ca84a4cc25f9fc37c929af5473f42450047b4e84942c90168f51fea4c9951553ae9d7c644a0b5cb9f3ea651a444da7d0e08720691e216c3f7f96deb3b76d9d599027d690174751d52c47ea58ad292b9b8b29859fa792bdf17c834c0c0b827be5df51d91509d7721f47d19e4093c36a47605db96d6fd5cbf746fd2c5df0ea4a4f65d20639f516a8bd3742621797dd88cd17faef4d404fd77d0cf21333bb508b360f35186818d7874557dcb4440206c5a5b000c57b64ed81a0dffbd08d8cfa6f494b7393d10ee4a95f3d3271c42d51b8692122b07db954dd11477d1a5bb78fcfad40ea5dcfab8df26838c384cdb435130020d4fe2767634873bb81d17e14a51dc1ecf41b8a6c8ffb3c6b79bc13eb8637a4691996805d7641d65b29a9138f357f116163861923451c764d7bb69de40850c32dee8e03c762e6f5cb7360b502e2e4bf585d9f4b638e0795ac4588477752487e346fd3a7bda721569afe04d427ec6e7934907c7667417c28257ee9181f76447d7057254c1b69071149c189044f756c445daf47e2be766e0d3fa80187b75b553c76934dfd797ee83860a668359c0f242dfd950a9cb7f97ee0937fc0c373ecca319480f3e746af428949ef1f31db9a78cc7f62d84696710f95cfa49a6a8c7ade1208eac03b2218ada747116f95e4297bb38e59aeda627b8ff396830c723019613e4965c377608f5499f4f07d4bef48ca58f4b48ddaddb2d7be74f6ddb5fe3afad805b6ca8056686994f357d0992bc54a4f3d4115de504d7ff9a02d3c6b9066f38873f04d1466908b11f2f9f7add3a9b91a2b61568b41205e5c8e21fdd70994aee96b9dfdf83d9cdd56769b6e88da71931e7e3de679c463e9e21cad03707f5f7293c1e8ff1a7b5d020e28e3c6e7f0add8691c0a7472d048415ea0499022e50816f4b1f13efd4671df011df250800173c20fee4d6e73993b761b050ef5fce05e9a0d54efd7e797c6a31a96fe71dd972144aa96b91e6cc2678efd92fd21244df33bdb3e779e7c9a3a2509b8d2c6b5ba2626521edb136d896ea64fe11898c9ae82de735910d537d3bc249c7505cb7c61933740cb4356a2a01579c4f1c8c05c73a21caec799471acca684b0b50eb03a74592e5f171edac0da37c78416c8a74c2572a6be20d82dcd97f17e43b2486af602a1133009254a0bbe3b8e057eefa1d4bca7631dac6cad534862d4aceb52f8d5b92c110afd865de66331a5ecc22772de2559c9b84ef58a9de130d1e5fbe654caef0268bdcdee51324b2c7f79d197963edabb62aec06f3b9edac6fb9f8b926a7f8608522eb83e08ee00fa2627f64d1db2b386caa97457d875fed88a725ef57f74a211a230fcc7b8a92b4a544f53553e6b8e7682fb431d99842a4f7e77a92b5976aa0d3247faccf29380833b24088ca9ea377b7e84bd3d90e075aab7c8d8aed11ac79ab63cbdc27b24bf6e4219094d24e52bbe6419776f3a441ccc71936fc0a4f9c36c43b5c08f8fee8a099f20ab77070ce45942b2db48163847dd99e95a3a9774969e0956264a59d5f07078d44332149b7dfefd38dc0309da70941fb71c93884b347b862e33af5f94c7c5bb4fdf19e7ccdd77932116123d143f7b3a773c983ec41a066b23dfa6dab422c7e1828f0cc49a29e9b26bbbe83279cf616df45e528b7431d17eb8a16361cd27f266fc80811e1bd6e47ac8e9b17c1417f7c198223da88de36878f49533d55d32e5cd7904e89d99196289a7e42;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h456a016947e8f5dd6eca3edc933a664dc85173b7dd7572e5385db83a71e20a8713bc018bb6d27e5dd18908c587a234576487be525409144ed0ef8818b1a3c153c7608116313fb980ba94bb5e841b0fec228761dc7d5061315633c5def58a7b65d170d0838b1f4a3c0a017477e0240cf698c5852a5b663d5260bc1c5049445c97064f1eda22b09e083f75ac8b4304cc4e08452fa31f53587ba4278e01a4efd5738e7b1f5be35cd3e2948b9f14859c5fda146d5b131e1a854dfe0228c2691e7c03e55de1cc76c22cee407214f60e213e647242c2ad91aa00b2fb405650e09eb05542f4bde31dd8ddca9cbb4a8d0d1ed60a2782f41f076096d7f9709d92e64b754bc3afb7669429d18d749b9b79cf84d4c6dafd1cc86e21f38faac90ea7527a2cac4c7359e89bd17b0c9af6a495059783af30c4370935656d00b9f99810bf74b859100131c34076364b0157713aa3fdb672a692b3ac7e56926953bb20603a73b24c82ba44d15dc6710eea723f503a6d36c239b6c6bd5043c7a1a8c5f1d90221323687fe8ec33a783c6c3fbc540913b4b705f7e31b0579b8ad73e39d41c986489f45625bfc46c5105eff33af3449f4f83b34c56c16ec91fe1237abc34531968c8a371939566a5afc9019653509a6308b89caac637ba216a78749aa4cd8d6ea16186eff7771549c11495b725485ed877b02a610d0e2f79e95329ecb7e75606ea754d9258387abdbfe556ce65a3cec6eb53f4dccaf224ab220e61a380a732d3f457df913a6b6d171f2540a46d9011a8f753b52a8d173cb22c426b86ddc501e9cef7c6ae8e3993b73a80170358fefb731d1c0bd041dd37d1ab043030e7d37ffb29190aab191a3af54907b4d267fc5262912b803a19615bfc2dd78cafe0fa11dba92e78e843ac40886f8a58f0cfaec6aef4046ba91a4fd1c992d7278954b839c5d31ab745fc1fe763a1b5e3d2ebc6149f082a1ccdb5a8dbb73692c6c0fde6018bde33823cacf2e2938eb636384dff771cbe7000446fa45b33297d896b32bce3d10a55e0e68b8b3621e8629dc47e200e18c72bb31896e8273aac2f6f3950c6e19811d3f3a7b7aaaf69c292eb17ade4e6f67003270c07f4a4d88749eb76aae2cc76cb05952ac7ee7737558bfb5516777c26863c9521b304a126f124eaa5cb225e38db3c38b3310a39e45b4782edd5477b396b2f8bc4f6541e9412a156b59dc301bd45db76eb7a75d75d37379db07018293292f1320b2dc265fc5e57d4582cbeca5129e6321f3e68d6bf9f672361595e0e4ce30253d029fda3b397c9b1d55a67d56941ed4f540d47750eaccfbe0acd5b81d23c5d0479ee446d7559e1c72d5cec51a8698bd87f23d6cc58501a9b7e77504875812abb1527152fb803a070c17492e9a74c87691a47dd601384cc054cd6adafd45a623f4347a4077b0972fc636ec8c525223a5a10c5106f1d45b3e88f4c1b6bfbb63673817db0b8854d55ee623a3e51b9eedeba9ca454a46ce3bf4e6edcb1f088206577235514abdc1a078f230252f575b64cc76bc25e2461a4a10952bc2288c0230599e2b480a4d197105163fa7ab698f8694bc54643e193905bf6f95202e6c7792761e55d8cada474ee670abd192fe99974e0962aee2ebf5355ddadafde4b3a575fdb42aa0b4c2d25dbe445a65f8ff1953bf12602caf9425d042655953306ffa53b31dcb5c7d88a7e7a7ea9c2b8dddaf196206c79ee2298e4a133618bf03192c838f7f35623328033ad695c378f0d86058bb50e6a623786e55adddca271c30a33369e632f40561dfb5a3506dce8e37b1f6485a9dc31974e606bdd0bd1f0afd6494b364a886f40253723965ebac1ead06698e1a072825478c5bb6f6c055bdce46f7565303d43d653a07682723cd93404c6956c194edd04da60e108862220ad6613cab3816c875473b2ecb21e0505d5ef6e3732b63b5c9f53b88d26f35088b0bc79a662e8c4175192c602b5820a56f76bd57e77edd985d5d6a2831348be18e7c05bde4b31dba3781b400218e3774d8b6f8eaeaa37f3c38c9a9c1f7d750d7b5d2b3b1253e9da1e965fa1e79b128d042e141f375313aa75264509d47483abb8fdf29793752ad42aa921e68afa7d43eb96e46e8c4b464939452f227dae93f0096edf8ac77bdee625a95832dda121638cbd582c4fb8b2d7514ab7404dae784096beba01e9c1e6edcb188d62a079728b1402cd00cadeb00f45c7e38d479ca74ed392d1706825e8c48cdaafac4b28333606a53de42c2d0f2d95b7c4f8426e7e982ad19ffadc7b710bb92f81ab0bf3011eadca74f48892d438af498b20e27f8b46d6fe5255fa6aea0112b0df05980a3f961b9806cfa756714c965590d7db7185738a9682840a5edfd7127c3a5cc1bd802459a7dfad84eae086ce2609d657b7148d497f45ae2edad81a49d315f13956ebee07da2c007208634bb0221eea8d82e0d7a853b1c0f29db805464bc1ec9a44d1f204f43f3f04eac8abc629a69a58fe3a6f417e11284f741840b69c5d1f7f80ef94f3c94bb131057c77f417ae5e7986e9d16eee3a9c306406d91fbb74053c0ca4b020ff4a749d77481ca4a19a420f600bc038108ae76db7a1ef7965075972572de36a38982f2682f8165c20309508eaac037d5e726d72f06e589303f552af54a3f8d1c17c15bca0c551e808720a54bab4b1e7261c339571d176f2b7a2fdc6e09e3c7aec221862cf38e8db50e48ba947b9355e69f9ca63bdfc301b41c2062c1f3161dd8e6fc79f03ec2c5bee47ee61ba23149ee2215d189b9b25e6dbdcf1791c5c9565de67fea1a8db209c73cff50e9b9defe08246aeadf0d9549aff5fde067d7a8ad248ec2c4566c11e1155ad55cbfa83b10f368f6f303cb7b31cd52d848a93ba1a414b09f453038c640f7215c2009d30dd145d61a7fb4526759c74abc7329b93207088e83aa12359fac1a4779eca3519eaddd14a022c7323c02090eef63286577007a39d9c7a03f0f77e0308ea9266c17460c4e46aadb4fe1636f9e59f3da277e57ef3630c7b0b58ec73f24979f945758408c3bddd87a734bbcf9c998521674b75ffa2e3cbce3c55b4552810ae976b15d591c53784244ee80fbc8329638857de8400d15dd67813fd4b07911c849547186394bfa7353acd579ef8a05654bffd281e8fc912e6198288a55901e0c04729c1cddde7a271c7b1bd00f897667640de59cfba2fcaf3c25473fa96ed44dec0732d26a3ee2321cbc799141ce67ca4a3cff9d3e06da0f6bb10af852ed244dbdfdb4fb8d8f533ac23b67b89797df1b31b84a1a8762ae5c6ec1380c8f389e6d5661ea48e3555cf96f7a997af2ee4500b7294324622119f8e90a199197e7481d8cc9029f7cba5fd34a8751a797e149abaab40afb663b93c7c063fce90d13435845e0e71ca4ed926bf9c34001165fa6094478b7f8d92be97ac8bab9a9013e9f9d98749bd9c65d81c3ba0b7d2175c44d3b60ce22ff86a55c16213b6924743bbadc2da3b2a4982c6cc6d22827609f110c3ccaa79e04c6073875f29278181440f239e6253245e39f134f7fa2fc1a19792f175891ab340e36bebe022537473914525cffad48c1084afdd65c1133532ab4c6750fc77959ca34a35bc99417ba46025343a10c1ac755fb826880c59c5c228d6c0d7aaef59f42bb02340c8094904b9ea4e3efa1c096e75d1428297ffc04e35476e20a46401c6427986c37fc4c162e8dadf9b1ee66fe85464ae796393724543fe5f0489c5389acc31c181fc1784dc4f15b71cc3238d5038e1416724c402fcd77e88240e39b29a0ba9969f0737d21f42aff5152bb14d9b60f27dbf884bfc1d4f74454626fd6e67f6db286c90cfa18441cb08eab172b0d381a4168ed229c00c172bdf50762726b0e157a5743b08a729ee07d2733fb46c4f581acd99da105c502167013e1b9e3c93de44ea47e3d77bd2f4a169ea8845d5363be70e29625d477b20a50057dc6cb3f22fb3e2179f366f92a2c0601581d2d7190aaf3121d5f89e99ede2e9edfe03b3c35c2dfa201d0397b758109bef89fce4abfd19597270fa69752acada0a9cdcac8cf7f28a65cda6daf19a3e58ed17719019ce6a98fa988100fc2dfc39450559b39e103f246676de5584619c687e3fe629d1446a5bf81e02ba0def758ed673fdeba679f0d3ce91a9c6f28477f6fe3307bc932321b432fe60b9a9f1ac5c147c65373fc94a88afdb22eb5656ce6244543618a6a095532c1daf215c9986122ef322b8c4a77e9032926761023b9e368e4f9502b6de2cd8774313e72fa340468ebd32a46abfd343a1193501a6df1ec27943cd179a3874eafc58307c9e61770e6276896f4b9a9ef7408c98e23cd68c2f412c157a4d2006400091df95b9bded54012d796d163be0dddf3624771b062a458801a61c89bb10d06364fdf443dd60a89bd8b8c5d5230c1b5717771d18501efc3de207637d809a309dc9acc9c4524e28caf3049c0f72ae0f0911a053a51f192c0324eb778d06868c61f67ce3968d8a21a6cc2c88a36635b09046adec75fcdc95ee4128c3f9c9835de943b5297868c734bd02afff7ab36ca34fd5246fc0a156b08a89261dd151a3d211a063649982125ef1b5c7d02027f25b2f44a9650b01664f5d60a9357104cee7db722ea9613ae35c2e6a4b0c71385ba91d0b307d03230fbd01947e584e0108b65e6784ae8650c4997ab4cfde3531442ba9acc30cefa826a62c747020a1851a3744a3dd2337896f63866e8c69ae7ff724b0b6c3ac4039912254fd481fc7bc3d4efd3cb90313b0f6f6cdba2a431d213a666eae36c4100b2635cc1c51cac035e986e210aef21223c88bc4c916ea8706fe804e4cfaf18681d667ddc911a9de00c1c3880245b47ae6f66226d81a69fa09fffb9cbd993285fa343fc42bc36a48bb4a0d2adf5d1fddcfbe0040179871f2c9040fc15471eb6650ed4a7f5e84f2c1e8b4820a1c34c457f71c39a03f26a754e1814799bdc538b141dd382e1a763e6de72a6761bc5bb67771050f3a707b8748940f52213fa31fc8d71a7ea442f76284719827d7800626c337dc5c8fa084b8b51d8bcec35b1ee694383103941cbe5e3eca4957499f0b1a38b07a01bebc217e15bbf2619a8df84cabf245d4019b11c594d7806745c2f8e37991ed146070d2349e68564de7eaf855523e25e7932fd8cf7f77eb05ec13f5b495987a8540efb9b2120f63bb23bdf567c897d0f9f56ce583770caae7aa73d8b964a046ee3f1f7de94207e37d3e6ad2e5c83d876e815415e79676cb2e45bccfe5302284f7f1b2d38843bd9c7aaa85502f76f8e143562696bbfb8325b1d509c2bbb2de690a2b121327378e01b89cf7294265208af3b70ae5d2bbd70e686d553ade7b47ae5a01a0dcd42852bc8bb08ecc9a6c1d31e09820f577fafa860d8f8296dba9a4cefd9edc82778d8d688afa98ebe4e49616ea72d249dce7a6f750150052fe68cc318869a4021437f919bc3c772af8f1f9721fa950eedc3e005c3864ad233;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h64fb9961d54ba8075d47b7031fff20749da32f404707ab05be504a1ed9150545f16c19b7b398c18a08fdc23aa5d40230fbe8d1189b50bbc7296fbdc8309294e781bac547708d7033fcc7658f88faea0d5124cd861a431785575724f52402aeca1d041fd42bbcfa4a32c332f7fcfc61f51cbb137a731570e2873d53ef4d1640f9e9b962e30fd266257ffa9ae4150597aa3c814907a2a3441938df65f2f387075b0a643edf5944701251fae05ea61dbc9c8148c6fc5f3179ed6d1c264c06bad9cec151956a832581245f89b3fdb32e44bb9b0f5f204cfebf12264f07f6fb11761cd6cb8b8139cbe6f879eb4a1e51f71fa1e7e594c1c4887710c2722131cb84b69b91e2fe9342272da539884d7fa14898ff626e7ed04e5d737594bc176eeb69332062def4057b7008a0686611c2af0afed756d11c4f4e8f89ee97530dd956d83d5ed58fdfade559a6ae57b5ea2e78d6c126d1b45695cac36cea6343d09942cacc0c5999bf82b4193af6f3ad199def02323a5912a4d36e94528359ed81a1752bbbdddb8c858f055a259a38360a32d5b0a2e248ac27032348c661b70404ac0b7a58e78c53c68565d5acae29eaa4e63828361b204659ee0ea49fd467ff9bc00b1b688622bad949288a29276102724c237a8ee08bfe2cadaedcb2ab009d7505d0ec5b3635f3276442e75e4a0f9c94f3c6732fbe1081eefc6bd532b82e478d71a0a095202ada752696335bc4df9bdccd2fea2f64e97079a2a916240b0c997535594b647c14d8dbc61f166392c78b7ee910e5fa778fd47f6c92cd549c4279e3390f108852dae85129aac639a8f173c0b9259e06d8fcebcbadff6f16e2df838469ad5e659697b8f234a98837c16774619117f429ca0206e3f01bb2d554ab47a4dc76f78b074d39a8319df87a5aa51819f6a277e5b520844e3d4ca524a0ede60f049172ff68a58cd14ec631bf9bd68995ac0b44549de995741617a8e91cd606be564f3ac3daa86158921c753808de601374d12fc8ac684b7daf852cf2516988efaea6586923d49b8ba455381464b5a8c7dc4f74b1a0ae3d4fc81a49f666e1a745f0d4bf7b17dc7c27a62a0770d2df22eb39f9e5534c1158107e054dd21d9b61621448a910377b5382add7c77b7cc930a95142a959b9262fe2485e60e865dd19089d220e17deea3e86656fdfe4b52d8ec8e8dc29b2a4f46e7d931cf6d309f6481fdbe65a5cff1dd062e809ee7befae335512e9a9e2df6dd35198a16948c722f48bef91e799bb642b8fdd424d89551147fded5eebb6a5a2878899a1003e474633b95b44d1029de51a8fb4970338db04009d53d19370d2eab58c781e9acd53f4cf1eb3158135526e251bd33d0660e7252ade764cd67017832faf773394e797b0e80715a1a37cf99b7c0444bd6fec1776328d1381a9f090533513ada613f162ab792a004a37fb1f9884e22b1ad8e5bf12d6343e9b95e7e55931f6f0c25a1faca6b19bd0e865311f9ef862265bd1efbe540a35ecbdc8e1671f50da059f58eaec0dfa01e87d3863a25328672287ad9ffc0e3811fa78f2fbbd9080f02ff8ed42201f3bd2c15ffe5c10ec9f0b9489f73daaff077f2f1956d2e612225bac8de93355943f2cc3a785e1085e462cf18ae1e19e8fc6803495bf1d9188b135a8c11daac091caa572ce1715a02da58d9d363f07e38b00038361d585ed205cbe8e857bd475cfde0d8378d0371cd1138ab13e595666a04808360fee5d4b94584ef46d602a0338f00cca19b2fcc10bf32bb255424beb0644a269b921470bb674043bd32b5d601eb51d4ddbca0047bdfbb320ea5edfc5c60a84303452bd7a2100fa1d993e4388cd8db2dfff43ba78cd3fd24e77c364be96e0d7491a1ac1d7c51df682d7754e64b7c94e2a8556219e70380dca94ec9ae47c988123acb1e8d529798111ffd0be717f6e1eeefa7f5bde3e6bd3f2a9b86ee681cdc1e49718f4c666bc74de23531a6ca777f16c123341c6ba485ac761ac4df7acd766de03cb7cff40d73578376bd7bd01c4820c92f9fb93a5c410f2403251d6ffdb58bf12211f697fea8b8a4d376ec54f621f77e8eb4089909fb58a55990b664cdadd2d46e90823082bd7daa800a9b05c442f4f629b93e21303235403b7e470a4dee9853810dad1f269a572eb50273307f8b1d6cf978988fe287032ab3a1a0c15092b424ac5b895e4800370dc20612ac388f806ac8504dc5b23ad75c400f313d0c1dd8048c39077658940c3f67e8ce6e26c0eaf2355b518a7e5258ffbe890f246b0050bb17b52dd158d5c5f2d476b41976ca0072b9acf7bde10106f917d7a71548ae2bfb284810b8c4de771c2558ef2f2727691bcab69824c7a7004907c0698c91ca0bfdcf75dd5fc4b9095f0fbe13ee0449960d9079ddc1dccc130705bc1e04f84aabd4233829de56877adbe4b859947fecc0ca344ca8feb91a3c2a7a71cbd38b7b8ff12d6efb91eff3d053184b5f6e6658b1b8c310b68396b0bb913ea685e2c3a455edf80a08b2e8892f3b3d644a7226ec11ef136fbd82f6b33b1d77b014c4ae1d8ab6c40d0fb020075dea1daa7812e678e67b946f7364b013c32d1114a2c5a0250d78171e95c49f7c3e42ebea726ffe0b75ff9c71e799ee13e43392adc49113f59c8259d2e3fc2d0d391f30a153c691eb02257a9c3d41c53661d39a6e76d88170e1770bdf6a32193c25ccb63ee9c802727d5520d6e88741c144b6eb19a3c075dfb8aa8cbb4642c75fe04d9361fafee3b2f2aeef15d206a0df20391167b3294f2da00cdd23520b5d5a1cc6807aa828abda89f47de65deb16adc79f6222649c7c9a41abd87bef5a1f4991679e58998f2ee751c9254d5f2be3e3469594e898bf827cfa4665d7cabe6278ee8360a8d59491a9c440a4c8a4f2ecd0f2cd3d8a8aada268db547f3a64b3b8702b7d21a95459214a4453f2635723dd9ad3b5447e14581bd6cbaf79c0afa5877b5d8fa9a9553ff926af8bdcf1610f29479689e2233768ab56ceba68ef3fdfd90abee88ad8624a86a9c72063bafb316790f87c12da2436af76f2f09b7684da3d819148b6577a69927edada94a5a560ac5b2fa761933960a22769be9607622a318a76fb84cd13aa881d65399577a01ccaeb9577a982958f3117a27fe9b87648521b3cb3e2b3b433a2f87cbf466bae080218bb8a58e9d58dcdec1ba463b280ce4771ba5086de20b5222ee72a4d1834fbb2b700472e6a9cc1e1a9c97573604b526b18ebd4f39f117f9de1054bdcea528c7e6842a1116f82dbdae31f24673fbb76ac16ead441061b79955948406c8d6a97ee8062be113e18b4ebf687f2cfc7066300e0ac652fb09c7972cef8cf3f88b166d00fc956b837fa844b5e0b9b799aa764766a02ce8163de087d5eb573fce268abe937b9e9d3eadf79a75d02dd476b43261c0fb5292c0514f7c499ec272f56fe36906c40c07d29b71b44920646c6805c0b374a6d143c211e035974156da339f588be59aff851e6681099be008e61687ea3566281d1be5404d1806d5e3f4403f9015609603879cff5e136621728c24158a4ccb5accc7a1b258528d99054f908bd12971e7bc457997ad0fe6537303200c7b91c4b4f0df03362b064d867e55a4f16c2dce0738e52cf1c0faee8390415550e9f640d00d4caafc60f684828a71320481c000fd992145e413145ea93ffc88653c10dffd6d6ce0f3f85e8501dc54624c1146e89173fd9628b7ea2d0b37cbfb6aaf375af684d3c31a6ffefd3a04904c702757bc93590a6a6aae62173e1e65e36f7d275d1856fe6f21a3bfa2c852f97fe7b3532c1d0f5e3ec4942876e8711ade6aaf942ee5248e22b2ec013e2223f60a688225b9cc328bce61658927557a0824982a86ba890aa94ee75623991f8bedac0d52dde7a93a216521ec51e85ea1f01bb548e660842690eafd60cfc9389396df8ef090e90471831f2da60bee562ade574620f300cd31eab8a054a33cf1578c4e527dfa39cc3b34b3081cb899f46d426a92a2b044d2b83405d2e5329dd338cab390e2b41b60b9a9446be9dfd768d20e504a4291c7f6813eed01b83f35eb9450ae102f7261a0ba023c3bfe0c7c1d7b10bfe52f36d8e053ddbb573b57aeef684f55f5c750598939a8fb21f52a1ef4947a97ef5ff5a11f1a9912bd84b6a304a38eff7e11a72e504cb1fe917e5f04f1458d070574842adb632cd3a1f264befd08f2fbd20f8833849a3e20cf4267df87d16ae4b4079095e787a43c9465865da35151fe0ac4ddbf63f7e39c127f7bab302cc3955ac283eb6573a8496f1296b6ec6366d0618514bc25f3808a46a508ef8678401476d06d30395b0877fad22dabeae22e9f9e21e2f49f3cc5a57dd06ba777b92906a666f8a769e1accbf688de97d84394cea8ac5749d64437058e845924d6e5a47e83275fc64c6330e65935b4c3e6c5f891a4007a23c3f2bb5671f1a6f6ea2535e2bf3ba5fe6285c6e7b765f8a1b8336207e5463c7712713fcbbd0f523cacfeec4805fc8dab626a74d16e1830d3b652dcaca6b8d3085111a9f138167268556d24340e5e202af37a3b6ed80c5d3a320d59d57bb71544a4d2da3eceacdacaf5c0a23565c15c29da57dd0bf0ec66a4033adc4171a1528d6f8a76626f7a96a09eb22bfc2707429ab33de3cc5394dd4ce3c2fec84be3eb004034fe944f08d71c9f14a5fd4056e348ae645655689833dd54e9282124d728fe1a5daedfa49cc2b076f4b3257683df5ea4ebe56bae93787cf1ecbde4da0548caf1ab44c2f4a8009e12475053f7e663e13807169cc93480a89e888f39c2a563043ae23f774b58edbc132c6b9b50cac94551a8bd38da23474b233d341763f25e486f8500b5d80bbb7327fe3e7d7ba41a5ec919ad9ea87221c8e2991e464b957ecc6627d93709c9a443789efa1e0f839511cab255433a87e03da91a1901056e33e86e93fcdf9e13be4ba3def57d4f1bf8e654ff22282384831a4c58f192d0dcd04e08336b1cc1949dfe4f24ed72748e9eb512d9a7121b40ef15e930ee08741aeb19c1332f97c23f0bd948af5196dc86282b8a2baac5a88dd83487165284cbcb695d1fbc6ac8630abf5f551a89c000a02c4ebd682cdfae8adbc1007426b9ca221093e7c9dd8b06089abfc15feed56cc4925cbd765a6cce29e051edad331a257bc899dc47b60d489c93796ea225338ba00a11da03b42e97a3fbd378868d8f29b1786d64c80e27a464f59f2c6fffcab994b3edaf37cac6ed2462f0bc606b80f837896ea13d97b6e5a8872528f88c4df3ade8f76daaa5a5f2950c11a6fb8396cc39a17b4cffa242a50cef083e9f452e008e0beab32b852cb82a408237ed1a90e57ebb95e300d742bbe67c3e1e35bb17fb562e8bef55f20d1286fb2b73dd547d868ae129a651729fa856a1fe255d6beaa20370c256b0b0ae83fe0280cd3fe2d3492b3f06b51c30f9020721239adc1387151b55da037289826972d318fbf47bff94df3fcf91c110112b8b267b5459159fe133;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h7b33f6194f357b4b98c37982f0c33b4ea36610b3f9e4685e667da9c546026ef17cfe37964bd0e23fbbfce607fcc18f1d66a4efd47ee7b291abc83352d15c16329e87ef3d5cc5d94fb8c43405dcc56fda15a8b584f335e44c2861996ecd599f0dcbf6dddbf50a4e24018b4ec0823e07c6f7d07a0f3668983ca22e3fb774f2c4d010e9c478dda17a97aeb04fe7fd852fa76d905681c3f007d5bc4ef9e5a245547b22d3e03a219eb152e75a315b59b646b8a3eea572cedad85b7335b79c5caed0b8df21015c6895b4c9255e9a534b8fc449c318ac22262a2085eb3b359912422bd5c8e2a541f2501a40382632f6695a2a9fd0b5aeb6fa8d60337974b2692765f8926bad2e0d969cd14b94cfab8a01212078f32aa0f29c7abd1b95ca01e90f37fec4421e8f05a856340cbbd5bdee1f940ec12fa0ab5ae9c047a689aa1713ca7049aeb560388c9240740e29fc5c80b2d5c309c74c1d0ab0cb337cc1777201bb4ecfd3274afbab1818998bf19d590f6eec3a6f7dcf0d417a3f765f13b021139a27dc023399084359ae6d50fe8cc23f60e7d78acf5b4df27143e584075f91d40d66f9d3405f9690b597bdf3f88e977b95a3ab097da71514764bf1f9521e2b2b0c9fc25790bc8e20a7f77c85fd38ce4ce0288efd936aa3de6f5081f53e208f37d0cda2d57e5a5c90f1b667d3754acbc59e8e60124a287f4771f0251746cb9f4cfcf1adbade211a09dbb5ba87913a7f460c598de862a8b6c9078a2dd9d83949e3b16f2d5a90d97d0f0fff42428735523a6f3fee8b4cb4ff240f337a8da6612507c4ed649539682055f356a7b27b30e78ebf8c99f236eab6d571d901ee53ed7dec59ff22e8f5032300c22161d7956faf564c6b716a0ac8a45705e25ca75858e806901c79ed5bf2efd86f40fbd511eb3f4a8fb86e80600d04995e8c74e77be06c9458a0d17be1019ac3124da585a30331c61a08d3f9226b37623a34c38d7e01d5dac7ac2bab71b60747e2713ae004879ca4f2e87cb0288aba3d87502ba195bf2b6fc50ca177b5721584b39fb416b51511753e7ef1ff54ffc0a4123220bcdd71a35db681322f7fc49940ce4fdd3297c939b78ae1b43806180253678d441e8008384fce2f76cd8bc5dfa61fcb30df915c843f03b7f1a9c8fa4c4e51f0889e165f9fe5ba37fb8b413a1b6f0eff40935b8b4fa4fe29e59aba4e3a4c44489bb1124ad17421a8c91006c4bb9f5c7fd5b7ecc89e6d7bc850b7ae89c998c4fd533bd2f565c70a03f4894547a7fe01bcfbcc6728c23aeb43711bd6d9eabc75864170ec34968560ed401cbdfc0ffa9a3581d1b7f939087e3474dead5356dd58716b27597d1e136532b41920989eadbc3d4f22dad079e61bc8aebe570faf28831f56db005bd70355a7f03fa3e7ca4b5e6da7214b34cd4884826bcd3bfaf2111a7ca8e4448aa15ae7c60e4c8828704de50826c1d4de0446b0621a35237d22e1015f4f266cf798a6f662ce455d5716942d42c2f7ab037d5e570487f91b572fad1a67c1afffb76606bbd33fe7f2b66f0db9cb5947dd2e26b8f2a31986717825258c8217c10930df7bd88845146d0bcf48184dcbb9d04fa576820d2c562314b4a0432fdc81fdc728c7472b4d34fd46403055a9f6f8202d492ff6f4ae3dcfd7b7daed01aa1e0898d27d4f2eed55b785d10fc43e382b35dc39795d8cf7ab785f34bab5eff01ad6976c552a71e6ae8e7976fe397ebef018b97b3455d72dc490f225a88bcdc92983fddda829884d41976ff1e7e1e6a51bd02a620d2753f7b2c8e6377c396a3787399a70235dc662e0671c862007f20f6876c3df3e232897ce804143ffb2b3c1bdc3279470840ad401f4bd1fb5215294e34eeef6fccc790b47b2de30dee7c924ce259894fdadcd05e96c69d44dff38cfe0ddf2e70dec80a6ff7fc94fcd9c8ba2035f296b6bbc251abba4fc7f3cf7e983cc6f58fac143f9b6a6151307f517e04c1cbb05857aed4a420b3c8de788934c02328032bf8383d05edc320517a7bc91322c4f0f2c294c83d2157a6ac4ddf106804034ea4b9062bcbd541c1be7756e36cbf8ac942f497964e04c71486c8bf7cc73fb4a323b27637cc97f8d4295fdf8c1e549c4b930bd94c7cd4594c9697cb45a7d8e1658df9bf2b3c7efdd4da0af69dd3dadda14bd27539f30a54973fcd29e67294fcfcc0d2e6bf05695e52608be69cfebdd37fc8d31a38394736ff9f34314891cb7daa2f0909a020fd7feac7ec1a3d16e95fd4a5142c24e1ec994236d868677f03a749b63c082475e8013b112a292108ffe151e68c32f799b907f3c84f7d160262b5425161d8cf6654b3bf98b812c71ce98aa12ccf30268e738c450b3e31b344575fdc3b30d8cfa9673002d9f26dc7c0cb8ab925e5401df5ce38a8bd182ebba0eafee63aac8c00904df32e7087b88dd55883e4bc412bcbbd5b31a92383dc4646ac9a6527d103343919592b701ff293275406366115d544c7c4cf0153319afed898e5752f2052e2c1c02a44f6819630df2661aea284729ee27271c5ef0a4a44ece04cad8ff4a7d324b07b84adc3d8f1290a0e12ee8726bf1f4e7abf383a311cb6dcb0512ffec3d4af7f2d330974da25399e9399e631b27dea7aacb10d7d4298b3762bd3b5c18fbe345eab5ef086c003339f83f0178385474bc1fe6152e8e915423bba4e030fa745b2a7a1829463154381545e1340e149892129f0f81b3c07c5bcc3d384bb583440f5c710827cb3604fdfae3a98724bb1c1e1815d9f31d7faf47fb0b15fe92a5a40749dcf5514ecdf0ae9edb88c2cb7925bedba4991b74bb63bb18b6b561aef249d92a6a11363a75e2eb0e77f1acfe064f195debb3244832d7edc602bf6bea6f2d7f1bdb5034fb3026aa446b1d9c8f4dd711f7683c255ae66cde0f66ac6d790716e440df1f1bb0045e6d6d0cbb66b6e86bfd49b2beed47953ac782df01da33a29a85fec90b822a42bc412403d70a20863c90319c3c31a857ff8dfaf2e4831e3c936aad007fe7fad213397580251d5010bfafad2faad82dc7c86dd5d41350c4503d73b3ad8079db045204fbc1f3c112528d27243668ebe36ed9b72a413054c045c9751886dcf98e4d6099c7e6cfa47f61be2aebba743d709c70c16b5a731f4fa24f9a2725f68080dff55716deb19245ad2167ffaab741a6d4484a61ed710ed16738d355b119cc832d4ead82358f584a44b9e43f2cc7e62a72f3798910faf5397853e97ce2fd3eedcbee785a535bb3bdaa91749d6b0b52b4f2908d7a7782cf37493b5df79c88cc029ef2fefa6d32c89ef8104d4d70bf1beb4e138050fc1beb3d30bd353448e96837f0c6cbad20a0f572c6d9ff9c4c532a4d572f76c02c27ab90bee2531ddb8ac0f128736cdd1edec80bd821febb0b258f2436a48bf4f28e00bae620e43fdda9d9b04292806187117a60ce01cb269e97649394d06cc7f6185d91b47df522b788a5fd4a395a6f114d803058cffae6ab6ff21b0fa48da64e0e69bce8b72b622e9b6444488347bc3eaa909ca32178377145a1f6705e1833c0f1dd9b9bcc0d590b73e1302ee17177c2c714e5cbe69a44d361b6237b591a5d5213c9953037c7f0b22cbb3cfa1ef19e347cee76d445fe00df05d79a4c7a398d4cf067d964d70626b17e06d8660a348d157ab42311b1f44f79b92938d9baa4d58959fd899c155ea75a7405f3c32d6542346af5d2061b4a621fd91cb8c557471ab6d89eaa0fa98d6e9262769d4d703b90bf9afc0057112b2035a60fc019fab19ada48eb59d46a86da86a092f22c271eb29d91a28bbb22edf6dc855d1d79550d3b08acf225067a0713a4435008cd40868f493fc83020c4d3aeed30be6b5e6704aa3947c0a48fc90e3c1b06c15041915b7a88f52fb695323243d20ad3c3a0c21a6cc9e39d33311d9d0338d1449287200268ff9ba254740af9d5b8f9d1840fbb7ec82be9f128c746f6083c23a788962eafd207ae3d6ccc809a9b6d14ddceb1b1609480fb8e70351ca62a5c665bfd72f59eda8923d8866a6eb89811d916a847807aa8f5becfe20348f4fe7be046066c472aac1ca328d9c014a313ebc079b2a5275542dc4049af157031a9c33804910faf5e82bfb36f39524177b7e1aafe2b522bab02a31228d9ff8385693cbedf32dc315b1152fdbdff7eaebbf79cdf0d9ddf9b770e88faf69b83880a96fc9e5f9d52ae3a5f9cca9eac45fb7dae63316356553283c1c7cf9a82609ec09e194feb70fbe9569278161e961420d9e5f649697443d852ba95b02a3d31d030b821eb5ecd3c958429aaa7808d3794bd1eabe8b7b3301282a236b47be7cf7b4b4178bbeaa54b2d989d48645a609d2783dd3f9552b441674ce62488eaacac327352b933d51e4a55670e54dd3570f84c60390d3b4fa014d6245e34c47a5328b49a687be0d38f17f84d1d1ed6b523d090fd8724cbcf639613570be9b27a744c4356bad4e9903785d999fb064f8afa34b1f08846d808ed68fe9501f9392b939c9c18a642b825af94682054f220ff0060adbf398b7ac60454b36359352696d8b9c6e1c3090605ea9adb28fd2c93132205828514ee4b21c0c7ea0e1a79fb1a9de87065a27805330fc2bbb4db0dc77087aa38b7f247c64f399859abd83c6997ee05f40a4201585271bd51ab27e0f578e461d4704f9a6701760da185d4cfab6ffc40cb5b520c578cc987cc9271f2fe2edd9cf510129f995df339cd483547e78f0ecb2a70711d6c964848475f8e63e61e5f50dcd02c69b9238b0c77d078000068796aae99d7eb01d1181a3cdf8aed9ef142459d6c6101bbf0b5659eb30516ecd9fed20ab0f18ea066eb96146b3c78c5a214e4f30a4e1a37753e7428bf4ab84e8eb4fd6a4b6d3af8fac6fad5d4176ce662650c191fc47538bebeda6747358e9c604be21d2a499821113a793c91d5d2995c2ced7ad40c9b9839c68dcfe4257699ff0c04e2669b22d1c7b0d439401bf63c033f58436dfc232f071e382f6cd41303df618befae79323e89d6d45d471341aa690206f27b85b58eee0e552bc6e93e6d7c1cbd4131d42a936344cf833dc33b2ff9178c37f26284b8c1563951b0601048a91f2de413e63ae05282a1d7c0a2edd5615b5e6d147bcb98b713911c687d411de975845345c3d168326b550a5705481d8af8a6a801be1da587b253cb9515901f0342b171a4b33fbd5ecea4b7cd470bbce3ffac1966cd55fabd9cb04a259621639218effefde58600c2ce44eca1636b10ebb8e7668a79c5de661c103114446c28f62bf1794c2be04291e2736b7cb7ef76673156fe84a73be4568d645f58c54b5bd2146f017b5db88adfaaa5a701670145c523f3c51c00adaea127e799ee56e705f24df65c6d0324e20fbb06d04fc0b5eaba77f08361b679cf2fdb483acc38b90a31523e6b5d57e33bbe798c7f91a32c5b4e083dd894ae13d32bcdb8a087a3ec154924c8a014c050e436cd4a372f749476428affb690ca1377c87617e31fe3f2358e0d5f9a9a313a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3b7bf32559a779b9234a2a59239945b3ee701a5d2c1b692549b3906afd6ee277389d2cb0432fe87867cda4282398c32ab737b406d8d98537a1ac6d5e2c22c87169dce675d611b4766eaacaf7ef7ac050b36a6e49caddb016cc922dd0255423b72819545e9238151ac39e94e6a4447ae3cfa2ca497a8b1ac26ad00b5e8accfa3100f45bc150a8ddeb9faec2131cf9ac7e51117bf8b0543bda73e639a1588e50da83b1d9cdd7a2b808f64a94e4e773aee2484067ab3670cbec1bcf6ba4fb6f5629db1342bc6098e9f671d597070ba756deda95c6aa9f397cc863637fc7c52848f67fbafd65967ffb7290fb694b8af359e817fd35e642fc3a7ed61c301f4bf025ff700d1125048a7c5e5a0792ec312086539bd47857aac406aa31f2e9f633666e46623552978791f02ccc0f536efcc06c049c84eaac41d4db6e3032083870e581da5dbceb86c89d597300c8d2d1d8668b32fc8efaaafd0820abf5b2d0b7af9c1ad4879759b941496061e216088a803f962c63f25fff1a52cee535a647e77ce35ffe32db7e0198397bb7d480da78657dfd38afd4655d976814898ae74074efaf71a0f973a1b4f822ddfb165a839326bbb6be266e933833340b2bb76f3297e3c9a4586d4226489d5646ed38cc9ac428f04ef56ba951532aaf666e42350d8f6fb4b5cf0edc5ad1858d36ed84d49f8b0d965a3759f9597b578102fc418bc1188f24fac4f60dc25761de1f62b96eb4c80cc40ce173e9f66f59a1eea8652cfc0b12a383a39ddd207076c3281e0103db7f3165a32b8c547c05d8343c0d7ac1021ee29edc05774b88a3e65d896978bd221ebd04cf34f3003933c2248bd62dd981823e3ec336816db42026b480deb69c75687c90411f6405eb06ced0fb40492d77705ac61350c5d42027ef59ea61daab7ba50066331c55f1e9351397d83b221f6d699a2a9545772087c5efce0877f9fc0e5bad44f2a9506f02fc18a1e0d8718f654cea9b2afbcd99664a6d3a8e250e288c4a7bdefb0b8fc1b35370ba29e5193217d4b77cb4911f2a25eb80fad87658be2409cd9d0f9efe7b54f2bc8853c1155d97ec7ba6738e755187d1ac804a507d9eb965e8d5c087c23e788382d15ef8d26a64bd75af82ab111ba2adf5039bb79d74f94136622de494a3c2113dc1770633ac6cd98884ca6d99c264c147828e9931bd97afc7dae5025bf80b90cadd8f63ed11131f5ef9d81135d85a158c56cb475790831280e0dea46078586056ce6e98275b5f9e94e596f6e123a1442ff7ddc5105af25e1414c8bfd57e048aabd8f3f2461038cad1cdf6a8dae3febfa4e5301ea76669da427c3869be1d74b921a900c523c7afebcec55c1b1030af911b11db59185194dd41adc9888fe22b3edf76f82df6a1e225f5e3d4d52500302cc6ec259bc87d689825cf83e8e388ac5f15ca05d94bf5083b561bcbdf5d47b5b3b0307eac5a20547dced6c94ec9fd09d85195f5b72d3999297ea68e2d26adca011d523cbdab881287fc15172d88670fddb5b7eb5ad28315255df4f594a658e259a66d0fa15859d87e8f70ecac16c147ac2b96e11bbfd1ab774d40ac3310c73a5ee8bbf42b5f5fcc190b02ee4dc67a84f98c54853785c4373ad31c147090b83d5adb65da4e381f860d22b59284d3b6b641b4ca2ec727a63183529ce5b8902e6d73200a081281cb0e1f18aa357f6e3cc019d23fbc2f4ea4e4dd1bc3fc18cb59bbd73f8d798c36d086789fd6d4e63e39caf3b26bc033a44478b6bfae6cb7073f3073d488f19cda248c8159e1a54fdf3094c4adc205c1c84b8da1cef649b64811f9764b2cd12d53d63e18a4dd6fe5d260f5fd01354b754a94098ffb80b1a4c08b09fbfea3d865583452d21422fd517feb59cd60fbc5d7c08efbfebc587f81779b8afb16e41a9720c44ec7723736e653f42e6e7c120c07cc5243763b49511090e4b45937936465f1685dc7537e88d15dc318b78790f3d6b48767e8cb42fa62671fb79bcedb4853fa4a0a60e26b5430acfb89f7706b8d0bf8942d199d2f20bec101b954b46e76d374c75be1acdd7a295fdb0302479ada6aee52e7fe803cd66511a34ec1a8b3b7cf003b3c4f46bb547e307c12e3cc0766d9e885c14e202c625ed54f6f9d3ff58752906f836c6af11225a55b16574687b778793e0df4e731ae17a4af5b5445499c6a4c460bfabed03636c0a4c8a78de95877e437633bab561dda93c9e01c4c2409ea1fffbe4821ffb2c92111364e3248400f944aa22f70866b7af39d0f53d51860dab2f6cddc52ac6bada382f283434f9c53078155f189aecd6d090b50d902fbb74f86548da55af3406a3020ef4942aa7c840822cdc81bbc2d1ca01b4e9de53c4f40f6f2c55ed86f666c18f7a2c0c5deb77d5b28faa0681de110607333261442fc828a0f04246304c7276f5e9bab1c1dab7f93c7b212767b1b39fe703daa03f3795875bf03fc8e149decb82d2b49a327541f76e0dceb427180397e49426fd1b1b097985fe4f34c8fb1a12fad7f2499134d0745ac1865915760e14890d81dff7295b8c8da192083d696303fc71fe9f79993180c3c0029ba3c249ee13b5e7aeb5d9ab1f00518d93ee53b4594c71f7a07f19cf94eb039d82be2e14f0fc095a18b145a98abf1bc5ad7d3acb58f90f1b241d582cdf065c01852cbd1d17f60141993660976b28ccfddce966c2e2963deda748d5472ad18eb5bf7cc22176287c1ce87ef9e2d6b4aee2c95a726cd71c45d574d927020d2ab51aabd4b182056bda4052cdc062f79fb00e2fc39854d602619016809c6dd2bc712cd6027352e60619c6d46e5d199f6e65d7ef0e0415b656eee0e77c3724cebdbba99f04e97f54ccbde8e59e131b9646bbf5fe54bd62e6bd085a61bec7ffa22b2ee64c6756cf905e4f12af3f2ca435477a1f0d81b227a8dc95659992a74cc098f4b636e9dd181800edbc610fb7cd4b3620ab3a2b40eeae702d058e98dd6616bea48368c5e148127e72eb1b636c2ea9ac3e2ee2a3f733fec9f52a8174b86d80f5148f87d0536614e70fd49a3ac038438d281d84cf06371894ac716314becafeec2257176eb33b5d375a1323196e35d1c01990ec4beb8eb5ad7a820feaae045cc11fd0b41ead72fd3ccc9bcaeaafda323b12371ddd276f30ba661f932c527cfbcf4562d13527355b8a2c729a78a2d981152e506112cf9bbdfd3b9b7f3f7a426199c0e62bfec073ec869bf966f443ac26cf612a198c1d9ce0512624eef9f453dd79d0694f35343bcbea05642fd1533be74da09be769dd2fc7dea13f3fd5a40f739da8fe1102a788a781cf094c5c6230d5fd5cecd47798b9ac172fef6ca4f073da147900d9bc12b999ceaab92629cd02cb163f1cdf77176d699b930dd7110ebeb1749d49b7c5956c748553d8d58870c7ea56a403ec7b7963ceefe99c910d7c407fc21c2a6fc7fa9fc80d94d13f08eb11b64b0a9986c51d3a5f70f3a507a0e29db305768defe83a898609f98e09766b7082cd5e195c3aa646a1ac64ef1782d0ff55e1e2654dbd8567a8afb1ebb07ed36f9051911772a03a5864c986f711b8350a7ce49d8ec27adb53b2196be56bbd3452a787e57ba5fb7ea19fb565ff3fee65fc2ec7a19483975dcb21f802d958b25c6af26b481a87e06c8dd6c75ac948c3aaeb489766297c11968ff4644bbd0067959ef9a31fdceb99a518f21293c61dbb5494fd28fc96ad236cfa7faf9835cfb109687b2aab6f6df3dca9bacd7ebee1dbebb32c4faed21b3387ff12bab2aae56f4c3232b7e2681b325da7ef587a736c31abf24979641eae4fb7e0b5c72309f9b769efcc040217c4c8225f9f5a9269e4bb0d8dfb8c092c11a39da8f89f0844d9b2c1942a22d6abc96569dfabd62783684cf420d6be595c4bf0038e1d8c8a0b13c6569181460d1fb21021e07ce81a044b34fc6cb5788cd356a441130722a210fc6de1919e18fb8f0519be3871c535335290707c2ad4ea7171b336925b61028ec674b655275befd474b8c4751e92ebefe692cd1a44416bf763ac5b069ffefd0b9fd78430e0019ba06584264014eb7a490ce7d8941bd059b04755c64a02975a3f6ac4bcbcedcd9c9bd673ecb37e03dd83c87f812d8f4b23810d70c42bbaf16a850129c2253dcec9ebb757b401ffa86de7adb42a720452f8cc01af4a9686d2a85126613a6673ee086f212db2d6aa27879cd23fe90c55d6c4902ea24185f5397e46a8503f05fc3dafef10ddf7c1ebf05646442215dbe99487c8f1991e1b9bdb105f71382d3ebe679d975c293bb55bd889cc4883aee34683330808039ad166d7c49fe06df18c780669e23afc430303bf8169a1b96bd4415a294ae014781174a0a0693a9d891aecd372c4355f2a22607195afaee152f2c825c4623dba65e1532c4a1603d35636c06a42b91f2d69627c802be253d8297706e08218637ba356b9cef3c77ac808f3cc4c1db435031fbac8cd8a352840cee3427c8ad1ce11341354974c953b9882f1d549368aaf97ac526e84829beaffafbb0e7c7d2b9de0183c8ec7e251c98cd28a9f26e0671170223a2282a54aa85b1c5b8924ccf44cd6b539737fe7bf1cd57767fe351aeb34005c12c500010efde6a86ea89680951baa9726bd82e7d01b1802c6e13450849ff0d81f39e68fd749cc0f568465bfa78b1325654a378edcbd4b439f14af496b0993b75663e5b423a170d17d48aceee22906945a32d4d7615d00d93016be7e8957fed7d5baa0f82df8ba81ba527326a67150a86937931776ca996d03ca921ec40cfac034e0d81407fee089aeca6bf8800d126ebc3eb736fbb3854f65f9dd7ea53fd4c00ca2ee0cdc662c19bc60493cd2133e9851c1a175175b917ed6c18180b1a187def048037ade763eb667a5015d7346a3b5e1509ceddf8e711b003b9033cac4ffd20a84d042b28779be895805c65b3778eb02649bfb32d216877e801231544c5cab7dd636352788279fab2553d513f7ff424541f5b91e2e9bef8301c2c31c373aa5546bf4b06155eec51467cc8a02a7cb27ddfbc0732ddddaa0e0132a93c810f16db2f33daf15ef55a6f221201a8d621e5740c1f12b433e2bbab050967f551b6fc864b39fa0ae81c22c18223789286245733264c9e29927395e8582c5faeafc010a0053079e1c52482b8c4a8e8abbf1c3ee420d4b8be5377a260f2b156a20b9d9f766a75eb5d1bbe78668227a7a63e2d15ed354cdd882624eb2dfb437ab2c5ceba1a97622d1674035411ccf5d04122b966ff3782ce776c75ff8cf87a2d56f5324dbd18b86923da085df797665df0f8ae729870ae1ae954e00e0cd559d28ca906bf53b98c58bc9c6778b8d33adb3f948a8766f86ed75158edf85963fa1ff73a7f3fa3aac7a8dc3d87216ab7eaa82302c3b0d04c2ab6aa2cb74852984f9ea054f69ceec0f924cea3f7d7fb967cd674a20f8776207b3825246b7ebfbbef402e266139a4fe704c10276904c0b6b03310abb88f210a0affa68383d26f46d5e4db90ddc2f63;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hcc1e341a2a995c3daa8ac2885085f581312884a41b876e43cb089727a27c4103e45e9af2f181cc8fb722108701010597f910e0684e6be9d5e7b780e89ad100e59ea7ea374faac0c8d18a7662b49251a449ff7a595788f1caf5e71d624208e89804987e33e47e57e307899a98fdf2732cdde92bd8c0c5764f1418bd0d9b447a810c70969e4e0e4b0bd45455742505fb45cc5ed9641d7edd38e1bba9ffcb5192c3b0d8936a490ac99a97d342d1e5561eb00154281ebfda9b33d8532556113c15e31723af38955d885a9c1560b1efe0cb484fc6a45382e9449914c445eb1ed46fac7b911fd03b2d1505709066f948385a92fbabd53fc4eddee4bb0f8026472bf6a486cfc4445f157e04cdc8eb034a1e4f3ef637aad9c2794fe9ae152334a231cb4027ae444ebf12b99eb2a558e580de6a93b745033184ce9a1ab1667b3c84f86832219fd13cbf0ef02844b97ade453a42890504407474562d43b7038030d9a7ed2ed016221a6ad7b3ea68c903065a282406e526718053460218ecce5a68f2408d429b0c5ef421facf040520fd5de27ac3c3fd45d4735368541e577aa00aa428af2633729d9a0cb0bef6cd1dd8aab8840b67bbea21154b2314d1fb83a8f9087271ae14b8f8d33d950448919305d6c00b2f4f002b786740ba3eaed6a336416f5185796bf4913a94f92885378d8b269b355f321fc10d24d699a8a2b1a63af1b903a2c76ad9ba734ca7a4e5adb13f4bd007dc3a30762dee71d1d03de0a675ae6df26362161d6d87e8ed19d949f1973cd27c78f2a3d9c035473299cafa2593efe36bedd12138ed1b4d775e11c22cb7c863af4c22492d289bce02e2a782431c67013c21cb53a7cc9b8ca3514f089613dd8e5587c2e965f221c8c8101383fd7f1085ef64c34e3db2635ac726730a4ff0b06a0a97a2dd6bdd48f6047f1574c75bebe95b99586f3031c375d717c2e59b0f7938346762b36c6fa5995aef476e8a3a1081130515b6916febfff2f4225cca4b49cb34a9f966347b53680ed46a8bdd78bda5df09b4ebcd9cf8646eced7943af118a04c8341e07e1ef352a828367ef145eaa63e39d3b8c39f9190591a50aa017b07d61126a5d39f7bbd1877aebbe295a8588ec30db70a0fd0ad36ccd4bc35434d7b0d312ee56186bcf8b2cad1b05374c9797e54887b07c2ea074115ff675499ecd4e18f104201d74e9771e7c46178301e6d724e9edaea95a5023f8a2230f45eb8c179f80bf0e49e1582b5b1ef7f9bac7e949eaa874a351d779be34fffc7c9a4117abed1d3da90d4a6d68f4a699d2f70d443345a379975749dcdefeb2d81be2ad3f388de21fb9004c4e1791a2f470e4f3e8bfed1e3d171b7b24a45424061d04a502b22a138724b02bcd0c2473245040aadcedd44f4cf1d2cbb34156177d8a9c33adad0c15790a82282ccdc040d00dae6402ed0381ee32d3434188f4ef08563d4149b81da5e5770643a7bcfaad9b6a0de5c505ce3f477f851d62cfb8572aabbdc84629e4fa8e7e0ab851a64664c6e8a85e757f1e3a15819fc3186dbbde54e4179c2b49f032bcfb2f849a52d34b7d8602304b1d45a05393d6d5f666da54fe93102ee9ab04fad3a9b9e893eeafc23eb4d4152fbd686000c50410057804d96337792315ba90e2fc57bd55a99ffc8b0423c66568fe7a3e81548d9967eae16c04d3eaf9a3b446f03f4de1dbb6f2032460e54bf1642fabdd58c1d0de9183d305951428297e2a13fa5f5288cb9aa57019cfcf946db2cd0a8439756ee43c665501c8a326c72bebefbe5c446e9ef8a82287e86a37602e62952cc258e5aaa1a3d690b6bb62e8b0ccd7776d0fd2ae745bd6d39c5f5382921687b172c72b58c87fe18dfbf8fb08ab29eeeefea9b272251bf4a5d15374cccf8907a66385deb2e1a21f3d6578893862d76bfb20a3681d31129a7931042fbcd74426c0193af9301faf313a3e9e69d4f9cd9659255043cd62de6be3d588ec59234770d8fdfe46b1d7f5c8d8d2579bb2d098a73651300897a7bfc455847111ae540345b607f28b9a71472de52d22e8e05fdc67ab0f9ef5112e21a42379460671f50991cc25659d738cf9a8e90df1117c40d72b8fc1bd14fb96644b8b8921fb4486c36a121e563cec30c6d7ecbdf04dd0e3b22868a1bf5f16b6a40211a02e9e71b59ba92e0e72fef7827512d97ad9892210992ea3947b33f63d9dcff1dbf330d04bf9b8937851dbd9e1c7eec7d5a3b3f7e56dd52267f1c0117df8ac980443dd0e40688335fbce60972c8741abb03752513744dd13eaee7fd329ca99ceb6789b8762ea86a2b28386ebe78b7209b5901231af3ad0160d5ce8ff71d1c20d91c7aa36efa4bcb2308accaf56002d1c1d1c1d131243b4485d82cdaf7e21e1fc7315b26b775a0cb6d6835d61da03ccc9266b8fa8d33d2d9c99b46f4591a238656dbd25d1b0b8c529092f4a67d55729de0f1cd9f8224c83059bf4acd1b0556ff6eee77d20c1a62f0a3924a7a03dbc4b8be674adc6649cfdd1d6a4b5157ecebdacecfa74fd1454d2ade753da7c800874dde5f77d6e535e7d632aae9a783450a35a270e85015f82381f84218f1aea6764320510108138e14af6e364bd8e5a79646d3f428fa074e2f2b4c4ad70d9e77618ead283d951f98d48acd7d04c856dc118100748f1132c89e991e4023cc44d280db195856e197b1f8ca5f1f3848860987cd7fa51c1d53326ebb0ea2eec48526aae9d6092253e2142e4a86584a812940175835a20ee524e2e05ba21c9ccdcc5a50d3c505013048206e41d0b1f1ad4a3307ff56a3d9987d41961720b5eb4c4d5380a312a5fe0e15ffe4aa7bd545ad4f888ffb24964984ce9e0b04e183266ff21446dceaafd0ba59801b3eaf64b59f38645aba00396803864fc5927034ad17c2bd8387c445c7befb4d4234005d98977c46c81922f0be06c9ee7dc574c2b83fadd7e8626a8f66c0caa8310bbdf4d7970862af23d5e83a5a91dc7efdf4a77eced9222ce95ae857537f5cdf21cc2e73a70623006cfa23be9589f5de9897f70493c9cb51b6fd68bc445fa4deb15e963af4d5726db5ca2e5defaa4214b43ce429e9b063a590bf9b051ef6e9c638737f96c2393237a57abc303a784eaf705a1edae0a437ad57a0fefe72932da32221a80893c7d4a6f31256aa052e48721405065ed0e012a90124fa50ac5636e27a824428e7d2f2db24e576ac2123a871bb5ec445863618d886b2232c8a0947b1e20df93ae8866b33d97e48c4ea32dfb42fd8dba6a6570b044eeff05a7da8bdaf5944a7039457c97147ad388fec78acddd10674106a752578f4306fa607aea4589893b2eddd8e4c8a92e134d798391989ba53b139fe18a0c523a3e11f64954e14171475cf61307864a3767d5d03d4294548595017fb2495e3683fa0aa8ebf226fe23127058447f7f7544794a53bf0573d7f4d0f62e8dd3dc715fdfae080972d7af7398e885747a980e379e1a77dd99c3c2f5077bdc5994fa37b0aa2c154cf941848dfea97967a34c22b337e1730bd1435ca6b87e1c3e80123c6cea90500c63ed2f2d26dfb85dc85b9e9d3c78c29694191edcd293773c5d19b7a74c30d855a6d44b9bfaf6147bb13ec3cb8749c9da8e4428ec938bc66e7fc426d22207b3df657464bfe63c46d3127f465e03cb0b74d4db5d1468cb606fa635112cea1d76d6046e9589d498deb193ffca75301c27eaae33ca7fb6f83ee37ae7771b02743969c3008c14b5b1eb0b89365d01b52011897c362525045b27a09cfd34802f7bd1578633d72ed9968412468a04fcad5246eae05395c5b3b4fbef2d0b7a37a2bf82f6f1931b10a76c295218a62c86a8776d82823f361a5e231c1f7df1864c88a4e97d1d861f4bf9e7165736940f303a5c4e3f79a9673147e6d9f0a2e7e239219ad8deb2e0fa0a73b48483c7f410c4c230d54b76cd17fa359b81ca9e2b7b770e3851efb54b89085302980d284b6b057dda9fffce33b33a59c0285d976c7ba5f650593d610d597b366862d254f80d95aebd5a11d2d0e1f5a4d0741279cde3de2eceb3e38a158a1b35868ade5a12d64ab8dfebfa397529cd5d36d93b79dfac283b52b4485a60459ddb73f02278e6a5cd84d5a063ae48a1d60bab54d1dd7fef12769dfce753a514fa553dbcfd293bb15efb293bed38a51a58bcac8310134cb206b4d0c94e638cfc9632b9418b63abd35d644720c3cbc636f6f5e9af0e99d8a9277528418a8608995dbf531e2fca994bac501d515aa0448c8f5b510d98e9d575802b569e6b10362b7780b59c544054df2f6b81a9caaa6c86d03546fcfbd4816132d0c4b91c73e373ba579d014a26e75ff52589b99acf26da393bbfa1a2467847564f04d8d0e61eb376de491338aefb48d06cd641daf04b5b933ed98109fe661dbbe81a414b379e1248f3ff9358725739e4ee6353a9964e8ecb00a259426cd3a04ffd41f4755697bd27a8c6b46ad0c7eacecddb1acfb56f0a46ae063072783647d59cdc7e2cf500463d516b429f2bcb6e7115648102cdc7864d0339774feb433c0ae948f0dcd2bd0901b7d1f0d92c47be6ff5c798412916c04392ec77706ab9d815277a68f9fa3e3cb67cd9dab28f6af34cdb872d236acd6c58bf23b1519e196bdb64c07d37dcee6a82daa87e1a21e59aaa5bb428e632578fda02ab86da5cad45e98357818ab6ca4329cb335546e3b0be0b31cc62e55d11fe547f0ff720166231f2e00bca3742433772fc41e102fac7d0929126274a5e0794825b42f8830b780b6a8f31cb0a60f96577ca137667d2d99251aafc2b8a0ee3d938cf0ab1f8da44f8a9d2dfd111a40335a29542ec79f1bb8aed3058d46b2564cecae32e8feb1f9f2c4308980a7e642db8c7b30cf1854bf9b51e5f3ce8132907772c92ca2ce7e0de8dd30ff12e5f606f331e120c692dd4e79e5973d9198b4487a2c95bd644a94b636e30b53a5eb34c2705baf078c60db27691f2e0fa50b409893535aea610a183dd83254382c20c37d11f0773e6b1ea9ad6c9a6018fd15ca82e4cce601e315bcf0ed58ead7638e20d77d096fc3bd517a2863f70d8a20e33e016fdaf3fa13903ff246433815d8f804cd9dd691d434ac999e68ec97eb95449fd2b2322eb333b68cebadd90a6d8b8e7aaebe1698055efb5ee65290b628f72c2b47827c3ab1f4b4453900feb12c06bdaf7d0bda06480e5110d6c23fc01f8b46469a8869d07489c945ecc19f34145fff2db529b4358d143b07a9cfc5ce9cf6f476f83a901c5f9f1f8e7a1441e6f77a8dc0e5b824d1b9ace6fb1edf5f34b5ff375a4fe2afe63647dd3cd5b985122c11394a5aa173de2f347754b6ddb98e67c5816a4cd6ae3942e9943882f1554df16d263152a809301922df9195418bef6b04a1412e19217e5dec595a97a130deb6869f20160cbca2198306a81097f8c8cf6e72a0ea177db8abde2cda4bf9ef000479c9d178d1af975dcd774f5de5a642f9aba786a190cb4b1f62eecf4326fb62263ce729eb824497f4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h24899f2da302101b352c39d209d1758ff9efd4c1bf76508ad134b297ba9904ac599df5d4e73951960113f73b1a24a142b4b7525cb674ec212c10a503356fe7ba64c2335d8a2709f0b4546cda0269c1c55687b084c38e334719aeb2ab6aaafea8a090c4e48d9aad4a352f2cbd422cf9547d77eb8fcd157c4d219a852424f974b8d17ccd9c47723845fd2a2e7e9c7ac5d640187555f4bd527f1ba8ecfe7344aef72c548936a3805272fbf2725bd57fa7cfbfb39ebdd560dd8b3cb2ac81391d280bd640db1739255bd9edce859b2d9f1ac5b3c96d44ec1d0eb44983423f2df23689c909d2af2e766a243d693aa83496b012d250825e734a94ef972a580c15df36c86ee923c33e237aca3a6e71ac912311a30ad82aa1e7825a4587030fc08e6daa23a8333054bd9cf4bc86515dd0a099c71f086fbc7eac765aca28b3e746a85d7baea8ce98ea76d0976401e49fa2ac83e11d26f1992171ba06ac6ec692e35684b22614b2433f803d8849e601954f8c6553fc72e2ae20ad84cd8bc0066a99d4effa22c2f1e8ee02574d4d6a91f9386b7748f23df06b45e2ab61ed416813e5b7c837be002bca8a4052508da49d5b5e104357ebe28d248e1c322ef965fc9fc83f5194aa72b05c63eabb8b4819217f86452a6415c9c3be1df91b0f7512a8fd08512c95cac6c5644bb761f67a21a011387ef34ba0f9d893c6fa76770d52b795e69275a1dd04dc97751e208fa9997505ee3f3740ff57e6580f8799d745cf9afd1032777d699b890d7e6d530928f7f2373ec12c757439a9bd9491a4f7705ea21438aa5110120a693bc9c5650c53fe8be671987b50dcc7738866dc96e5f6a33fe0b174dc32e7c93a663ff1f7b9de159d59294d24e9047147f3b8490c20ebb3cd544b64c77732a53c991c705344ef3b82f203c388295046537bfed276f00f5e4122f822640219e741199c307235965fa7c616979cf16cd32601ea4ebf860c652750b287507d70d96590db0c2ea6755914335e5901eb8016457b3b1002abbb51dc255da9028ae9cad3ef47aa047f24aff39958dd2cfb883dd4687f7389a7ee4f58b45fa8f08d7f43d63f83dcd862bbf4ec2f9dc578a516ddbbc96e74d27c562e8334bcbf8b6cfac4897bf5e313a4a6cd5fdb45693c93083a4071ee30ec895ca21f1fb9b5526c14b9bb0e69577216150921da0c13b6cb2dcc3cb7ca3044c8a27d820e5ddc1042c6c96f7cc47b4a7c390fbfe3741c8594c5ed727918377bcdf1d98a6eebf5c59abeace13b415e82caea2477b35d3551653bf7b375ff9161c77ed066994ce7ba71d9e9e42d95b4345eaf1796aa0b3c6d473132a716a243742494cf8894f8500ae986b6dc008820eaa04d19aaf511da9e2906d2a05582632ee984a1e52277b972cdf55acc1e92881f35b5064cbf3ff1649495fd2ceedcbe7130a1cc36903f2b473a15a8df55124c5e1f5e5fc7893604bbb86f34458d1dfe9fc470768673aac67ae554dacbf454434440077cacaafd3b6b133761304711f9e543edf017abab0cff7ef09aa914e69dc05635857371d0851f8538320ea1c0fa50b5846c40261cb49ef3073b79bdfeca58390742967ce4920c123d6126385e879216450188760fdc7cc26747f1a79f6460a900a4c762f2d3507396574ac449ef1d26dece28d7f341888fd6d3dc9e42d461a1d8721c0392d33d0ed14c4733e0220a1833ee34510fefcb3ac8566bc9d12ffb22c118ef4b90c4098fb70eb9cb9d045eba71d9735e1152c5d8f27de01d795dc93387c4ccb413a736023142cef1de9c17d3eec571d8360cfa674beedd768b5f1250512664bac8bc0b1069b2a11e49829f8ca8a72f88ae7b5cfd4cde94806e1c1bfc80f6639a181564be335c947bdeff3c1c906f032afd2cdbe87f031f6d5347ca88bdc2a94a0c00a91e60c25c6e1bfb973a3fd06bf31dc3a948f113a7db1b30d17b9fed9d7dc20c746c14a4ff5dd256d0b9f9f23cc5aef7313f48398d49439ea50a5d9fd0d155c37cf6a9a97d72a2a2fa4388adea447b3d91c8159971fe3289a019e051105f2ecf6c1772bbeb1c1199405d53d41b7a02dbfdec622cd30a3b4b999e4f84f1d0ad938e81f807847d54465b32107d003f2a3e4250ac34e6bea2ac767837bb8763e0bcf42b30faab2e5edf359e83bda4f83c13b01603190453a1b17cada95facb11b2b3eda853cdcb09a5e1c63a310cc3c507022d03002435c168fcf57322200737e91322f51eebc73440c722a58513a0644da8e7b47e34d30ab9dad80b4b22a179b8be4dc5c48c4032d1e939f20fbe03395a86f24ecabd6c1d6fb6b14a9de4664566d20f4ebe48220b8a068beb41951c81878b1d959dfcf0114496358a08c1a10899dd4449ad601763dbc61cb0278fce4ec83be6d6e348bd6a0357a835b0358d3ca06204409c1c5dfe116bc35c93aeab7dba97fab401aa40c370bd76588b2a9535b038b2e9911be8514f7f09a5c9ffa70cfe19b73fdd2df0382dcaa55496fc3e58afaa2847f9aa95dade479a44fede008cc52c05de0768bea18f863a946b842fd91ad7be5aa0f512b7c7c299c399d80019d7d62512d18a2235c1dc026a26390b394203b0033a486fdb265c6cb12b80c49c2ec4724d7b27c9226e0136bab9e918cd9b7050f60ed2040ae0d30922423ead6abf0b4b7749c1d8957d3ecb4be13e81b0a97319f8e1e5501565173f954aa7955901aee0476b5ca59dc0ac4c82bb9ff6676d646f042c57f42c95f3df1452f4398ca621b90e667320acd5fefaa9eb7b5208c9adf2d898ec37905ae741efbc9b3ae178a668cff48a4d84245180e4d4131849e9d535cc11c6cf144e8cd408281c14e7f3e258a9f1bc41e6d5025a31430202f9b8c59582830be3cb99bbe72a15c6f22135904d23044aa5cbf2364907af9e917ac128051ac598320582aaed10ca65bba7c9ab5a847c2e316b59fe9495f577bdc1f93d1d8e3e2f87471b932449eb091b67021861c1c8cf81013b986ed636b8028081cb7ddef24cc010b641b48782700d709e6b8bd999bedc660972edee02019a51f8eefc52ab9176ddaf57593b04fabbc2500e1d27d20de873a3972bbf16830937b67dcc403bbb079806b7d99807618cd03aac91d81f32e7279d5e33d130d4d1ca2fb52fc9528497d8e7fd5e82ca48eb3f18a7731a342cc00ad4bb7ac92ae40b0997f731dc08f89c7d6fd8fd23ed460de6193730c0b8476682fa8be311605f158372db82cc298636c054b4b02faa524552fcb415f033fbe37ee15529edd487666a13716a53b44ace0b147c401d23c6d6289ba9af52b8e6471dcb52f7850e49eb79931ec3ccea616e503efd1a62f93e11e33d53c3b6d030caa7ad7a737e97f6e08fa8c9394aeafbafbe97715f74d4b2383be98d6e872db76c682aaa1ed6290b8bdb7d3c45e6957c89633aefcdbb4a12da6eb14d514adb5d84ea7287de41dac306aae4ac0ea1d79de0434df612cb17ec4e8f6d542a1fa27c35c79a1938c3c00edc50290b3bd47d13d514a736c407ea2abe7fa9795b925d2a97e29f611a97bcb712d8019e029f0a86da37e70ceed519dacafb04f5d5de5fcde0891808d944fafc87bd1cefb47d52ce7d1be1bb07a0cab63e0ff8ac081a9596b32efde22b59b2d7e2feeb2154a0fb4a35831834114b5a27554d225a08970faa6badf8d5615c318a8faf02dd0f2ca19dfac3ebce0c53d9a6a428ae59c3a63e79f7b4c857ef48a56982c331e697da8b5dbc49b624ccc047784e280dcc2a1bfa6ca29ad529cc540e18a089f2f346be2a95d846998b96bfe0c0f4d9045b27c1d8252e121d944a520cb94c1387c4ed12c81e85d4f73a861f7a89839cfc83a2e3ad5ee1ca61764d27fe3949742f3ad6a1dd54c136e0bdf434bd6abde4127984c11fb7b2eed02c8ee6f66a24b9f27474516c01ad1b4f252ea07cb2b3611f1d95de9f77e82986502b1aa3b365d2994f38082b5a48dc3ec05622a56623fbc7a710d57d040d2d6812b33a243d12495b1d52c5b2dc11ae54ef96b710585043cce45e0dde1df6232c42ca1c289e71ae6eef9ffe568d19f194607c10950c9c7303f1d7834b1b3088c797df16aa19f84f342f8de68b10779d8e7ec139ad66f8603760777c7300d5555a7a7cab63755694aa499b7ee7b8e7721be64e869939d3f57d141eb49d942e19777ef944133bf30de0db39901dd8dab60892bb7587a77b054a3774da946d784aa9c09d438d837d5f698502b6fc255fe67b7382ca3845dc4c617a7f69211a77d505e8e8728e908c9a5f42d2b849b7832c5155f95abbc57a3bb68e9d6c226925b0b4563d0c9e8e095cf07fd532a66bdaf83e5af9e193283090fa0d7582405ebda9625e64fc033096a00b2e200a7522bfd88a1c34ed83fe1f8c8fd2784a2c92fcbe5a7c2a062cf8f12c0f77ea64102dfe5b5131dbcdad2f2b549fef8660db539b1e2e048098fa2783a3c44850f85999c65dd8767e8989d01dc2e21e1ecc9eb7c391db755e7a3817ecfcf84e293b646d81292fd71c314c240ce7bfb902daa381467d2b7b54dd3f4c896fa060f5b2abba03fd82eb2e49fd310db0b7e6148aadd84161bbfbb0ee926640787c692e9c873476c07e3831302b9cdcfeb928ca41004e61dd8e4840f4a7815bba109bb646cf5d3a835c65fca24e8b71a258b146e6992de3153807083e710292555df2c491a72fe195e2a52691290526876f0cf3b59ea3cee79229617ecaaee094af9f299d3b7a22bf7d92e8a760a5ccef4d2e394a93c3db7450e415117cd4c4061d99353de9bf33bc56d15d76a2f74a9c0b7ad9970f326569f49f9f00a9f434b66b7b443a09b269b7eb2db36b861e71d76229d05974bd1ed17f8afafa3aedf7cf337584fcdace6ad4b4ec3cbda06fed5cce5a8bcd7a1059ee2c29667833ef97cdf0f7c472a02bc2510288dd5b503dd2145c749b614f654eef6599972bc408a1e34d49bc9923994ca4343c86ba23b9cb6fc89e6c607064fc63ef50804d89a1ea9b004b07975d9793573e09df47ad3f6cfb8682551385b7b828a4f06c1338eb3b201a3f41219face495ee1386b17f1d614dd2138c27d2cb47c8b33c0e10b83edc49a5751f76db5758245b91bab6432dbc451ebf8d350843ed4014f598b5ade23e1f77133b601b810ea6ca6f33ea1139674aac00d1ddd50c3387085640203bbb84cadc29d1c56cb9c544e6c8fd69bf42260e25c4c18d6bbed156403aaa8e5609071a30a1d800dbdd8f0cfc905e141f2e4899c139763e47a9cdfa9619b13dfed2e83b37df1e4678abaecd5a04e0fcc40868895016b59fbec61fc5ecc8e2db93dedb41d11d52936a7e03c346480e3aecc54880241b89aed53884c1022fb013052fa4271d996ef4048dfeecc4c40289e52fee5f93cb66e3965087865cf172964835fb835ba95f3bd29f7ceec4a882d35b0e1ff2a3a173a07c4db53d36b702db859654fbe54f4220abada5de7c3b1b2110677702eceb6fa022ee5a147f9349ad6812eed95e4d5525a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h91c7641f5c7c861fb557d13a1e5d8dcff6418aafd78d73ab908093ebf5d6f334394d9b9c80da51f1de1d5fc9436b111f39e3adacb1350ef2748db61926a091fdb4d587ae4c7b2ec3f78118011bf2f937d24fd3776ee38bb0f3b156a9479bd916058f6e17fe1130a0541891143ed5dcd6a971c1b49be0855a5c72e32015b109bb458713bd942ec9f209771cf5e9efadfdbb8c5746bb4d30f8a002484d83c7a5f48522c97ce1cf5a70ec983c243e4bb42172ca94840ef2f097ea58a91dafab4eb04ed73eadfb381fe06f68629311a1611cf83577a2adcd16402674aa534183bf38f7df838bc78c093f64257a21bae0f750c8f5ac713a0d4fd6df13fb28df2c80f02ffaeee35eac21d8a20818fc5d9eef5b9347737cbb1083eafcd9a4aaafa7ab6f9ba5966eb099706cb83dc5bce11517843ec2dc554735c37e27e91d3875e16ddb3ca84d53ba69c9ea93f42f1f030bb5fdd2ecdd28162b70164a480a1256d906f97393408bb8fd11359c5e210103f000fc95d8af270ddddcc17a1344ed48db28c2aa5221d285d49b7d4cdb3367fd2c1689c7c9c22291eb9dfa471e5d3ca0dc504c19b49220b093f7de71204c84c042b2e8a6fb9ecfdfeb6c1efe6eb78ccbfbd86f9daa282864ced6b6ecf70e895c889843153b31b518712fca24996d827f20ae691363e8e6169fc9ac1c67dd9ee156c312666aa0d3088dd7637210d5b5cb2a8376b9b6d9d201443e87564394843b70393035bc5eebd1af8de14057b5349e46254c2efee23545ba4bcbe804295a2437ced0620c3381a9762b2523ecab71702857a3f33307a0875d42a439057bcfd293202a33c99102f1ba95443ed2037495be024aa9e82f1615cbe03fafc8e2924feee147b854a4fb13f002e68e0447c9c580471df1d6d8d09ac16d56acc42348396feacf38a492c8ae4e5ce8eb92f098c34a55fba513af6593a4f7c55352683398b7ef33db30a72ec6b8706cc3247cb9f4d5b25d9a2b2516916519f453fc5f0d4ca58e3a075deeeba4f7c30aa2529e6fbc08f3d56599799340258d904a26cf0dd5050797793f8605e649536785cfa99e5c3e9274aa1d158b6aaeb9c1d50b0edbd52fdec94c1180418d290708460bf313654900d3c4bd5b9779c75ae95318392b3ca6b89c4e9492a181aafc7cbf8247e188df15a2ba8519be856d1427125f128f315a2555e2fa214403e4ac5eb5689b5d1053dd6d5929e833de6f9ed0d55b82996a493bd0556086b61f433d0e83ece970d6db91f496ccd11c716459f5008cc0b39a344ee947c7c7fe83f973613f7b454ae0042823af24ab63a582fc2fb548455258ac6942faba256ca9e2702a658b2167418323cbda9e94b384a849a298d3a1ebcdb6b76fc8abdba3b1fcbc477ff966bc4f784d6b00ffab7a9fdcc180d002c2bc8967d2c8ff31cf5e8cc6d4518abfd0c10e16e2f9581c7dc118a145c812e670a5fa4869b0d1eeafe0e490213affb42c4c0810f384121ba5806842b2dd84cd62b85a00edcf2565a6889ca747814f8f011e1c0e7dd1fe78d4cea7e5500230600820c1ceebe4f876ab08234416ed3a326e43ee9e0667b968b83a43f48f96b87a927ef52fb65116acc7f631d4e2c04e31fa522719acffc0d92c2a2049d0752857d133136873c50667492c5fde1aed4e213bd2469822db6bf150cb40d27e87f406145f49e18893b622c6101b5b2115db485e44cf5d9419e822fd4d0778435d0337d26be7f2e58b3e3939c4be890f6767704a814eb2a38050557e0f71594f8af8fb9f052354d0d50f32e931d309ef1e36434f0559ff677e9fc49c1d1a59e1676f1a10c22e61b53d1df534ad8373660f0c4dbffb0bd11acfbe167cf07810b63d18fc7376e38c3582a51b35023021af20aafef99f7c57e0c98dcbe2afc6da863244de3fe20849f6470d7e8079287884ad97c5c7c93565934a3fc1198b5f67572d3ade51a83d90ae8333b0630ab3935192ec23fb5d3045ae19ea1b77abd7ca7f685fcc95263a0e74e8cb7a3ac2f6280aeb7cab3336b7723225ac5b5d20f9aa74b8427c195b18cf8897f7242904b9162904a8109e1aaeded107fa6433700e5048bda731d20a28e0d9a6da7ab1868d216585c4013d4e9fcaa4a86cafdc21b5cabaa6b9e6e726d218d8cc985d36084df7f3cf7bab9aa13040b8f760ff181085259a6b05195c91018f8a90c459715b38818378cb9ae9105972a06b7e57ef00c391ee32af990d67cee40d676c988d24d1e2f40fefa74d681b99f2b06c272061ab93b9be3a0fbb266df3c1bd141175409fb8adb155432c332b8f2301cba909930a54e01448130eb7381a07ae2a850b7a009ab10724a71a091156d2bd0f84d3f7e772dd5ebb418f48d615db9c41e5bf7942438b0c2a69b0d9fdc62a1a87e661916dad3b9896d5e6e5d9972c8842c4dcd5b1de1dc8313d29b7db09c4f10cde190e2c3a0050663b8664ee015fa2fd019f656940178d025462b64f08725c6814f09a558cb026c79ff60fdf80b89340c2be4fe05cb816a1d29685a8f7cc62f89459a1ef79ed5cf177227022bf5086b0b6e51f0a760d747f79a73f151a474f79ab58fdd5b67d3d77f4d007d5f70f6d7ee1e072be11fbafde23a2f04e4e33ff23c094ab2a76a914b767deac2b0afd148041d0856ceceae4d628ea47c3a241890bf470c0c2b3550a0c2c2abb492afed4ab1b04c6d313e243a16a536ea903dc221a8762f9f96325c4e8f68598d5adac3b24a17d82ecb0c70c451648d9effab5e1215118d4f3c9b19a1c3eceaf1d9df80d4ca94dcf7df725c4d8601f51fc54b870350e4f6dfdcbc09e03511cd0c1fa2e39f97c218f021c58eef6e586618215f7a18e20e4979ed015f139a2d2a20e13ab67db08b7911ba695b4b888be0d78740bb805965b6c679438b599a07047d49d2543bdd3c89db36f255798064d65698c92b53b8607949fb568d59683bee736223eab20b2e18337963f49f5791c8dd3f7320a56923be67c813d20bf920c9d6c78c1cd565f493b176bc60305f70d7cde3f366c13924815db11ffcef209854d2b07d1d3ca251d204edc197ca0915240669c7874d88061f249e32feab52773eb0e542e5c25b0651298b3bc6cb5da96aa13581b9b34c4552723fbbc03dc74353efe4ed5c7cbe5f705301601c279ec0826c47d3750831ca655a8cdabcc5c24bca6a6c6555b23b7e65eb3219b067e5d787e67bede1d81c63e6e143aced8bab53e98100b5980ecd56ebde16d78e28640a7c97451c960318d27a6362890eb10682d15247866314c5896fe0171ab34ddb263994e2a970d80965a317e5e029cfd211203bc5761401801846955eae50278ba29f4480ef28bec6d36dfc219608f98db793e24924e9121ad3b9b52a87072c53de4235ce42a6764e3ada86956d20965164de6955f65d94fd7a9018788604acc72b086ed88d4c738707e601430cc54c4700ec0d3e6b734a16a4112a6c876e25e34ac4b57444c2a5f73859631d1e8a88d7d861d3faaa3e16498e503b40963c6d08f0eb21b7f3fd8dd0b51ceaf3984af8cb609a66994aecdb91541810a2447816799946405b176a13a305b07f875213691e097f801b8b802ff7e769a86ae775daabc9fbb753e59fc93b5dc4533e45dd94128774b69cfb9d12e84b43bf26a75ed32fd5b340db23eb557d03b8b0469f66c8adf8a3f078e84cbaf5eb80cf0df8b0eb6a7f42c896310b732b6806917d8ba1bc6d6f9e80f1ed11f08b2b6e4d626479ac70f36df458acc154e035a2424a30fee68b702300be90732b68ae65410ecc3c81de4a73c0e2e86075937c5ba76ac22415f1b44a3574b759ee9f9bfd87de447b2cafe2ccf342166d71c0690100e9c620f512725368578a6b40fc71370679958e329a928c2ea371c8965a02665eb8820ab937de613649a0007ea8c0e0300ad4175723f97bea413764eddb6e95be62eb2f9989b181a9d846437808f9adcb0b6412ea3ba8e7629185f49b348d7b53018f9484036dd5b0bc5e99c5f4dc94d713ed2f7ec752f7467f299b071bea7926e5209136811ed3d037fa67f0c589123941aa5a436e29ed9b82645dcdd0ffc72d4c11927502e77cd3d8fb3b55c5bb3fc393b054bdff17c8b427d0ac762ac4ec4d973319401347bfd37c4b52afa6ad07ae26937afb11fe44e77357862dc41eec4db0aa05e5dd577d42281b5705b2f2303d1882cc2ca975558726ede29ed047688f9aa639b803f27b95d6983cb1706bf08c07b1cc97d87f3216b92b2de49f1d6fb9384da99d0f6f35cefe339111b06422bf31d90a0fc4fd3b3ccbfb4606dd38c36312e3e7f06eca53dc2a721cd20f0009f703c8d5a548d9efd79d53d91564255d4bdfa8af871c38e622e0c9c563b5ef29700312624ff7cfab95883e66c26bcd21884ebc38d548be8df4090e5b7896dfc2228febdf84ffb8db9ce94bd0932595352cd5f98155f3b68192ace8d9eea79dfc3220c8b56985d6ad5e711333a7b85ddae73e2964a533c13e2c8c12a4b2f4054054992e52381181c5d938a2ccaaa70d84e3e55a5cf15a93d8a3a583a39490499ce4f46c1a4e967da107eba1495c8074885356b9682aa769b71b4c41275cb69241cafd018abe80810c420265830fa7b2f596e96b93de2ebb9aae7b51fb11bb4e438f2f8b9697d4e9863c853602cb30bc53a7e9a7583401c9e8e573f23b2f5231a97c48e2c9d1637aef27fd4000e8451d2a6454904cbc6abe478cfc4a339d7a8819ad4da5133bdfb60ceb57cc5ca124e3afb14c3c33e03466f256cdac154d5f4d548a8b29dbf1600f9cc0cc1d8bde6bfba12d37d53ac751bbdcd33ed2676eeac19bb12dac1bf73f97fcf296ea63c3b365a464219c351e6bf7c8d1861b8d6742a7b8a44f7aea42287531d1e2e6e8ed64f9c28df4adb53aeb2d732cb0feb139c060118a680f06872fb102615d7b2510bea0207c6cccac5d12c6112c630cced3f78723cac6c69ecf948dae04ba60657ebdd7d707e46547b9d11e3aa00cbc829eddcb04b0963764b389b3df48f44f788f8189945c7a1929f9d24e256dd12d62cb39788fa8eca0b02703f603104541ba95d887034b43c44ad0eb808309db1719cab0b3b05b87d62180b57ca40f2f721a889b0269d0d00e4bbc029d473a75e1d34b8bdffd63bf276f34701e5ec88c042c0e4b9afa045d87d316ff1bb1997f225a889cda23f0ca9ccfd8cee2add2e86e908e2992e1fd8c59047455d5fa68bf6703016021782833744f2e7fe60037f55d5eaf023c845f591878950fea5417403384155e59e028e41c43e7d430c0444d97ba786ab4b532f6fac3b0a4c45487a5322c893be55e02241168dfc4643d6d1e5b933595d0a4974537f1d5ceee4c996b26517feba43241d1be57f9e460ba1dc01e4c3640e830884ea5a26007b6d7593f5f87988a7b04e3cb8f1111a205d6e8e5a89eb30180de93d71a6eb12659be13d2335728771a8054527cb0710e73af453af990a7f6c4da26b708711b48ad8df79069876;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h397f6080366c18140db54c72da22e74557b56a1f0afc592c536968529077510890e0d73e0355573bd9de0a3bbeda40e907fe3c2cd00c4f8279ba2194c1057f28f3bbde016025591698ee49b39412e58e2fa9b5f077d9ecbb0a264486ec2e009b6f7fce4e5c729e1fa9389ea7f802e7e720886ee091097b4c881c72fc6a38c2484255a15b84634ba74e4996614f748f21731048d0513c23e270695789d86e59d7468445bd6488116a5be936d7d3f606de371c15750d44c2727ff8c938a5310a46bfcb55c50f2d771f5d48f13f2463e81524a536bda3e86ee8ea55c8b76363bb77467ad4fe6d2b1b5220e3ebdb171ca2b32ca149a3a7952f392734eef6481374e4e3dd8d3122bbff0be1d3b94060999122d7bcd4a8bbc47838e7b767f0651da41412f4c12fbea29f99bf6c4a9adb4a5e1400cfd0a0ad74197f94225725de3977edc5b6f6dd273e10cd0b55dfa0786ec2cf88765052eb888a546e4715f95aaae67ef618fd416be9b3ae16f857dc651521e4338e9b4ac39c5ad4dcc48b6abb1a74c15570ddef1d99d77c46465026640252a5eb427cd76f58305362bdee90e9e58309c7ced7ddd51c080c7995d57b56e42d4543bba10a99c6fb8d26fc01017f9353050b97fedfbd74c36e85240531fa0380aae0008417554a4764af5803c55f93743c69f0b752243fdd3c354eed693eb2e006df9757b35f548bd49f47bcba785808612f213fb137e084e7a2e28bc7001ca869f428c59f0b0c42b6e5de27aeae8ae82f0d633bdb2de5d81127ee6ddb5b3bc20cb7b9159eaa1df8a11a38c2bcd178591204f73f93e563c9bc6e01adc2411e69be4445645599b2fe372e1ff2184348edc99a1ba31eeb1450f69f478cba066b0b037b7b75fec37acbda80e284e2d90ff2396fcc8c029a56ad74c1aa763a3fc4a0a77db29aeadd68f9a88939c8859964cf2ac7102561bff4df321ff172dbffb089d5bfec007b9f00797c1be02e6ec4a15f76d04074a00d5f060f30746e6c8c8f09aca28372e7896c0fe6311b7e5882e8ab904fc9b29ff468d0b0acc0ff23cac37edc0685ccd9c5c380d9cde05ef6eaf3408b21d733659a78a95239ebe4c4ae314aac21dcd55f327662e76647264ce6c7cca420c1e22bbd8068510682831435a02fa5e66ed8531a6f8a4e741d590cf3159968dc0abb2c781ddc912d593f6dfbb4459f05f669410404db58de25afead121f6f01d332061fd2f0c48f232e45d19aea9c33d14e37928ec5a2857c39359538b3d6490938296483f434083563ee845ed53c5c2963b876c131be31ef8eceaac788ad1674d43107150ed1c23b10371084ee2ba21596b31567e9ae4d5a9133b4400c4418341dc5065aa964e9493af8adb2d2158213860daaaf8b76f15ce39a2c160b7d4d8e8240f5a9efed36c57091ead65f0f46370ffc82dd7cd3c784450d63687b4a863f964bdef63681a06e5c7997e05fca1016a5cc1bbf8607d0d9d30b65f4340652e9d1ee711cef350359c38993bedd98860b675e0c076b90a066c2150a407bbac7c6f8885aeb955893b23bd146d1cd9059156a27f875ea39000a7a799e5eda76d81be21d58672bbb1f7edf9ef913fd425fafcf25a94e97b6a79c1e641e4d7284d7f4309e68d346b748fb2b2b5f61b6d99c6134c7cee1ca00b30dbf708f9fec5cff17aab69f78cfa4f74c03b40bb809caa1955f352bf624c4602ffa179791c768f2b15badcd41e373f2be2f61dffbaeb15152950260ef459add157646c4789ee75a466bff0ca56ba2e1a43c601e4f399de840dfc0d6b93e91cbf6365ed3243b4132d4bc201ac35479dde3c65d6a04724e82600f4bcd3a23955639bf1acbad85684b339d069b682f6acf4bc2e7d5bb6df2063be574e8fa3f1a3040c3efd5492be239049a2502006cedb80bc9367473001f41ada1485db470c07fc6c103455785cfa46d5b0ef581ac609dee14d4b86aa20c6849eb1badf3f938ec5a802f719f91c959d14347a9252048f922f919d27d2297f70e86600733b8b087799b2beda0bd3ca7ba3afa672e1ccf2e3825279026593a85ac6d6658979bc7ef3b2afbcfa192e9dce98aff8939f3b4ab5ece989cba67d63b860e4b1e0696e8687a94c2028a54efc3a17f14a911e1d9afd2b445b817b03c295c0906dbd591fa0b878b6b9a64a286c344681db17c7af20cd7308b7187fad08f617c4b1ce5a8f0c10b435e5b7a42cb067f7cca66a93f5bcf7debe7c57feb6d3ffdc396abb35dc3b9b0ef02ded2a6dfd079dfe2366bfa4344e7e93d30d83516037b121d5cc5805e1c6fb26ee6619a875cc8d89129205092d3ee109317290b79ac45f7c189fa99d6944c13bcd0ad6d3b3595691541ef01d9aa9e1d942c520b32066d84049a76f52fe8825be4beeef3d85bcadd47f5784eb001c055d0961cd4135d83ac3b26fd651f779b430b8ad03c5f80c96ee4c02494e5eebe4a002569199478e9437f3faed0c57b453d216980434d46f8c471f5e4635b14c91e4d4afe6ecd5b1dc3868d97b3f825bf4a00b72c8f54db54248bd8e5860a74bafa70e3bf9f0930ef1ef4fc37f66032f8fed2bd216b9e0acf750e7cf1f856f16a6fed45472c2d59c2201b95d5148747b5a11ceb706d537fe2fedac1b5540d94cde9769c85ef0e1488d081a4edfd8d9e22ff6b9e0310fda9f4603f7ea2d3f45e927d15cc41813b9a71faf9acc5442cc1281ddf4eba1b5111bf4958e22e7fdf1ab728a63836f3d14b912964cf5fb4eadc4744ab7bb75aa2fc3c68f92665989f8fe5136d89305849bbbd3dd253d4aac518907a1aaa577ca7bf3a4ff8dae4dbacb8e02cec5be96f3ae3d5ad0b90d4cc00fc5313f0ae72dd53a82a1294c3e953515c2e0065cef335c49287bf2bfbe23003eb169155d9b24efea22bc3d7d5d9e2de640267b48ac3696b444cdc552e582237abace63dd5a083dfb043aea4688071128aabbaa65e8ec18d16cbb2f3a734ea73e1e82054684c5ca4aee7eb6877dddec488ec7749b5c2258b2bbe23afa123156847aee470030782d6d1f81d066053a9c9d0433a45fa0e30a6d8af63d42bf791a63752d0d388ce8d2fbaf8c5585aa94035e0e48cf2fda51b2a0d1c3ee63513d4c12f336e8398491da867983e830f89c0da0e4f3afa8bb571da77d4b905f7c98c3dde1172cd74728c7129a744d753b12b11f2d2995cbbcb15d4fbf5f5094c790a96755a78836e28cdb21add5357545fc3e6640d683d92208bb003c9dddd036d1ca8d6cf696efab76222792c0d2d979054122bc78e83cb8cb2fb3445ae021567216d55604862ecbe043e7fbed2b14bde9ce4c54084c20fd69fefa036ad47bddeef908c29a3f08b571a1dcd31ed38de2967a787e8bc417c37066326cbc2ba7ed4a755215e857bd90b36ae7cc22bdec896e70620e395c80907f9d596314b06925062aed26db137b8edb34fc527162883a91f7245554abde8bd8dc2186e9212804119a34e814e38e49083f59ba0031d8b505b0da488382b8b7f3bba61c70791d595cdc477d6fad229527ff985d3c039403e3049abdff20df2eb46dc45a7244bd2b80b2f21da4727904d20d6a70a07c3aecb3ee4252e88c27c48f7286c9e8de6b41b8c8c1ac0c809ee555ab2c22d450223a913397da431526091780fbd71f8bb66e6cdf7e8c5c6b21003c24779bf26953debe726e946e48c934729a182dbbe7660162bfab810b9c9d83be6fb2b3c1032ac673d77c689c8e6e51815131d4ae19f13acca441ccb6b549901dc958acd8e1bd95514da17938d39e4af99d807129eb23a5d47aa467d089cad45fb47c463e6d60b316ce106f00af3b43b3d16982b407fd9a471e9c24019ee4181705022cc08858d7f37d1b2499153ea5d99e8366a2d27cf16760dc3ebbd9dc8d75b16e253aa766e4d2b44433fad28a63e13d05d8234ff417a7070ad98ec0b7ac777f3fc94fe9ada7611c75389cff3487aee94e46facd5a543f07b73d6697462b318449eec3aafee087d76a55eb65217ce7dc89da66a127ea1207b05262b512e6813b78cae2800c125ebe31608c6d8a21071f06dadf1077db8abfe6c1a519c64475d389dbf32d22aa82b8b4059d2f387fd0d29e2a62e54e406f9aef9436305a15163983149d69e0165b852f0e616c8f38773b49c1e75e97ab06b59b4f10a6853b69d45f7579e1dfe88cad7f53b8d4f7d357ec3298a4cbe27ae9f6825fdded3353246ddf29af4aa51468766d23e303173c60c3e3093c452081ec45889b4f8111eba0e18df60619d818bd354ee15c04bac37931f6bff1768a265ee423bc216d20d798b310bdfdd395ce1fc7061bf3784a5c19cf424052f4650bd1ae4b80f0aa538592e3ad450dcfca77bf0653d95fcea3c13042ef2ac9b6087ce6be2f5e8d1136be52008f46b38571de467a39eede46595ebb7b011942234de690aeb292eaa90a3b00958d69c5cd49ea9f05338b0ce6ecbb401f7d66f2076fce35083833082132bd922ae49b80fbd6ed1d656444de8399dc2e76653c0735708737825617c9cbd6ca31c47e35cbdda3075e2adba5e56a556d157c2dd89b913e9d7a2abb74d525f234d7a90167381a16295124679c579824ae5b0a7966b5bf6f54af3168604ee01a783477ee00c71f5722705338fd0fa7878a2586a585ad21374adba8ce313dcbf4f612e12d5bc97ae899bb05021830063c953928bdeede40cf477a47500d334cf3b4ba653596b02bbea8be7481123c1f7cad08b711df727804de65801f834802c3081b4304908e729a0ff84b7639aa665730892736ee66aa65f83f2d3fc99fe920e31ad2f9d5b5f694a765ba0875a327846a97d52b51d3381d70713c76ac194f71c6924222e87deced65afea02e6cdd7d13f3f29edcd5db27dfb04277bc47208a38cbf4e51879792dfda6f1608c485a3e21604f905d868556609cf88dfd336f47ec8ded9a296aa50f80274153979a301893ca9d4e3f60cadf7a1f9546061a89906a7e70173c09d2db3f32c47bfa8ed91ae8d04190104fa616c72c0035c5cecd348ca1b42b2903cdfebafc21c19179c34562f597d0002c1044540a1608f0d72148c022286a264ab923bb3be4d6e51f8efe468aff70f292d3e8c40c649222669aaffb9173a28b76e60427a1808d12821715380b6e9a18e2f159c0508573196e90bdbaef214b1845c2235bb549840c289985383f28cfea2db6aacba3b2da0f4935340a56278f163f4249e9d3266651a69cfc20d7847a64be82e64c62f8eeb1327fa1ed4d9e9f1eaa22c5d7ce848f3aaad70aa32bf1c82ea4ad02ce0d14961db7443d4d623e4711b056849720ddedb17ba16df3b701cc3603599b0c5375fc2ea8b8b4c83b259a36efc16aa93b553f65bc84cfbaf28bc774bbf8cb42793f57e70716350babe8397ccf179ac90919276a16e2a7799168ea493ba17bb901ae6de8340c95d89556b1709f80bde2fb6177bef0ea11ee61deb648c12b8a8fa956fda9ba6b9eb14a6f8998ca5bdca07fcd378bfa38c152043dbde;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h940969ba76ce92ca96cb5bcc5a705b2277b54bfcf67b53719725fb11b5150e6948b43f0cff894cee70489724d57f34c6720c2d78cf965f207d91ff6612438da7100761bbc59c7172d1d959a3fcdbf499ef671e8adedbb37b51876cebc7fe4efefc1a50a8ac0a4f00de5b1499abe0df971b0aed7160705cf6ac92f39e935baa02995162eba3b723482cde524c3e917a076fe9394b9463a41b56f515901914f12aeaa6acb380083eaefb76f8466cf2a660f90c319ce4f31b5654f07fe6806343f1ace995c985954eadd4d137daafc18cbff9f609a588e63e148935f2d385a4b2eb499eeaaea8a2f2d8a13006a5d4b4b30c2e92d5ea1694ff6f7ff726b6806c625bf851bb9d760a0be02c454040d9e2e71fcee6e8ec6b310d6a1665b2f19a6f41f139042a48df028ce376e3b1ce57e6ca25b7563536593a9bf4a493527698f8ba06346999d33d900043c67ff55c835e227117923f73ed0fb2b13397bd9968e618a9d0e2049fa84e493de09f201b339e96243c05ea7872db9dcebd36e3ba5b68f0851c870718c22bef29c1e61381301d4fde6f81d1823d465245460f951865f0324ed697cf3f7ca750581531f126ea001732fb0309b2be69ca238303e4d7e73e34a68dde09325bfea046309a7a9648b221656eae7df0c68d844620bf5845b4a40da098ef5422fd84c754cb321c234865e0199613eb2b0f326e37d2a7f32e17e8373f3f7720ad7c70b70ce5289daeb5cdd8bcdef510f3e035d9a8d21b170e7a9bb8a0adfc585964252e7f3b49b1d957cd5293b8c066ddbfc2ccb4ec81877e4ad599f577beacead5ef698b4bd1e9f5791f70fc380195dd19dae18ed82898faeddd1f1c4bee76510ed792c0b545e817f2e26bfd293d6425534b6b81f578f80ba7682b5ef58b5a0ec1f2a1e271fdcc0b1a26ad822de49aee3fb40f02db08796501d47444a1b1c58c6d14546409475608aaaf26bf7c9ceea770f60d724f4fbdae17a6a49b21f6e92a1b2b6939912ba3e3762b7516001b9d45946ff7e2ec6f31571cf1b5a8a9c3f9913bcb309607ab8c18b98958094958981926604c127c6fa8a63889aa5def1c78fc3c7a0d9706365ff7263f8dbd26862aaa331a16707d271fb6fabe76e24e8d57b1c384c1b1e1fd587937518b2cbbfdeeddf7be5f45a3284f24c09306527efef72afa27ea1b9b61c6e674f8bf0aacc9a50ef69ef8be74b7627c877f109e0eaa7c5f6045a8481ee7cef6c78dd017d54a896173133b1f2288d5ee20628b0111db20337abe5de71c59fa20c63e545ee9d33e5eeebe0bd71efd2eb736b5c0b146d4ca7ff40c5760bac7b71a095edab8130961c232001ba1087e71e95755590ad1a29675f8acbe874f3946bce045c95e8ba6cb28d553332d745d9efb3aa3a08a6d60441d990ce2024537c5c32e2413318f2a949da4c33b0cf98c3b08067f635b12024944a6277a721bc5e4f5afc6d8b86c835e93fec4c1e6bb2233182ada552b629453a78e891c991abfbdaedf1e47a00077f3546779677cdb7abac684ef5a503cb819654475f4d9c18609080871b4faaad9c027f29ef515194f3469cb27c1f5b4b11c41b694782df9d41cc306934231e661c40425a5b87451f074e8ae0db56d1e9d0f2c8660b3b00c37004c83a82ed272d2c527f64c8db5fe7e5062f3d30ef54522cb52b25eea10ce427a93d278b7c46924180a48e6c7f2042818ec6a5cae69ca5598270d9e4ed7ad5184e319acefd1f09e47c7a6b95192d21c2cc40937e0222e7217cff75766c978ef035f90fda148255d7efd9b1328993d1e09eba39bb0a46d3a23fee48a67d09d60b731402e045ae4676ad94ce5876076192a713518c1bd2442d4b5fb6b209aa0e553d4084be75c0a7d1871fea45bbfc0f5c2c88534e3fefc5aea764d93a3900b2dfd6ae8f3170c123748b8ab31381aebf757ec4ec09bba8c5754b4a14f2d510664c6538f105dfdab55761e466a21eedc3da8592735164a511ac2abb9caea78a87ef329a53a29c4b0de83017f600157564bd38971363b7b0cc02cc9f1099c3d44a103a794d1ec42d9fa6919eecbc21e059efb38b0928e6263f9be7fcaa22fc89002f9351bf4fa0deeb38c2cdf6549b4bba9e11e8354ec2c88e567356cd8d0aaca074df0d77ea3683c108ee92fe0daad5c35acb60e6a9785921cf0497916af75758bc64bebbdc91c5679bc700bf191f321958fe55769cca3720565979c28c23212b77bb54c7f5e303760e2e7fe5e87bbcbe72f192d0f7c7ef8f91ef5601d63eaae8a5da8a8082e9f1601e5b57b441ed9b9b7f738c0a9dcfa1cb644b756f2c9c90922a20f46bcba5ee3f70c9441ca75e8aea748fa20a9af8b5c0d11ffe7a79e0a9364ee9f9c86c70542bb0d849bea5535518a415b4dbd5392365ac20fc5bae1f89228229592b0a1d4fd80cd88ba125b970df85c2af66b48e3eb8e7b3c991cf918ee40c1d56f361ba6e5daf806c18782ce5524a2ecdd5ff865292f346fb625c8be402951179b88c0b895c6658ac1c39eed6002ef052d8b13a25d2ae03fd6f689cf03fa3dd5139272d2b9b8b5971892788f27919458326c02fc1b74b66156329fd66d96f08b1112b40a47ed791763fb3270b6e8b07e32b9fbc4e21eeaf2bc9edadd64cc9f604f05a37f278b17df980974fa8e168e070ed0dcb40a9fd8c0ef62126d42119947c2877456870aaea51249f3f21d940cd18847b39cc5f11d3175b749a0c62fb5cc0b626ef81d6ed4c46c3a2669465a71ecf644e289f95bdc5f6e5d4a5b670ecfafcc19ce2d870b7a714027e6723a070f0558ac2fcd0359adf9d5e395e9c6f7fa936bbcda410738de88c3b1c320969d063ee16a4f8f27a8d0874a971673b0d0e51ef6f6d85f906abadae44ca879c91bdfcd44ac508aa8fb2d18fd7289cd5f6aa178d3b9b54bb171e84a5dcdb348d394e73c7e857b59194a87ffdfbd1355eca31086747e96956d8c66bc5bbff98533fb0e468298950cfbbe3286cb86cc853298bbb4ed6ae88efca2b930574689c482006160144fc625e5574d1bc4162b5880bb595ee36afdc6ebe3ef78a88be6cf9304b8b2f83a226df5899b866df44071bcd71e2a0da2b3687a64b5d13cc69a9b321b828bfc325a03c2e51bf6f604fca4102a993fd5c67bb101c0d5b2f9d500472c8ce4d547ed4415e3c4affc74e051d701f0fe7c6d8100f23ff5a59bfc28a9601d30f5275fca8f318bb3e6941758176881266f9bf034cd354f9f87bb034799d58da590e3a8dce33c37c48eb92240cc9d01efd27267cd9cbfa065367dbc498b661b5baf4694df19c935ffee311947bb9b34a63fe47ccbfd70d270865489462687b57f203a48c969a107f9c74b4ece6b655d1d11b82927cfc09cb44134497818cf45f4b0b4f9687e4f73560a705a00318d3ac94635b498ca97f898bcf8600e50edcc72ca176c9e1465b2e0c921aa50c7686a5805888bb6897b862694fe99c3566727d9981e32483fb544112d11726ccebdf4395b33fff026de1f34b41049333c90ecad6add883229e9684e6d86abd10fd3d2f305c54649e79b103e0e4853ccf4b4082e770e6b64487add069b43a5e5f87ba1569da0e6ee5ade25ed84d185eeb10c2dfa3bebb658cd5343f69b4a59b8e9307443858fd3a8da1ebb89a8d332d8353c021f57863602ca8422390f1d7e5c85eb2aaf9b96defa2468c1ca02332a17e5202cbe4a9847814615666e55bfa05406546c74c2daef4ee984f5d29842e58fee653c0946fd09688f8a4211635e8a4fdbdd891708d26e1ffbcbcec08acf02387f982505b4515774dde219a32df5a4d8e782fa01155c2f711b350ea2192c120f96b1b8b9056bdb68a14e82917b5b49be6cb539108a01a8ea725e3111e8c85547eb8f2581724cb1263207482644c5a244175117bd28ca216ec2e310c66f58e3a74a15b8359ad90ff5154e1217ef61cd99892dbbf6d299d8218705029f86bea7beec3360a78e1aa7afeb17fc989eb3fa6b377b3d1d6bb2cedf0b78275c0290549ad0db98f761c01087c6af66d4c182c63ebd42075aa82cf61d77ee97796f7a690f8769d379a0aa8700983016c20450e296cec0375a74aa45cfbd69a8a45b435d7d43c8f3a10d4d8379c76a737a2fe696300455c7e147676deeb0f4b6dfe53213b07c1544918d8c7f061018d01c491dc840abe9a8c8ce824ddfd7c64f85265fa9f15998ebb0c559a3e7e1826c7ed3c50172e56afdc7c4e9942ee7407f64c8cab41d221e508ef3c7a3093e03a93f440487fcfd25c1f43ef50f9bca2242a91c04a98f1d8ccff352e4fe1bdb24e3ba70d456d609ccc1b4cb387f3edbbdc3c1c25b5e5f1cdbb0b741f08d47398f1b9aa006290e2089d62ebf16f2cd3ae442a2547f6ec3b178be83b8bc676eedf5a903537cb177a54e340de4ef228b8c401c6cc039c9bebaa9fa1d5cf5ec947b24fb40471a0d7035bf68db3a1085f190b83ff1f539e2c3358895ac9b3bf91fb7dd20922126c717d130d14e1e9aa8c81750919b4f732a1d488e804107d540389b8d5ddb40e3613e7f1facfe00a278eae50ddda0cc8f3c14db7a9769107dca8823b0c635ad9976de945615709723d74e860b46c4566c76ab942983ceb5b25249f38fae2af4cf9d69b51d745ec63219def1903396bf8f531fdc15831add5db95a4485cad67cfff1e2776ae98998190e570801f24c026030bb7c78d0c79c5f740705c0526fa67df775f9cc9972956d346dcf163b32f18de64ce5411f938675719f760d7ce79661f6c62a02b6b5b858a21ae05dfc91fe6706943bda0a554ef4578db829dceffe4d065fd6bb52728451e077648f0c574a8afb95e84faceb96da8176ce7183426dc49718e38f9b0f449569376fb83107afc50887c63c32b819ace6dc85de39f91a7319a349606f29224b751a89e8b0d98c036f3b177519f7909ba269eff068222455832b36307d5588656863b682480256f317e77f993c57332f2261ab516ac34352289314ee1917902d0c12e777dd48eec2d7feb5c4f2081773a74994ae5786dce29a510c7be997b9a6b65e18d82f84a4f40dbd5a67b7770d5c9beda32e6c275f3766846cef26f3db44ee1f303d9cd5efb40356cd15e19e2d756a39caab9db371e983bb1f5715138179debb3fc2fde2d22a333119eda487b1bec4573a70270f15a06edf6d4fe4d5e2f27d85c5ac1fc9eceb66ca4f3bb13ece3afe7204ae45e677d3addb8faf5f904d07529e137822191bc07dd85072e959a4bc612473ad8495de7598f9104ebf1967725b55c64c1cfa2fd6255b1568f36823d4c609b23846e91489040ae20573fa6ef8103462b016d5e4d33a4864e6519cd6c74fd77a826d05f901c5c972e7511bc1d3442cb497970283fb96c2a921f7d1e757d32afa1712dfd3b6879e8367532cf9bc0c28151fbcfd282e5a194b9c972864bce66525438e0c4eba8cc470b6a8b23dab511045b83a93bacb0cf49c7e9443b2a5574840e765e963c1e5bb7dc62ccca05e20d223b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hbf491e55ba808a0d18765086070ca1a6c96cc4d9ed11449bf178af969d0b5fafd482cda77a135e133cd5f19389aecb0133ae1361934334378c3176cd9c344b3715a408fb2858fb081bd3707134702d113c2c32dff65d8c8a9c10e569158806b61448246f7b5e7c0c45c6e9f525e622907e78c4688f52a35e47b024500de0b0726c8692597d352cb24bf5f4774c23b650783e2a474047c4f8f93bdf6951a60e66fdc927d69894baeb56374ecfe88d44609d6ffb2eedd10764017e86cc0a6b51ae7cefa70e4b8aae9341c8ac150e0a0d46879f7f2d1c3077f511e6d3325949852b17e6cec23bc83352b6f43a3425710a202ba8f9b38a9df3ca9aafeb9282c10b9d183bbab83d057431728ec00c377c31b384f8a5dd4435bfb35fdfaa66137897d77f261dd84ebde5fd434ac5dd683361aa4bc6a68902d5669354b6be611fd7bebc65644bf0b897d83899609debb3eb7a77a9e9089e8ceab0ec4bdafeacfebd3d2514d6071c5cb225b65de7b3fead53710a3b88ec2474b30673d3e9839d856e2e932c2cc3169f6db9ca41b7b2d297c141e0a8ffbee72ac5ed1974fc25ae615c64ef1ccdb9af6668356abe2b5610b37efeb6177ff73d97dfdeb65f181479854cef6c2fe6820044c6489d650c099d49460d8c3aebd4628b931a889b0ed3ec2fa237bafddc4ce2df4c29f38f25eaaf1ecb55f5196346a3751eca03d4cc0b3c5ab912f7037426e0f078240316121aeb19377981b3f76a7ec919f6c1fd07475672a094ac0dc3f6f31f40a9bd94a4ab5af9a8ab3ff329d406c69db95dba6d040b259e98cb50fdf2bb0d9f81823cf9f0338d94cd90403ee0bbe61abc6816bd8a103090cb4eda2f961cf927e86c4625c75562b6ce7eec98ad3f63e2cb6293d3f2e2daff658df36c808d717effc94e595c20c30f7e9f3d192f642d8e782a075df47577792eb4877296f7f7c0252ccd89bef9aaeb9b4c8ed847bad1f64a72ec8af8b4d1bcace19abd64c0930640cb41fd1efe60e9d632281b0232e1368ab4103e9820c6f0914b85140e239e20e58ee3db84047cfc5867685eb971a4b185a2e739d9dcc11713185b8212083ea358a5940e1d1a791651d935621fb57f816ea2d22403c33f142e78e9eb3ea321492ef9e9625b82db419c7bb98f622f7b5e2cb33e427ea67673399b7af6b60009b62c51c1dc8b078b5caa40449f0555c0454cc2e74c5b99efe077c4d22ac4b90111e2eec30dbf399f747d73d40402a58dd71dc1d397194b3c3b053d4a934e9eb8ffcc47a846e54a5d71a44f0d7ff67a2432ed4c5ff452da8b2ffee1f7e5679c544ed5d8c28a836315270aa5b869f631011b392678276744725120e0a8d814d5ff37b0925de95a68fdfc7a5a88affaa932348f4e4e8e121cbb658c3dbdcd536f538fc5a0b2f63c0c7b8a84848b1e721bfa3b24c9db6c86cae8aac4466ed73915b8c2419d7971ddea0a80b8a8b9097538d7053de0a6f9db4114c6b8fbc966b1e4a3cf4ac5ff94fbfb08d9faa448b6e683411edcaae4975014d8857d2ce157cac4b7fcd645b12352d708d316a7417bfe1224d504e8d3b5aae305eaccfca35abfd7fa3e989c092d7051f677c4c3b5ed5c9fd4d2f20e1389b0473a81e7036d74f37b0dc450bddc6adaa57decaa571f719f1500280bcc4e8cbc3b854730508b8b537a8aacd207a9f195087e6f442b198b0ed5e7c77c70730ca5ef458d36207ad9ff71c66fe9b2e9090790425634febaa0b6a02fc2bdc2b169d2d90b766ad9741f18a7061227cbc0b43e46f3051554e793d538b535fa80e3bd5999595eb27378c1259e4dcb90be4001739f51c3b633963546e24b05b74d1a933e4fe9bfb77b8005a0311f31004dba364a1308ce67d310199e8ff27620cc70a6aaea4253d452bbbc257276217387cd91062b3d303ba7af52629237258d6c9be7d0dbb7e52244b7b159d9fc5102ab861908cc6d10483a9632175bc2a8f34014b5a24e5c693a41e58f1afd22e266016204a6322e7040d36c7ec778cdacc4c49df9189ebd4a38475b0492c19f2e7971ce7457ab5613513cc5f08cb9c75949ec85ece082e3015bb15f93d8c9d3ef9b9254a473ed4477bb71ab5e3287900af0f80aaea339cc6c69436b7285f130086d78e37b8f6e1cd5f80417213dfc49794d28404bc343e634d7c66530c8835f3b2b2b2b6cff5078258f7037f893b9e412089bae982d1a2ab30c14d105b423a411c31890e8805ed8e89e6f533a23cdff1ec8e252d5bcb1edb6706227f074efa4afc7790e4c8a1cb3f3c1585612158182703dd670341af1d398ebf1ab4aa5357acfba4e3eff5d8692b0d69b0cb4f9868840c931b13e2e13971caeaefb747583148ce8c2120f1087051c44f4ca836882870055d5a8f43df642ad4f98067f512426640c197023430a8e02d02627f242100641ec55d71b633565106356236dd629782af91f8ebfa1adff15cd02844d540626e0564f106eb6e493c53f2456b98203f849861fadda200cfd5dcd1ea0b08c62921b6e138bfd55a6efe2165302ae8588b323633bda4f454731d7a05a4e10913b56a194049d87e04fbe733d6a7f4e0248d5da6c9eb20ccd8e74e375fe910d480b99f0e83972e0e5a982fc281172127ffbe2dbec48182b403f03c7140759ba740abeea39fdde34fb64b209b823a9390db5eed9e4938baa9a01689eceb600acfff0753ad0cbd8d8006094adfbd1e3bbc5ba4b1bf9d91d5ffcacc236248617e3dabad307a0cf3ad4a190b0107b38d7bcfdb551d90e8c5088d094191a529e4c2106046844aec6a0be32132907d5a4bb02385572b7f292f23ce2b4d7d59e741cda4cc059d8d80566acc4a9c8de1ba4ab1ab0a3735d51507d4e23aabcbc2a9af7620a99acafdc0cc1fd8080d07d094b60f285e423463f96cbbe6d60e8444ec4f68104ddc49dbd151a6a971af08e6be26c712c22f1c2f943d98f1108d64a6d8abfaefb76c917acc2decf448b78688330c1bc3ab221c389cb81f4f682f7d31e344bcfbc624a311e6aa10ae0eff89ea4fe9cb9ed0101ff070c08f171d3eb32d27c059f6925908ef503311d81dd9a17aa802189b88d7bd9d30a8cac517ede31f776d1c11358115290033bd4c0fb1574d42fcc7c1b1e811599f7be169b47e5b318dc58f578486f8788424bac799d852186ec1fef28ba187d221ce4f4244db6b3af02e77de9e0cca945bc0439b7782cfd22dfacbaa678a8d627ba0a209fdc43ba5ffb2478f41bdc8f45909ace2c17c57935478b80882ac1c3b0369fd0b4bbd18e44b7a0bdd2371744edb391ba568fed1a17c29e5be866ca5daa71a5a610724b559d9cf1ff675e66bd1701db34945dc6b490403fa699e0b71989f5e588fd505e44d7a0b80b03b7ebbe1ce7aefd26ea07ba79c0254dc724144596f1d4a0e91ed08e839c1d00b3035d63b7ddfd5cf6b9aa85e13c5341ea49b93ebe931555eca121d0c06db258a17d8eccd0a3a57f3315c1246acd5b2afdcd1c88652854ead5500a4be4dfe409f70f4fa06ec84359d9fe8c96d51e18e22d28679044c038878624c15dae14d082c554bdbe0ae8985f984ff7e138af524efe79968b68af9981a5afcd27ed27d0f50ba7bf530069a46120daff229d27a0d2e38dcfa99be71039967993d72a14d1424cc003600c05b8db8aef0acc8c96b195a8f9fb59b850a1be848c668ec81667757708082427aa124e5d6a526c027baa98faac9c1bd150e472b55214a3942c23a195d2739ee8d620564624e3b4a9132e64bb599c9923f92b2256ad1b6a33b833d990f493bc77bdd32a449c01f898a064d9675f1655dce14d21f85d1ba7687194ed124aef8c8153cd6b121d3265eac13da9b4705138e53b57ee40db5cbbbb48998bfc663313402e55f6694aa347c2f662e285583bd549a60356b42e779eb7b18cdcdce94599518e984de47bb712bf07be89b3e9bde2e77750711b086ceee55e562a18da76521a5e62370abbb7a5617e4dca5e584bc008f2287b50832e7e7e5f6fad4507dfa651d0d3312f9c0acaedcacaa2afb6682dd58c8ff07dac22ba67eb30f35f4c2fae493ce09f509af907d36faddbab0bd6e2885f8fd98292dc8cccbbb5b87a5eec4936a083963228b50be3ba3d5b9aa43ef7ecb9668a7af636cb22e9ab0c706817566eb5a8dbac571c7c0ca90226cb5dde3a8fea210ac32e668952e9346b2f3a0f0861f1682e28ba2e9142e0b9ad67967856830da0d9e2ff6c6060d9f9590de21ba97614a115b710f199f791bf47dda457fa67ec2777c29663282967880fc39fc50d368b7a6897edece8815f6d7c948e50e45239ac2749428ecd0dc9bd3d90f2f9dd4c85faeadb7945fb03bd5a1312ee77f35a8041150e98f48980fa0de5166dcc28cc125da82cdef8f22370b44e03a3fd40e517035bea408c6a81be4fd3a5cc1463a3fec22827ebd028c5d5b51fe4f6ab2e7f993ad91c65c69985818bf96f29bd92aa99578e52ec0a6e4667ec4e3f2c9d4068ad836ee13fafcd9567604006a9532e8fc2ef3098ce5bc06175673539c0b38440f6caeb5352a766470d0d2500e78367e06ea68665af753a15ff1fd45f2e45b0edcabbc0a4f8bb6af5c4f0084030ed1b30b3d47fe13f58052c252f9abab804b3f2a6f6465ebe87d46049dd000db299be89fb2c33ae613d691a25e3274254183ae623246aca38aff37e53fee6178657e0f92cbdca816b3f3fa2a9e6cd45f26368b14600081cd229c555adac30e4624cd964b8af8584ffd8a048dc0aa10c73cd40319d27a42186a652960b82a627152f84165b5f4a871c00297120e16cbad5dfafba97d7b307044108eff72da0c04c8f7132d086e0f87731ae4a2dac61719f6067000270c0eb584aabb221b8cc018cb6f826cba2441d92978ee048adb14a1a3bd6695f019ddbff947d7d4a198415021ab521991950b94a05fc3af7413ed57fb77ac4a56a76116f11c6592e5ae74b1eb257f31b4d7c0b71cb8f1727e4bd33f1a8035ee21c97e7edbe8316becb0a2a27aa061819b8a0a4d0749a31ff68a6ce5d170cad51165609da0d3bfd4a6425d5f98dac44e56f7503b151b3d5deea211210888bab7b573f97ed3f66b874ea20ce6a514dbac08c0059ed6b9d8f8f2d5c18e0239dbb1cc19482a605d34b86b5527a11256a8f0c7f075b189fb76d0bff3adb2d16e5ac31099380aede10c287a77dcbbdf572c30a2a5d6f50fea2ec29a8e0d35aecd96842a7cb9370fa1f0c3ce1fefec71f8b06df51782c3559307251c18f068156a724530f287bd402ec549839a90cc2b35d2f37bd90733395d88cc44c82063a77ef68ecc79bf2795503eee1845ecdd25304a4c6f93163ae5176d1e6d296fe7ef9cf19e397615751d7c8abdba93b38d5f336846c7bd7dc4a251dca474de83092f22c086343d29f59de3f87c66a126ca400408602bd1d2eaa7a3adc7a906a0be822acd698f1cf20c8c18b30bc1da86f0d59dfc8acce077fd25f36418d505d2f6327b0c71e1e150da35c5bd318;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hd6c445883795d87444816927ec9a9ae80055354a513eabb2fbb77f4423861fe7f65f1dfe72f76ec8398c65a73ec9d6b5483e64a2937494b54f40bbd086f6c4ab5d3a7d92fd28f1b3549a7f57fc41dd83d3f74c940a8f0935899535b4722012483a604be59602c6fa061ca638178eef61c04d2ea374ab88f687dd3c842797a81338801ae2f37a5654851ecef9abb31bc7abda0ed30c01274e514f5ae4a91ab2987c95d47fb48330bc083e9b6beeff0b26204582195284a14528f1ddafb40bde97954ca4f447e86425315eb285dc7742b75112e5da7d6172bca072c14b992f4479485bfede845e08d91b982b2d7bfd30d870046107eb618e48d8cdff215666105517baeebdc70881b4936ac9fb4d6667ea39de795a850761686f8e965813f1fa3de6acca2cbcac15ddeb1234a91eb3fbac2d798a7b25882bb208366891bb7fb7b3b2ac82f7df2f0d6edd61e53103cd2d60dc909e253eddf5debb049749aed2727c2c1e8810cba2e8628443f94e23fb06c09d9e82ef0f99e85f60b2e412eab6cf6552a711c2d48e786db97f40bd746bc0e1189b010b41d2c77735073aa6cfff1c959ab14309c6364311671584c91a604e076fdefe7aec3079b2ada66461579ac14cb90c7537370e5c6bbd1aa093e42aa64a069b6ce2e46b32d90edd6f6a76cccfd36858620f56f30cd946dee47d9f41700305ab8232f10b987e6fa4c6c016446d324d96dfe03033857888847257459bf132c9823415bd083b35048e006105859249ca1e7476ddc9edd99e29f83214e700be12e1448aa3a841191aca1deaa6aa6abf810aedb1887513b0dfae24694cda2bb8e025309f3220e7134839ad7a0b51b1265c08877d5ba3d8524be114fa7b755093475d677b3e0ca624373950fa2c5e7296dcb28b17a85be0df7c9180c9171ee0ca911fe5a6c233b55a3f8bfbd14abe49eeb207d83feb650cbd6aeb3fc7376f3cda0d3c782123ed967ab726a00fa409144e7d5cbe0a0f381da24e1100706dbd11e7f63c13857e73a07e281518ec39807856e0115b7115c1ac7ac7685ea9c75703134350cc4215989428e4cd8a2d5dbd7e87bcfd3cd0493b162b4ab794fd1a1c35353bf7fb0e40a90cf9de270f8d4d762103e2d89d7c6be6cdd8d7ae7918ab3d056d178f6c3bf2158f3f10cdb88f92dba9eb9deda8f186b5fcb1f05a6a1951acfa38750cf3990201ba28fc955ac13bfda8831e6ba24942b567c8ea7a6b8dc562e4a12a1e80a27769932eb9b5f16fb633c03deab121f10fa082eab9f8a4bf29fbed1a5b18c414132d818c5ea8c08e0e0251c0998a2e104d7b7b7344a46a5d41b29409a68e33c24b9a9928f5b0afe9cad4cbcc74c85ddd6c5f1982b5c6a87fe30d36199b50b9d3e9ea3ff75adade047bf90cf042b4fa13d4f4ca5560e670114e207963c48bebae4fe11c5b70b484ea9e56ca73096fad48edc3d5ee17da9e0e2536b68df54df7e2e857cf87581c0f1b92d84336234f681cd70a024a50f89bdf41760eafe3bedefa0352a0f86ed85a03f0496fc131a5e7754ad6b885db7d97e31b61a12966c2c7861cf7a8fbe75e093a07603d49312a80388b4a7c32577ea070b6e5c843d8f3bafbc16099c0f0476e7324393714eff1b7712e0eb1e4dc9c13b2d6a380228f22f906acca72d0a5f87a7b99fa39edbb5fc05fc9bed1a862dc9f9dd9efb4c14bdc80f7ccb5609b7c9048939d71afcf6ce8753fcf219cab65c5d874256996d97ded882dbd641f0f3a92272e097fe1f78bc053d6ca1bf5042928fb33fd348bc5a7826fa78ce7aee8f08e76d944a0529752b29a0f9fa923e5c2e6d82874d82dc649fa0f7250864ea4649258b19228d30234c3ce79f57b9094ea87e181054b916348feb2fd08d5855f885956c872b7538b910387706a29f945cb4046bc40567d56f6a6221bba166025c4bf014c65fa734e4a00ead0cada47c1f5535e46ed20700c8d12f405474223a5d15838cbdfe248bb17102474d0d6938d961b442d76ca186866f44a6e612d99cf72625b8ad6db455357851a576cb756f67dda158bf1b75bd4bb2e4c27ab68ebb63a865948a264b5a8e5a33c477e8e5647cbb48bc578eecfbafdfd53a5732068eca85ea642928a991123256026525b26f3103e3f25dd4b13c170757d14382ab70050a61e8dd0f4e8b6a39d105053b5dc5ca8c6f6cc40552a52f37b1a8d96226a334c0d1970905ada845d060f8420b06262bd4a96eb1ef25ccd7013797e4eb3eff925ddf4763d82095e7d04f8c5509225cae19d740b040e8f5a8aa079541cb511ea7166694a32e1baa4ae5c7a736b06922b715fe3cb8913dd59a6b169fdd0fd274f8d0af7e01885c713d1edb16bfbf6d31aa7d44efedcb1e8236e9f4c0327f4a154dce8ec1006fecb1d88199d6c336385876be66445a8f758698fcfc58ae41fbb5d51c3fcf4ff6ab4a07d72a88e8a83d5eda816a89b8409eb0463231aa70ad1ebb8b0e85cedfc501d49aa9da7c8839bbe2b93fa6993545102bb61a9a4b57594e209e19c2893d93c22d37539d04e056950249593e475c4411c7f2a663274cd03545469668d6a6d15ddfe542230efc264ebc4aebe9ea702dac32c0b1baaea253efba97e754eb4751d70b4d502b69a93ee6185b99be5a8c179f876c283ad4543ec0fe4c02f1a6d75197eb90874cb8ab7b87d262b88f07a249e6a57348ede9218fc4d7d35fd2fcd87352f6a4d3fbaf88d325327c290b0f92967ea2a9755abb24a9a91e54e8bbfe70abaf0193f406854fee5663d72189882346816d4b99b3ad095333357ba737791acb7a142284f81d6263ad46947df6f2ce92715f0254f2d2daf088d5816afe5ffaa3b84962d421d320ad634008ae9e1a3de4ddac0966ea2247699c8d14f182b8744a7f8246742782a60a28b69e63b5b58458d9d2a60f235568c0be8a4d44dd1aa0ddb70de6c242f7bdc9711c776fe1fd250eaa636b938b6732898f12eea66455114de3b3ea3b5b15f5023e69dfe1880f4eddf7ff2d9d25b334e685bf5abc85c20ff52f219f76133ef6334d8832995cae620c2b20c0d76bd30281772cdf89cbcd74c035d2a9bd5b6619a6712bf99710b931abc44acf20295efd54b67389f7112a95c10591f4853c2240f668f7fe0a113dfdfe8d0793503ba789e64b4fcdd819cd2a32120f1245be65be5bbb251a6c319e0b566d913fc38dffd1ebaf31efb8b25229c89d02c277f7b90c27492883ab5f9e7ef64fd1840f0b1e216a7b7d16dc6d54245f7aeac184c8108580216d75dab333ff548e6266cf600be6be520939eaa1d16375867e19784d41aed6fd4836927cf27ab3326e0630dac6495ff40c7ce6810d9130e9c8f86bb0f16c2220528a3a25d9f0c64697dbdaf57c9a79dfb2579fd7230d243d5757f46ca565567f4f2014e4d04a5dac992e30a4713a8dad42edf3a73981207c71fbf2d5a8d31dccb265c0b0fb6da27ddfb52005a9d9059f2cf86793ca44990782dbd224c344b4d68bbc34bb1a7b2581c3b84bcc480c1cd8ff9b114ed3c8bf7d547158cc8e5bd8af6709df94338f004693f0c2404852fb8d8674922b82de8b37ab50d25a072e1e4917efaa02b2d6991d54d7a2c9f966d383c774ceba8985848dc9f15193fa91cc8204b8a86d76211ee33b5334be603977fcd2ce3f41d2daff6e6d1db70b7b11a702db736d428be8c5597386a9147a86236f544d8532b9a3aa8393c62d1e343cdde2fae851ba13b5a84b06a785896147cd335d8a8a9dc478238404c1d609ad82c135287b562e781b330a76999ed001976e8c57d42d7ff75ba2c3027e60e644262a549133e232515492f03d4fa020cbfcf700ca1af2b9d715e3e376ade149784d6808d94e380016a25d1f4ded57bbf77b6c15949d708aef117fae1cdde685aea440058959c4ada7e83664ba55ae2096840ffd7d4faa4a6fe0f7a58252b64ca26ff63bc7d48b576c28f02822d3414c52e00529378e3a86138b9241676c22318efac5237f89781d7402ae5d5792202b60df004ca940bb2011cb1193beacc7e20178c25e00469be53e7fd6c2326129bb781098743038c78c02dd20444360ffae17a8904a90eb7f97fa3a487e96bda78540ad0d2cafc596cd7dc67c162d80c389ea1e2750d42f99687663cca1277b259658a850e585fda70d68221e5b40484adc40ce0c94bd801ddfd314d966d8de625cdaff0f7c67a195d16b3581ca93cba60f1422e04dc6d809bbfa9403973382d3f88d64014f42709457bd315274c76951db38801e6320fc5853ded45610feae66d2c0a570df6e24bc8134b563e1f1f97caf56f3596e0cde43b9440b9cd17f44bc9705996c438482ac1474be29e724394966c4ab47a40d3de4466341a4cae4b054b77ba70f6f48dd7249febf958dc1cf6ec324f58bf603f3f4b0f15cb06a69ca8847b12dd6a7ec28b59102e3e6018f2f98c1ec56d75e9f190eae354709bf2d3e45af3a2c94894bb01325eaff35128cba955f5fb74ed876b29d6f1e779afd75962326b07d71165159daf86b956c04b39cb64297860cea1d425ab8ece991e67780acebf2df0b58baaf3e185ace44d69c3031f097157cc6e743938c195c649c9c91c47163f89eee689f2a3217d289d73667bd8f8745d6e33a947623bfb0d11cff599dd58052737b07ba836514868052fbcf93e04ff680ccd4278fbb2f39f0e231519d6662434fb884e551c4940558016f9b0ab614da3e1d5feb0dd913f33d8f5eb44295e1686461d5133bf4bcdaebe544407772c287cd0dbd92d3508d6509d10d4eef04c54d14633baa1d3b2a64e712eeb58846d6de6b4d095d7d806583b75ac9d439892347bf79c9dcd41b5c0580a0a4064111887ac37aaa8e2c7daa857e70b4f3b200ee05377c0aad89b035bede1697765bd570eb022ea39a48bbb4981fb218ee280d9064f3c3a28ee81780d291bd35b664c19a0730a30971e364ebef8a73dfeab7e156593615d01b091afc0c6a3ac7b5937cdac2df9629ae0aa1ea1e52b28d43a2d38a7a4fe300f29162e5efdbe48ecf5fb22905d89de967a7789f1b2688eefd5216808842428bec7b300ef9b66ed80797948c22c5bc5c8b758839c297ba3909abc96f4f9ef09d86e2b6c9a193e658ce19751dbae0551226186fb0477757f5ae347ca15451930817aeb0c31bae8ef32cb2195d2416e1eaff0a94ede21665b07cbf879de663891c18ff58193247e3017ba2223fd85eefb3f5b359e2970bdcdbc72b6eb37d3415c94fd8152b163a9aef924a7ad6157056d1570e31f1b17f0ab4b6dbe86add1ca4468226ae54d715b90621c349f52231849363b681aab988edff9d817ae1d284d4c391696a945d0ee6ee976944476951248a1f4d6373fda16032ab89c695ebcd865431bd945081c6c848ffdf2f898a6f11ba40c911431d5111f33b8ae5d654796ecb53129e3347cd0cbc0a77e172643b9c9d7e34cd6d517d40f9e0c7811413dc5599d0672227bd8cb39038e8da3f17ab7d6f86ebc81d358aa578b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h54529c33413e1652f3b103afa18cdb6a9adbd486972a0e5c726b9968ebff1dae9cd98456eafdaeaf06b1d0833d0786214ab873561b224062c3de3137b2671ab74d2d9dafb633434b6cb9569f9530c337ef89e874a81ab7724440acdf3b929762254c6f45641331d7988733cc8f28cbc2e64bc027451c49d7cc432f30b0ff3fde98830e079b112121bab893520c2710f5ca849cb208639cbb276a425338746afe60b6a9d58ac67cea6ced3cddffd50b5412595d11664bab2e4573e64304bdfffc0fc5a76686b5ad42b91af50f68361d1ec542dcd15b19d0d7578bfa1b380336120de614920f6438a969157e48319e52f40ead4b5ab6b2e105de70a4f224f91402a45ac064587799288bd4dc4d2588c2f2b8709d227da83e268af9457ca625652bd01f059f2719509167c5e203189e44f48d0dd23844e31ace9f95d2764d475a8ee97324d0ee5cc017f3400b0f52ad76938c70a5d9033136e4fb037760b7bcacfbc6d9f3644b72c763867984d35b9e820f89d155db8f0f53c6745df2b2f174d449ff33458787ee2c8a05959e563a95ef0a8a46c1c9f6d46b5e7018beb56da76d281697ebfc7e895dc50161bc0dea7844190c5f6a41715cc55d14b80bcde58d4f43cd5f7ebc31558c644c473c061ef74a1dc96496b5ab60a92c6ab54ad2631454bcb7e2ff7c1c56d4a3aaae7641f35390faa88b673ea41ffd9f1a3974e57c0d39d5469c923ecd65b5f73b41706b1ccbf10595d5afe2d055c622079d28c8d7b38d5ad2e0b5e05a7b7fe961cea4e8e3d71ed2aa82980fe9e52ab86e02115332e3dc6952d4e70102030952c721185a7ce4708a79d9c7be9feca1e5ff7526f356b06f8fb4ea35e35ae14f28ced956778f2d674815f2396095b5c60c72804af8600a44ba88c306e7afd82a3a45b404ddfe0cc0a772d51b851969eaa7b8ee1d09fb290e7598fb1a8fb8fa039f6f8b6a4c000dd161b10df32a5022212c6e61eccd7f2c766c5425e73f803bd9ed810a7a2e2ac6610e718e0b95ff674a1a6eabdc0b22c34a6f6286622fd703e11017e6cbaf6e78c0bc3e456db7a4085c160f05d10fb018dfc4b4dc897034734dca9ac3ca0577d103019ef74946ca1f139e5573459b604a53c2e7b53feff3b4edb0ea66b56fbafe8109f2b63bc214a299c8a9de085e033dd2a237f49bd06e5630f1d1fed6bed202f6e60b567dfe4de172549d6eb5f97d6c5e89b8edd6a678fee06476221533bb3432bc21ab751fbb1d5962439ed43bd9d2027dbb9e70c9a1236635594e924abe94127a92f769fb1fef712304e25fff96a80bfba535942c593a1cf858f6002f0936dca952c85a9d3a91898aecdf6d8f58b7bbd2b7ec1c07084416b801330ec852ba3b23817fc79a476dec762867871863e6ad6d15ee8722223b2b47a66a014c5d87054c264897caab84cc51f25753027c23f8d6e5ab91cdc875f4e1ec9399946d782ce128765705436c749ac20dad248fb48b20e07a465752dfe86b2bb304bd3d67470b9ef5bea4a7a3a3958614c8e7084fcc44976ad41f652187740d96d9b8538b8734ad9119fffaa1c2cc2c36a5634102cd222c13f5d21a100c5abcb6401c61df8240be3e4d83bd2361fe17317eae9fec9d079ef124447a23ab758ad9a14a7afa9be751456c99f2fde60b0fafbe5fde6dca72e58525add65b31d24a5f98268ec656a41fd439ff278de47523f876d784566cef3fa3480ce9fa2225790a153ca160873ae8e49405b0aeefe990dff9f0d860842ad7641abc92cc80969bedd69161b78e9061a3533abc7dd39a9631aa54cc51534ff80e83d1d271cefc08ef7047525205548166f84173e07ebc9ff04edadf4052bd2963c8964d212b6333c330e99c17c58bc4526e31b35944636f759a43bd33534dd49bd340a00dbe9b8ead5faaaad6bc4a9a53fef26fc80c6d71c13ed6c5ee3b826fa03b70a56edc187f7448d322b1c8d8e902c51d13ad8fa270cb770ec0aa14245a463628cbf3a70ca9ae1502fd29fc01d7d47539a1e6b2c8be997f7b8ce8568832a0cf09be91b225ea626b5ac1cd85ac9f4fe0ba7036da1561104b8fda768b320093f8508065a43f628a3eca60fadf1e31f1bfd295c4f78f55a30a1ddb02c94928a464214ba1938a692cbd23f3bdc430c78a4fbb1b28365b93b085e054c0349fb1a1a2afce2ce2b3ab3775724866539caf4164519eb7e0fb8f0ff2178ea6b4587f10c05ccfbca3190609bb43cc99b923f6b53a47f559ec44894759c91589103e5baaafacac38aafe8e463d78c1cab50fe4403aa33f8f203bce538ad663bb99de7817885e5cc7a1179021011ef2398d12e7a9820367f6147c7434dbf49829d4c93d98f2469ab7518b85dea29ced206609c5abcc430b259c681b4dd32379188fa3f930dd328a931448451b3cb51224f0d21f6d0d4bd8f570219371105312f82526c723e7241cb963cb41795b73f827b79efa95577fdb8e7c7308bdb66fc665873e231ab4c6e7ae9ae2ee99467481d9f49012a3513ff33d6416ae60b47838d5cf91195de47bb750d77fa8bf85d9a261c16479e0282699bd574ecbd1694875234fc1868abbf4538b2bb95764026987eb9d3a899c3a97a7dfa1305ff525bbfd1b8e59f7b79de38bb570d806b02698ebdce42ea3ed3e492ab1877c33b49a832b4ebddbf5e3167ba407e089ecdabbf0d0c10efe8d2b623dfaede6481affa0e07cc67c155a6d82aabe69104bf6a9e8555bb48a70b3e4535d2a7dafbad666d1098dbbd266c051ba4a93af64caf51342a5ee0e61178389d4259f440df1914f47dd1ae5ecdcacac7d716b9876bab86d1c3285dfda754fb542bb8174d2ba3e62b37e781fb5854b4204bb86caaf927099fd60c3e7459100fbd3a627c4313f17928861b6fc6ce98b435c6fdf887044d41079c95d50176aa5106c31041fd9f05e3dcab0d94cab0ebacc1959881ae8d7334d5b3f6d6902bd4315d01b43c3ba01ddb0dc2f7879513113014de7788629b758ee5761811771de39ac9af833ba7546efe995500526b7329bc90d680ce62b24cce00fdfabdc8078f53e1199dbdccf00d12d10c8a8194cab15f5edac415f3fd9e204bab56b58849fbfc4c44dc377dba2102bebca500b569b2b02894e4d65384932e4fcdd266baf5df4832d1632bf7b7480983e6de3485879c20ebdfa28f99a321bce870c4cb42d1e32db0e5d4b552e6bb6e12680514a7a6c0bc4062d8011ea9b0efe3ebb635d652d7df65d5258e539e325df6be8584ac20b0ec7692fb159065ae58f280779543be34b88c520de903ca45fc6f5b9762e895ed9504d7fef4731ac6edfc817938543abc315c3886621a3834f1e699d79764cdb27cea673dc50202b1c408ac9d6b25f1abfef81deaf201d809fc310c536ac2e10ec15ff28ffdf1f0b01414d89717548ebacec1e8ff1cb2aae73daac44eca10c025a40c7e3852425d771cde1d78a6fa49e2e07059659971fb4484e8f0bb6bb2db83f8a27c0f8589ed6ef62c7bcacccb20cc0fda76bbf2b3fe3d3f9884a2be59b88430c5df4737294ea8bf7b3614f234a0a58b94841f1a762609447e705f05d240c82f52fc30a734c8d555e11f4667e6103ecba8782c75b9196bfd6f4a15a34de4c652c6a5ce9d542ccd237fb6a3ef8c13b29209d12f8e100348bd110d50b3c51b9b4aa282fbd1c736f54926288415ac780159d5688da86380aec7988bcb609e9a1d712f9bf43d2f99d7968baffe3cd8c5c181d2d52b49f920ccdbc540bcfcd6a2688868d373f902cc1e715c1436229e72a2b9e7515a5b13b39123c4612c6389e0ce69a565d6c399f47641ad1ef93d54520f9416fcd73d1753bf75b5383377bce66feb8f556a1752538eaba004c53d81a7e35b4215dea506433a005d500f20d2c478acdb4497b8d3d69e97af697c41b9cbb497ee9defa81183eb1d45040962aa5113cd57b9c3a8442e8a5f6aa8927e412695171fd6b87e732e84d0ab781eabed060fd8f4f89d19226cc394f0a2cb1215534f181a4e95a6bcc90e28ca05f3b160d1ae0cc0ffa0c047810a2b94d5c5bb3aa176222b335da8c5c29ce8c0ce1fe6ce30cf5c97ea09e1d2e6969e061794ec9aed8e05cd2cf25c8c7d01e33a8ae3296468ac917295336922777f3a35bda9fa9bdd65ae6006119b5cd1a929091e67813b8ad2fde68591ed59db6f75ae15b5f46b9e8891a6f0c3c381e65c742f43efb5188a663422a064a76fdc8a4c0d607f6979e9205474892a83ffeb8956f4e36b9cf1e451d25e90c1992a763ad68ef1ce1df673d312f9e74af848b2fde64f6e3324b058f810366fd9602d38650e617e1c34b4dc1720dfce95fac1812993bf23c1868ffb35399181eb400d04a06fc2233a612a4066314b97bdbb54ef484543390029dc22a13c961f29011bd363f91cf7b3de2071ea9f930a0f51d5387da0fd09e8d2cbb6ee45d0f9ec645765d0522aca8e9d039641df5e3a486d5a6bcf51f53bb5a56a86ffc97c3a0776e87b07dabb09e092e443238b0177a9756e99ff959f9d95fc351f45d70d0ef88d91acc56a7c953509a98384c7a2f3dd18db77eeddbdef7a32dacefa7bc4e1c6be3ced78d4243e6d24974d937864e9ae3eaf83915704c8f808bd02e76ec7e56150b92799bb931e4f7a5d9d5206a0c46f48d39e728f306e8329f3194ce2fcd118b295b9f28d38546cd2a0d258af9ddb5a7d66cec34d97fb6e30bde24e37f6431d051b5b68bef8f257dcc67784208e1c94c7e5bc8b479360db165ecbcbd20d3c31c7cc55a2e391dac08092aa05eae56aa103a8be0f00570ffe5998443cd930331b8289f69ac9b6772fc724b8270a14fb5ef4903f99378361c418b5133bc4e491ee32037714bf169394264bdea1c78695e64ab7aa29c261a0d7ed560ff9fdcb840f7556b7dd9ef26bded09b04a3807095d1aafe5aaa30e1067181a07ba355e72aac61813df3d2076bf8d75a124da32d28ead6ec9d7c5139794c8a3034fea1f10b6294814782944649d684831a0c6261525d4f46f22e007be59b8f75d15cbc5dad4a4bdf35f1c8beb0838bbf3c5cec9287dd6a466c67fc8fe1da54f1c4f56d482f31eea6dced4413863d366fcf82f7954c07a86143dd6526d5d94f788c0036293478dc9949f98ccbb5792ba389b1c7cee8c44a1cb32c34d6db1e7e79f66654b7042c4e56fbd537ba58099509f6d9659a52af2395057bca1fa22deb5f5e8673069eb95ff46ecbfbb41429a1d065fc5ed4998b5d5e699f7d3e726804594fce2e5e9a8e6420ebd56a9bd290e56f09ad714dee7c049012787856dca107be5ca4077727aa7fe23c5f81b207bbece0fcceba321d283ff32d218b24a6001525ce3a691b18e6ab3ab2bb1c7d0f0930b1041581c7c80832896270781a2f2f40f1f029fe8ee41c3fa65fb8a0cf91a131ef15a27c70a69f0adee9dbd664d3769cf7b58fa2be56c8ad9fb5a220e131e075b35661f6d81cf874d482084d837cc2b1bb19029ee6fb01ae544022b8447246ce00db0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hfac079255b65a03a03659374d54184e17d92beb692b2844a489c6a626a0b015029549b5a1de8f9c97e8f60e0d03f8e24dc1ebc370610f39d6d0e9c2ea4ee9579d81243c0d777282d2e9d58b039740d473c1f521ddce8f583f7afc01a04ecd747eec54e9602b70ad101959af681bac8731370ad3c2618206456a64045b0d3f380c4aba52aa5e023b3f27733ff55593969c8995dd978fc037fcf2b30811e553bedafd251f221b4884fed0a3552167eb7d217421c7d8eb4f22f0bda3058b247dfc3bebba3e480e7e2dc128fc060c48071c269ab5f765e14310f957cbcc2e82e50415fde698a14838937aab378fce2c40901ae8ec8601d7384d632da33f0264213d677c375e2edbc9dc4f3942e944d7f73f8029a729f7e777bb5560398d3b20c87dd1e628395a9836e0f0bc1266e810239a6c5b4b455dd2dcff9c55d93b4832f860cd5f3906ec1752b9fa4d50d86534e0735042552ccaca6f3fbb75b853adc2e3f110f4b5af3099a2676c5341127d3fa952bfce69fb860ce6ca77181316eb6470c994283f5c0fe9563be4f21e3744ff3377ee5d046c5b9abb4cbeb3f876507289685e5120beb41da458b34a7c1a01a494f512c86610bd19e2335e663889e2deece5875ce2b5ae948f4083820f8f32b71c7dd8c3fc8a8185a4d8271edca0452021fa090e91ad10e8ce1a415ea6a37dcb19787baaac2be293a927a3e1f45fee505cf6375e7f04d20813f6b5533222c2c272601bbe6de075627c63e021ec081b03ba23b93775489cf4ef98a305ea120e11972bb393776f8d01bf5345748d5f9f97cf500d5b6f8f085fd5812284ae2f9bfa975af114ef8b9cb797a677252220f8d7fe0707989dfb48e50ef1b394b39b56e1024de396300db6c7f7dd1471465e56fbe6dca57a0b6826b3d09462067c4f82c1a78e43aab8e567d2f56d046753f049b0b0763d073a5f8728345f14238ff4d612b68c2d591acddc89ca7e36e007344a43a06d9a86c0beeb8efb70eefb2ee79f443e12d2cdec536c316362fb52b4117472fa89d110ce1e6f71c70eb5c99fc0173fd24d354882c9708076f0e517362fc1eda289cbc472fdb84a0baf8f7c8cfea77dc3e4bbb34bd157eb76fb937553592cc2d247083655df270e45e7d00f8e5bc148c148c4bf6a86c3593355088d2ebfc8e6fc907f5f70f44120dcc98a8ea9c852d7db63690947c8923df753114173bf2fb57dbd2609d7dc5826815d8325ab8ab34d8ffaff6d02bf6588973b8bc00d5ee5cc83d380adedbf13c37173e50ab2b0ee55680db869c86b9a491582f471eeeda80c254c744681b473a9129f4d0ac72ab08b85b45fa6d750294697ab7bd4ddfd3a531116173e85d281be86bc43535f1665db64d2d9eb6a649c13463b62ff1b97dece0a71f2e214060786d1df7ff9c9a53b7983a22c8a40fdb2d9307ffe5e1d47affe27d9f7eab669591028fd3a3c7cf8cd5d18d0efd9a2dce09155975f9ff7446372acbb450c1a08b54c3e9ea9bca5c3c59830de915766eb53a49df5432d4c2139215b390a68a9b1734510316280768e9fb3bb73ba6ebd0be0d6a1ab99a9d370dc38b02cb44276cfe5b0d0ef460b227b522bcb85e0148e0feb5aebc16708115e1d824222144773060f674a4106b0e746699e77b4f1b2bb71addde9cad29f9213749f029a5926765a096b27d836cd39a21cbcaeebfc24a99b061387b98673a27af83093330866aa145cb5477fc3239c4615b5572219899f5525bb15ddd24b789fc4af00d21237ae3ca1577ded28e079fa97f726ae4d419ea66046fa9aa9066b3adef57662267514ab1534ece63d39dfa532fb6a7acfc40faed811f1b0842eca84704664ce6d24196832d57bbdb3cfa1f4c667ee653135133f6180ff73c4ca9276f948320273998846bd6e5934c2bee562cae219244c423f56dd5757091272b323fb91bb06b374ce53d7f3ad35302353a848d3f3adb0a9f442dd04b3d3273ba0b08f78ace51ff419ace3252d97e67faee715ccbe79c50295ba2c2185738453bb897411a730f39c5b2c1f995809f3e48f10983f0ac10b0571de9271803e5659acd9ea6caa1ad47e948ce081f64081459e7aec8bdb1c10962da65cd3be196df6b7037abb2ebc3e2c901881bcea835c4fb2d1d00df1ff692033da7fa777c189412e88426f795efb863a88686247f7812833a5acb07cf23dfd6ddbeb9d47284dbee3893b9ba65db8e25ed712e2a1527383ef74938b9cddb096c9831daa152b2faa35ba741874cd406fd748325acb68f665263acca88ab955a1598b896d64b32c2997e94a279b4e2df50ed737ea1cdfe35906732e77eebd181aa3a9de01bb02201cdc113f9515a63a408946ddf99f50db850e96b55fe185a6fe31dcddfd33fab2231051982400b576ba49a56cbae9c6a74864b6a493a647c6f5087a8988567db4fb8f1d705c907769eddee524960e4a1317c068407e0ad0172c07b6d54500d8b61a9a0aef8b23dbf971d40c396e9947b6d38edc9aff19d9086afaf472cda0fed8b8c35c7a0670e2b6cf7841ddeb1c14181fd794f1b9c7baebcc56731f05fe3dae912d6f308e8cee311e7be8cdb0b5dbc82b0a483f445f8c127cd89435e3a71e93a91cb556f3be9d872af48e8d93595e59e6ffd06eea598c5cec08386fe505561b59aa3b4f88715672fccfa920c78c5d2823413de4210ff503a33586e01775012ee03001b1dc278c9519304db665a6a407d5fda9b958dc8cfa1a8771c32c6181880faabeccbe1a308889b93d5e6a8bd1a7d251aa2aad000a561daef55e89bc20a232f9be4949a97b3644ba4d4aeb293d190bd57ca7e393bb3c9fe8eaebfa2a487f00a8ed0de983038f4697da98786014cc8f47554178bf9215e4f5675ac54e5a5f2add8b53eeb002696ec94aca81696b83bbaa069c57911b3856214770fd9b560a796fdb59e38de05c5c24a33cb55b12267e9a2a968e263f0d2a0786555902ff8c1c0dc442d5a411ee00dae80bee60aa851dbb2bcb20c58b785facb9e9188934fb4596f786bf6cfc5246e53f74af9052233986ee6d8f179f96fc47938d22b9911fb1f9a4279ef7b529fe2e6681cea1615932876cd9caad32525a44a2c14ab82db258c02a756fc813eec9aa0b64bc90ed20172c85249c8cd2eca713e59f862693147fc43083b3a33e9a65fc2ed5e6b82eff9cf8f14479feff64cdc24d756837cbfdd79e370a36ffde35bea2aa46e231000220f45b80dfd31330b36336e827a5f58132893b152da42c5fe36672890f7cbc1a9172af1e1cb720de023216f9cb4f0f3eaa9ba4fc3c0c121467b91c8c5e0c458d9d74e7df563d5f6f32bcbc906a76687b7167fb5fa087f9e987d6be25b173c4f42bfeb5a28146ce0297cf6e4ff4f8469cf8076fd4909c5582321f7533e0fabacb4c2b9ff122bee0678f711b64e49be2b60770f94e5a8a65df33f7ab3938054b3d15672b51120a12800157f4379b7535ecaf408cefad9b1798809810be3bec7328b88a7f39d2a03c1a67770694061045d82091729c63035a9a03e72f5889b45eb67014f8ba2d2406c88fc2fdb3d6943e24dbf985969d9eabef9861d261215cccb57cdc8370d449ff9da0f1a15066f06bcc02a5959696cc5d286606a22b41ec45e9b423d7444732a66a853e937e19a3e4f8c2b6f891cffc26bceabb5244e153795aa8bd80e5497c1aa0a1d99affcf33843bc2374080dce2106c5d181a1472588ff747ad393f8876ca2fa22756d81d2adc44f782c336cebb0372eab16bfda815b8d5449e4d76310de269f293136aa3efb56cf68c9bd809a1058de5f4246a6dfb376a391a1678c431f69e9aa75905cfdbeea8619ba339e8d323a2f9b8a0271f733a6d57ab43dfeffbb69374c582ea4404c14ad99c2b34a6c58d3b3e4f98e61cc23b722a516e750c467709a739eadb8cc9fd8d700aa561f40f75092dc543e7cead9aac5611e45f171dbc86f320297dc79328ae804ced05af814e0d09b17cb3d4931453d219a261645a6b3e0da9d3bb1fa293936c234c78f3d81ee86c0c4c2ac396139fb8cb321b3b2c792889a1c45b1a579152f9d6c9fb3aa1f2957e9c4b735488aa7aa656865fca572a628b6c9492ac430f91f3db034c70f48050db89dd024d1a3caf851240b1ba271b28360a2f45e8a4bc5d0e694433e1b714c9cffebd38ebe955342366ef7bd952de3d3b46b8bcd4b8704dfd2fc27de4682ee2b2829c3e24d7edbafef8ce0a7715681b02b1fcc804d0cb4a872004601b5c24afce2adfe74af0584740a2632408c67df127259922a7e0f67c4d87a6a523755fde183eeab0af95c177664c3806162301f9ab71420997c2985f0e80c75dc90584314f8748db600eae63d3bff8ccf1c094de825b91c0da5fad32ba6df63ab7b057163bf1bbf131e8c82ad9c77410be9765886fed28dac674c295a03bfac420625101d425546883712acbe925e31e3af67f8ad93c6a2ef3908b574e9cff481b3765d115139221e182aa6266142048e82c22a7daf269b835dae16bf4aef0c9ceb94bef50b78c0e3ab5c4f9eccebbec2250e60c045418bc8bfc5b87898db357da938aed2f6c00b18012015f8aae72085537bc24df8b02cce6f900d0b426069d5e8452561a421318cd514bbc095a6640957e9eab27e85da0b068edff0b1ed5ff762b2eaa721adb81dc337016bbc0c510f7c08e6eacaeb82fdc0f093b4724d813f2bf24a290af4ddf5f6222e9d97662ca37546b036c6feb4a4fb0552739ebbe769c7376dd1f1e92044d4f16b7aa68f41124e14f233d343808b53da400644dd64e9989aea72360f6ac7b2faac4c10007615fdf2e2a11426aa6cadd0edf42e67a8e393aefede8d98639a7967433aaece8c9b535e4b8c92def8d24bd950923a32fdde522b7ab6199f9662668c3627f851c9a811dd4034dfd2821e5d451ed79d1b8ed31b443fb9b68ef0e5daca93d7ccb6cced0274d664f362e6fa23d3a1ab166d01eb7c63ea79a1962373c4484a597ad98f6d0c26e0a0ffbe381d2793dab18fbac80a9ef6614d191e262c468f47bcbcff705bb23e0530d7b72625d1dcd1653520adea2f9f9bcf5a66e285b9f1606890cf6a242a0dace546db706294f92a0b3dcbdd890910ab9454c736cf61788ab04f8d5f5073fafdcdaa193fac4739e9fc6402d566abe918a55bd212132d07ad72e16cf5ecb8701984f5990fa677c2603edae7b16cea1bd85195bcb2c57b4fcd6c1fe1e6f5a8f2ad758f26c9014f25a0179d57977dc0feb537e51bea33143141919590c3e3d67cecc2224ab30ae286b0c438d334f4a3250b4be241e68d8a33851de0fe9089119f57540d05521c831116991daa35d76a729cf1557e3ec6fc62b41e662a80e324e2b0df124ee85fc4e55a2c0a1272e9f80be01740d55568ea4f8c0cbfe2d89d06b24ba0c7be290d121237cc1a5854e391ab4e6514c97c2fe2a868a931701a1004ffbb65ab1b5d60ac81d1893b96e38121378d7194bf8b8454e10a1e52125907b13a8c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h2ac5150a01cea685a1851530cec21dbfe693043018a3ee72ab1e0b124d40541993d14d8049f96a361770232b6ecf845eb1cf71ab84de80caf4d9a0f409f2707c4042746f3ecbe3c529f99a7f2aae5cb0b4ff60d8d615110460129a50d1b7f1e33540e917d4b54565e6de61d6d589215406f500777cd315b93a88e201181f1f26c78e61c805284de0c3744967be37d9d99361d75617d92eaf808e4602a892a07812ac28a7ee213145122a839c6be4e6d1f53757d57a879d23f7033429b658dc991d1626a2da44938d57507bde3a66a6f1f2acc0a41a5bebb3ba000e5b3f43768cf652e843230270a2495e190f615a0fbc8c78629a174ebb26e44c8ff9c73e4ec471c39a2b90f748c050b2bee5fbcd2b8ba2d17533e763e05af71515e811204763702f77e94f51c624051d0928a3ac380951e1191bc639acb781475f999f2d7c6d53bfb8bceac71c3ca84e3c1fb3ad6b7192e527e7e72f45c8d0793bbc095a06e6fa17ab32659716b34b857907d8ca94d89b8421033dfb092941311dc1b88dbc4cc5c88bfb7d8be0e747870912de42ab44bd18f53899d06d23aa5f27c3e49c75286a84a4bdaf731cf87680bd0f874d93ea844acb2bfbf49ffa080a8d13c0a61873ea6d8baa3833dc02e49bc030dbce992fb3f3b928b44ac8b91d990e29bb7532ea90b065272491e66bc087a44260c9629a6ba183cb0987eb865cef31473e5cb75988a7a941a0165ac14caa612cd1c1ce9db60d805ab874535ef4cf71c727eba2841c67fd754a12df5d9a9ef6c949c8742d5ee93486671e2c935023d5ceb2738de0bba730d3323839404b7cc3984be858c684dc8aa3fd59139846b9c0597ddef30b32955356dc830d37a195eef483f3859a798dd8256b7a234e5e2dc7009338376a78e5169b0414ca55efb5f82e5d95546753b9046ed912c1b0d0093892215322accfca82ba7ccd32e290e75ad36b2ffe7a3222bea2d7d93cb5d71bedad18608189f1bfc61b6eb7f72d032b15e98527398aa1c4a02996b290ed01943e35a44e26630441a448b1a1897699d0ad7ac1c7ffcc807d06936525e9948b335c767b2c0e6f8cd5062aa70ed839300eddad203b97f828cdd86783bc5e71747bf9b047bb3e46956152bc61a7b1064453ce490c1b3aae36257db0135b595b238922787822ab759ece60521251afca83cda892d35be9df90ab49232579fdfd41b6910400224df8a5dfc758fd537eb68b8f8a4b4fa5b1203652bd2ba527a43d1776c19d70e28fe9bb7e20214a016c62974146ba6b2732b9e5619bd7b3ece184afba61765bc9bb96e71d7ad0ce60fa246f851425f422445570321f54ff8756cc44825e8c1aef8bc08349f0d23dfdc4c0c793d3a71f47dab4eed2728f693a8d1ff03fc9cab43edacedf581e0a3b74e5423a985ea843c18bbecf2c13e2d6bbbc966b06cf16b4a12fc01a7ca302bc59ad261156cdbc1871803d27a9cbd233692809e39a2de4a9ced84b01528f496a3cdb9a41e54d952f32f77cf203a298947af38d3059c327e3b479a6899288c49c201006c181644c636f7bb817f7703a01f264b28e09c35443f9bd4bdd162e3a5a04b1aa4652251ee216ec5e65dcd0993aaf91d56f86f2084ff7478ab28082735eb4c5aedac11c8c094ec2934b8eb33b2ac9663c5eebc433b00355ca94c4a301ee474196d989399301273f980b761838e7b6d9f690fd48973d4b863961c0efc0673189408070b2de4f9b60e5f4ad729dd91c8c3090e27c53173091ecfcb2b4b538769d071a44d4c0c559739317c3353e34036fe061a0e35a1e8f7599d922f1c5f4e60bacfccbe6ec90666d11e0ebae337646333814583004f0ce48a008d45f8378644fd9dca01f8b7c881d2c32422071d73a2a12db33d65c99c3cbe3932092da655be2e35029be4e9d0ccc130fd94cf7b86283dd788814f33957fa020a6bdae0d4fe92a67ce6e29c94f6e951d2059a2d913745bb179821c643d1968fc29bc2f09b15fb0e7d2c796d6d3d37d29bef3affea24be05050cf0e8fd1dc07bd835c9d13f1356b7e356803441c5f9f9c8d13d66266d0ed6c41318ba1f70193affe5e589497175527bd59d209c8899459086fafe232d96db3e7250c07d60a267e98cfadaf1fc667e8ddb0b1434f78d5b54bbf6fca8fad23e56e2d7c8c99d9e88f513f98428922fe6400bdf894a88cb8be2f46634db41b9c3be6e7c504155e68bf970e856db2876cefa9715fe1469a9d54ee4611e11d92ba2c29120410cd3ca376c28b5dcb9115ed4827f984e8cdc540fd00084ffa73df96640c31cf07df0ce3ea2bc096565e4ba4046e482a69baa67b90a2514a48776cab693f51e6255e9888c6f63a834cf2883d2046193c937c36b33cc6863a63ad526283ee62df0bd8879afb655f8b70f991f193e74be4bae72d8450a3575af45f59a1ae8bfb7cfa04b14f4669f5838c6b917f47ab01dc19c24457f1dab0dec3fbef36567b5bb7191f0865c36c8bfc3036d7f993840095dd684fab9b4bf75b07acf4b11e8ed10d22475bdf192a02cf3e8562dc2face5a0dad38c88d6c704f39f430bd2eef4995462d544a1c3c6bc38c04f8e1a15d376f93638343981c25c0158ffc5bbcea3899dbc0048417cb40cbd17fccaa1b7375f21df7e1ee8de06b8816442427584d9b931bbcb4f670200308347d49252ebcf026f6746893b034ce946589e0c979831329c27e33529023457d2015c1f433c07e9ce41d25396fd38b5ca9e67e35991077bd2524b369f32d057126e8c8909061c60f3e819bbbe1970687415de9d1a958c94d90ceeb1218b5dd2df013aed5834a564cf84910f05169479c8052d493fb6474d241e8a368d0e27118615eb535baf626e42b2a0628d351f48e5eda10638a531c5acd148fa89d499e0a88a23883665d4a932f1052095d32276beac7c5832cb2b0047c6becec7bb775ac52d33e1187dc7de81c8c5597c5fd29b4872a29894a1d018b3289b43f8eb8419b9b942a18e4a8bebebbf76fc811081c2c3588b966423d0cda48792d56e98f2e17e2a2b23c9648add380c83d3952ed3634412e4d1f73f39de0181c595dbfb313b76ec5f7f4a87b8fb1608e672f83cd2adb6f3c5dffc1794fbf05437fc9bd18a9afba93dcb761495a35553a3944b3c5af2de2b5ae4a9e3ff235f9fe79ab63687a3009f80678f728d1ea852ed5db2f0dac699b08bf550e8b34e310bf561dca15d716f1c0e1afaa36fb539f3b0ccdbe4cf8e511386a96eaa47865905140e2fc1cb5d5b8cfb4e275e490ebb6e8355f27c5ef5bc1f2283d57a49e8abec2ae4d5e0621b58e80fc4a310e03708810a0d1784846172703141e0ed47a2ce32e56dbeca94cf3691dcda18a8291bb5591fed6ff7e8e86b1d6e4cdef929f0115d6efef8dcd089006d0a6100c3ce62f2ea7d1f4baeb656ce7c1fe8383fabf9f835f94bac8850d503be60069b2b00bcdcba346cab9edc92197395409f56c84714af9d5b08dbb9874ef9cf61b04fa0e1982f6b2a811854490d9ed0e0ff174625628b2d96bb2ac71b9fd16fdcf62e956e0faaa4298e2bd36d345a80113d2e646a18b1ecded73e4b6df8c13f441c8abfc286e478393a6ba92b45e44d0444f6441fa9606756928a9ec4bf0a825173b571d887bb506181edbf596d5bd32b75b895b89d710aa73384ee2527abfb0374df078bd4e69aa3e2e4ccc3e000bf3afc9eb9f53f62b02cfc72155877111f257ae3d699bf6b3bbfe91ae9440bf55416b38a75c55a4a5d6539f2091708e3620af03c861aeb821436fe544bf0278681767d82755e0939d1541dfa9a9d05d4be3a46388d00948345377f23856df330c1dfce71e832d9eac634292d9c1dd68df525e8beee8272eb9987601568e17ef7fffdc3e477808b0d580a3d7d9770d17b4316282ec89c7414d5c924c15580832034ded94d5487667316174ace9db355c4867b2f152d8a6a3f1aa5fe8ea5ee6044c898d2bbf4cbe890aaa8f98f1cd36168d5f8020fd1a712537463a3ec1b6264aa9b0c88e321ea3566b2ca53cd62730aa74b96e31ae2f2328d16e07eba1bd715ada653b3baa0c8c609f0aa2d3765b259d714f49f4fbe0cce61b55320f9c3b085e51723d7434a70fe39d7f4dfaaf553ecd9483a847ae70a74f59afd0ad276cb6f12371220627e6745731f53a2db0b8fe238b93bbd08225e312320daf96c1b61acfdaa9b987e5056865410be98c624d9bc711c5fedab91d7844ce5f36b50c1f6676b0b08b51d2e961eb49364f351821789bb8802a278bd8767a0e57a4cdc8ea4f9682c96b2eb7e411c7cb44f519a749a7c40b610f9e1e859a707758bce39e74ba47da7ad09c15f0692e03b399d7852a05fab4930318d9307c0dcc0556c5e31d13a82e6e8de5cca6c28792f6e905a6e1db32817a4c7c22e3b787ecccc76129b7a04c12d727a6581a66caf2e2f73cd7fe24dfa1ac61cbdc3a5f9caaf3bc0001aab917f3f156c73a0a2ec409675944d8b399529f72bf214719a9efa05e77457ee02281d10c7d27a70a17c37fcf4deaa5e46a06073700d95e5ebc10abc1e156f5307c49b479feccba689e57752d5edca01c9ef351ec35309df48cab38b0614ada1c01e544d64de3b14bd9391097380ff9585d48e30579a7071141baadb4584c04efeec28165017ac16215b797af9410abed5f619c06b575f7c67ef38fe18255707955a8ae24f288bf51537584627936dd89ac5368ebfbff5168faf14d3f241ded8307d7f9aa0a2ff6eff253a614d86ae914f13effabcf7fc29100e4c298eb818385813eed838f4ee1545e19c435527768e76f25cd38de4ce499d46ffe593a9b389264771180b0fcf8004ce6da158e48c779ef8d7244f01e0a69be8ad55711487674765746eda5b2527d8bfa83c0d71aa08eecc499799cfb9da085d939df4c3a61b7d7261825a07be2274f9ffd1703a98f2feccb195ffbc8311e0345017d08a7f3f2ef7d324db6a821fea44a90da4bd212bc48cbc77cb212cab4d51e8fd7053bcecc3edbc2668ccad3b70d82f9888dd75033a135c3d7bd8b6dc14754061ca7e054ecca813466e8abec7544422f33c83454964e883af9cafb42c9fbcc3112f9bb0dd038938de9e7f81dff1fc3b0dcf36d013f11cd5213349fd4d551974335eb7e4d406e61f5ac38e83bd2c772847c9f3842131ac5086e31ca572ab6f972ccea03f3cd67f1ae1f870576451982c042b55159b33ff8a3c5811227bf4d288cd22fb9c25d68a41f5b84c831604c27a3005634a431ee70c13e540040a0372b11441af82bd82fd808244b2a03b0a07b26e8aba0b7706462c9d78e177e347aea5ad6217b330fb4575aaf6bf7fc3edeef040985ad23cd0512a3407241542d9f36ac453dd418b0d24d417ddd572d9f5f54510030d71c5e5485d30af86ef14ac7c50d5b6b6eef7a1b48e80d14cfe7d56223be826a312ec88b2be18923292adc56ad7924fef4028fbda08005c9063edc4ac9b0bbfa3367b96b91c51b497e2cf88b68353ddedd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h43de17db8448944a8670093791a38dd8b6e0b16ff5b6fe1c63d2e7c3dd72203edc3a2f228c1062060a53445473e54d4fbfea57419e66ab5127b605f7f7f92a9b3cf9bde236a3ab13b76f9922007eb2ef9090df137e3556d75d8c5da68140aa118ca5d7a53c971f75a50b7fcaf644dd48a3fbe2ef7ac4ae2638d33b0c62e1b719ccab7717d4ab09e3892020757b2cf1d3e36c729cf50eb21cad2c66c8f1ac7565a16dcd01c2da89b1d5e1e5e211d94c16f706687b31763c3047486ba6f729c8b5692c9c7e41d7c2f4520472411131b238c5a4f536bd6baab3dee7c14aa97fd5b9f9539dd3c8ff55d4149d85f7cf6d2a4221ba6350e429b9f335b301a6123d3da9851732da760775714fbfc623dc237db8edcf8fa50c188c45f633c04a922478f06f6335a10a4d39b7ba960baf2b2adcef15f29d558d9b9b5196878298d12bf64144861250f8c1a3fdc9a1007adf8fb964b8a01ad61a8dcbe9c7c9cfaff47d3a33b8ca892bab182b12f01a237f9ff7be0e75ac359300cf85ac203f584fb06c2efe5d9d1692468dfccb6841886fd8bbd81b5b159855129a4f3c911be6c5fa3fb47cb05c2d642b4cd78ded17ce7ea2de2df0925e713697bab5c53968d001db750846dbcac9995e946f59a5cf66f82f4a81266ed2a1357c94ba1adc9b358d6a240e2fe73e11a2a0d3e14d91f1e796d7050c2f39211ba1106a649b7271a183b245775919a6334ff432234ed861fff08da87592b3c94277f7fa9c2ea7978c1eb0e0efb834e660b9cb7dbe5859f57f6df256d298d66bbb15be887018538e109db112a2c635824aa3777196db53c9a006ee2bb25b1653851eb276b798dc6e2471e46b63b958b1bf7cf779e7ee6ab1733c1127d6922a38ad48bb52c8287da39b1fc4c6598095f357bff02ccfc7d1670a40415cfb07470ec7ab05bf4ec505027b7381a4aec9b42e5e8110335c7b1f3abbe99bf219fec644b57b4ef18ac42bd9abb5c516d61d8d143557408c9e6ebcc691c2d233e1c90091c41bc54d788fd11660dc41cbebb81ae1aea175dfacded4bf38b2f9cc6b7234d8df3bb08821704339bdc96a7822d44fa849b4a190a09c3a7683f72b3c00ba695ea2c5ae36f856d465b939ea80b5b22667cdd57e918939e8fd6037652aea28e3b2a842c8c5c83438f86982d6421e0fc74b93e85b48f70c91575923051931c7c3e89ade85e94497569ab2f027923b67e9f30eb32ef07e18a9366f32504f4850c70e38644ab99627429d665c1eb978d8f44b3a0fdd0b03b32c3d1bbf41111906122a2bf6bc2af5033418e9cf615a726ef049254bbcee39801f488af19c7408a8ff92950fa163af0567ef04583e31173180f9f94d3d87f8c1aecfdcb2573c9a4878a4958c590e77809a5196b10054afeb58d453bd3a328abfe3fc790e1e99cc7a18f74defbb2810179211e9e0a123ebad9790b44c1f131d514955628db025ecee236d16bfcff8aad144c364b779df81aacebd7584fa28f2cb6a385bddc661a245cedfe73b7014a9d46451cb95ae7a9545ea11a9fc15fc7704964f0179ae0eccfd1d742c73d4ff7c54c7b599c2c432cae15189fe708e43888462e00ccfeae1b0df8964b4a8bb7bdd2dc97c8abbd9a5ab2c60645af933b36e74c3af68beec466e21d5c3f5ac7b90cd042c33c4de4c1463145e5e9a44a11c4c1ba116d0e4405a2067903f9e84910004dc58f02db54b149593d264ea87c914698ad19b92f6bac9f42caaa5497d0b690c37a4cd1588ef1d2f2877f89047a55ff5cf858988f197df010ca04e15860d79e74a3ffc14137cee83e7dad6f4f49cc3af97d1c87c497a4954216dcbff6d516b06a802e124d8317538820ab27a11c6c890d327b4fb8d312c3aad2d6b87cea36e7851a16a8d56701d94bc61414c472a34003f54fb706df6578504449c57c69fa9ce1e80bae3ec584dc67e3abc582188695c97f900155e14bf0db315e1641e38c751c4250b15acaec5c4f41510933d6bbaaa2e093f217bd3bdec33e2bcd1703f7faa2a13b8eba96356e0cc024ecd04d1b5920eb684aef9538e356ee17454c6c42ae0c772d4ee8237055867619b5b80abf9dff5a2e41d68c8c64fa85a210df48ef52da4f7467a8127ec1f5a1f5589d066b31ea5a3f130ac20356592a5ac2eaf42f8937ad56921797e47f676411ee53cb3082fc1513d07f58a05b4e5efecde3e6edcd9fb6201ff5ad36a653f7fa4a0114da4cddd377e811c5a21922d17d210add496fb37d2edee5c20616a9ca6aacbbc62b341f47ebb784cc373404f7c5fb8440c3096fb2453fb85bb3a4496a859826412cd88e3f28eba7266cd253dba23eb080ce27e40f86deab877fcec34574e527f2746ab7c772a4faa726376f04c26c96d5f9d614dcc850adb6b7acac562a583bc95ca06bcfbee76aa230ba092337b2be3fbc59cc4437c18584d33fc5b9eeaf76f702dc82b730fa52cce59fac5356fba3b64362aecd61b7fa13f68b94299be5427b06e2c00a3c29c1168927aa9de358430c8b43645301f63b5a7f9a75a4580bc50317adc0dc9b8b0bfa257da84365ba8a26fed2c0f25a575ae3a11a7af4c14435cd0d2101b55bbac8a3710a0bc95dbd65034c881cdf2e5e7803131c38ce3a4fb8dc85039f96ca0430ef57da3bc4ca9ca6d57ac5d0a24c2b06a41a2d6063a7d1191a5c6496c68f2d71dc5149f43c4e70eda0d74d3188dc23ed9dc9539da094d4f1b4e7414db4bcb204884ac2dc1194c87222da17839b4256045848a892ce0f0d2526653e19a07926829b15d693a148fbba364c540360c284b6ad9368ea4d3e8bff3470f23aa811e314d1db6c8033099fc2899ba17d952c2da471d855bba29cf2f1803934eed483df3890364bca87ecd005485a555034f1dd1307b91275cb40516726a63a7601d81c8f14314aeb4f18b8e3185aabe0cf8426445df7201f4bf153c0f8ff93a15f557ff41e6d314dcefc04219f7270cded7610c35372e619d775373f0a67441e680e0cc934fe205627bfb64a03f108770511d30cefb4972e081085472ae8f90ba6202f0ae40142080cba33602bb3983c5d8fb0eab7079094f16a118c77a4837a33a6251ac25d15b01b5b98460fcaed1c5e201f7149d33907df3b8d3fb9dcdbe31ba1d88f9d60747d6b3af799541bc7e01a8faa09d7c3beec5ea1dd41287d91a6e77d46b316ad8365d38692862895e13710eb571d246a1b9aafe42fd97f4edb4c9ee294e600d7319b8afd3669420be5c9bee0f9dd37fbbee98090ce85827bf1e8947f40f562625f7dcc089d4516259b69cec4beb10132e1f27b51a2ca61198eb582e60e56128f241a46b98746c2dcf1a0f1097749d7d01ef8c576c261b14e9176d630e8d79b02c37503a429612661d84afde70c9cca46ff7d822b1d5aaa9a5e0a3dfa7cca7fa3b94f603ffb48630b321367e960315edf194b4e96635ee29205f14f4d6e4a99383b5f1258cd7f291960af5a8ebad68ae3d882e7d00ff5866cf72cdac870ec702331f3f9c7fe54cc24e971c19fd9ef3a5c45fad909530ec079746a18cfe404cb468c8d710e398e97ef227b778528885b6345bbfc31eed06de4ace3aecc0329b0923a3d603b4901a605d5563b4faeee52760a8efbe930c8bcc99a352b3691be23fe78cf92b33a2fa062b6e66279e4d159c0c09a337255b5fdb5154eceb0258ba4947922b17f19f916b9f0fae87f1668f34f0bd1a49d71dbd920463b6c5e67c54c58a63c45a77f47569ecb86d7713b76ddb49bbcf9a079505a5f74b795fd14336524923d15b2fc1e16441e19c5cbac6176f0d71468f4e981f0b0c7614fcc2d8075aedb8ccd4d9f2d31839bd529e38823e6154ab9513fe9fd8082e47cc6f8fa01926c51e4747f06f5c2381e557ea716869f0389ad16f42001ac516159ccb8039b6c19699f8ca8ca70276e6d71fa45db8a7698d4de197dc6eba38cdf40c093a1205c6e1975578067bd2eb1131a9a88af8146c11c3da76861b01926a266446f94d47ca8ae380f678cf78cb7b55476ab41f4198dea061ec0882800f2b1c102a7ef6b2a85601cf5e784222ca7be05082b10c034e4da48d15e98706507e7f16506551b3833f9fd0c3b2f5a265c43cb525a4ebce10447a3bda105f109ff03e8dc020d80c783adda864afa95330d6af75e5104655bdd739926aa8ff113bd0da195215d7faac021659be069af094d2fff9dc8793426c5548e407cbca4d0bb7a1d342785a1ffde56221fa6a48f8974c656d0a980b5ed0fa76d933029968a694689f83cf680c5e80c10a0a297a1726489623c8946b95200819995f7fcfe728b44105161e07f33051134681d923dd855f323c7ef8d90b6901576689989a8300851cfb31f8f3eeb5b5aa3b61423250a13ce389064194e47464bc15deaf7cc27d54f86fe4622ffbc9cd6c22e9bd7d7296a43852f7ff23fa98fcafe34708b45180246ab0aea0b83d8ca646a14655a3b014eb4f3424d18d60a2020ecd832ff384c1a86581bf9b852cca719440663fe640457b7a68b9e2f69e31dda3e7576f3e75618c4eea2403f53ab3a193a7b547448c102bfc98148707044d784a63c30071130dede0234311b180cbddd468ac2527678013f6433f7d9298c3b4628125d7575e34f73a3cdf6b38d7acf4f3aef5386653c1c2e6bfe7bc177aa8a0ea10e9b5f92df0cd754976fae8e6420db563e5d9dfc5cc70af37ffcb6b12d63f69cf28141df86ef3f6005991223b0708803b257a079501f6e4f4a1a7462c3033851aa6b45f8c88215035d2f7414c85cecfe793ce4e8100b7e57d38e5d677b0b6ada7eec63a2887234cd2756b94c238b1d103e8da1d04a2702843303810a5ddf09d2dff248ee0951cfeff2e1b6a9edd1b35824a1623f7437476c00f4bfaf7a74c3672c3aa0e242704f593d35400ee79d6ce62d1f9e3f74ad4e9d6d615c8a95cef4aa6867ce5ada711ba2dd72368a3e2ab7862532ae2e0322ed9dcae2f1235b58836f5ddffe03667d374f58d9b13307352799206f0263ec9b9207c69ffe65ffe6518874afeb63d0efa63972b5f84ad42914a7d1577c3fe88910b75f62d3329fdeff6c5255bfcbc62d5881cdbd30f7418a1fb505654cd14256be7974a90cd72f90c7185f6ab27cd297653e62ba80b4b2ef4ff3cf4ad2caac991434fd4ff2305f0e2b788b708a4c640dd2dd0ea9cc56deca045d3a5458305150d10312337ed46dde54d8e0dcb6a8aca21136569cdf2d9575c82ff83be059f804a75f69d14893efb0d2fcb68992b967ac5016ba44f46bce209e6dc832e8cf07fc3b2b4298bb2e075b15f95ecebf9deb528bc7a05525309e14ea9dbe0a8524ebf237061eba236aa69b86915d0485e40fe392324d3479d9f7849f1dc7101848eaf7f739baca64cf9d383a8a63e257c3651bc45604b09ab487d5a3ee8ecbabf031863abb1d17933a0cab958c4ce67c39fec9e62cdbc8b50fe8c9d9d60ed641f3e4909d5b0eb6f72d5ef63aa9e7f98113c68064fd431eefaf044124237;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h882a85ffac91ad47e39e6d8baae7a2b8bc9f69ac9b65e2f9d6f31e017596eb85828f7a8a6db6d8d4677acb553ad2bbd6c926f931a4fd3b500e7cae96dfd99d859175d0fcccb326a86f8de876818c0f722440e0561194c34d83bac4a89df83431d0be5410e752d7089d2ac58cb2f5eac0f6b1441af2b40d0a779b432d252621ad64760a5a7ae4ccad841956195a843b1d9e909fdf3cd8fb20163cace3e361f4bff65f6bd89b81ac7eefe5109896d7a010bdbbf388550c207fb1edf156fc1fc1ddb121f78148839d75dd0827db06127e9c38747c20f546edac3e94da2b3cfc8634e6866d5517d742b36b34bb51735b6d64c5103b68fc384826f2c59365daf76bd6cdaa1c67069ee7a17673509a6c53c99570e0320bdba7241d6b8ce12d8358e832c11d4aa6684215596ceadad4e11ccf9984edcba3e2d75f62af99ef56a4720311956a9e29e44cd3562c3c6cf819c2ac22b9bd4d45e813623d919d70e3bc5f2902aa5b5359dc42794dfd253ef32aee497bb9465a963ea2eef3e121fc6c328835afb939ce8388acc376c84e168b2c3572b9a1357bc2399dac780175eca07efdfe4103becb5a9dd5d5adc7bafd888bec28eedb64fd1645fac37e9724d852ed433e0f64c08cea63c211ca6badbdf16e605b55802f1e492ceab7eb2f0dbbc320fcf068dee5933d79740768d7e0b1b85d78bf33e00cbc117b5e0711e6e53812de629d39f12ab88e551c67034ebd4a51f9304e7b7257be64d3a72a03417293830d34321a06527b31b6eaeee4c1536d0ef868abf3ae12c293bd30f6af30dc22e3654d8a2e21bab8043ce3a470cfe2107590d1b96868118c5222148d8f97deb20a22a7ca3734461def0dbacf1ca10c1ae36d9895acd1e651db80aa83330f512c63576456602561fbdfc259f8b5581d5d9c7d821abd113da9d004ef2327d3658cd8900738b834e7af67b694e750ce859d5b9e96bc9c8eae15058282daed9aa56015351bd540ca5929c8b1ae2264ea51bccba06ed67107303668f58d131edf03eb523858484cf6a6ce65240977b3f93ecad52b7951eb18b619a6575892e97ce5de5da275085090ad20a54afafda68f98462ec42eaf5c41b5e50e7e0182465737d1ff3d9cd1a8d4c53d9dbf1e6a0acdcfc5caf510814723c87cbd84ec81d0b04b0282eb4082dc61424b30e98f82b7c2a09fd9ecf06f4a7904b6e279644350fa538d1165d6a870fb7f9e650f1333b7ea44e3b91bb4eb8ede9b89ef6868921333d0c9e717a23989fbb429becb9acfe1936b30ae85f6cd0584ebcf486ee9068098474d031ea2a257e8dc720203c6f71b1ddd7fa2e26e1f9295ed7c9b3de4b037253674437f3374394d8e3c1488630ad5c47b85baad68c79f9b85d7d8a95fc34e734cb3ec4ee98c0be624380fb4831e883c6eaabec160c639ac5c6a07354c7206cf3c14592be5cf071aa9dffdbb06b2a1fcb5b1618ea1368f49e003cb32a2ac7e3fe3651f6a956c871b8b850889e5f15ede2b706314d61447fa015dd670f28cd8dceffd4e0ff598446eab588a93729693173b7888a3196009d33a3ebbf399c897516999c081944f6221f8f6189f9df3fe35216aa8e4e02f0323673b9eb388c3e7f99c28ee6ea741bbb998f3bedcea3a25cbbc48a2e60e4a54d2a44e8de958a9dc3fa0f65d60bdc4356a1add0bfa85c3e2dce1df23c58449d221337ac03aa8f307cc02b695e9273375edd81be40c4b1b78c50a428c439a8cd5e356224bce444c3be072698ffd0bbf0b4364565a5d137e96ee33de32de914a73711a014379970d63f667acbb85fcc19bf45f4c30fd980655140565a709e25135106f4256667271d2f3958ccb03c1854f8ecaf22446334cbdb57e03d894f6126438e8ef3bff0897103dbf3679f08edf8b74e4b7f056f7ee9e58f587b0d5dfcb273d9e01219912d7c14178850f738aaa8b40ee426ab771b208829c491dd3127197a912a47e25c160efa6074d0ca685c87fa6ceda797fc27e2204f1cab3564116571f0964c10e834d8f9f682c46887d07b295a18c821999d6d91f046e178d634e8d530236872c14b06ae2322a8f6651b340175c20ad454f28005306870ca7c40f907b0f8078a202e5f77e65f5fecdf06a058f8260d0616c89e57b14f9f6e1ae7ced729bd9d11da70de0b588b3502213dce653a559af252db9dc6fd0a05fda3a836e270d125e2ee6cfb533274d4c8ed27fb0ccf68f45164bba4cc35f62e82786dca61960db6be0c548b7716706f567e0130519fe66be20ed24b93295e5ad30e1eeaff079b73c3bd8b07eb77ff21f778ddbc62cbd01868d06897c19ae60b50b9ab0740d59e57b91e0b74b838651f6916286fdfcda8ce52b94a46081538ae21d31b778823dd950ec79be7b3afb58ad2c1877421f52654164e8afc1938658b9b5925a7da7ca2f264ac6c1e16ba754ca562fdf1aeff880d69eea409b5abedb0edf68c9aa95de0d2a712a7b976256595341ad9c7b11d5223765b41e7f8057d7be0278cd6192b4b800b750a9fc8707beb89c7e3b67e5dfcd7d93c3db0e3b14fda3dc45a318edf077f160927dd692d2dcff4df55d24b32f963169c7ccf27c16c55976f5a7ff6ca095aafba7bf20f28fdb0648441695304aa6c4d2e1a9eb5bd62cfcff838c1b96c5fa805d4d38d1a389dd01097503eccc1dcd3a2fd4c29a1fe0d5eb95c753adf65c5d11691ca85c5b36ace52e3214f506726d66b3740a8f0052fd281ca9ac06863cdc91ac73b77f092e1c3b241bea52eeb023f0820f9867822b8f230059b80e999dde5957b02c8ca91712c8221b70b8fc04449a4ff9db1ebaff06f1637fe5b51036f2bafe79e4bd0cb92fa7049605bac2af30be90c7610e77c33c3812a0d2e08e4437a5602556e995858ca4a2a1c63faec09d71764202aac914ad4b7d289ac5ca02b3f72bc7c0bfec3654aca275c0a6420464ca476692c030c04f37e01e40e7e17276a916c7c3129d6e5670bc94e606e8e82fba975605ff2bcbb5b7d9be82caa3115828e9cd396ddea26f465107b4c9372bdf0a7b70d73dae022c5a80031681976f569dd9f7412d79f7d4ee40443d9a457759a4ebb6b46280fb21aa89597da0efc825121f8c21ba694886fd44c665dc85104cd36e903d2bbcc5e6fcd8c5dd1e3d713ccd58315bfe47a715136a04ac4deb1d214b7583d92939ae6555a6136be5b63d3f04619feceb835eba40d36a75a3fd447dd2fa97c89454b20019c281f92a4a006c3da2a3bc017a48daf2586d7977e789c9e209f6f92fa91a107d2f94e4ba8a8dfba996c6b5952fa9c09cff989bf7a665e1ce0961d99bfe257a2508283880170e102718075f4af555f3ad7980ebe3a9f963e37f53e1b9a4c45c7836f03bb384e47d12a421aa9edd1f3442616d678b05076c1fc8a1d6405e37d2dc623005b176c53d6a95d8d6442f1ec783efe9fd5843dd85eefec7fb94a273a7932cb7bf7cdf126196eeba41af4d4294df2976a2881bf472bf7d7a2dbfa8d39e3ab34a5c6717bd0601e0aff9006ba4eed83bd3f3fd94a30798b85b8fa92e043d35cb4b843a2a50e02cf0bd5781bd43823af6418442273be47c1d889de89d95df3cc1701bd44d9e71d6c93bf9c62282660e4b7a421608229161f1e88162eecf116e4d13ee38842b06d734694847b447aa449ee75105fe65a880634b30f4533dbc19aad11a24994b07b2b752e091faa8b868faaa52eb4b2cd5175eeff12904445426836406781d7973b5eb0c05d417cb98ee8e8a14d8858a5960078f77e9d2831813014655ef4081870bedbfe4b8184599a81f3323419cd06e6716ec477874957aa04e8a135720312da84080000eb1e6f93d23a5a5e5b9d44777b1a0a85af32449bf41d7e99b4771b43c7816738080472fcf04e5011f9f733d98c31f055e20210df255575886b4441d71233d6fc6172b5c2729605cfc07b1d8f45185ccf40f254fcdbba549a1712d3053ba582e31fdd5ace08d842de1358bb7d4ba2cc7b0e576eccceedf1ef08613c5e3828d6b9d03c08f34613b6b6dc00bada1d168a9a3c3e6142ea854c2c1081039efefd552db7f73e499ba97c9241ae358199f2e6c67d24f3da751fd889efbf5b3fcf006f48a7268187b7a5e6c5c5fb6695fb950573cbe14ca0218d1d6e95080acb26a19cc641e8c9f9582f71e3b9af05044f313e9e9842912322572d19832da3224702bf0305e1d5d5d174d957dfd079a5fe05edbbab5ab54aa466a1202b55df14f5db22e9e3d48e70e06e6ef2d42f8f1b11ea87908d3e98bbff44d6b2a3a79601f807185cfb8a09e2a8f267d29837d7bedb77b50357ffffaaa1244c096e696ba84714753cd8f9692045980d265388975d7beeb08cf089257d3a7ae7f27f4378bf884158d11b29e4e7c13d8d406b335dcd48c5d99d7ea8b8041b07cec8ceef53c03e65a44c5c81bd0221e206ac79df73a80c1713c7232e5bf1a0161f8ef2f275780057136706b41664efd9d2bc728bee722cad9f6cf7c330da7ab8de25664e5a4a07949933db0d527bb6b3ac3cee6379a56b5f00fd2664cf0c75e3c969efaa3c4923817abc9a52b8b515791aeca2cfda207d704d3125b9c602222243bc62f7c8a8629b1d73ca724a5adc613e271afaf26f766d8927ef45c8e0d133ed6921c112a23d0029892fd87694fd1fd99067fc36350055d4096021fc4c73152c8fbefea4f7c5235d5fc5714d79f7a6154b8ebd871762b59330fcb58a937735305a12d8c36f529ce134e83af64a4b91d565f79d2fedb80cbf9210b48fc67683bef6cc9d84970df3d48873a4c708ecd1a0ce1355c87d1b5804ced7169e4ae5f749f98dda9b8eadff55d5ef669824e46f106d34ca08979726e95314acf3beb8c16f94ccd148075a8b4500516865e5915a4d7e3cbd2469e099875b8a3903829f77a37dd5ac018799ba3d95b66442054fdfc8bcbb1f0a02073ae8997de74660fdce30178d3f238a23877ae0787fbf169df194ba279bdc50156e5f9f4cfccf6dcc1e2d5a5ef5bc0c28cac67bf4af3aa2bc271d6ea46ebbd1a0e39940e753c3530049f3c65701331fa280b7d3bf1504ba98ad31420e2c049403886c0f85691fcba4ce587fefcbed4758b9d92adeec38ebcc9de48aae2c8727a809f1134b0f1a9c07b3e16fd44d062bc9e9964d34488e00956f27693a9c95a23b0a2ac3d8181099f91caf85ff0bad1bf8b571c1f7984da48e446cd59c13a863174839b43756ff5f92be156a64a6d6b401913763a597183aebd5bb4b9b3867fed86fe101f125eb73e5a917088d8f506680be0230f2c7274a838acec2f441fd73c3230a043700e519835658556460eddfc2c2a1d50a7d8f8847a1f71b7afa154dc9dc8d10d86035c44d022f148c6fb009e2fcf0730ff0ed52795550ab51a471843176e3231160041c69340c24a3ca250066964587557b4f5d2ec64215aa7e9522bb070671e87b4ab633c8549cd7f3818d1fa59fb45e6ba44059e014b3619b84eaf12d96d903390de106c7ae8a1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h43b6c526f95094fc45ba0fa71f510a39d47371ee0d7258948aa15cbb57499ce5b4d5bba81bb82d463608365ca8b99927e60e1c7dc14256ec6acea0b01f405d7284bec5115c7cf45bf73393b743712ce2676486783018340f70696bc28b7d18884aefa26e265e261e8cbd7dd302fd049c850dfa5404ccdf8377d42b36e2a53b5d3ad05a97703853700384e45e87fad7ed57aa876fc9c01289342e1dd7b7879d783b37cd8081116faf0d60029f62e22fb780fdc657f82f33cbe48d285e340fb712b6df4010626a6cf0fe7eb2159da2d72e90c41c44f04d9176e7b37ffda71e1a21b1ff000e1462f6e222ad6fa6d34b006ba873d87cea8dc06f033e2117f9644af0958623158bb6d648d725fa23f7911215ab22b63a0a4b1d2f15476f2789eacab89803c1be0455406f93f54a4663a607db197e0faa01d23a4e47ebf5ff1e9220893407c193246662f0b1beaa714388802f16f4d5100243613601ad48914da719409a8e98d08bbe863ea014687adafc391584439aa4ae515afdaa9d1c00e835d7a495c2541e68a79eb102d8c6959309c37249c5d9bc7c3a460ec9b366dcc3e71613f45ce85f61c5b4d6990d1ce0b5f0c1b8f07621f4327eb42b9a7cbebc5f72aa8df2e20271789549fd39665eaaecedde9137b4d8de6a61f86c9fe483009db71bba54e3acb03d70cfd7656b410719235c6e8b1bd9f285a6a649620c7e62f38438efec16801f0066e5ff2483950d20bce4cd14156fbf3aec6869adde0ec8cb07c59174f4188ddfc0f8e25444b197a6d2c09bac022e2ba4bd75bc594b50fca13e0051d2c5af839ca0c11cca91c1e826cedd17b408fba9403e5ee8d0df8ba5c66e3beb7a2084867d98532be12acf2076fa6581818ba01fd5dacfdd60a6fbf04c52d7a6c821d7e803faf7b35e447b6c44be7d4b2fafded0837aa2015f7c22258dc85b4a65d39cc12bee47794ac0afce6ddbb0892df33542a554df9b378aa97da3e97d221f9357354434a8849124f61be773a5ec03c2d895136b51362eb1543371d4e0b6e8d2743a1a0c44d1c5c6a05d48f78b7a86a8b6c6c6fe1188c312fe7e034d5c8b025076c03b772578757237dad86e643a622bcc0d40db9d5b9a270e7e6950a1feb1ab5ada25489930c82c27347e3161b20b34d7b7bb65cf5f28cdb9fb3016687d283afef3a31ac2ccc5b6cbe9f50a0fafad8002320294f0f02da7ae8a40d7c7207102325d21eeed17ffe9fdd6f608b0e31065d1c60a85427a5918ab30b8cd9c2d3c726a7280c3ae8f1143ab9739e89ab8bb913e91c71c7deda88c977fa57b14139d912916c338ed8da737f155f52c59f7cf544b8f67c378a6304ad76fcde173325a255875c3df5bd82915e643287ef265a0da5ffbbdfe177839e903fd9fa2d3b4203dbccb183378911560eab10fd214de2662aba2397314f70bdabbd52785d268ab173bb63d739d1657e8c326b00b3ea574fe9db1ba2f928deb6f5705aea05a62e900ddec3fc76de387f24691812f1d6fcadc5dbd4a230fe0e8763aabdd47a826ec86778aa9bab996a6674f376988f42d1561117bd379dd9241d7f91789bc7ec2eee0eee7184da6759f99764c7d964dfac8d1487d9e7428226d88bbf88b9d94504f9635e97a18da9dcf4f7327e377c0ee512c70e2726a24f1960cb847830fabc86c1c6eab2726b254a660365dd6bc01da00c98bd637a20a66f719e24249b9148253464a1a65a03b47730d3bb6deb2a530dad01af4377ca3614746bad6ada7e6dbff25616a0aca7d7ea49cd9eef23a06e45e82798932596fbaeab48b59d6a430a31ceebaffe3b54c6ff47529749d77ea6c613529dced6ea7f9782722b6f109a7424ffcf8184f4bf7bdc5cfdd54504673647a92c12f340c5f213bb8a5b325d31a46f89c752a888daddd1b113c6b326ad9a320b43e1f9f41d852486f0b333045cb3217959058398b18f9e621b2a32738d0e5f288863a2ccc37a568062b4eb18ab0f6dfd01c00ca3804263cef139757604c92b217926c05a10746b0ff720667759acbb29c269c3d3dbf645020d7c7a35b95ab50eab8d95a7878123a7cd95a3a033269215a78da788d5125a26766d5361d2df13f2665b93aa05aa2d1dc5a410e139ee0ecaf115cc2d52414eb454053c0c3d39a0ad24e0e47554f85bc58a14068d6a860786bbac943d14e1519c91753be2221f995e6be7dedf5e6c7580849923be4ba73faf1dc85ac7a65f3864c620efa110eb2563d830ccf061adddfe2d908c05e0dd67d7fbb68dfd183bce3719237a732c0e00383e4c054739eb23931d5c545e56a37d2f953d5268a7dbd58cc4a99aa22978a6c6db5b468870c97061a5c36e9abe8889c51280304423102ff62c46a317a7b0059be7f20f2534775e6f39030c1af59707d04c53c2f49311dc3d97cdaed269e27dd3b34e87a95d811396aa3908e13d5d320bad570a3441b1e41691934ac63dc17ceeed91f166cce798c0147b4588b06c929f602df891af3521ddd97c5c1a4609a6c38836d19b3c8d8651d38f4ca39fbb19634bb23d4e0f9aca2d3a6de7ce130e3cc8aa8f56aaa50c5e8e2bf7832ffb16f7c6c9b850cbf557723b71547957982a654a60fa353ea8e3a53706a5ab06664a9541a82f5ea0a87c5a69dea39af4fafa65aa927666680b299f097c8b8609669234450e6d16a88a76611f98fd22b8451a657db62d1d04d7fa7020e40686716ce7abab6f1516e2beaba52706b507eee07dca3cee88ea855e57455608a873aa04732f3244f159504b11d4430f40b547c901a8c15083bb9bca97980f645b9a26b9e087cdd162f3109e631b1bfe2933a634322984111b4665d933a55f139a5ac53aec287a5529a6f7cdce9aa3cb2221bf419f9944565e8e04df3050c89098f958391172dcb53cfd4229021d220692fe29e70ba0c892405606e825bb8fa6650a82d9954364f518c2c3903327c9613a3da1399e52e890c29ae5df4e410e5eecc4555bf418e36f55031ff38c469b814100224e03363020dcd5c98bf71245127fe8e5af839103f915caedf5f931ae813127fc831b87afbee90b8fead48cf1e98c56da60084b8e849b00e3f9db368e80c4f6dc737b861eb8714788082db06d53e36a5d1e61cb78d7cfb433882b08f60cccee16d34e57ba3748a73b995819cb795488e99c9e39d8cf1813f8af00c416c8b0569ac0d1e8dc25ee4c0095776dc8cb296bf71a2ecf3f866d2c8d82875606276a58f6a5cfe5231f61425aa82d99ce77b666968427552bae7eb7fa529b7ba1ddba6e64c5e7926dd5addf657dd2a738a8f3bea4c9de4d01f9fc11e5a8479c6ba064b0dadf8faf713a89ebb3a584cf41f67fa2ca6f5af9ff7bc15cdbff4894cfb35433d975346728802edac54e5751f482869909a707422f91a4fa00365d3299ae3081ad63a1bee847a2686d4ebae6c47d4b0a148897f1c8de832019adcbbbcd212ae95ff72a17eaf8a40d2e424242aa9b1c0903709dfdf23ca02f33f5bde46a899cca9bd7624538ba013fbb6a8ceac94290fb8c746b11898490e3879abcbd0bc075e7dfed701592b64ac10e4718a77d5f63950b432fd7cca4a5774ca20a334c6add91aea7dd215ee157a697f9007b1788205678461e84f953376a0641ff245cc4b80d93098b623c358eb1474d6166886684eacd11f4b21ff20190e0a58ad83dc39e4264e92af5b96a9709ab7663edd34d68fd6555b0feb89558364ca91c160000508b90c404fa31577ee6dbc34f3bd0813b920d91de4126a24589a0c34dda1907e16e46d33366b2b100f35186adeb30baebc7b149206af1d41c796382e83090d7399587f643d0fc3aa1698bc7ad2d422b99066e80ee7951266b0958046048de6cb2ce8bd8313b533544dfdbbb769bf59fd7f91a278f5afde607ddfccbae2948bf0c9cdd26507a5a90f5b5ebabcea2ee36637a906a5454a671d24290e69294d3d20a240b1f48c099cba85ec3afec8fe8504834730a7d07103d90143a4e1287aa2a33c008bc28e08df9eaf884f1d6c2fe07daa1da1965a689214c742cfe687f7fb1b42d5b5f2116cb7ab777a375855ecf108bccbd1914a419df3f44dbca76d25645754e704d15b7a7f1851b60f173d2a9dd6bc10d9d94ca1658512d51586d5b418bbb5abd06cc3adce9693b4cd381b60ddedcbcd6114b8529b5e6187bb8e8dbe735419b4157ab7074026c37afd18fa035597ac67a3983cc8b536999f53c65189017e819c4648d0fc89b60b8e0329014084836578cd8a931a6c3b851730d1d93a3930b9a8ed51639eeff47af0c3879928131ba894147e8c94e493db1fd0fa72e8d1cef3d87087196993ba4921d0b324a423d4bf557640c66f1943cfca153e09b117cbe07a0fa10eb04675b063b7fd0a22d378c220a65be0c5e120854c76187a654a7f126fc657206e7adf6edf20162a9346ffe4e9109ff4e6674b18bdc18efe67ebed01a326da2abb740d119509237f270f3c9a0ed4082124273e0bbe2c06dd841f438bd7232a258b9afe95e86448b7fe7011684c087aeb1611f4c5f915162f9cabf2ca685694d130310911f5b1897f302ac6cb3fcde16ae37b98243a999b13bb1dd4a8961c249b3cdd1264f82e08483e65aa4dc55a3942ad9c443254d0547b6c70a6559786a54bccfa8d1e54d00944af754650c5a22f468b40a64b774ad256755029afeff2d427ccc692007d819cef4ad8da1bc247a6e794e68ee4b6d62d7989ce57c155fa5f8dc1d0d189d53bcc3293d288ba18761140e8b12821a2bca91ec4bad9996e0ba151e6a77443e2c239f52c18036fa4a68dc2a36d09183ebb6c7f53a1d67e92695ed09206667b67b0acf7027a2250fcefe6ae29f5cc6eee018423dde6398c251a8213f457f15fbdbad99b3a5eba2cec59a785016ed69d59a02316bdb336b1a5526fc2380b5386f6719e1ac3923f853172b3c85879dcf84de382c20f2ced49bc4cc598690d436c27200a6f2ea8e1b20ca201814ba805054ce61943cddf510634bd8f867c5d5aa32aa57b2c67f97964d4f3bafc43f8aaa6318454055ea206e8aa7301ac790f25b0b35fb85d407eb888e00aab20cadf228e4fc348f6101670bbeae568d2da67b9e7f03230a4e5e2d26b81000c649beffcc50742efbbda9bd7501fafa116fbdff161d2756fe810aca118bc4301a06ce8865123a46e134a00c82982b21ed20f2ebba28963f1a8fe1c5a8e7f2480408b6948f67e292c67db406842e5abe1990efb72184c637e66a6b7c91b7696f3d51e624bdc5dda48a0c1b13a801248e3de519d692f87f53c3adcd19d001c268f5a0435fc486b5d24b8eca212eb182c2d835dc3dfae266e9e8aa1b19681bb78e6564c912c7dd1a9b74eec276cec9971a2aedb9d1712fd8b2361c6e4cb149e7c533eaf19bedc62d49a2580f79a9c907c85029305ed411145fda5c2942b6e1e68c76ab4a1a3fc2beaeacda36762d20fb977ea3319ed9a67b0f4bbc2d69a1b1243c8238cd34832e44aa022d01c2d7d9c33d162;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h24ff59bd065ed4e5af31a3b56510bf484b0f17e8c0d0f13207944ddb1442ee20d5c069d8de3ec45a7bde6de96c900b9c3c919c629abc2a8a90c18f91958e6ec79f677e375542520a42dbd1152523d2bcae4a28d3ae55cd71bbf52a4039ac53f87c1a418d56af3c484c1518125c7d9aafcb74ec4db089c56e8b38ea6b91e8884af4da79e7f328d9c0536b7826fad9054d32ca815826623729bb462e77f0242cd7094ec4c468e7e5d78f2b619c9f3442487628e134164d61a473696576278cd348787e8c54a4f8aecde05da4517b6298931f7374aa54c8ecd61db140b5bbbf0714333dc265685ad2b715353920cc5e7991b026b195eae6e30f27aaeedf9dc20d6f250880a72db1d341c32e7ebcea537ddf11ce70a5219aebab13a1f36389b5e9680a818caf8bb2710f734d04a6c730dd61a04ca0c7f36bd6301f9ef1be548b00058cf1975695fdb6b09e69a1889c86429fe49e06d54a1c89b5b8ce394f418d8d6049259fd51e1e9f7405a79c41a88d6b51851ecba4b17037f68968ad080418f0a507b0021b0c45bd43e6df55d1f3cb0ecff5db27b136c1acd41080adee34d77316f8bdac23aa2e911cc04d5268247548355a35e48ac851c11bfa39ba406472138211ed7a4c4f12b005db34a157e26fa4700d29febfce888c499420317701bdaba3eb6cb3bc23c72a5eb7e31f920bf2fd791cf3ffb45386cc83bdd03b239fd5f1faaffe9de53ab710e7b34d8cf5f1c30b0f31022f02a9eee9bdcd1319fed3d5729398016f05f591b6ec424d7f5b5d0f0cc08b10f31acf056d70537c3d11a8d856caf9afbaa7cecdf174ca46ef6cbeaf896656c66026cc2f1003e25c009ea0e5361ef9783a6ef41240eebaa523bde4b039e253cd86d3d9d6fb7359e11e01802e76702ded1db878bb54c468607bd7e751dbea829ba7c6ba3627f828c17208a9e1db483ae7bade67dab8f59745c9ab84e42c203ab1867f493c2535d1e6bf88be4ea6524f1e94ba85761dc85ece28e3bac360eb320c4544a69ff9681a5dddeac5ccc625a2f391b5ce3c25ba2f2821e5436762489eac97a255e7917bd098da7bb0b52f965fb180b54f2acf11d1ce3f73d3a0a55b1d42eca45cbc8ab274e4eabce6ba4ea4d2d94fef882a0da43e750c26fbbfd1729178700617505553f561d05514019fdccdb0450a6891ef3975b6a692b951be93398c3839b785f44e794c737f6de000cf0b4b4773d80fc37e82c76d54a9860eb040087d8d00a6862199a2610e3be5c6a4cbce9c585d223118f8613432ca4c3d0f64277d81c5bdde220b9985d57b1ba75b3085ba45b03035e3608ea84d0e5d7e558d0fe578b8c9f2344e72a9fe4015c593dc9f74343fbc4852bf60633ad1e12a9d36820b9b880c4f1dce9821d8c61919400bd3131a4ef4dcf3f0f18f5f1bc523df275ed6c7b8a16f2d53d1462dae21151cabf2b21b3209db1c17b4a46450cf26bb192cac2d038f32c1eac020c73e5fa7f33a21ad58f63142fb26821a46dec2868f4c298d11ec2d21e8b015980eb649a974b5cc284cb93bbe1db9c4072cc4c34ee3db4589cdb3fe228d787bf514b68cc921cb315a8042f0a261ea0128f94fa3babc5a95d65406f7fb4e447b37740e1576d98ccc3926c891dfda6b8e5b53d5aac1225caad2bd3b0f16a8258fe8d7e3713953b8eb494748329b6fd8334f2a90b731cee4c3fadc76bfc1ca656c1787ee77c2a67ea1eafdde397c3838e2ea149dfd39abee9f75ac3ed1adfd18fc94281de1550f64420a8c2bf8f6ee511801aece1881a86a137d3b4308c0c9b469f98131bd305636adb8965f980f4eef2f753640284b3395a6ea81be1de66d6a8d4f6d14e674f029b8e8748728a8aba788e58f87190e108f13579973b428f65967b4e6676f87853ced2b7139a3ede909d9a125c6488e2955ad849750f11f320cca9bd5ef5c69f5e4e7669b27a34a73ce622947380bc49cd53f7e591ac57d7f8f44c3f1b35aafe09ab382b2da3b723fcd7b50852b5117dc6ccfb52aa51fc195f5b5e85d92818339ff33ec0a535b8d32b689c90898c9b5aadb404c574d1899b26e40950700ef2c0eb00cd96a01e5413d1847f335de954e84c00a8e68512c3027ec920bb01e196e04f302e978dd4ca9a4de871472faa3631af8170f0c8d20bafdf52fe559a5b8a838459f46219f284062fb881b61cf77eb5c9085d0fe722308e1b424ff9c12b141ac21ef84ad48b6d5484af9c53f1d24338ba35fcf4fca8b318c70e01d43db9e3865d3826f93c213b6f0ff6e31cb881cb400667900d9a0167ff09f567dc7fb4eb49b8e7b1a231acee90b5b85e2a02670ea659d2293fb37f2ea7037497392b93b4448b8c4e54aa84ed077608e8ebdfe05d07ed2c529d2500a78deb761e0eadb3048ebdfa02fef276d344fccb0efe094b875d2b231a96f8eb8197b2217ad718acf841fc332b7de1bde8413a0e63245f227b8b91e37bb3348350d3235928d65b6b1218bef665b5ef65a2e89248da75d1774b3d6fa34efafe2b42abdcd0ff0c71fce2ff5a7afbd537d57bd06b6a91017a7b90630e6133c7ae1c5d3244a16ea540b748f04f1930eae36fb3bd3cf8658d0caee09e53ec80f63b21331c354c9ae2eb2aa10f1e5b188bc7f765f7af267fa59133d6c61fd507b78aa71bcf27385edcdfd3ebf614482b64ba7643f6e3ff71962e3a1397d1ffea0a0d9b52d71671725244b48bce00b175c0ba9f7dfd02fca4f6503101e697cd1588701e37adabc9e78b961d7792fd02630ff68f7ff9f93bd4e0704e25ac50d72f29642378d3f6ea9592a8b5fe02b34821a08185ab939ff055519ece2fedf5cfabb99b16f03659f42725f5748d61b33312e4b3837c602719652dfc29c5fa81e802914fe37acaf5840e08194e94c5658083192b778de37c3b62cb0f7e24db9047ffa024101a9bc1af76fa72462845a58c43b6111700c9bd3eae52835d2fcbac9252163578378aa0381dd20cc2b964af8231117120a85895bc5c9e49c2e1a767ee58cc581e52747eb968d886b9115e4a9886e6bf187b8e8af8e01d3182e9373f525875dc43138e8b1285618a6eb009ae3101377427f2fbcae28146706e1e06e746813ff304675d898316cde2c78e7dfc834d476d8a4466c1567ded5676cf47b70e2084ba046cbc6dfd77a158bbcc875e0a2e3b994f66edf1e56354f42939777ab0480ba6ef960d0edbf8789c160d7f16b6e99b4e5aa560944210277c1bbda61c0d9dd2210a4944b787f50aa92440f1d10966d0b4047ca143f7f24f41e5b69e57bb085ebfba6c3cb29dd9fd270d129e403539414514dda242367d29492409f3990a8d1430de45de521cd85b5084ad01d6d45413df6eaccb23777d4030f6b1d4efa1aec5d0ff7f149ce8376c54f1a6240b85a77d8f0f714caa69c17a1fc7378dac962067e6e66b001965cee343e02e0613fd0bff2ec07e1c25d643979c8001ad916393def40dc7db6102c05ff6eb007547564d53cab81bdda02dc6fcb35a105d4021ebda53028e5f61b81c4c2c39bf7c91e3afde8537ceab797ecdc85b1f88401de3bd859db8cccc07a96f21939b3452afeffdd702fa02ecb02bb8f9b9fbb19dc0050acf97593dd5c523d3b10529611b32de70ba8b4074d7bb179354afc146b0b5c37f398eec1dfd7db8f1b82dcb982f679a2e31ce83abc2a4fd144a7cf2c90510eefa87faea8aedc0e9742c49f65717854f780777ad279896b4ed1cb5f00d65d6713c206011aae6509e75f1a51873022ed7c8934fc2bdcf226ea43b59dbe8f5e44c9b831b3ace706e5544faa30134fb5c72348051ca070d2c3962be6a6abf6c3e448d1d02f5082cfd2a9a2bd3ef1595346ce5113669f0e9b71d54e3f19e0746ac79795a3da1f0b02e5d1a6395f1ba68f968bc744eb1a8efe985310ea98617638f140e6a2604e0dc37608b9564c31cc558edaeb3a09f19add084937f0862fcac704b9664339527d1882da2ab36bc0969f20361096026df03eb8ba8b6fd9ed8fe33de3b4242ca6d6630b021b847e4cd276d1d4e17f67d820b02d414903b35d5be22fea26465cfbc2ca6e553fa8f03e4712e1f8610af1adfff29d3a9ba862f3a7321cbcfb52265900dbba9100b9a4d4eb9288d614335ea6dbe87387c84e345c0ca5351a01dfc479579376ab0730c8473909c8d2efcf64cfb01bf0b55fa7e61d3529bb23275a9e1268cdc10dc1e40bb59f8d4bfb9b1e320c3f4a39e810308bcb0c9d015280ac1fd444b87139a7678b2d666e7d53acf240f471d56fa47764edcd69c5b21d6f942d185468ae32c507375da1ed2f5d62481b249723fbcb045b055591831198e8c543fb2878a0848082506ae5d38e8190688a82a39151f3e1ce6acdd08aa9c814019fecf39520a08341530346d7922bbd5f72df1474da235fb172e848d78774364e2a81e71103977c064094adb2a8d9e7dd4e57394b3a5444c388f2a5efbdd264a0914783ebec6324e8ce1713cfaf37de691ba98842cbb92bb8af3c95fff7946c768ed95aaf0a855c0337ad368d283893aa7b00ee0b16e2e4abb9fcc172d0eb94de92356f95d610a02bf6467871e31fff4a14c4de64682f31ba154659dd9f6923ba8593d384f9e3b5b31abd3671dcd30c44c5f026c47ef1c4ad9f235f6e6323897d68347c3cb3d0daea818535b9119b99fc7113670a752b038b40f86644b84190bb56d6a3672428cb5949eac7446429ca5f1294ee3641c4f37ccf21dda0a6eb73ea65ca569527632bcbecf6157a0e7bf333f532f32780105c3c111486d6bf02ba210ce81b4346ad1aea37d89d0f1eeb8974d4a70cd7d04d138913e0644971dba4f9490c49ecbe772244582a55ec22fe00c3e483caf35a634124eccccce055961cc9da4ee18b75e66954915f293ea9183ce57d7f22c6c461a78ad1eda9d071cd799955d736752964afebab2af1bdccb4720f3937a5b3cc3a4b11c5b992b8fce64b2e583928e65f930370d068111c6ddaf13ffcc641f5d8738d2374fbb3c77e81c19a172cc8f3317e625402dc3a7f730f38b9c8981d9ddade895bbf2af58539633d5cd32961911314812bfc1166b4bcb6a6c5f127b01db03e20362109c3fb882a0a61ce28f401285966e7fd2b915ecc69e2c8c5048b6518b59b3516554fafef39620854d1bd3254b646aefe7cbb3784ad0cfe6e94c02e240a02347df7bc45178bb706034d21b4121c1eaf22f516dbdb04a8408fcf00b9471841121bb86337a807b6f5ef1b776860a91de4ecf4e07eb2003486769aaa10eb7b50ac47657b5d8787ad618aac95979c7c14109e8dcaea92eea8b3951a15dfd03ddc76149de00abc5d60e604f60ddffadd8a8d7552df032fcf8d7a275134af00bc4878bd50c006e9e6745b6ca85bbd6cf38e377e05d967f264772fce11b5623e099a7c998958ecc50764555c9f1c1c1fe0bd62725142a6e5a7338eb0cd2549b095900df62e00a0b648bfc288e54d3199367df774015f5ac9b807e2355121afc533921ac67f09b8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h6b6cf3598af280f070d19c381b755f5cee8bad87bb563ca5f84f022a6360d9bd8e149cb93ed9c5765502fc1fe4e1b029178f9193b762778db9fe8364dd592c3312260149d37fab1f9a9236fdc664cd8ae9a80b27af3254d4c431fb5b68f39a449c8e68a67d0ebe374d628513f85351f17b0fcd6c169b81da53a33fa9d9d8705dd1db30f693a6537cbc85902c6d34a37c65acf806a05df21ed93c72c35d2c5bb43748cf293f8445fe46de8d8b49f76ee263a53aa239037d45fa47acfc6fa25d0133bb516b9e2aec375367ecfe758312fa6c92ce59fb57f6f9513611828e524b5a3eb26a6a35649b956557e6470cc5c32b81fde0559aad3cd265d46fb6847f16163a1e49a7a322207a1c229c1ef62e96d8e6c3ab17def942c8193dcea7418746fba2a3d12a7924745671467678e4af3a701a60733072a905398a411dbe4ebf7642bf0cf35a6c57330a78a7312049cf26f38da81924aa36857c5d99fd187ff383cfb23dd852449f21be49588ff45bcc2d651f9734c110695d42ce0d5d0740af5a734abebdf124920e3e09ad7c3e8698245020033f9a6dbd6cce13835acc3275c8e146819d012e1c2bd53141c4b2340d7479b66d96c9d5a9e6e92b934a165a2565197dc59681be60137c104352102be4ae42f9bb847f68927a8f6d372c33ba27053835d532690e004f10ba597c9ce12e616fd0e76ad5a5e04dd05393d694ea6ec9040f2a151c84a72857c2f8bc4bdc80e664b680980658162075a78f90d72651af7b1efc23671dfb2b2df260974e77ec586fa6014ecde7ca23859aaacb484681278f8d783c1da9a732081d0d4a01b3bc2a460acd4f2b627e090498b4f945325240089175fd7a848e3bdaf15ab9629f4c2ca831c826a6d881c33048671efbbdb603bda9acfb6ef5b2245379d591013f00fb96ad4cea32323a2fe1f335075bc17f21ebf2ff11171ad990f2036ab95789b02138f5764492c649a2aaac94e2e9cc7a474fabc379bbc6742f750dc95c298880d38352142eb89e10bfb98e29c37fc80fe5ea5ba2d1b5747b5f2402bb17b975682de9aeb5373a42a726f2567dc9b28734c92d8bbe2cddc82ac8c4de5ba1c1d8409008e9006916ca1489b11552b5b286bcb6d5e4d75b67d211284e475cad13d13d3ca54791c04874d77a37379a9414b86809cddc6f42738adbcd99cba56347342a20e1a3d97db1f122014948f3695a6e510eaef0433ca30dc8269eddbe5c89d2f581a7fb15a2b32d1915e3745fa4e2d5db1da70b638bf1139501997e4bc598feff09e24816665710525a965e59743bf765af6bc6f7e622637c71222eb5a45a26d2988db0420bab2d239a8b94e24692a282a7bf52febc9ff109a98f2a20e2331d676096a3938a44c875c6a5c9f0f5b10c66207e099a6b57327b81b8679ba19ca7329e76feb6c567a1b400d4ad8e3a5249d52a6c4543a49ae8a47577a2cdbdc5c3965c71127f6c0a0c5847f82314767397787aa8c299da5992a681971222eab043adbf5a396f7d491185c018c0c91e0c768b3d0ca7e97295bf23d9f0b875959053a3168f6fbec30e7a3eb531be3ed818a9b578694750b6b965d14e760363a5e1ff28b1a03aa482d35055df0060740ca44229b1f20f87d915fb9d5319d9ab11909be55354a635e45133843ebda18eeb0036c678ce8005afabf6cbaadcfa630a0d24d7e4cae51569df46311027a12963da936e75a17adab02ba230fb328337425425ba1cdee45113cf746da26379daeac8d4cfbf74d7974480895d4dd6d94333e856914496de68912303cc13ebac4ebfbe1f1b4b3e6341cc25183d6e53e46b71982d5190c549de6773ef8588158171f096ca6c3ea120205fbf181f55a119ba4707f72034e326064fcbb29d9697b7426efaa36e9468daf3d7f5fb7ca8665c3d37ee51edfb2d8612889ed6a93281a56131e2cebbc8bb4357a3316c534a8ff4c9fd1305862a1006a41c4a385d76d4772ea381728ae0f52bd3955e448442f77ab2d39a2c975f6d7e3929a2ce5a6cf79eeb397657a64e71dd277cfbda7f9d2cf8e3d8f2251160c4532e97952d5dd8201fa2380766a6e4633386a1178a3c9ff2e7dd406b3f45e4795ebae9dbae88bb9b0e832259f67f31483c6d5ace6015f21c444dd0e6a6634298c368644b599a84917f0343cbb4a3f6c105e5ce8ef76198ac81300464b1d2ced0a0ccc809945f7480124dba61b7a47b5987b18cecf0c622458c02a38eee305b518afdc61f7237797eb1d2628d9c74d226b4b08bb2b72fdde33a7637745293e8a9f89c148181c47fe0b3a28a050de1e20d79aa07d19b8ae282a2ffc3ce6f01917deb8bbeeeb70dd285bf334f746c5a10efef9a2fc88d69756d9ba535727e592ea6064ff1e84497989b6907107195bf797759167409ab8e51513aad9aa5da5f51100c4e599f20ed00a03a71ee344bffd11eddd4c2022474737532a61eb4e008eadcb5325d3cfe71095544f3c37821f209ceb3221b5ef1b8fa8350f6b56f1e714e5b8e4b0eedb5686372d27cb585928b961198d41d675fd2bca9af1c5b7feb738e481df53ed0c60b97e44d3a5355d615111304b01cf4e0648d5fc7a2b3188f848a5302804a14cc3426d682057f87de86b572cc9dbd80f970c551354925bed7efa89989b21120985ff67a1bdebb48e10faf0bcb3b9e8536ef57a4bd140c7b3eaad03b114c00ea15df0ab9f67e052b6273e80c7d8c99398f63e88f7e1a2e59156e4e3ddc84aea352d7770f879f20c3ea657aaaf7fb08eb2473238f9a2a3b1c93b58d08072693f8f58d767b56bbea51d094e0a47d0afbbcf679ce87989c7ee33adc4419fb1535cf28baad0504528ef2cdb232aa8c585b96f68b158b731c6f89f25f2f65d11f363ea3bb3ba69f5b60687c407be77fce29142d4f4f9aaf7e7f37263137d7a1a73a3d889112924826ede9c0c1c73fcc0ec4dba5e66af8e6acbd8699d2351b2d010dc4d9086dd41c0fb80eeb2c5543fc69f1dd199b1a55837fc5294895a95a4c549412efb074065869ccc697aed98f2cfd6274defd317da50b3e71a45df1aa80a2e090cfc641d7a11560058469f34d20686717a94f8f4429174c9540313d98086b2a1e6de6f7bfd9fb46dc6f64bb6e5c05373c23bd7967ca10184c56f963974e1817ca26a5e15f7e12e3f1aa785551dc21ffcf87b3da59d9bdf394a6f341968f08542c0d48251379cc80c4d221d4652f7e7e9658abd9cf1aa6372f625c1bf00f9765dbe8177f2cb031b80dab43c9642e721b0bf0b90aa562c60796b07d4bc93f250e19417ae2745219b4841633cd7669c57c88debefa7edb2441fbb482cfd4419c4ac108c27cd9e8547cc7744403df43398f6b53652b089d4c78fddca4e787b72a004dce603be4ff661e033dfaab5ceab715d4ceebe88f135d1178b8309b9216aa9022cf666c2df28b274d3978e294ce40fb7fa34d97b9b64fc47fc060a1d86e637fd1ce18fc922d4dfaef3a9ec74ecaaf8b9a79a8135a888b27ac1cf91e951665686f3f51dc856e53e49237fde9c01834d322151d325b9ad319ff9cfd5e02536e97166d8513fa716b30ec1978db54516a56bfaf7e42e7ec5eb6723223b24515d9109c4b7bd261162a5b257c6c508459ac0cabaa2b82c9eea1f507d4c23be51588803004a71d59090513d724c7424ff06e3167a83cc6f8f89e130e823026f3fc92eec91803362d09b77d562fbacb4716e63b3853fee3ab17d78b7a3c13e8b3384dfe6d74176c619bff2071eb47c9567acd863b537665578caca7692ecc6ff89aaa1c7e6c3c02a59c2cded0379133b2dd344974e9c9e75344c7682bef60af39bbaa31e9dc12db1f3ca5e746e5ee25b16a35fe73b145a44cc352d90022da98932ad9822d4b4e9da904cd30c65a5a7a8c0665e1c47c23079c8987a1126fc46f5247853c59ac5d7508387641037260cd622f927f6fac8c7ea68092fab27f9de750088d66be97700fefb104522857f12eaedc5cf21ec1f2820c4e75a9e1c7d4bb7504572c3d8653516a7a58459366f339e30afb0efe7e94db43a0bfcdd85b603160408922f94c78c6ae0c96dc91f3741ec24f518efb4a62cb48163cf4e427bedeafbfaf1ed47495efa3b24bb7b8a9bec868920cf032507d40a89759626589924c27e73df54877457ac67e472b601b66699501ffd183fe5a36c0ccffca3d4410938da905475e069bcefed7bd724ebbd98cbe4cca425504a41d3a8ddce439c2d22dd1aa15de81da2db74619005212a9743561ecad741deba26e5261386ccc61809d0f74a347bf4a955739d7037718d6c2f70054b4a1a58d3d901e8b322dbb333a59521c6d69989cf29d0261d9d703f8c1bce6e3f887c51d6625bcd7bd485cba0d040e36dbacb8a8a6b14aa7f7daaeb39feb28a763be1be8065606d78aeb0259cc2e1a896a3415b72fec66b1b7a68ea61c6f44f0ba2cb64c93cde2198a332a2fa21659afcddcac4737db9b26f511c9dabd3ed7dcdf516d7246bdfff41c8f5d14a68fd21fc4ce3cea46a95926a749cafd972368445d50195c14dc91c75ed54b04009c028e37a281a2e27092a188c952a60252403ce7b1d40b7a60ee4cdf5bb31b632196176dd32235d060d2ed9d3610734f03c4b71a092d8d407582c9a74239f9746a4032bea54cfd4e9a695b626030dd230e70ba1f8318177ed572f7fbaffbe6b7b7a583d7f59ee24406b6eaf69ba81ce9fad70149e5ec2eb945f27daea8a73d92d70f039206cac42d411dca6732c8fac3bf4b019402433cd68e28b2c12722db882ae9ed3c032028e1e47b8e127ad77e885dd8a82402ab46e881e35b0bdb5d4d5672dd028adc974a56b7505fcc7577c5a907a28714aed6fa7f62468392648951e136a8d19f09bc4c00625d2786569598b36d3af86411083cccac9f3863caf8f150bf05954ee7342429e0ae829f9a879655e854eee13386b2fdf3d7ab245dc61b332bea9d8719a7f57e8880a7ccf8fe798428abba495bab385d2b8f67c111023fb19f32eda8a31df35a359cf2433a43a746b564f0aad9b5c86b585ab585a4ee53e62bcc7f1b3edb90505e4964b7e0eaad5d2a47b9fc8589d1d8af3a8a67389b1f8b16acf9d3a28961967e8b1d2c0fdfdc1226299e467667310591a30f4023eaa5d292fc03b66a9b2bc1b903adcb50d3f430bc41631e4d12326c6a82ea1be71c76fd588b37410659e1d3dbb0b3f79c590a2b7a81e63c934880707d1a0245346680444c35f04ea9596045f7c5fb0bdf5b3a88c766c2a7c3c8b3b88508fc58aa5cf182c90de2504460db33aab5519d5e0e89b9a9def017db775197024a5e5a5772e6683a4615ec6c51d26cedefe6f3667eb0e65c692c07b0a21c2f0f02a4002ff45454eee1dd2a3a4aca4c51044f29cfbc2fccd2cfd0f312fbd6d17d0b8b5f926b8aab3332cacaa45cff5d55e9c29a8a36b5c3dc378dfc5143e559f784c345d10006538269cf7bd68880e836970a0ee73772021d957bdb332eb5024c43dabc5b5ca3390760;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h23287c3105a34aa69a9cea511fb009d7c9b6ed280259f1541fc9d96c5c1aa2a2d3b249c085ae949aed385af864084f32b2c9bcf9cc5b2a4b0d09a12f26f551ae566546545335d13d052ba7cde57b267c5d58b549f1925e3f47573d924f76fa9c68e7a8d0fb1fb1727f3829bf717e323fdebd9ba4a7da22d713e4aa1028588ad604d415d64f70a690e6c4a34647638c8b2c0c6640e55e6283cfaa0af9579b0edff2f86533298098287e05234552c0ce5f4eef367d02bf2659ddae3456b3b6a739789ce07c4caf941e815110f0d68f8fc0705be61291c6c18c68cc7ef9c3fbf3ede1e33998b613100c2c914542e9fa4e4e6a6fb1f21608145d6eb7b25d7e419d9b4080c29d5a7883d7f886df8ae28fea77e94e9729b0e5a82cd780568e4e0de444b43338a2d66bb8722b7d7211abcadeca3936ed83436e5099cbf1288bf1d5c28711c498560038818ac08064026cd1a1f98f20c7ab6b609face8d205b3e8b1f13a0c156694cc5f9ae7da64fce501763d6cc905f78b9d504b9736b0d6f8feb7da7a10e907e7e4b21f1b242745238ff6ccbb30a8b518a784e3f804e3b79a9446095fbd56f2315eaf5b1ba3285a77ad786a7e118e81b4a1ea1e85b96704abd764268138c6d9ed43c6884f451c9dae353a6a2d5337f9abf43d45c8a585769ad648289eab7e5f3282ad535524c4435c407a81e3ce65370e014b713781768f27776d4307b66943535c08d6e35fd9f99aba1a47ab2274beb998a9c370a4236735a6e3b8403d53f0381c6d1a8d64de053c20ede969ae0829726d920bb99aaac50ef9b7e55c8b14c1935bbfd761c821755523e382bf667798ca1cebafcd4c4403e5f6e1d09d1f1f17acb4ce480f0cd1b4ccc8f08e10cffbb6ee0723391b9a5c99930be76d116eebbf326434bd394d00cd09b7769487479f886988baf26fab7f58a65ce9df2e6b9d64e3444da464e65717c3c8447a8292ef910e07933a10852f7f0f461180ba265afc90f549c4df82de2b0ae4be7e673bbcad925a107ba71699b90d9f7d66c4c9bfae882832b6ccf2c7320072bedc9dbfc6f04e8851dc9cb1ff2caee1eb6ca18026588ae350bba0aba20e19306d8a95e266b515e25a3121eaf5dea35c39ba8a8d69459bd97b0a76ae8dbf03fe25545de45c83901bd974b8e13ccd9d00af92c4fb52f4c128442efe2c43ba2a126e2fab21026aa710733c205eb547e0162b0b1d9fff62f9b96dd46ee057d677d67954d0e7c7ac4818b291d7fb6b3cf3a5e668ef0564c470466d22e27f731ab6b2a698280f2d855268548a4be9d0664ee4da9dc34368a00800a825467e908b8fb57692a2fe93f8bf60d0fe4f9c32f36d798b2b25a412319cbbd4d751921100faf52724fe063c0b858142e25b0ec4ba41b6274a857cb1097705abd874afa580562f382816e429b9d96b9f3060775ab88d89ed9aa1bfe2fafe20acdfb580ab59fb060896075dfaab54b04d342c86086b854944f14b6a45d9dafa7fd6ae9476839e1f7e8d315f90922d3ca890252559ffa5045ae18180ce364ac8ea900ec139ce98c5143facb424c2658fc32952a0d080df6c47af73e9beb55588de2bbb46c36067c3373d45776037cabcde0580dfcc791fde932f67a88aa4b0bd378ae9642278461ec12210b8b063caa88f0c285171cb77d9e42131103023e6c4c9adcc49919663c3d47081e2c1a07f9b5185512e9b32b707b7da8329906abaa16fcc4a72495da67c34abdff06b44c9ffd3a555025753fc110765c54efb36e7f3dd20f4aed91a969a580400f962b851a4151ee409e3d8b6e881ab13e2a4df7874d76b0e3d868e16deb76fb0e1bca4198fed0ae4272f2116ccf0990d8c1916615e8aa7e5a1a282fa7789d8c2190e11cd114472a6018b5ca933c7d1a70e667b157cba9d11730abfaede11f4aae745683fa26ee1ca44aacd207d6a0a425b7bcbce237f655fb147c12ae54735cc03d8edf7fc388019a4f6bd1e36cd54f248829a21a5e33e2bddb454b865ceb47998c4b0723f5cf4eb969428bd21342c9b53ed92adf2619ba4918ad5418d7c659a32e19355e7ecff78d12cd171e49892f3c83df5ba93d19cb47303e294565bd63a4d83e5e9031d1784fdd89b31efabc475fc8328fb739996aadb893cf21fff405d61b5f7fcebdf5148b1b96364dccda6c520a0b79eea9cee4cc62445e67c1ba90f0ab32aa3e78e3c8703de467c27ea3bcff6436ac2fc14b0ed79531d72b0944da3647ee5a29b533302674eee577f90558df1ee29807f3de204d80283ee9caa7346ac5c30d77a9e9342a9eab64413aaa8302c0a6c65b046815ccf01e6716efe68c39d9bcbe883fdbd6c20d1e465714ccc80558874307a34c8ee45821d3c6135d00352b6cffd5b0a8702307360551d00e71bd407e3cf9ec8b7e2db5edd5dfa5d6f7f1156bcd27e7fbcf531c10c445c8e7a4d730ffc2f1e5f76363628bc58f31baccf8b20fc9e6b6e69f18612a87f5adc1a95be15bd255331fbe7eb8bbb9266be23a1b6c169601945f0109463dc69e3485f34b930710c9949e3a06c6197f50fd5b0843a9438f0ddd2e1960e55a2d347e2a7ecba49b34160a152b73ac3fef5af95c632017925f90b51cc7b69cc4eecb13e46bca999afd3d8b2ac80446f19c2a83fc64b815f17393ebdc0d8e60a24d4420e8e24f99665d70613e8e3c3c398e76331592a7bccef5cc41df98ddb8ce69dda58568bb024fcbd60ffb39d44ac8487af14427270bd533e2156f0e543ca7c60add8b8a0dae5f88d525e4bfcc786caaf6e466c5b8b679341e40ffb2f7461483346be5c842ebbed56d08914f56121a4f6fff55c816f86894dcd93c293ac896de5466d08d5fc8407ce4950b9bb041454d269f975de0bbc02ad1ebe54329a6c6010fbe7a2c3e0d225b5bf380a6e5292ab3e5e782965c1b84f8faa357e7dc7dfb32a96491a25ab7cb3b8cc35b32e44b1204151b0efb7c6f361d2603f28e1cb5ffebb870563dca07b6390c6f82afcca19fac8e53ea1f157851c470117accafcb94d0ba83d9e78092c54e26e7c0699ad82329d323b8f1f25b99ea91a57ad2a48289891611450c0effb2cc352121d9f532c390e40d2531fc6e9c3dac0bdba5fc2b2c23aae76a8694018d19c40f7057e9fbdfe0c2449a737e68991c5c6fbdb9f653714decfa2f1c29d27c6f007ec1d77cdf50f7d0c159a22958258d80f46b371426bd8a797775fdd6128dd90f20b2262a81b1522fa807f06f5e6a6effaf02c51b6e87cc09f624c8d7b7a16b07d6bb3b084c7d471faa2134b8b336ceb2e3bf34e7cce2b6739783d3a86df1e7b46dc505338d8ec1ebf5e3a7d89ed34535c45cf716d1eeca10e635faa30632dcc9ee7e7096e324a515059b397b68e6c61b27b812ebfdfcf6b386778bb653309e1dbb975951515bfb4d8c80b780ebb6939f8ce11e4f99033067fa957ee99354d55064a8a822168f96975722fa830bb37aaebb3bc1a4f9548bdbf38071c088bdb27b84d174f848aa471e0f758516a50e53b1c538e0d8e470accaea4b24e7c9b5609bb2f5c889c1002870aa8454b8332b2ec48567463ecea73a5cafc878b80b34ceb1959404d985290a536ad4fb3fb427c5a7e8182219b603783499afc92ccfe35d8c10d12c993aed8dd387917382972e2ddf9410d632b1f16a9f298cc56bf3a53025bbfbe91c770ff381c831c1047f70eb331620db60cb0039c22eb6c76885652d96c1fd6973b83f0c98659e4a5004e49bf5fa9972ffd169d22accf6ef57e53520429a506ff42bd3384da080e339ceb2e37ecc29331f368d4de823373e8b40d4723aab13fb39945e852b33ed2037f42895eefb5c0725841b3986de06ba85a1bc0a10d9df8d6bea7e18394c7e8e429ddfd6c83b30bd6d5673252459c054e725f86c9614737906e667be676275b6c4f152fba515018e6d3581356b3733efab0c2a5ff399773f3458c4122aa859873b1c0f5c966bce470fc1f828b75503d3fb4450cbfd071aa1a352d7e03308964ec8acbcbe8f19998fcb3b3ea80ea5c37184975573d431bf2fc3d76d831dd678439d6ab310fcec2e17dc5f13b2fe45b2d85f25aea86b77056377b9ee9430922a7cf6d519f293db100b50f76b57624ee79b3914ca8ae637539dbc5db0232fbb5ed7d3c39037a08171a1e561a267c991f9eb0ccf0920eae0b7b601f9d9835ee85b15dd32b2ce5d4bdc94b92fd375103f5e10e92d601d9ae74d87a0e42d2adae06422da654d8cf9a609cd9881ad1950b7aa54b54ce18f676a904983df87695d7d3e29110e4ca2148822231663c83b8f15405141a309a697079210ec86d31d8d136a4957ef0ba7fc551050e539cbfac5cb0acd853def9788bc1fb5ebb5272d4c16766dadc0e02c98450cf771ad21acd33ff897e8f6b1f80bf8b54ed60b1dce1d99d9e390c348fd4c63e8d518f1417cb979762753795ae128dc13cab75a5b34ac0455c67b575b0fa9bd4af454680d6d74244ad950e385a1aa228df0b09548c68abd70dcc0600d69edddb7be9ddb5cdde56385e497d97127ed8c962828b5c85a95b4d490fcad3052f91ece536f5b3be384a39d639511cfe5adb8051366e38a0c9b94c588b6ff9fecbc7664d2fd4b7e430592c5d43f38cacab1342bc202378fdc2772a95e5957362aefe409d0c8294a6b99290e3f6b4266cc5f079fa99754f4901e9da9f36aebfac6a9411de6320f2f746a579e6757cc2b0d081bcd75c85072fd75718894c34e1c08182985ff8748761efefaacd7b270a761b0f11f31071eb97045db12853666cd0fee7dfed41f9d55f838c5a97a652ba3677bee863b9e12050c626c50239ad055a4823c167a96d6602b820d9502f2b3c40d8b4821828bde2faabde638448521b7a880fc8d7e988a2c314ef730ae519ea32fd19f5596fab9e4225b8ad2ef0e96530aa278bd85e820325378f3fd6277f2e7f2817371135bcac09f5969d2e3b6b323e382c650c799ca40f4431fe270e3eed352424cc89e27e277aa7a46c8ee3262c4d0f1e43265ba3732b67b3e3447bdc4bce53c208d2dc450c8cdaf95f4d129a63c5e459e59a31bf995d262fc260fabaf4d70c5fc0a83373c3c5bff65290c39195eaecd10032485bb087146c4623b76b9ac3fb1c8409b57434080bae276fd9077e5d32c384aef87b5ceaf7b719a49508cf77b9c814e3f85c62c370a4421c33306879508837f78ff7e9b3a3d5725fac68d67006e5f5392e9e1f27b7bacb4916b9eb756c9a64b13fad1c2d86836db01b4ad499496d07fbb6079dff0978e927f3e400ca0314dc726828b6035e935ec2d5c47e858478d3308b4a5dcb0cd8b523b4d107ce6b0463f7b2252d82260bd7b1010bf7d14b3eb49aa318e558ae6275c68ab41bfd0c189ae79bf05f6aa0e5f34df865a16a3b6e30a96b2418c873534d1f9b8a7a25904aeb32a6fff0cc432e49e345edd7c7faa694c63df591db5127bdd7a10fb172e927aa052d2f6904b11546edafbf55d1f945ee1f441f88dfadb13170e4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h34e31cd1b5cfefa6ed07bc4754a1d8738ae33b8f2105c0bb1d5a35ed7577c57bb128359b9c1db827cbed93baa1773e4750e9b4dc8d4251c0289e47e5a4082bd7d9fab224c44128b1f68c61605e2dcdf39151d26750459b2fa189eebbc27edfae9b0c18d31d60d5008c1a429d2cefd2f1d3385e89da57f603cd841a09763075a8441ea0ccf8ad9e898149ccae64883f6c93cd230fce3b66860a31b6472230aca1224b8ccad2ae37dbb58ce670b919c17a6371dbd7ca77411d90c504e099b7965665663d1a0c622d2874b3d978a1cc6077aaf89346aba7bda3d28101ffec45d2e613a2a82b8be1afade3177ded09fbf3a607baeaa1098daf7d6788962e8e86df6636a9f8538c46e37770e6ef839e4280977f4e11d9e82f4bbc50f267c4038b1789cfcf2d90308736f50fab09c3801cbc8f4fa8bd864a41a38ee1faf08acc4dcc0b3c6a47a0d136bb16e08dfd32535c4399c6a73af54d5c864e75d13e4ad8a3e093a668865cb14f122344c5b4f7fc8ee45430f8975bbc8e4369aa622bc945973b3e72f9d30021f02a3631e858ada368744bb65d142ec82ed2ba0a959caa0e984ce1fc5810b39915d07c76b9c03c72d6e8f8042aae89873904de94b35b283908b8bfe176e75bec9f4792d0d933294d510545460ecf7a68c33eaaf4bd04d9cfa2fcd576cf9acb78b4fb1ca1d2914a4c7a631710910b9fff5c9b679dd10763eda5e91931cdae87b82b9bedabdd2e2065f6044c73dd5e65c10fd90ae9387e4330c5bf95d646763df378a5f8a9e50b673242d134b5c171abddb59346914dce3690ecea5fc343f59fa6ec1cbc15f1c11daf360ea9e8943eb8c47bfcf9cad03e1b7cf6ba79f47cc54f3c1d0d83de965515d104342b21816aeb69295c204721c41c16e1ee4aa6fa3b270938267692a367e441353f7e76a0aa9e5190e5ac758a2eb09a0e7a14a7b94a7caad0455b1867e02625fa984de7a49f74f168d0bd25683994ff941e4772f1812e9bc641e6ff7ab7c3cbb559c125ff8306fc2d4dc985df441da28a88a1e4dd7e35b889cf81b4a86adb7a78464486b3dec5d6b5952c120aadb209b2b53f2feb982dc6c2710e59052f5f0750f8fd775acae4270094768128b4c723d05cdcd6588c80cf8d5991e15172856ca229264ea5f1c96df39863e2385d386e5cc39ed8d17e31068ba42ca94ca51718f658a5e5f9d6190bb8b2a4eeeb07f44e3c38b8e0e28f4f9e47f18921b5997d8c9a35a5d59be3faf0e3f6e0a3f022f4e58abf35d15cc7e6077fb9bbc61c88a88df170669af6c33b6cc330deff38525f41f7b98634591a306e6eb713c282b14ada6ba9beac98b4f667e2ac8a122e45eccb78697d1c1fb16868b37c8b58afb3b1588bc1c15ba433b0fad02d488ef5512f918db7289f0e7013ae8c1cad655bf4fc87eb72eacd156a8ca86a7c1821d25cd9e856222c2366f23f762531f217f11dd3c8bd24ab546d99a42fcbfde114509867eebd393c0b9a37751db534cc784cd640e8f3ec4a8477ff57966036d7d310a6c9ffee627c433fe1831936ad62653f0ce0955c047d5da473dc63d442ad3888f721f36ed1908c2c229b65a5fbb7d035a5a91c0bd499b99d8caf650c5be05f678496348922d0898d5f476e33af10379616b3cea6a6f0e4fe385ccd42b5d3d405474d293b0411885459eada2e911b767e797730ad62a594686113cca79c25ab596c75f25bdac95ffd2097de06d0c82992999dae4b2a28f45f9d152aab9174893f9048723ee121899c616c0710c8bf4615352d3357ef8e18c2d956c1492fcef326f94c1f7efa97958964a8e6b4eb661f09cf00b89f798952cc695bc244d5b76cb2ef929fa114c55b68afe9bcc0fbfdf0b189b87997788cbae5d4dd0e6600c0caefa3519620a1c68b7a427160153aab0df28515368bd03ea1b671263d77f587b88c907428df7be30109cc2ce2746a0070d2dd88bdeb4ef267db7feea223ba7919fabc8d9c9aa983f7e1cbebf354da57081359930357113899d1d602fac827051637ef135a0289e750c9c3ee0a6349dce5399aeeee6b5c12400a297a25f8c30a6190732e03b83da162538e2c800d0526da0200848d273774651d770814d687c2687ef2afc75aae5de4785664728fa8293790b2b60621deca3024d9df6707e6b4b621f5f6eab05b13a1db1825063e0d3485e393910e0ae5d96b22a3dc14cffef708612ffc7914a6118d31bb97d82131ecaabf09498ce97175ce494de55a99be73610d4ee04eedf68f1d2570fddd0601ec0de99f3a47e25fd1fd717779727e78dd1e14720a9ca8a31b659d3f2dd2c532f161e06106af773ade9d42a05409c7f3d560d2f71d8c564dbd05513d46e0b8cb52163f5c051283bd08ff287bb516b5b614b1450cec226389e99922abb9c660831719c6072ff8ea5d0e44239debf3f3491f7a56be621eb4f9ab62ab019d3667486b4cb1fdb737cf29cc1c0a2ed05ba45132b557101af984d5680523f0a1f98a13f837aa0490e759db9c4a008ccdcd9942156cb9731f55df032b53ae15deb5db4db168e3e432d9c0cedd0dc17f190f1bb85dcde9c1966a2c71ba718ce65457ca9218c1f3bd119cbded68e34b0714f268c6bbe780d9c518a08a18ed61340f026eef09944c5bf1c918494b309da2576754fd6793ff5c3bf506dd5eb8d632f26a1216e3d2c200d8ca98849bb98058103a0529a8e5e29224d369591093a272278bb0b2b1f35e45981141efe459f001c80474aa29a5e421dda96d507cca70f3c01a7cb559ae1269b64daa9ba2a41cda09063ef20a7dc544c4c7c9231c622460312bfc7acbf25429ad3ea0e2245a556c35aaf8ce632d6aa01503571b7ad4c8276401d8ca7f017b00134d7ab362887bd71ed262b5d3ce4515435146f9f665d4a6f33a0690177f768c79fb42f1a0b9c116c3971d052227cb221b8d9c4bc7ec575037ecb2c6949bc938f53a2609b0a8138af67b655de65f877250274718e1b09821143c2ea25434ae441ce299399fc5fe2086005ff8216699788680ec1f1be705168b6e870ffdee8d138a480d995349455225dd356bd86cc3b7b1af5d3d2a990009358ac9a3c3e316bf96ac122dc09cc08c1ef6f44859394ea0c2c95d356ab45275fff9eec2c568f98f6e4125645709f99f699816108bdca365f4eb90d9b195ee9279496fe9c9c1079e22d8272adfb80b4574e8be4a3f31c72f5cae7cb8b6b9f3413de9a56823480bc0ee2a6f96cd0b18a60f79e0b16f156637abb25fba660245c11729df2d87128e8c67bc53318b773f99934482a399f93b5e859bd3ab1298f51c94793e7e35e4920dc60e760f3bff84266947720cebcd043f9b5f323f8ba2aa70e46e17667aca1cfb22941c63a2841ff57b006e4ec93daccde8d541204e6561ffd6534055d9add2e501c51d7d1495921249e59d4ef4e675a5a30a2ba60bb78becfba8673f666cf070bd3e90c0d3629f87abfea702f3fe14ce9900505b235111e31e2327a54de2b7a45d0abf3012d5f8d0c687c469583151eaacf1e6ca1e1c23f93c6be1aba93daae7ede2b2f227d246303a37ff82183cb674b575a4021126ed9bc9ac6fd36e17cd311a62744c042c61f967c95de68ebf42c95d9b6eb8286c55f9f6d32211b6ce38eb492dc0b901602e2045a25efbabead424831aeadc3b839c45575aaf030bfa0aa4dee3a2a695475215b53d63f5ecbb6c454cd35ad25b1f38c675e88a647dbf5de0ad916ac584a95b93f20a5366403575ccb28cc9cefc931ec7217595f55ca34100204290c62e509dd9bf7fb9f2933b65d5f18afcc16d030c9448952072c26f8c997f0cea995c954dd266706ad18a8d42007788dde794ee107d3f8ebc27b9aa8afc0d6fbfab95b3f8d599a4560f34f86283291d990535b1164cdd27a05a1b625579034b7ac3744d0d2cc00b46a19355af927eee28b3d1d2c1f319ca5abacf04e27dfc1d2424aea688345d77a71801e01a80c4291298440dcde7d22dc6fdef55c87572b3b2509ab8c79015a8d45cace0382cba2111eb6dd529e5e718904b026a06d5e4bbb44bb71bddbee4c6f30c093bd1d2c6ae9d0b069f6e3a9f53e906995a4bedcc130fe2f87f294ddd865f15006a56df2080259982a968ebe0e9d2af7058739dc0a0b836353aabdd46921637501994f74debe4a54cdadfe45843b9aae569d908fa10ac90e3955267af692c271cd0d34b25708a42d17153b387a91c36d9461f7ef218491eaf0da8852cf878c127caff42f0b7d9d2c4c160aafb9b3e7c8e7d39db91c22bfa6099df29cf03d9b4f6971f665dff7e5797c79b2b5a32b2d36bdedfb0ea2d253bf3e03e4ea82e95d525055af28521cbd8963aaef0ba6cef6704ea2212b2ce9f178b69eb46c1211fd98caf9e0d4ac26b0f2ca025d42c44b76b26d7bcf6d43f955a1fc1bb068efaa167f7736d567fa230601bd82d24537e42851237dd384a962e594f7db05ecbc1d7090a1c8608c3cc1c093cb2c9f49146e666ece44c4520f34e92818afea48b95ada93fbc8db66658f98a484def1c0cdb5456781fc419b753412353c338115f2fed84bcd2097f78676757c8c9c7bf2caf3b96e50eb31f4a8aec23ab964f0fb5d928ca531c44e0313789c18ef11074c6b204795db59c6d5c701310910f71834127e6477c613ac0a2423786c9b9f9f2ddb27260f8b382130196247fc40afd1e6eadde2bff31fcf3dad7a1b40e9a4b662ae24fb22cdb57c1683ee06de53fa4af2e5f6587629f90aa7efeae2c50495e53fdbf4c6f8716704af8ee7e190c4fb08e25a0a8b635652e30f11b74086479a51ff2ff1e8a2e69e4c8076c6335f7a7a4b04834ac41cec77eeaf303aa383b06a20e27fe3a83992c62741a9870e1dcc20086582e3527e6f03bd41ea009d0c699dfe4d9f65df455755fe0987ea4b4b76f96be12da9dd9dfc879df580526c880a106d0bd1788f076f32f8453494ef9d4d51c7d5c96815c401572b531fa5c4eb24d142f5a7952807145416e82809e360413dca1699efc4bd58e9e83e5d9cb97c479ddb4a8ab61ec67231c335265ce432841ddd70bb575502f1c5dcefb2a8d90309e498f0da1edb81e98edd3f1092b856d4fd1eafbc3de5c62ecfa802146d1faec8441b73e328725ed72653f0bb7cb3b3ffde207a0474a53e1a799034a78ef2a936a3fa9d17fb45b8babffe71edd76a7dbc3dfcab5183be96777a8655a9b257e56e83c56cb90375b319bda8b0911861792f441436c4f833c18ae747edfac8bf51267c54491f924a2d7f2da6703ddc648266769e0738c6cd7bea1e180f76d0a33667e658687e25b12ff5e72522845f1994a2b8961a23e8a764aa56e466d519bf3e864efe8e249cd4a3ff55d74a88a75e5a57cd52daf2ab81aae844994697f132c9ea49b038175f6625abe7b9566f33abfacceeb808da99be585cd55ad9dff523e265a305dbd94d653d49e6debf9127091ca9e2474acef1c196f6762043a48c08ac1ccad8f02bf29ba8fc7a38e0f1fa58f3b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h1ccc065ccee52f45c4822455ab22b71eb5bf35355da0f422820e8d694e0de5ae7a7111a25430a150fcdb136672563f2292e62a5fe878ec9eb5ffe309611e4fb6adeaa86c6f36903cb7a4de66bea96b151700eba3d01fb7c090c3c7e8c624d09359bd68be7dd0d326292bb96daf4bd092ba89e6fe213101aa2b1578852b516344e361ca2f084aa9e029785bd9c7c78a22aa81f6cb4b72872a3b4b09314f2b102e92f90aa9b8e3291a7fa3c73b41e5f791bc1346c0d5760fbb942854d90659980c3e4de1d39e6bb3528d061947931b0e671d24e1b0ac293c9829a0f1e12383ea10102159c93ec46b7efc4a773494fcb217bbd34a433193fe57556a5af6c7c470df2c2063ba46bfd9797968f71d36739a20c87331816dd5169e13563ce23771b1e9d68945fa013cb1e8225f0d3a8932d1b791ac03c9c0afa35c2d5a6cf7d15c57cfbf905fd1d18711c09ee04fcc7d7fb5154b929471dc4d27477fb55e454ab6c1af300c991c9feeb9c7c6b837871314fb2ee6931e5bc344770adb20fee54031e8f1613d0677c0482e195933793c1b906597dc9eebea0eea639ac4b903c68812a49185411c6f5a06b6c71be1c933c1b372c5b3ac259dd94d32b2d8a7630cbf89e161805f4d187f3b48d08629f2508bd156914c21ef796f72da46503184592b29490902bdf2cb610625d9810ed4ff74c3e773ca6fbb29e7f27b97a8953a265d943f221395371011070e8fb68f1de709daf388b3c92cb85051e74638525918cf25ff0ae41bde615a9da430db7120fc6062420e79dd8db54c4cb62c0ea550c377d823578bde4b864c7b24b0743f18bf3e5a6f7a9b0c648226b6d77541393953da4996663647e52d3cdcb5657897c878f768b3b94eda05784f92921ffb2db8b728bb724b00a3062bcc9a62244f6053d6e757261e63f58ca1ce38f69bb4b9eb2107264b0385e28d70e7dda4ef610d3c7cf8c0ec2a20f6c3e53e6f08faefec9b9dbf79eb197704c556b525e7eb93f136f5a765e0fc869d0baabaca1a223fffa125fa8d7053daf200187e4f9aeacace21630ec3498a32d22999164cd675c3c5401abed0489e0378be4d417aacc7caebde95aee921039cbf12a7ea9ff536cc85661c3fdd561647e8ce0faa282880a0636152d3918be21214cc3ed2c2ebbf2ab009fcbf29af76f41f8b14881f52d14f0a80db445301f5c5c0c99ddb55eab1c4fc27ef7ca9b6b2cd900d9f91b16b0273a1ff049bf968d268d15bfc89b44ec49086a3f0baa3882c9429d08e72d142eaa8df71619e63d7c2098c78325a097e4e2c904152dc17a4f0e32cda2f08eb30779166fd2110ff23f593906914dd9241096b2e8b6203c718a605b0f43e1c9bd077f8834237a8271b25504d425bedb6bbfc1f31c1670c9bc7f46f0a52e948738cb43a390a30d65c73adab582e62bbc60b922d560b0ebaad08b18b29999a63b7433186ec6204659009a012ada4d098bfecc81b7c52bb4d10550a945eba66746b3683fca433c91894579bf1c29d3ebdb3a870a22def7397af4996c1dfa69f1acd6afcc164faa25032997413629f1b2f27de557338bde208db74b48abb8c89e022f6d436074e8728b3dede2421055459fd2e7f7681af594c6ed565aed01219e8345363b6aa81d57e693317c570e9032d724148a558bd621d3474986196c21aa2e0c842353ec4c152c03e9950f066f742fd63824e0b21f5574108bad3df4901f59ebee612916cde8a07ea021f016e96570b91ead947ccdb532dde6d1339f36a6d24725c558a137a7e65965754c9eb54ac76b9a68d5495e118a1aeeda3d7deb1ab39da72b0ffc1f1cce7c4d167f1e89f2848ed48ca4a5a3ff8089e6c55a937e637e9f89b305b1a641fb75f59afcfd006ade82e61589d0e1a3fa449daf7e25838774946df43880cba183e7effcb40eb0edc1df74019e281340263e864c062cf5b506dc7ceaf817bfca4ee5afd1ebceb5b894f0cb5869f99404fbc89cfde743734b7bb8e29ca596bca918dc3e0a78c84e95a815e7060236cda564a44f5257253e41be867b348c23f9273687d812f3de72f7a540db6e1735a8ba8be411446de3f6ea6321eddfb619aa49d5a7be7d069f6b3d945121a823213b3bc29eae081049b7fd5cbb73f74df57d1569adaff2db6f17174f2a31373a4361a2e04776bb5579729ae258a37e8566daad07cdeadf924d2c5651f2830cf38a71480e76e4256a845616258caac60f8fba2327e247865761bd71b2da016037283ddaac63ee95684bdc6c8b3be72a0a8c1d1cc01270e4be689b61dbf961f7bd280e72b38714210c5f2c7432c6a117693eb9e08c192287c851421d0876faa99a51ffa3a7cb64d962954b56c4037198fdecd004402ecc1be4e13aa1ec952423935007d3e8ea96d0460324154b8cf94a40879c419b9d2e452538c5399fde0f22024e04e940b9993c9e997232ae2b3594f8e57627ed82ff316b7b9ba9ef6e4791fa563cf2791dafc3a3cfc0c25894b841ded26eb20e0bc97d6d0dcbed395009fbf2a567a984b8ff72b805866730774a31db06c5aabf8e78b563139bf6788eeb462b4e76089373afa9e95a17e411b569d16ca487e23a9d5c0094d5a6651db7adbd5978e416b8a903308934cfb33679c3883b77e8329b16c5671c4dbfb7c449804ac3c1cda9a8ee62a340fc21ea9f8eeb935e3987f7f6a94c767b86fc8f7cb4137c3a33f39780b9f23f9f457f946d8fad4665cf4a536a15a6b92bbf910695330b3f1e6ac98d9d97a5ac9a075c8e553f0635db3aef0c06f86e1ed7842d60e0ecb618a06e8a14632c4601cb56408c56f342362e1fa369f18b928391dc1c66a4d489ff3e472623b033d71ac5bdf1f7864656fe43cbc5bc3ee16eb11f57db2c302b1f1a4bacf513c5b5e583cdcdf8b88b39ed49f3a55c62d6ec95b9abc5c5938f159b4c5a2dfdc8f040badb3cd249ab8f02ef28faad26c78246b1e04eaf231bca96ea9cc224e33d02a238b8df8ffb18ec0d029e056b92b658e66889f1f2c421f138eb1afcaf72eed79d0de094bf5990b1d593d4ac08521b8e592834910741551c6e4cdb00a3e8537c6f488936c6f59b717c59460a48f4bbc67a9f41d2c0115ef5a65858a0cfa7fc855f4d6e4ad1fd9fea85323ff545b6102434278490a132114330e0e70fe57c61bbb84d1bf854d1e45293e7215f1a4be44c43a2badfaa5145200c17e1178a6f2bf5d4fb7d58386e84f44445cf8ee265fc24535df9cdec193e8ad5353b79b51d6facb047e4048e4548fd99eecf25987d54d1e91ed6385294bc6685cd488411d6ede525a4a24c9a471f90ec77000f10382b3bcd6b7a10813cfa4efed6aa96d56485190aee5b0752b142ef5ea8eabb485468f75e6ecaa85398579ad6dcec417e7ab4db126e9e843d0ca7f25e2b7453a7cc12ef5c48ec4e9fa5b4e085d87a874208f96e14659ee666dede56b1b8cb19d7d151d6ba311db2095d14f85baa046f1118aef741df401a19f00bd26b8f6c634224e3c085e80be7c9272b4284fd36cedea1cd0af67c0279d8eae2019a9e6f571321cf66862d71a46afcdaf5d3799733293e73d6cae32dbca0eb91d5e0aac2b6817f593d63897b055da2383add2b6dbffe0a1b55210b26b88fb83a7edb6d4c9312664109660471f9019ae27b3e09e1de80fa0219b71a34a43615c3a9f622f76721338032f9ec685a49597fd68f4e3bb63b214c7b6251914e57838526821499766aa25b214da5d158a13ed39cd4f15ee4a251b2f85bea0b17b0807115d935b6fb04bcc79074fa127295b574435d126d3ea73b9f975a3bf768888358a8e0405676c64d2d7968d8171855e0bebb08146447ba0739400e7f49f8f86d675bbbc31e10e22e1c2873c337ad9130b958aaae6083909ac66182af818522e8743d785d26fedf77915a2adf8c1d30fddd3b1ccf71224d47effe519082f328607936059f8e56f32435e01c9820245dc12375a86854fd8e6b3b30def2e9e2dae761c58e4bd92d726a7dbe81d9cf82a62f98ade4a4ca184fb460bb1095d9820bc3d286cd22cd30e7dfcd9887184736e0777df2534f89e5abef09f62476b4a4ba442c64e68d4ec1d95a8d86d8f4ef57d7395448ef4a340f631e09a16e6935f0093278be4044a48ab5490742321101aae6568fd840bb06a2a872f20ff3b5387a3fce90af43c87f7cb72a08c1c031d407f57be4e0f7790983939a3ac12e9d2cd9e9a2d848dcf97281f4c5c7313ca721ef92329627dbf1751c30ed49727ff258684cd3a2a9b089df20c7d49986d4ed32e9ed1e1978088ebe06f1b5807bf3516be310371846bcb8e9d6574c8bd2ba73952d082eabd333f290ebf6f15d12c9fcbcb743841f3ad670ec142c4f6e8367dc9a602004c0562646a5cb8b2984cb95e76013da9419a4fe764c75a8be5cb3ba514c73845c04b369f494347f67628ec814a18a094272302133299b8c25f9100501de26bc9a7fcf1c5c4c47852a1ca44335c5b41bb7597f4a12a8e5d79b2e075071d5de14b74ef3138af9a2d27e05d24f4e9ec0af1d858b68acc2fdff4094c3dd21e52ea91e4c2e398b8e3138350cfb8a585435df5a45abb3e8a9860e8cb80c7604ea7905645adab133cc8361b25af419c673229adca9f0c6c6eab302ade5e6173952c60591a1aed1ab5dd288685709b92cbe78c266adaab6aa5b2be432d18b3a7eaa0d3ed8bb61569e7848710dabb2e13f51322bfd89793becca8ade3374b52343e6e934679dcecadd6c0624b9ad4e17111adb707a5bdd87149988ed19a8f7e3917bd359b00cbf5de9b08612bfd6a521a76bb2c2311bdcb77f3f3cf534fe3e37ca6e86816a6d69e05fd4e9475c47b60abc58b97ed87be8f1109776cad14b85662c5f4879dd79b290fc8e0280df9611f56166e9702811bbdf26a21491fb326136587d69d412d469e7dfec860c0b2a3839e8cbbf97563eebd534a0b8799a5a5d450cd29a2f027bf4623313648d0507ee7d59fc5a83c3c5c029d31e68afbfbffa8575762b9c1208c3ea93b5d9659d2a67b129b6b114cf566539311d06b992636d646f12e1219e58e22459bc10b5e253f2b7ed5ae38c50148d1505b407ff458f6467ce78abf131787b7cf59a75a7fe8728edc5f37ee93ce2e2e5ff62bee66602555c2e30fc80999b847d081bb2857b43576b09517fbd9dd2ae2edc436fc535f411b43a17a15006cc0fc80d86048ac269fea72b8f47308edf044c6182475d6ab22de88a2763db06be189513f559c1e5d8f7ebee552030488784c349f97e7b5d50544b5ee0fc5e4a5a6d51b55c3eb5a877cf69301ca2c6c03f6ed7072e713c6d72833fca0a0f923cde912e68e404b2fce8d6b889a3aaa62fc28e7740308e24c1029cba6a0fcd71465c9d01a3c615428f2a553ea8fc7e1db7dd4947fc5851ecedd9b317c4b49195e9dc76bbd42710fa2a1a5566e60e5a170a6ec130a480a91ee1cba45e7ed2682a53e916aa7cb08677ba8dde34a624835ea7d3c781d5744acfc46d7a7a199;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hea8126f758960ec93b68ccd3444dd02fa1d1a726ad3038da483e2117b1d5a037e9b63f83f30022be11a1bf117a207c88230da356deea2b1d0506375a020e72270343d0b02edc2432d4afa964dc05d2849041dd2313c45c92987b91ebdf55a5720d0e3333d8069b9b054e3ca8a577ff4b65477f496026712a410dd438b8f4eac0bf1f58d514b4b3571222fecfc7c9722b59e3c90ea0ccdf330a17900992a9367ad4f0b49eda20d4b3727b2d58f013bd38e80acf79c3c2193ec2ead94b909cffe47d350794652df84904a6e4b496efc9fafe7b0875e55ff28ff5df90fd69b800564174758fbc6d1d5ee362f982f123feb269006d616d240103146134e5dee55cd308a5ef7cda56c04eaef511ed29a91dae9184f4c7cd2b21b1e79babd699668503fb296cf3bd8da2be5aedd322bc58b0e4f181df8427909be90f4a7eafb8d56498992553be22fa3ae208b5d3886b1590069de5ecf98705021de5d973dddf16ef50d239810edae7350c235019620f92b0b168ce4bc3d97cebd8db4b195197f5f09c39b5b6884550f899bd19d412b14033629c8dbc8fe03e579f9d9a756528d287cd0e3647605bb118b21dca62061daca548f86f55c5146b85d4755ae04ac8d9a96960c3ca403678b83005deb8bbfb9f20f34aecd1f258267adfc644348829276f658a409e081d31d10bb685a308128adb0297ee001ca84a4444042dc5436e38e9f0cff11620505ed915d3c1c8f76b127a280c14c682a2552e1753f7342fba24f3a2273c10729801f1a3b934e4108d11cee9e6b9ae2425a01099a4bc60a6edb2553de49ef19245158009e7106753b5bb70fc6aabef1f7ef9626db2eac8a17da0fd29186ca91ca7c36538ef8251502976c0066e4c45adafd78efb5db4a0dae2f60c636b60e3034dfdca906af9b33a8ea482309e3046883993a55c54482f2561b6a69e36a50460d5ed98878a1583beb5309cba3fb0b5f6c17b64261304340f0229937b21038d3792995318e89d08b3b390f62070cde1403d100de730a69a2609805214fc0b7dba7637f0d606feef3c1ebc318fe87876235108cdacb1a223d7f4b6e3615c8e3fa1c5c11c82e17e4b10657e2451178d44badf2ee9599e33959d66fcd62510508767b92257db3e5cac35cde85761e73f3538212eafb30d63638601a5d5d62116dc30881ef5d38b030eada2ebc987ae0901b7421cb5cbdd97e20cede9ca21c989c21d88a1ca38a1b8aab776a669f445a84be88fc95684c0da8505d8d4e95ece806f1cd7deef94e2c96bcb857c6ef1f6aa3ad43ca71c98a4e6f51e1b50602414955891ce16e0e5f65c0e7fe54ce22ba98506a7a5466d8f39bf4b6dc28dbc4e5a6612108ffa154b018ea9dd7511434fc468a9d4c045d596673bda7364fc2f575d6835763b5466c843d94ac7dd8170bd5d9e6210d83385180f9a0d124a50950c471cfdb08c3919e507297eefd3c0eff56cc50919eeb5a2326a1b3fd341b3cb004dcf8ead04799f29e51276d14c093b4eebaa670a84493917ef172d9b42297c051b95c5db29737cbc10a93a2a39a08a6a83ea46a6d86e5bfda0345ea72e31ca4614c8ee8bc2c59d05cf1da928113ddf372368e8ae61c19507573a6dc78188d5e5d13965895e5ea1aef0e51754e3c93090e37da57754586b935c80e414e038c5124d7ecbeacc78245eb0b09d2685f9b623ba326576bc079867c90077ed6e48e879ed801ff8ef91fcd7f46d883aa7c2b526b832bf84aebea4711a3b6fed65c02a0799c3c708cbf7173b73ca2d43aef7bd53810fb4fc939755650bd10de7aabdb326f8daa18e884679cd19dc1097bb4c049a929937f846ea4934d3d83ce259487237c2c6394cb529150e652be0143ffea3ce1f09aceb2ec8a314785977cbee3825ac0d0a4552c0aceb366d8a1d2262d17b55491ea97d4aa72915f7c1a2aea70166eeaaaf7dc2206fe22db4ee44ffa9d1429ef818cd72a10cbe7f86d24abe3fb3c975f720c1d9a53dedb6f21aa21a6e5354d48e02a478de7ba402a6a9944a4f2d99ce9df56520801c893067c2976b1543d330861f0bf9cb7591afb06db591611031d18000575b1a6bf37f56150c46c12c481087f280a44651d28f72dfb42aa2a37432021e6fb7d32dd368be7b450ccd167d22ec864fff2f3cfb5e0d1fc51f6a227213b0a9d9e431513fbd6956e9314213db6fdd3afa8118160fcfb44c6cb163a52df1f5855b37ce1b01a783a9440c48d13fafbeeff20a543c64c5c4bb3a1651e4e1d6e5705657b8e77d6539cf6954e7c448c20acad2716dc1bf90dc03d777ebcc1bff09564b0fba3840a09555bb07fbea2da691114dbba6c455c5a0e23a8343d0d4b99a5d24f5f606d40dfb9c915dfe21dc72b488cc3be8824402c72f9b4a11da5e93685d1af02b4802ad856d09171b923bc9e3a325f155f7d7f7bc296f3b8e387f7d6937e9af0da9ef1d3f5688f1382996eb2400474c2c6d8917d1ad2e9bea2eea619b922d122b82001f3d88a71700826591674aaae6919ad439eb595685be89934cb5c5d854878ae3c390e9da63257cd63c3bf65a47c823c7ec5f7ec3e6d55ba918e4434a79f68bbf5311d0d78bb79b5fa3b65c949e4e7168e92ba6d20372ad404fa1db88ddb50ef59412e08371f97fef649f624e805e99a5c103d6435ad390b27ef92e83acdc098ed9cf8704e99b5687e0f7525a9d8862cb96092d95b3f6993522a83530438dc817b3da7d254d2b5e8e01abe88fea7b49123375407c512fae4935be747efb087f78c5662de100dfeb047c4f48f1abdaade4b1b4b277d0d6dce4d59d2a0cae9c6f5a06bd18b15b31236cd15c423a6dcd03c15f158f1b0e8629ffad718838a48cfbb4846580dc1e4eb07908213e75a065df38e10b416a8af8694a4aa9555e6079058cbaf92e3899b37be96fd2b0b7da67ce08aaca73ade3e40332ac20b1bf8e09a8dac71914e79ce5092c5cc56d4ae1c42d8363c96efb6348032eaf2ed777088630cf80064081965432fc00f17a68b360bcf341004330018cb897ae2d00ed91a5c42cdd9c606ab9e78d4bab8f71d6acebf529052cb80ad101445e553845b762e4d486c475b7e5ce1d9ae5ed8ab58cef202954fb8de3280f2b592e9f0d5897195209c7c979a7a12b8c624b52d423411609fa3d1bc259a77c7b8637e2b1a7fc4f116d433a373bc28262c3d2963a9a90085d9c54f486968a2aebb18c5e2ea5e4a8049942dda70316b15c322a25d0266445797f59d440a1d08fca4181a2f1c0f3f97855d04424250fc7e06ccab868c011dc16add06c4133bbc23844913840aeee9b90f9f332e702b0187a399a781f8d0d235919ca01cea07ddb25fdd181c334f56f9d689ac9236cea76431e056ae1ee949e3f5dfbf578bcb5d6e4abd7e1f4ec377637a6989638fb2b3697e9e0c00d548f683bb4f8a820e200ccb902a5b96d25e7c3d6864267c652f5d810a5c484208b3d0b546a90f41fe7c959fc483d3868cc671ee3879b10672beb31de5f68fa6249829b90e33afa9af3aff56881a7400d7eaefa52746c7f153bc76b113175087b4ca016068adac0d99e80a1e64475ae6866c769d3de8b2ba15864d341cf459012461e4cd2e69f64b24f80a7236fff8c80d385a2d51f6dc478046af02b462cf5e6b606331fe033baf21b3faa3e01aa48170abe0bbac63bfd0dc9503733b82cfd4c862a9ac0fa3e0d8e978c1513feacc252326d3b3e1210b5b92b084139aa1c5e1e3808b335a14c8c32b27726fd3ae500f6587a334bc602f68b0f6e86a947e9b973cf3913aae7859b0c9d8b2033560d706b722d73feb8b74bd99e0b23d0d61ae58cce827065cd409dc16e01677ca9c8ffeb9b2f84688e2bf85276716830a4c8f7dbf6a8e7713bd3479535455093d83e8b9ce4025e5839ad360b373b2d88a5a04e02a5de35d6242c7aef5b2c657502949be94e760e543a8b71978829cecd4c984d246216a0df3e6ac1cf09445bb62f5e48d546c16bbacc6945ae9a2f74605ef9eafb3a7895be437bd8d399c62f761552cb0e9b2733edbcc9821e165e9bc99c3886aed214cafa476e3c1724e0d8d6ffb866bb31c86b373ef3e95e661b543263ba8ba7480c89b5c43a7e2bf3a320adbd2256c020ea740113496109a56f957b716e37f0d96b0b0558ccd5b49aef8a34221c39b6c8a01b95443223bd140443b11dd70853ec58040a0a144e747d8f5d5735cf29a853b0e0b2256fb07b3cbe09fe85835d4757f65b4ab022ce5f322c0805df2f5c5db678183639aaab0498d02d60d366235cdac58828f01b644d9c0486cd77f5e784c5830a027c7940a54e621df30eb8ee8c9d37e164d709ed2bdf14c098acce6518be7686b59b9eff5b94146957efeca56deb3e2eacd29444a1656affa272e94fae1f2ab8511ae21786e3d92c96cf0aea68ec7b3a57c147cd7cbc49c9c19664843c7d64cdcb065b4e347f76694432a1b51bd095ba38a40c05171843ff599e0cc30c0f490b0dc3d3929d9efbe8fe6c91f1b453cb6097131372881c7ab8b0ab84a2dbf8e29634bd514661845e0748c951cc6a00f4726f8d4aa19bfd98b35e6537c38a598b5fd1e76216db0664f7535174b547504d5e42ff6fd96dc1690ee613d7f56e59e9c17160ef825e2933947df29004bb3363265e99097a8fa25dd602ef2607df9f17e07edd967543b872bae71e994e229fd9010dba502fe5dfe4d35b7a1ff62a71a1ac0c29be49de21891290b18a137827f9fc367d2032346bf6d440ea9234428686e93391087a0157595a7fccd838b1cbff5517d6f9d196bf3659502748b7d4d97105df9a004ea1870c4f78047bf3d7134f67743b11b1cc0cb18f44b83f4d3e3832dd7971f5f4d431c33b8732e388c68f08c88c002ab9038a362b14c27fc6bfe8f9a18da24d5b167dfdc4b303237bcf61800be9f1cfa3d5e65738c846ceb1b818602f07c95d8c5f99162deca8b3cce19453435804d3eabc514d01548386f0f9de19920af025b571860b7aded464d82eb8804fdf0283dec2de14798471252d0aefd3344fa523762a165f6439eb95ff0976041e8b4237d72e017c255238135275feb3c4de8f341ca081f77f7f9ef702533bc59ddeafe50ad6c1ef4a7cdae79e1d297cfc298ee6822b2c2d1d2d57039c2aecd9ad34ea494c8f5a77eefd83650dc6d1f3393336482483bd97d53ae922b20711300baeec65896a3b01175882c565d24017644578759a68aa47611f96384f282fc6bd92815263eaacb4711f610cf04589ec5f5768624441b50a62499b336546d248aa75e3ecf584260ea5ea8d2cc3540f066f779290f7735ba3f42e49a5e452c095c4a8ceca653fcd84b43766443ed72a2764988d4093ebd7219a2876f73331a1d46b7f9a11ca311d1988380d9d7ecd5ef1629929113cc3177f604de65ebf6dae6aeabab7a8c620aea3e4db727f22f3ea841ded0d80f6c891c8f88ca1d32bf08dacd85ac2ede959ba2d514efde4adfe1a52e07f6febd796aadfa266f0dbb1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h1add15d92e76645a4b35a1335191a9e991b07bd707aa432b4031728d2c83115413844b956b6003c215e18fe97e6e134bcd4c240f3285a6b96467c65eaa8341776d7cd84fa508c9d9a00939e78b53a80da148ea4de97708df7cf94bcb798f32e7b6866d567d6f3a10f03db69041ccc82af14aa99973720fc6cd5f0170ae6d0c90c85c944e89db5d08eb36534310a839ad4a2a02b543368c25c46d61d8839515141c7e10cec761ee8db9e9dd96402bbdc5d322280812ae75b8c991487cc6e902aff4155af86f6e3f69281b9fb92cb78514ba5e570d24931c453ac8d7c6ded0aad1ba32e2e89d0c7f28ae9d01d53ade814ef64ab2dff2df4603938b1cb48b6289dd2020899267afcd4ac4d75fdd9dababe79c67c1509632af70fec4b141b5128ae0baa6e40de658875acf396f1da0e6bc0450470361155bd9f47f8730d9df49073735be096e8053bf81794e23f448fae0e6c8633d0b09cccdb7544b2540c39111dd76d6dec3d5d61b369930db5cd4ef51bc274a5a6b66ac85068aa0dd9df85d6d5cce931a4b0bd1eede293259946a764bfddec0ee8dab2da77e2fe8b3817697618c7cd7622ed8679d3756f05e073f14d67687007657efbb07de2e32abebc508ce7aa87d08ccd8c16c4616ff0009b9147ba104bb842b77284ea037cbf765968e8fa5a40e3158e886da4b313f20427fdbf6a259aed29fc05f5870e5850a263c43c5acc10008e8a8e046b937a844532e7b7a73e12f76262720b6cd818dfa95421ddf73e10d1d2fd9b9e23c438b0ce921ddfcce82caad3ea439f6f935e34bf54f2d2c7a2e431f92ae69b160cd18341f88ac135e17ea286c0e59f85fcbd837e9c2ba6f14eaef50acc6249c27b2b62991461b9854254e9e5f137165d8d64b09eab600b9655bc63981ea6296f7189c9c11a1c74e0a1d3405d93dc051d0a7e6f99f190c5c3d54df1ba6e029a91d92482706913d01e571286e0e1a14c21b92796baa2f1931a06a041b15ac34568b373e74815435feb789cd58e88e57af9a460792bd8a63b6910ca6466b6a8ae066c504b14927371c2cd33b323cf453f7d3fe2e9768f561409566f37e6f856ca105d2ccd7eee9a81c00562ecdd06610b348005fe34789cc42e3de0b1ed16a29e6d30f48f5b2388adb2e45049aa6729a627190e0cd060a90c9f891b2d851649792bff65b6e8bbd2bbafcc7361393197b467b4bb0069d8a3e25754446a65bba952e42f4446939eed022ece4526fcbf4b9008fd3b772794ecaffe6493a08413fb1603d5f4adae6ca9f8095c59e6961b8e695c69b4695579a7a2b02ab432c1f02c7953ecbe973863a4243ea332b84d4dbc567aa9911d0de5d64601ce8872b6effbb2274c4f05c84714d3c3510fbe82f0af2b507bba21c84cfc092513596ce6eb72cd6ef4db67c559bbed9c86c9b18b433b60e0899c7b24f9b8834b561a38dd65f3cc993b74a7de926595cef1fbe97d7b66ef0c70b67ddc3ce69d383c918314c763cb47d91d46ec4d57aa75cf45cbdfb3c52a4de8cfaf53699d4e87a9cb64acba0b248fa8d85d69c4feea96b2e07e65ede52b03cce69b6e2b1755eacf5cad407ba860dc315836da7e7bfd7544aa3181307ac8969e0d7d7834300aacbf725564e28aae2b53fe44648a3a5ee9b03a239aab68d19442b8eb43ef5d521f7af03354065557b912263baf067624199fd664830413d8101d134f6e7679c8dea1636a02cc1259d673a220556e5c4db2d6cde427025796e025ef7a728f723a3cee1a2e3842be5336380614020fadb23dcd4d073f0f73cf678b73deaef693153e47a6bcc7528a9acd08059f04965cec1417a4064a24aff963a6e0b4debd72c88b50b8e7536cefc88abdf854755f65e54f557af853a26f9f15a5e5b395b12ac7e099ed3f8e8a016f38397cf1473ebfe1c6383984cde78609bb9a23e9495b25fb6e73292d708160738976de664c92e286eccbbcf50a82562c1793d24a8ba66056f9589ca107b1a662ba6ab496608df217b51c00e58e77d604b65d9c1c757973dc56c50967f4ce9eb5762acb0304d7ea7e87097093e8061065c620c24d172d1e6e723c50a9971165ed5e2013935da7ad66525bd118ea36a9ea93ec85e7391352a82b4dbde6a2ecafdcfb2a307da8abc5c97c3abea07f3a806cb2165f77e897afc7fac8642c4bf3b729db9ba63fb13609fb5ea59ece97fb82cf5a9bb5fbdc35b5d32f957cf73c5d9f3445a2faf825cf9c51bb53ce55eab3b08ab3b990dfaa53eca2824a2c01870626deabd586a8769e16ec26ff17051cd21759d13dac90d4fdd1142204699cae3463dbc14473a4bed7f3b30fc6f64dcd1e99c4446cd0fc587fd63c5577512e991d615f0bdad1bb1ffb2a8e57c7d7475644798d5b13f0e35a381ce1ddb18d7815acdb51b06a09435faab14492b1a2935efede40b62eec7043dc0bb5660bde64c267afba0005d6c04b09286ab865911e3f6248e5001fe18a1501509a89e1549ed053f5fbe1f6d7cd3a9063c4bdda697ceec617292652c5eacc3db70a76a2bbc8a5b1629aebb2ce24943f06826179936e4fac61e3d0912f98a68210b27a821559aabe90707bfb677b3bb84d9a5b97e5843c8869e9754f38f401ea7b84d8b17c7205aae1b47af3309f54ebf1ecfb41877241b1a082c4d41203df6b4149c811a438024f0ff4a688c9eabf06f3d97809c63c0079dcb7ffb00ca4ab847e419f05415ac24ea23e666fa4bc6807dcddc22090402112d71bc95ffc8e5ea825fe7c8463c87d06b23cd80a4a0cca9ed68a883aae421ce19c3523b320cc76a01911ed030e19b6f634446581c7e5d5b9eb6cdbe5c4390aed051ac4258c02b97c1968426b53cbcef8fd86a187a91aaf935b50d409e4bf296d54e3c20f6f4e52c0429fed2f153f0a75d96b376d84cc993018036ca4be7f7c3c9624ad9bf7cceebb616edfdff9ed333577e3b3183588b70160a6ba9822de65440086cf16b90a8cd142aae1a121c998a8711de6da9c79b8e8498f30fc50f79b40917dacd79d7bd23d9d6580e220473bfbdfb70f5fc6857ee3c77afa197e5f70ac19c17a04f23ed9ae9f8f4bb1f7c00fa09b060d9bf7ccc5ecfce52d86878b78a68178d5ce9f2b42e65a029f658f158d20b1db75ce4d3d3efeebb4a55e42b801ebe05c5c95e91863e7169b534a3ba70ecf84323706d48a788db13b8625c87b4a44e891f44b7579838e95bc61dc9421ed81b9a6efc784e1864949eb36c54347495ba855f328a94f9fb55f9f6c95a0aa780c53b2d5657fd569d175e769a20e25dd040c7cfc2875bd44d0a9537cdb9e0ace4ad7c74469a6501cc7e78d50b48eb4e227fa6414b1631f5c623c1f936513f9577bbaad9e86ca39ef062a64f7d554d76a4dce847be41e1aa50eb36c8d9faea98f94b55576b22f7b50efc9721c1e724ff0661a78867368de926ab9f0c5a12f64feac1a4a894b6ca0b1c18b0afe05b3da54f7d6d78eb27564ad134e9cf31d5db86f5b37f979a51beb8d58a03add5845fdeafd0d16eb78648b4782a0e73a9e58374f10026918a77248a5e4e0614cf512ff5443a208987d0d88aa75ed21929ab306bd74d176ed15636c88be24b02b349f7b7523125d0f3bc7cc8c138e6d9c625bc9a7bff7a4af0fe037f6bb66e5066006fea889e0f29a009d95e1d0e15aca4075015e7290960375c906c6bbf2adb60c450ff4fc0ca7056057adfbfc39c953526bd95a2c120e8ffb8d4911c18a5c4e46daca53d9903652219a6b8e93f8f57c47505f8201583f43f2740bddf229485a922b440c6a4bfb5215ad173e520d8387e47a809231e10b02b0dcbb7627898e371bdc7c75991bfc2c2ecd172f1bda43156faf9288c1b53b3347c0b770e73b234e15036856b45389a4e853d5427ea425d40e21ae353b3cd707f53dd43c5ce2cee8f6bcc2999b857c67d55eaf6e20d494798b40afc5bb681af1b5a72a8b2ac9cb7ce5e3866095c1701a8becf8157404d0528bfaa13dc80078d6549313c440c01b0abe69439749d10fc556d977bf52303ac790109b1de63ee56346e077fcfc181f651b92f93dc583b8d837e0909aa6117a2ff789c4904b84359aacd32b45e7c8977b75e77835d05b6ecb3d6bc3595ccdae245003e0c70901afaabf442ca7ecb5bba2eea1af7cc8ce8b5f8e4207f6bcfdcf0e8a4c80fae331afc7ad98c7c8c15aba912e4c089afef4db5d10f7079a34603112851e0fa09a793c93d0568bf95ac77aedd0124de95ea791dfc85b42c33674123a1bd18c60d6973c2470e9caba103f8f4f0d1d297bf8f50c51bc878e9a6a532de3593c2c9427ee1e4fb1123e85effa93355b9a562f230c4bad2feb88a65c14c7df6daebba12bb9ee47490f1d5c94f0a5c8086cc1c01b229ceae629f32459542a0c5d4b874739dae94406e588648ee8f4c1ce0ad9b7d373ca9e6322f87c5f57f01a498826b772b201961647c7bd2e4a8ce5e069b8118715b18d65c3c9a0fb473c9241f19874db8698b410caada20c4924880ced381895bf81d4889b0865548a545e8c51a82e92bf3d2fcca6b5195826244660c71841a07651c84bea9997f4cedd4495943c6dbaf3e1d8e142601d160fefb57b6e4431cdedcb701b236f1f767e4a7e03d745b800535264a960617142e27b3ee57686d1d7c5b3260854a10ccc145ff38c609977b08c37547470c27d0a097da774ea0a0b807622e59bc2bad64bb56d2606393af26c7649ea70176761cee69a61f35f04c0a6e37697ee03acd84b03aad2ddb9830a950f9391cdd35c2d4be7a2bdeedefd0518bc9d8b8a3abdfb4fb115fd3c5290907fff706086a1fe0dd9e422048dc96e427c9db56862c45966577c23a637aefdc98a4a2ae252d386b406d6a5bbfc22029e9fb205bbd554341433ee8b6d11db0e0d57c9101d98b75827e504abeb953dcfd68523027fa857962a19012fa0d2eb3eb483ff9328f2ab62b657460112e10c0d0ab2d6f296904c077a987e18435ba299a92561128607ea7e06be3b3163125817f75e9ca78d6362dfd295173667b19b621744a64d5ec7f85a4a5dad352040e290022f70a4e52fa68be1fae9555cefa7cfb5cb8b5bde9e3cb851d807e0ba66a335d0e6fc273cf719139bd8124c96bfd1ad299641d097c98ac607f44047b55208d12d2dfb5e2359312a4539c2557c1cff96a26d32c66ab39336152da57fe60ce0253f520239b6e50c839e8e84b9357a71bfaf040aaf50f1789b9b3224149624a94c9a2d64baf06fc37e5fa718318e2805ad1b7d879c2b298cfcd34d03862761ebc5d6b4d33d7f1c4a12e4d82da8697bcbd107cad60dfa6c97aafbcb426df189f604f6e50582daeefc0a5b13edccb2c2d0b140c75da917aa42ce54a536b4a91cf934cb307f85709f8cdd3ebee977e6bd009531197ba8b0588144867fc7277e36852da4afc7b12d653d1e004f029066c0d90706223aa10a748c3c5d20f45d0b6865eb957e75d9156e052e009cf8ecb2df29b6c2862e7c46dd10150f12ec2bb7b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc69aa439f0252925eb901b97cfcdbf6f3c25fbfb452775e8eab1457719d8d41eafbdd0f2dbb202b89c75a4bcf47d0e50878bd5befa6be9f3cd862a1bcf17207db5ccd43fcc5942ea83fa8aeefaa0828c583300687a44c0ba8ea57ae7ca73733b37447d3d00920e34a26efc7818c5fe6ca3c0700469824a9670a6580f45edd0b6b480726db3ce74ccb58329891dd12c844782cbcdecf3ae0c7889041a7db5e1df63afea1d95c6e01a3ea04b94d2b0302c84dbec45a6cef2dde8d8ca06c12ec2d861f1f198e4031945fc485b6c6cb8282a64e307fd0190c6f37fadd514bd3c1692ea96bb9da12c7023496dd75e9b0752e106d2a6fd5ea2ba4e2e94c8b776cdc7d9fc854322e60b878e5e14cddaeb9326562bd687f4570713375ead3eb688b012c5dd447a1dcd0dc3bdb0191a4dcd06e661af9355c703860744579a7ee8780ce373e512fc69fe2c8ce64c60bb7c552846447af72175ec050bb71cf27ad244beb09a4132c785d6ec7f47cdf5fbe5b611e0e3a388d54e17a2a368ff1e48b2872021edf35710b41e9e9ee1a4559adf5f0403563abb627b9212df57b2615b4fdaeb93f497c9498942e6172a9866f20b700b22d8b1899ea4eab4352933c0f91bc923c3f49309dceb64e2df7dec94312160409961142f3367834ccbeb57182dda6e937d6efb0665481c87fedf1bcbdbb572a39285115db64f93ac3d1643ca6fd6b3e86888171f998fb31a6ec1440e96612237a622c47d49d87535e5ea7d794962bf82558cc686047051f072be6a05e91e9639b4ded6dbc0e0e74fe5f88e3741fc302cc054611c7907a498b090b490955c97541de751779b10f8d71cf1ef7cf0fd0720404a369c5513abc7d932b1495b3e2def1f866a3976159afa31080e4bd705e2bdefe81aceff1a88f384ef44aa6d14415d077be71bbf265a76245262ec797967842ce7229687442872b66a6a9c05ec001d47f1ae884095ce1644e3b98a37f407064670c40246782b93193a36b99745c654407237a6185f68fdaf5ab0b4cc6617b37ac13f0c6e6cd8a4532064f24260e3d3d7846a1df91b8a73a04a088b98080fbc25ddd844435b0bd4f3f36ef461209ab9d046e2d9df1912c2e11afa6fdc13696b983164f1d2b971cc300b6ae605ba92c1a25925dc7c52f4acba19bacd8fc4291d30125d762236459ef495ec0cb87ba104c5d947b527a71869c98a470a0f767e69db82efe9ad39c1d8bf16ced2012b3318f59a415b41e06ee6ed379f218e18f3eed0ade40ba4bb7231a46d645b3da34bfc2a5ab636befcf192cd03c621086a0c2bc7951af8946b33e47f335cb30f8efa57275c1375cf165da36dfcdd60a530db23672301ac74fe80a69e374d411749e49d7bcf522d838ebc63617b1bd2bcd09e4e9aa11001a4bd6c4292bda222fc7b173cbe187a23435708ed9097be7f98aee0a668d2ee30cf91827eaa7707531ce59669de7eb478a814255d72394d8a40418f8e9910cb7637f524690e98ba751f63f37bea1ad8e14a95989b2195b227ba9ab6aeed1aa30df54c10bb221f1449c2c9582879b70105413f00997e5ede3d68e46c3329bc8d78a11ab5917fc36197b20102cdd05733509ef455fd2272fdb85cb554806b53461b36fb2305521ab7dfd05c01d87414648590760e5dd453f230e91e8bf52cb40cb8a25e346d69bdf2fb14105fdafc1a93b347545119b948a1f4d7328888b4490062d544f6cb8f9bef44fcb46c8aeadfbb9c7baf8c20b0619db065f810a6f19090db9248f709bf6008a0f20d8242c9793c19544cef72e127ab01cc57e380a06a795ccc2b2f7919ea8e9312f486f1dbb09aa6696aa132913cda279f4471d26ae44d8f0015ed7eb824e1af7e2493aa5a920278a415e2233acd0ce8c0b250c590011e267010ae232f9d47270c102093bc9ce32e1277a7e03b7a3e3e8d789b0a6ecddbaed63e4595c0bb7c6d6f2e6f4259b0abec49cd08df59e13132d17bb1e2d21dfa51342f7b8df5a45b7fe8c99f6aecdf24465c6aa20bd61eb885e37002f20ec10fa3f7982ff0f2f124ccdb00cb1024bbfaaf10a22b40df052dbb80d91ff60cc7e3f4d231799e9d3439262c85c85b98d9d786240759a23c6ef4d4fbf630ccdd831befb0cc81d8a7b63464e30c5b2a48490e10cb6ea9f6ad4baad00f38166c51509c46b1e7c360369684afc844e4b795f251b0d52066ca80ddbc778211bbbeeb00155c12db5cae59b92c7122ab479efa74994149f314962cd4da32689bd0b01a883d68019fdfc92355019f675280cf581e77ae39782b466fc60338e9dfc3e2a6d19bdf617a285aae52098bac1643883821011e8b6cfed46acc2e5ec1f410afea3b619746758a923c553f716d6dfc393d592623e9dc1384647668b372f364cc54c41798928ae0ae1e31e96c0c25fa856c40ea5637806a4426931b8a0de5b7fa055349725e7265a66cb409f2b508c5a324da441f5111383e96162a4e0c6d11aca3f6452a449de30332491bd59b228f249387cab39656ff23fc4940853e53aacd84eb76095fded8952ae8f142e364dbd57654d8aff8a6e27472d8ced0b3b34a9bb9d5c642b3ea56aeeecd8d4a374a044448431aa22842586c26ea81721399199f678fef819a2b5ec23f956a79cce2ea3fdba68dcc55abd5f3b3a88d00eca6bc069bf830a840ef215f758ecdeca806264bb483c000b48a77530e9a2c69a347af93c7c33216d4b225eef8956bd3321abc2041f994f2ca94ca1e5a0281ec4f9960f841f6e4de1cad57b927c214f49f230702f5584a122090b965e710b7beddd2599812e79445723eaf4f6bab1382e3baa907c0e78c0a80586aea0756078d585d3ff0988e0c78d36cc5b48bacd1879141818b3de230f46530ec78c85f1cd7ff812a5c5636d40abf16a390bad088fea1abcf84d494362e9031346a76ee00249fa2593db16a69e71fc807894af3ce84d0453738e893295987d77aa819a8e82be0e7ac7349a3abffc5e51bfed58d3f6f59347f6ca6eb55ec74b9c2b1007efbc4295770a765966d6eac9417abd9940c68eafd78a647bf270b0c2448eebd3d368e022c5fe11bfc3512ae43a63b78dda0f70b1420c343ea0df6cc734327b8c029ca502e3afc57311c76f2d7e08551a6817a7604b231873e680c9862fbc40fa97e5b576ae5b8cce245cbb3b10965f94cdfee3d75aa4aaba2fcca05f49a837a3e0d6a0ac3af428333755372ae54cffeca76195d027de3dd285450eaaec3af9748a82662a4310d9a5de1ea6c4cfc8ae76b922abccc13097f4f97d9847e4b465a939207dea44c66f7624152abbbb3c74e53c70477b1065534ed62ee0697c6f8686ae7eb2bc098e0431b2761e96fc4a64a5f40266fbe4dd1280a32b95ed1ecef5d3833101fca4b586143fbd6a3b12262f3e078ab2dff4829b1fb148f0fc69b96079ca9c8ecb5336e74e2c09044571ec24550f65e8b63443ed2be08c08e34daf82f4758becc84906988be14245ade23732f31cfbeb9a3bea1b8d230e710c5de5220438f9a41751b0005264dffc644840591a82cf31b419ca0aef2882cddf0d9c9dc4344894eb643f505d40382874cfb0d7da9962ea757b040376d9ab39954b282617b18df6be77583caa9b8419ae2b7851686e0e03438aec92f9fac5b27a871eabdaf6bb760c4afc865974d0b9c4eb76b0957696cec83c5e5c9f5266848de005c34985d755624c68c3263fd5e572eb85ad2181654a7b2df362cf0d2570c24e48ab85601d9d66f0669186c4a7da313464ffe1fd50a60770e1bb990a812464783530dd695e6076830ccba13af4531356fb02de0a557799875a3d7913aa1b79c06920a0782db3ec4a1ba535704b5dd3c23ea87f959432134194ced3415ed0b4d2ebf71bc00800e2331dd9e277841c8342ebf688abea0fefbc30b7e52d1fe9ae1700abcf52af39aa049fe9c2caac82dac14d1f23f1ebddbe3e3acc368bb05f2b294213446f830dba7eb048361c3623e8154db893f62d9c291316369ba3ff5caecc2cf862b448b41111873394f011ff238916b800ed65092f501c18b2f21d4190ccd9d5bf6c2d6a35f3fc54aaa1842c988c8c09dc53c6d2f2ee142cddab49bddedcb17739d1a39418c58b3d239af51756500aa1c16e7b191c935ae92879f6f2d73c91e48a85ebd2ee4cb57d9e42f71abafc5ba8262f309dadde6bc2669b7bf3026efce4964bad11bd812b33dec1b2c98c92aed161835cbd25500f661464df877732609c24442e86761c77256c790f072c414836f4ed40a08fefb2469bd5caa5d0560f7f75fd723be76d642d8cc5430cf9a84474496c06105c50bc4f53ab99020aa459692321f54aae0f241a08e446d51bb499c2f887ba5920b7c59b8ff57a74f0f940e5ec747d83e4a16faba511ae5baf82711b3f159ce8591e37d7b6c0979405fa32cb7eb721c48d7cc03887e3a2cda34ac2530ab64254dc8dd6359555db29e6b7ab0108da67e21fd6991c393dbf7c057a73efe3aad691a0a75f685dadfa984bf2352a3b64602d009c0b99c97e575fdd4c8605672f37c9c20edf044d0942928da5ea177246cbd609d71a385a39c53d9d174d8a0fdd55b8f63b12cbf5306381911a4e97b8cc7fbd8eb1db513c5cf4b20e447ee2fef11c38b1e07a06ecad3d61379ff62476e5dfbee54aee979f3df989c3c63a4dfebd46aa7545e0424105156f97e448d12f68a5b9955341615366290d07fd45381c53950d90a9ef1571264e28d24b92ddca370b6e432ec851c2870e8d18f5b7a8d70592192950cf075f367b9a2cb7981ed5abacd49e5cdb591dc69449e08672a342af32bef8e692868cf17fb1956e6b85fb51011a60a2eabbfa468d88076e35cbbf07d764345f227cbcfb99b43d8590ec84b61c467cdac88dbc85d702742b1a960f0d39647ea178dd989fb23fa1678648b7166ee9e25108c97fa37e5d7a4ab8cff8a0843cc17f30da7b271cff1d7375fb8fb4d1a72edf22de153093c88cfedee609233ea45645eb00fbaf61270edf66f179616082d58ce3e037d266793271983c48f047235eebdcef7aac5e008c1e34b7f85ed457c15c6bcf67cd1e9d5ac8995258a495b9ec26004df0a9da971ff5729749eadcaf7c06cb3e42572f4c168e0a948f2b8e34d8b9acdbab17817fd372d18e00aa3acd3b73c638708e98355a26356ac7803159ed65e16396117f550965fe529ffa7acb8a2b5980c3c718b6dadd739a10494a5a5381c02868ff19ca84f3a0b8c6a8828409054d3c67e7a36b1c9654dc5bc61770feb303745f087eacab6427dc7ca08d66089bb747a9f00014e09db4a2b154418dcd97e5d98184aac1953ca019d899c1d73c0c33da102f705bd346ba5f1dafd472f70987cc30433922f90d4ac9c2daa89c2a4a75d985f2b5d71f0ec6046362a71840616a547b42604a99eb2412738da1d91fb5c31d35e192428ef767d3f832e57d0567f07c0feb8e9cfd9f3cce46edce82dade32a7cc0a0be1466247457a38c047f9b04abc37a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'heb3259985a5d934fc6069b73073e077cc13c230a740da7b6ed4a0ba34679b4710c9252dac22e295813a30dcd8d9fb7dca4965adebe1aad3c1dd31bd79f0bf9816a6c7a6bcc2781a3c53084f5c14d5b1b9c945ef7c7a6e136da5ac32128f9cb72ebccdf48e6afd8bd111feb6b4c6dbe02e01cbc0bbe3467208830213b4bf95dcd397ffd9aca4565251ee224fac2e4bf689ad8182e61c14534f081e14e6d02ef922d29ded302a1ee54e8c5156e4de90764798873eb7386996f95c6a362c7c5612535ccc9db149e195551a8550fb2404565e75f1c5e942f12633a6a13a2081d08b4d0787d80a24c141d7a67e534fe8c0aa49b25e313e5ff07239be70339725acadaabfa4269eab139ba25ae4633b1782b31824a743f99c95c29f90dc9c5bfe826c279f1cb155037d10e7dda59a6de0e60cd174804218b4eca7c39d13baade63846b4fd749695d459f39990b815202f1ae09233f8a831eae69ceddc17acc698d473714b7440d2f58637617373710f5c9f21de1da0b47f138556ed86e30785d12e3a2230a561aaf620ec3469b30e18dc62c74806f2d75019f9e3c1d8c89183657943520b28be8fded12a8ff7ac0d70082201f0c6af363ee9a841b281092a0d5d8b9ccdbd490f0f36b2c1b08d8e132fff47ab70a1dcbf090978f6a81dba63a35d93b636762e589b63a8dbaa2551f4b45682a2be576c575e17104460912a54b18274f5d9d06f6555a892c6a6f0562cc81170315bcf7b01311ff9b42c741928de0a78867518ef2f24bc608fce728a29619e24aaaa9bb1d66dcd2a3dafb360a33850eb67654ba7eb21bbef8e6d16b5ac58bf6237033968151c1eeb39df1ae7154cdd3758c281112e22c85b4f0040d4ccaf25cddb23debc3ae68f2087a809fa9a8114d566c64906bb37e285692ad77c19df0ca504cb1053b24d0fc56d1a3d8bbae5535cd2d35cb35dc1deb0e047dccee94e9b0900241ea6e33ef0d031078d4c7559aaf5d7f1392414adfc62ce0d4cd1c886781faf9577ea958497d6c860aa51d4cd07bfa6462a457dfb8c6ad4c26d73ff1e306b915ca45e0c22b41e3dfcd0dfac27c3d10685b615bfacbdb4e6161d132c29a632bcdf92478ee529441b0e63d400c996ff40c3d5801de574400d8dc5d6371b9e08b5e9890335bf344a71589769da6be14a42766d27bcc2b64ec558c50cca18b9d2359f1a24e6243a039cbbb3494667db0dbb7b92a4727ce9532b6e01f3215928945c9d639bac9a7f394ce3cf008a17fd49e8d99eb513e0387f0a86e2db2ff82804ba097a1ef4f3b3664f4481c5ccc1153864725fffaea20cf1a2654c276f04163afa4d7582a4cd9e9c994ce3481d4cf3564029356dc70a34cbfdca74d0a1ff85c3a06ca384a13ccb34083e0bb3c23f2dc8a7172e50f4e31c8f74324ee91abc0589370f91a87526281fb87964215ff2373e7948e731b80b5233ce54c9fbf8681cc6c001fa151e1aefb253c05697dccb101cd43edf2b2945ff3cb65207ff1c9c3c6001232beb961ac4b8670524a7929c4c07604ac03543fdc407b1117a421908377e6aa78030d3471ed23bb41750620b912649c2d69b947e573f04f044681bfced2db43296d6f420f4be128f6c84772a6f659babdaec4a4e2441bfd94c0f256d721e4a25c702fdd0bb2c8d1f0f091cbfb5004a24682dca395c0f7fa0290f0114ae83c1deacd3d2ac2cf2d0f391f06d17c96f8b766915224b6d067ea9288dccbe0e900627db35c96e2958b58d537875c5e8a9d4cee88099f42ad6341a8ba166844ed202ddb8f71562b2d395b4aecf4635b2da6163959752137006198dcb6be1621babe28191028748679bffcbad9b2da975eafa61de2e688506ce91830074d85c6341e0c37f1b187f2336e862aeaf24ab518ff8914e5c970446ba03e3fc7ba0d7cfa21afaece4cd41dc13fc7d498d1d087de632b894cf191293f9fb662391612681de5662fa215c843a8e9d490b1afd8f605ff88b0aa04239cb2aa27c111cd0a1af9575e4d654aee67e934e63e10c0b2653a6fc247760fe108de18accb7efd9932652fca37aca2d2656030876ae44709b2b467b2f607744dcae0d4e122d62c840c44430cd503526f99edec0e5d0b738bf5b4d05de12cf8aca3f6d10abcecf051c4191e756c269d86e90e5b4446cec169a4b138a98423213b2e08a24f16834c3e9ba24e9f98b8f11ea4ae46d3aeb1e6fdada6ff914096f6d58c156ad83cf241aed852b75eb9842505293e7fea90620658df881f238c7b345e078368a18079fd67ef720fba04e4a5875953ea56dfaeb03bf550571b415926e0402d2aabb89d49ab3b2723562836e06cc36ae8f2ce8d0dfb7220c6cb43a2d1e8765ba39c10336cb165da448dea50ee7a23fa4691a4f9baa444cb0eb7e925b2e7f91d0c2fc9ed52a38b84efc94b36d7f20bbf82cb0178eb93a31b52fef3818ecd12ebb2e3ccfc7f6017ec7866b6bed4838ecdf1025f6c8f0392dad31af55250af82cde3d6e31167f4733776ad67c53352b243566e2146d160e69b54639abfa1fcde16132724b142e100f03260b35ba27d9db732db2bf37b8905794525fa1f11ed03eac6b5b4714bf501b80400962c89b5dab3c86a4e018d216b50d926ebcd88d5fd597c387667191fa4ab0e9f28375cfc9cc3b29c04a5392891c068668b786f61fc74e503fbad75b2c545bcbee8ba40a3f4205230627e66a9f83aaa78ca0b637c4e953d29cf8746ff17b277f8804544ee9303c85a44a6901e960a04896c0a6c6d9c2205dd9b53ef8a85f4d39a76f73092b3b9e3f5648366ee855bf7cc736c76e449b799ab50685aee12501a8dd305c530e16e18d1a66ca7b7048bf7e2b2d964d1d2c88317f1436b2f6086915f434b3db0dba029317542ea2d0523649435e6862e85283d02d053ce2c368f11c510ab5c0beb8e65d81ef5793afa151ee8b35554169c171c7fab52c588ef7c3c71ef7a5373597ef5c91fa14893adb1e1736f55ab259b5b9248006fdcfbdb30c3f052f0198d7141fe64f3a1d468f99104b18658bfdcf4ac5f5df814bbde6e20fc2b98e8a09c06cdd37b4de2380902a894c36e15c8a5d8196d0c748525b4ee7a9830138e54256a8e2852b95c9225d04b7019fd631062394b16efb40f69c775f7ae431ab0e65fb46ad1d1525635c302a676d7cdcc362a73583c99475798e52a2e023f8cfecc8c5ec9404bee6c887b54a74d6742ee81188536761fc13bdeee84de6aa0d9e38ff62eab10dd016f3803520b29be12d2e9c3e3ced84a49a1a5b019cfb2b47c53a75d5b45b2642f9b74c2168dd59f2350d5edd4a3fac629bc69e60500b4d80b289416a35cd97f357acbd0cef899f45e49ab6d389ecea37a44269f516fabc124a1409dcbe5575ae95db465d8955bc45f94b2cfa6939f187ff8cd5ae6e1c76fd1521e7dc60e221349ee5f8f5915a076825eaf8b326af27c30cc256002d59674a594e323b7e090a1ea67475abc9fabbf3e578279788b03a0f4ce4b9ff13b7cedb4bae928b437e48aec13bfdf5dc3344ad062516753bfdef83808e673b4dd5d1a2da4b929f6cdfbe9c5ad16b43d62b2cec6d397352dd8ce72cd309c095e726ff423c1045c1ec4dbfae137c8d22633c2dcccbd144131f6f142ab18354c72d5929dcb7cff9cb8d5d22ae39530cf5357a3fdaf3899ca8ca6b0bea40961ee8feeb573f73eed2c0078bf2ac308067487f68f030fe35a910d0698c1535e524a698eddc7692f1b925f6667b63b5977cdd142e7b7508bf3d4ef76e5b40aa6d0e3546c79e026abcd49b2b8c918918d872ae71f046af99b017851c9ab2bbf025851753e126cbe19d46cec1e5b42fd6bb260f51ef5070080a00e99dac7d81b1eda49ea4f08290ad2d98130b9ca65ce6a1b4fe6bc50c773703872980aaedbc76dfcebdf79d2fa27485c7176a25fb046fa8836b00d111e144c7934ef81862bbb6a496a13ae4abb9f41ca8eeb76455cf57f537838fb6824a2bf2d0ac94311995fc88eba3b38bd8ada54d6258dbe0dc3a41cf923b996fc882afda68630a8c7b0f4b85dc1121488cfea50cd3a95624a2e1b57c77cc8e81a15a9ddf4b3f561e29331a3c3bae4a9ac140000d4560bbc9c9eb016dfdf2f0ef15aeac2d2f35665cc9fe9b8a362193192330b7976a43f96dce5444c219f160da4abed6c76171c06e0f5b8e5d5c097ee7a3f2e5af38ce5bf4c9739db157739be388e05556dfc8abf5f6f1803660a5142c9935bc7cec425305dc527a0184ee048aae942814e4ded4c02715c9ecef8d10e26144624f11965facb60c83da78d0f26295e60f14254bd33494a514e5497c6f85a11674ae285d62fb3447d817968b31c7a44ad9e58b9fcc0ff76a839c3144693333e8b1425c7d4c99423b29aee91604305a8378f464c34dbfd38722d67e7ce863b910262d5f3d9eb57ed97ab50bb0074d5ddd139201e92bb16de5eee9d77b8dbb08d83285164ec0b8f898599fe82ac53b85d66d00780a0140192fc4c66ddc42b77884fed3cceaba8883a93b223a5030b484121083f8e2712f8247551fed510e2023a51310c81f513d5dd10efa5d798aa8af887dceb4ec2f4e7760c8897a8d19a34c737cfb57f6906fed69f66326d6eba631cae0ce1628ffeb34d4258051be18ca827690ef926138ef8b49a4c2b1fa1b90f2e21a79a051e348e9bf4eacb6db907505d8a817be0dd9fe5b1cf49c528faa86060c5e0ae38364e771a35563e0b05e7a8b4a7ec78ca8f3b79412b2a350f73f693e79c37a3fff0335646fda1155da2276f0c8268b5d92062f5e7350ba928993eb4feb09e33629ab4fe3a2f66ce33e95e9c7dc0230abd550ae75923d858907cd2e8509b2df19d2042530fd48fcd0b6efea8fd2c505805ba9e1c5b08286d197448d0a0541e0fe86b8e75b164c67111acbd2aab30e2609969fe56cb26ae8a8659ae51c9f2e987435d0233037609f7a3a59172b3c90e6d6303285e8d405c152996ceb9a3f5ba854bfaf6054aa681f3a9abd7a56390a9dd6246a70dbd380887b823551659ad2b7a26b1d36bfd07a555a0ea5dcf2c73c74bca5053216f4ff7a36efc94dfe86fbf900f46026be7261f21a33992561eb9dee2b8e0a0c00a06641956c97ca799ae32717dc4ac9f57888df4a57c5c5f9d56e6ef62afb86e7f2572c5b02fbbcdbc1e955b2cb4b687849151128e9571df96af06d7afe4071d9a99b8c5a8d1c6ebb90230b4d1e2b9defbeb0942e8e5ef2077d74d274bfe062c82c5d035110e9ca5cc816d261792b9aa07d43a2f2cdf4d0d9e6b7c7230b3f56f33adf88414f21b0d3b0154c15f1e223306407ba4426f13647c48b600dff58d944651aa2fe9198bee519026c7b4311fb152118c208afeef335fe4190337af0610f16977b6372c83072ecdbcf88f50d6c6b8ad1265ea29887c7ba93857e8a45cc0fb7eb7b0407ef88cd62bfca4d12ead4ea1e7a9d2088b8d96a2bf2f6d62d73df28726f329c5c552b36c0a0ea96d20592bd33a9a5a46786e4023;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3a9b4feba5d5d3ba534f65ef46fbbc94f9128c4b25bdfa10cfe4c071565f1c98e5813ff4ce019731e2b14ab9a6a2dca3e7cb09694ab4a5698fc316eb72aa4af356566aa51d5742e5e64524472b7f0a414a22247e76be8aab82e8ce7e9ddf96fd430058ce40ab13db5c54425bfc6c3ff2f789873db13e684809db2810ea3abba951e67ffeadcb4b22842265ce084b4f6ed4662509724b329006a670da698df8b2c59d7c068f6338a836357cb3529b1c1a7d0f65a88561ae6ef7e7a7a6a5644c4dd3885cd52834942b97af0a509ac70a7f75232fb39bf12b6664f62b43961ef194782e6accbac66407bf1a40cf21a2c1df8b910623aaf0b74b6123551eb095b3091ac26a36093c1fa03e38c03a8b99dc7a4da0929201f821eb9aedaaa02cc91525342ed317d027660e26e8dc44734eeabe0e747ea01a255d317188567c5591ab9e9b2126943b663b1091fff9d24d688c685b4175d7c3ab029f4858eac2a87d4903877c6c7021453647d391792aaad2f3d1d8e6b666e5f390e51495a15ac436ac87843bc812fcd9f70d3f0524ba306f07aa1c80f182022b2ab4f7de2f4a686edc9b54f0cb0113edc06809eb3af802d54f13e91312c5b3a83570f867f2b1a75b62383cd01bd8406cbc0c62ef88cb8eadddafc606d14bcdd797b15ed0705967c258c3283ced8363f01dd3a9da96e624378fae6f8001c0ee467a56701c02a4f40149094d936d2c789dbab60ad1595c6bfd0f2f67ee42e96397b6f57b69f08d039fb461de129b9c5807c959e27bf9477e7decb62c13248c3258d556d5d7b5ea65ba27ff18728528c8a8c6836bb5c046d8ef5fb86823a79aba55c6137599763ab56b9b669d9dd2adcc1847395fed0e61aab6c75969090e2528acb2365a98e70dfca5ba22db8130f775d31c24602beb706cde110928d898b86c62ea03bc4743df1cd5b0b97b5a8e9c31b1773149baf431626ca8bece990e71805c8cf58108baa6b95d48f03dc5757678f7bf771c7130d59942089bd17928f68119df939ab4cc9872506239752ea8794b417550a28339e10a879c6baffeca690f1173368c67a7f9790c387ddd395933ac9e5a887a03db9d71fb3701d9dce34627000a2142cc008fe7c65e93a4b1debb7d21671175ba1d56ca4ca58d94e82bdc3cb92bf97bfa3cfeda8b30542f465908335607e19d3dc44d65a716b736d668f03ee826df984a1c1b26149681fa595f9e68f308429b96476574be1d3a035b48c8f270a217c118c28e4e47a606075ea9fe27f7d782390de3370fed50855244358f4af4ad73d24d10b6d4325eb610e814494ebe023c7ea7bd2e6a37cf83aebe7d6ed229e5b69fe07a235b30be8351f28a3428c60ca326990836cb0017c695ce1343490e9e68505368bd5aa539f4beba090961e2a5f8392da8a9c4997a0b59d5a9412ac3cc06d7b94c63fea3269e9865eec293e073e5248d784518b110bc1b4a159728d2616a906ff1acf1597e8f60cd3e5227425eb1d28b9c2a0645efc043d4b4865e8247e1a9fe8e561be2f701e49facbb327a6468f7faa86450d3509ea948502eff3433166c06f81ef1e9a7f4faf3889188d764c1d173fe8e88e320a58361eb3cd92c9db7d71ceac360268c81f46992b8f879ee724dd5d0925cf454444a3da153844b6ee90440f27cc46fd86d29a01559b2e03c0ce7588b1ee2082b59b68392355655ea98ff9842c929067984ce1902054a249171928d887a43fdbd2c4a9f0eceb9b7e8b7c130b9d605a6994a644732b8a4b77fb5b3ead4d13c1e8025335452ba2056c757d9051fb2f7542718c60db29d36e10b222c86ba782604b7c6db0509f78b499df83594cb3d542ed6c59742ca1c1c39d4c6e77d0acb46bacfbc04d5bd3a78e10b0cf67a0aac2eabf8ec6eb3b9459b3ea9235434cff22203dd11f9ffd1d4d59e76bad805da372e523d5c8b12a20d69760b4f6ca2f7f748d5b0e0557beeb97b9127274cd2e900c45a15da8abf8dac6e739a52013d1390b4a48c429e78bce46608cbe906b9ab2e2eb722df1830e997ff19165bfe9bf4f9306e163fc882fca71c3f5edd7ebacf0e0459bd0836bf81c87eec0c302f1acd7ed0046418e99caf774e78eccd7f1cbc62951ea581eb5d9e681fb899bf45fb476f87c921fdcf9570b794688a3e4d806bf41bc3f44435b74f8245b4214d588a0a634d21444b9cf6db89d265554dbd25bb1dcee1c720d66c4c7445621bbb008b5974cabd715ba68eba1fcc3c4846bbd70b451e423aecaec32561c1d897d44ecb4bc897fd5ac9cdc84cdaf007972245a6092e7a2f7524444f442dd8c7203066bf3418f82931a5a94a2d4c20b6a35169be128cbeeba0df6a0ea4b1cef96a9cb8e85d7fad7e52b9c0f0daf1a95c3952615c36400d19a514904f7eba4c21a8169724cedd3c1c30809bd5a0356dc03c2a395b946116b8c01fd19b4ffde01e724955d09b7603544394c56e3abf5f97c48126f43b41416e91687eaf9720be4d986b1ab6bf27ef5af992d04e2ccb931420cb83d27e4b0ecdd84f18c1f262bb58d933fddc83d55e80f3dc56e7bb6232dc4e18fef6227d8acd9def68b618acf3660277a0990f3d5e0722412a7228a29a7f157e28eab367df83f27a2887d560efe941def5e0b65dfc6199c1a2e794cac49ec649c9588b1021e062f5d30c5c4fc4e3eaff4b4a158b9df359250decb46b8289f7013874e6f8d1ce1cc680262b871c344a8f59d8e76b0ed592dea86b617c598b85a52790f3f4537a9efd65b410bde386a9ced71cca0851810e22830da7422203ff1afc48f56d36a5c32c553ea59977f793c5f5a406cbecda1bff0642e1910f09f586e4be06a36cfd24772358dfb5da65c93fb00fec2965386786db877ec77e89a48445fdc03cab38eafd1549bb7f3c88e506b1f29d39a4fe921052baec6bb8e759c3c63feba4935e1747d65337a4ac0ccc66dbaf3b1c1a6946d6561e5f62503faba10b21efc3a35fba77a07517520d0ca842aa9f30317fc771fdc3d804e7f3e8dc6b74726a6b8c03327e15558c802f6600a6cb71d99c0aa11bf49e62590b32266b1a2808576239bf03a8420e57b9ec0e5fc1f0407518610deb1ba549c983bfb0745ce5977f868b2c61dc91dbdc2a3443c4aeecea7288bd90dd489c7596088877148415a97243fae159b8517bf0693bd6b499d804094cbd5d54b2218695c19c4be17d3a456bcab2cd448a2f9116e01ba18f20dc4eda6e1174d1ed19814d5743cfe5d17504f17ee4e3a21e0e5351fb8bd6bc6bc160a278fd62f9a2fe00b1d7322db2ffec3a9f36d6ee7fb05eea9bafd1821ed6cbd196e6f6723fd5e91ad5460a2cace986208338c38978f4ce50b5a7dca0ebf000059883ab2bb0317958e87905368f9c3f0a227402f377fe4fa288548a316a7d1bbc3322a0fee75f3a2ff75f77d408e2257ff10fd14fce136845ab25da3933f1c9c4061ff499eba14ec03038e547cb1556d2bd15225a965c1abffcdb0cad39f30fb63d0b2bce443a8e4473b428e2f0a33930bbb6bf99db93f2f3da9f753172a8e254c219c481b34aedc7f569695b45e1bf6a9358607325285cf8e0cd236a849b1ce5861884e7c091f447851afbf6506e195983d70109e5bceab53ebee5bc0007adfe6011bbd03623af1c089254e39022594b33106fa0be2f00ae5bb2b08490c2ee7dcac5b20e61421fffc6c6c87b507ae0687a0ae248513d9ea250823588ca5223301149f5b2d17f6c698b4eceee6d9f1c804a1325361c3eebd9c7719f37fda1757f5575e5993dc31255f85396c7e9e350437f8da1a90b4387c3b34458f153efe2a0951967c2d988f7b779830028639f15b91affd757e0f3f7fa0ec868a9e241505d69620136c8414465c72127086aa5ef5ac9c1af616cb4c852be619c39ec1150019cf37845249b06d4dcfdca8120fe91d926c8873c9ad3846f683fc1d81611b0581b81225b8e7569d67503344b7c5f710df8971a03569e0e92f0e40742c4bf68b89fff8caff563bf33a7e6f2404b9a4d0af5befcfed0b76f3941ae02c38da81b9d75cb8290e4934e0e450cea491ed9f631543912f4718a3ba60ae0bebab51fa6d8b877a5742b04683200fb98f83646e5f421c7cd5a9808704c752b2dc5810e302e6da230f3f8b2ce62d5eccde2f571b11f9f65569c0dcfb26a1363ffc8d23a9ea5525f6defb57fc232f1177af6884358e9a5e202ed309b30d85ab56cb6a198e36cd274a17bde14a42057934547c68b051e1ceb024e7ec6ffc748b5df9644f042bd3e8ea175cf0f7b77f559c9eb776fc847f731c03607e795233e6407e0d9fdacd506b5ab20fc761fefec2767372f64c9fd6b2d64611642646380f826e2bac943a5a6a5410e3aeb643f5b6e8fab407103dd692c80bae9b7f8e2b963c396840bd29e1d744e338d2aec453cf53160e7dc50b60faabf009de8212f138399c3a92c375a38906e44c53cb6faafc43f05090973d71b411fc11a8c2dcfbbb1125b2c3b88447b2821cf41b7193a92ba1c215c16fd6378f19e43ff603a9e327023f7db294d17954ea1fd26e389131c133374a727bd77f0fbabe34643ac7870a37fc7d20a951cc306802bedffa93b774f7c9c0531565244e3f4a36a0dc3cf64b61310d36626566bc4ffcf59267592e7f495b951abe48353cc300b8c22fd01db72938208248da690ba61d43ec8e4ebacb1b601d48e5140962aa0dff01486d79306bec14eeeba77154bec178168ee06f14e6f8b71819a8982ada98c47693b38b982702e5d179d35538bc6d897e0d239dbae9cafe7e30801c2f8599f3c5f9000654891fe43daae2c0cf707a21cfe396fbf44fcd80120e6d2817793685cbcff74710672e35c744fbb7bda1c02992495d4c08fe05f6ffad48e1976e496590723447f819ac2525fb8b5562c7233ffe53754848880ec67752aae5a22b22b04e43a0c8b228be801f93600e1820bf32c7f5c93b55441a0f3f70849794453877413236ba8be760a9a52b37775dd05c4322f57f25ae00e9a1217f6fd551231d9b4233d782d8ddc469b355897176a84d00659b89bfc087b05b871b5a4014d672fa261ed543a29133f7a6052a8c0e60c6eb9f2c8c53d41d9b9558e7b9c092e30f09f64eba6f54dafc43898ed94254b74c73a8c8d0e59e1e34c72122ff76a74be016c89f0dd27f7929dd59d096201efb12c07c0a9eafa6d26a7cb29bdc28461904a63e811cb0242ec3f20d0af270669614cf33947f4b06ad894d3ebc16752ecd891e1a825f66c3de3c2e86034a87b71e6feb091b41e3898f87d5ad5435c1511ebdb4d8eb7e395fd7936faaf3f7fe9da647d755ce8ad525a2f75432d124f818bf7c5fcefc45c55132491b57770a02e73f75107853e95905ac90fac9cd93239260107b892a483d6895c3b76076a7e90fa85407f5da8974b2392f40793852251ccb7c197696d9b14edc94df8e1cd04fbc65fc4e94767d6fdc662c54adf5c1ef2ffea4469e2983e33c4c7b11805154f1194c3d0b0f7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h836beb7ac899a1f9d5ae0606d34a852a72fe6d0ffae9b8b74df52842d2f4803d8111ce352facc51c06938a044571b197e0696b7ef54c1606f855943069a197c9d9677615bf44f5192c47b790519d4fe51323cc0c02d715f1edc77203e6c49f8c743ec6671f673651412d51402df5bfddf5707f4b0113fc398196a365415ddcecce58f19e272e79ab6530a635edd275475c823a8d86e1551241649fbb6b1e3b6158f6b483d09e114a39fbb79659fcbf15e273bc09f67bdc3c45e8d61c905f2fb03197fb024bd1f227bb84875004f792be0b02721da3373b6cdb0978552697cfcbd6dd1ff25eacbb8888d650ef1f37d358357fa70f5a066d2902d19a01fb79a6124e15ab61843176437cbacce7a5ba6d126f3df8ee632674f6454eb4f4c70ebc3e1f16a9fbd812d0db5bd76189f1b90ae4334ba267440285ead3b5380017867617ca3848e3b12c01633180df59e64a778775f48c4dc3232eb74caf1dbf9a94a9771e70bff1fd6ec6da113d3b725bcae524518bd4c711a16cdf34d47824395a89fbacb99527ae7a535f3fce7c190def5b64c1cb5f3cf34a2fe4045ef0670259b874d4480bf2123c3f6bb1ecb79b202a68b8724fd05d71cc13ca2d2e60682795f0e613be381c39cc4da799a2b144c4212be6a017afcf1c6c33d9e7cd21999bc3220fddeee7d30c4be836a578a8dc2a1887129bb2ba41c1eef0b750b54800e4035bd2a0d9d5a2b24a10d54f8dc2f2693d931ca53dc056209920dacd6f1ddef3be756a736eca2d3765855c1e451e0f3263ca2c481ba107287b144c014ea8c1c9df9a0305e57834c55759f98d3d9afbe1e22aeb8ddcb3249df6fda73a50acb20d7b659c3720592fd32ae9b904c55312ff5950a14a0edbae922a4a5b8922eb981b1aebd9a739deabf2e16654ed3ac88cd45ac8ae04ca23e874f2c4e3c791ddb759af2cdd8deeb1a6d36fc97622df777749a2c12bed898e14bfd6c76e432e311f7853a6d73c689efb668f8b6a75550ea74471e0dcac650e59ebaacc5510fdcbf59262c053608a4658fdb1d4f6dae41b4ce13c58d47e9c8b57e41477daa5a42a68198edd30667d61e1ab0da0a748360c9427e13be93c865df0262819218c97a16813fcf1e2eba896ba77d570af464fabf4e48fc988bb455e32e2ebab6cd50729f7cbc570fc76cfe13155d5dde3f0608e1752cc3029c44efd95f6b8eb29e6bbb6f54b700156591d7657036047893d225f7e61e72038fd1660e3053f9501b810d4468ef6abb08cf4a5017ece73621df3565cb88cdd246d9c35c6576c91f7b66ac17cb600f2733d21250653e76d9f44ec9e9c246c0f4ca5ba1f66edc21cb2d9c27d25e440f721eefffec0f367aefdd012f1ff23a9442336cb48ee9658d242e5cfc7de0a3847ecaa9d4ae2bf3f1781c71743a7c7f80be2956014c8fb10978fbcc636f0b346e2967a815017faac27348d11d7b65ade708ddcf17bab8c435e6c3097c7eeb04a7e7cd430327250b3c2b957ba6e70b5905286b5675163a0a7558dc912fac5b635e706958215248a1b44d6e456edf47e9980f295ff66440dd97ca3e508fe132ec80e08054067ebfae0e1a551976dd25d6f9aa65db22fa4a0acc3ebdd6389f8e332099642b90df80ac9388b69c89a722caabbb17c6bdf7bc5dbdc2bc973ab3bf715cef4bba96cbf08c6fdcd99a7877972d7374c2a84e9041475e4d29117d8337f7b4379ff28834466632e39f665f46ed41e0cfc0b394c880468e61ae2e470986c788bfa1eb26a6ed03e63b309cc65e75ed857223a9b06bb186f9d6034c760553610a968d2ac1f56d9e45918743eedd0e8c059bf70762ac3ba9440b5c66d92b22f5d4ddc8490d788118bd29491e3341b06b58ee9a39f0b58f1bcbef051dd2aeeb7643d95cba54155ef9b909aa8a1acfa91eeade68e1640e2f6140a2c4189b459be5ea097dd3f33e2f32bc9126a6d8ca607b66ee961ec87deb3c9fa495d23f631fba211106d71e5620f8f58cd2dbc90eedab5f3e7a5e0d9e559c5ffea7be5f5ee58e05e98acaad9ad1cb7278b42c4491231e5a084a49e190f01308bd8bb53d6926976d4bf6c663395a25edcd7ea87160fb833dec25570a763c914226042d59c32a714e0cf91e9438f5c22868e3e84e30f75c2e83e07497233ff2584d5d10bdbcfb5d0450ad2db62846399cc8dbaf8c88b5eb2fe3fc79c99bbf88ead70548e7b3f5d1090ff75446b675fc325d87266fa7c2aa6e9d837a77280df4995edcf05e68bfffc0c19461ae3c6d838df26ffdde779a03ca9d73eb02c16c148423f6ddc698200fdf3821688b94d5e841da73d257de86717c0cb422e4d71e9b5c69a7544fb626ed21b062a72b90aa5b398a17c604fc6ed3bc833ad62aeb5e2413cb0ca7c1d5820d6eefc2eb73761f5aab39b99418ef944bf0a72907fab3c1d318dcd7da28fcdf8e031b79f523cc4e7b76e4f9695b408342493d82f697541d17b17a50c83cf3de6df0b6b06823369910bc6a72fac6dfa2cc50422cd1e6a97694ff854779ab5e9df3d51ffa249abb3c6b26b13e34a17df8fac488fb0d80a1116400406b794f1d58692141d4dfa2570d0d21853434efb913f33fd8bbe29bcfbbc7e227dd41888cacd68d7fd10f356ff9a8e3b3cffdac56df990ed5d9d64b3ba554329fde6e48343411775f98a4018a613b7ff35f97ab30d8ec511ca0f4aa7b4cd8bd0b3d743fddcceb5bade7a85cd35b8ab6dab9157d70c0686f6fe97e1ba29765648270e1ceddc4fd89164bc4f2c77970a7882266cd92d1d1f528b204c21d962d1b2d851526fe1ebdcef1df174fc99de0a92b7640b6e471ccc3429e478aca2e01fd0674990e7a5d4f2e07d024e0693d80527e205505f43974a91ac9dcf17baa21c4efe80387014434f3d98ffd2224ed50fd51139796cee078afa2b9d79c13a0e2632df06609b878b095af6bd6e0bd6cd17cdf315e1f58e1f369d52769ea1fb5b173a2adbc0846eb5d4fc104f7714d086fa69ed9cc8887a06a27c8664325dd29dff2a20d3316fd250292bbc177ab0302e7e20541d14792b7627fc1ffb3bb7ab4856aaac3f87a42f8fdd7ec8512f2dff7e8f9059b74eec4b85bc67144a22cb9eac4d5ace48cda6557b820e6b6ba9e4c21e33ad9e9c93af7ae6f382433ee2041d700b414270a7477dd8229a4868ff00fcee5e9cb8bb3249cb3ffddc63d07bf4d9ced84e67ca44d7231ba5c20d3f0317e805ecfc5c9f4bef243cd249aa51c0723cdaaced0fc8e9200a7610ad58d968ffc10578e4883e1bccd956dccb5e9410e03fe0530e1b8699b5da781af75f3faed67ee18fa07723ec9e433b68b55e4a99fd0cc45a21715931451a5aa3d8cd5d7656ec7aee9565527914a44dac15c5331c5d4867fcc6e3e2cdc2ff3d902e702f23a3a8c9994e2f39e51acb2b05c35ad0a368d3ad90da2c440332c4166ffac994566213c103abced9362f52e6bca9378d230c9dbbd01180fc5d41054d942a09cd54452eca42827c212f5e48540b962ba431b27a31849a7859797f346f3c4900587116e0fd86f3f0551ab57a48bcee3b6a37810b56a848997125aa95e099ca6aa734c020d0326d5a77ee33d4f787d6ca911dd213e884cb23dd28fd7f77ff66676a4bb5ba9f59036fabb8a822d6618cd42a70611f9d7b9eb4bb7d5d614bfda09619e57ddbfd4bafd2e5938227848e0a908eacef2ccbeb1cc4ea83e021867b5b7be5af50173b370b46fd64af3b6436a58b746549a2d37c75316bf3f51e62d5fa0d97c727cdbe468c9bae3283db8321c5669756078b1d2214b6f4b2a2b37dbe7c097886d263f3aff0231da87cce18956c7978238d2f9bdd8f62fae91808f50dca3331f74eab655c527064af1f523e62501edd44002c50fabe35d099ae2c2f0783ade9af3e378741af6a0fbe41ca82b7731fbb741809668e76941aea36e1fba215f44266606d266474ec83b62e062ba49fde526424d0f1276143be80b9b15bb96050d2149859198fb4022fff54847d58cc7fa26995f3847ebb4f0374f1c395adad18d0d74f0d11246d57a4fac5490e79611f0214cc114cd7344707ae9d8ef6f504b1f5355960d75997b00090a7dabf6bdfc20c8f52176dccd67fa3321b5cd03c94549d98cc515d89bd8f1124139e74512610a9d1306dc11208e90c2bce3a1fdb072ac6a120ddd13a17d63db523c77a3ba609f0afd4e6e84c30649c5fc093e82e8ec16e5d9007dcba20dd63dea82db2c19b9ba318a7227f55f14161dd3950ad01e36ee05f7b22f1fec76b87d0a5fd5cf00edcceb97c58ccd1ef61dba63424714f00d738ec357280426d174da1ff1ed23cacc8f4e7e917b32647ec0d5cb371f2984fb33a9da88107142075f76b11f2a11c4374ca3280403e84c8e16c1404ce85de2836c6e1fe1d32c806df151c9da092f8d68a37e77cad610b7ba6ecca0766a700e62cbd2c19b9852f927a750ef9995911bd8623725d9cc5d81593ab0541e6be5b075c81668643e2e7f8c6ca86b7b3e1ffa5dec0b13d085e317ef543a019f3ced3c9d56edd8a516c63a035949b924c494ea53bd444f1b1d7eb76e36a623f5f202f766262ac77f9d6b1952968a9bf7a9d3c2e59e6650a8afd0392d8634106ca7d1f8ac0adb15eec6f6217aa093cebe300997016f32fe416bb85ec8a6cd9734d0387e77aadb9169ce179d8819c64ed841c7291c41fd6b76a6b209ce06aa11de86dd36f408b91c7fe1367d7b0be9a9e3a7149ba67e3f8d971280a6bffd402c5b78e567e1224df56265d2bc228b2b54631ba83ac9f31d1aab955b92d94df5d79d7a87ecb3df57e5ab367340a205b7198a1c4501fa5820f66c7c5a1b16ad6df0e47d84e6c933098281b51e550f379577263eadcd7fa2971024df3c25b646c0ed8d6b03f21907490532bb4d18d197e6d407c096fc009dd274e0c0624fae2aab268dd73fe8283d9b326bd08bb124810b0931faf5939103323c16539cafaf2fa185eba0b239918fcd179a871ef1efbe5e2ab2843706ec57a87990353b132fac8b68c0f66ab6d5c1155216ab2721eea8ab59a107a479d313e3476dfc0445bf8fff0ed73352532672dab04b2b7d1366461b2dcc734e638de26deab9c24fa75c8635be59fbcd5cb3e259c65dc3b5cfbca288eb1fe83db6be32b60ff3fc3291c3dce887ef7a02a9d27f35e3efff0486f2c1b03b05ab2758d3732dc2c850e9bfe96c0cd172f31961463b61769d602eb60c5804a924e4c77d50f7f9473f3dad89c6e5f999bb93bb24ebf54bb6b42152d241b8159e78f6ce76bcadf3a7893d8ad786d2ba35d7d7a2f56a24d74947d5fad00b168919690577dfe881b986beaffff6042ae88914ac15669d8509ce8da10026796d774909ddbabc8d215c07e13d3729daa05ae2f530a004b2682054927a64610d7d4d6ee06fde15b070d3c086589b2c09247463447423613de527ef8681801738770090ccea37607c8bb7d134f13d6ae4c242c7466a7181e219630f1b7c41ab3b5057da824ef509c26;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc422d621c7261d6d0ee7c693209c62d1ce0e7ed67a983dec4336b9f5695f9708d05945af60d84e7e09393da86adc4c6496e48d30a5b795ea0acc7e0d7f3905f319e938cff2fb7298194f0e5cc5360bf5e176cfe04cdb53e6879b50dfdc25914a20130ab7f25836f4b952b1b9896a37396750ab16e4162f36a111510828a2f2ca30164eaa1e4d789e62f088f1488bdf7ee34d8173edac87b4a86e131500284707cd28410845ab12f05a6a19602dcb4683db15618642725fef28e8e7da8c98dc58ff7deaad269723f7c57a8ccf9d8bd3ec9e6bdc6c5ca21d48c5fb9a244b16a4e2778302f428b07704995820a485cb44450edff3167d9831dcdf10679f751d057684fc628d74f0a71010fd11f7293901c879047bdac6e7ebc9a02d08fc79a227b03a6a5f1a3f1a6d93989d5357e81e715a4e3d121f83e5e4ce41c762f678967db82a8855780bc69780a4f1d73172459bcbc27e4171640664d0e7379a6b046667fb655c77e54e34c948138780c1e77cb103c5f4b89765bb193ca6219c0215a1a00c1c61452ec71bffc4d6247f588c0333871f7661aa42eeb22b443bc8e4562eacdb058e029618b47633a23191ea8449e2f979f1f7882db80ddcb9bfd6e607517cf4e863ecd135325dc11a7eed2cbbd28c4c32453b2e17968b13ca1f79f662c65aeb422b0880cd90941e521d51c1e7fd66698556e4aacc468ef3e93bab0763c607afd2bc94ae39d1d99423d480b63464268fc4f94e77e8ff18c0d9c9b785237578e0ac53756b3eb8572c5449b81152fa5ca48f3e596c4aa0cac5b036c3e8281df4e3caa5fa9378bc8db43feb651d78501479e27485f0c8719ae3d428c584eec889d38526506a0bdbd84c33bea63c25008d4f22f97b5badb19f816e94bfd04a8338acbfaeab39fd73dc392023e639d6a00316196ae4a7410c4976a1d43ae48e683aa65b32edbcdc65793837315376f8bda1d767aeb28d3b41b9ff4e204fea115383d6457e0b41d8999d66527409007f8c0e9c921bd3585572edf0a3e9c885fe12a775f1013c34165145a8be77edfcd5f2f318df634196aad6f0786d97f1cb7d4153ec4b964a8da3bec4a23dab6f729526f0961edfe31aae06291660588b0ed886f8b16c682528314927c5b327f24b0d26423551d796dda959f698de2da978c786795ac81e3164d4530a32363f1e332ee32f7d61a83ad20928eeb7412a9aecdbceeb0d3b81513bfbffc044c77c34125eb839abb4ca844536a45b9dfac5b4c5b60d886b68d48c353d57a16476ddf626a7e5fea1ddd74fb65774590e1055412506816d1ada3f6c5c72cfda39e57d304c6142a16155e6bb82382a2e3afc50c705292f1a087563f831428a59f91847c8d9894ae938c0254f1e8d493d493a1a52ac14a9d7c2e6172f1724a0071e09c5fb81bec5b519ce475b2b55e038c95008729cbf890241ba6d30a5a235d93b26fae3a0b0584d30baf5779c41f75546309bace5d96366668e66f6de77d2cc00ac9e7a58186890574459926699203936a79bd216528155f5a10e84ef963879a8481edca8c6825db3acddf0c5c733434cb3697a512e7ff7965541611db213858a55c22c19afb49af598eaceab668c0e36f2b7c81fb7d71046fdc3f35faea0ffa7a3fd55820a4f96fb546d1e8bffb8cc5ed79d6a675106b2aa1f947621a6052ae9e640c3acef4faac295abd66b9dd3e16a53d1b153a96fe251ac8e181d7a192c7d0b96f3265a03545e488bac6eab1077580b16a4d22e6e2bff659a731607817cf779480c790363e5bfc8112c1a0a3ad25f67d190010fbb44ce98ae62f77d4d028d6130733e4fdc14200e6e12e98b813a716c7a2c7238a31660685e8c46a1c63a236ac63b89f1080425702df70cc6a6a9c98ff7557489c6e291712ce88f01661d8d9ac88919d5813fb3b5ebc8dca25b55024b10de1f32f823c455e8e72cb4ce2e3624c061205b956034c3742df6e373730c63041e52f398b7405f96b9366fee8879237916998ad1ba585afeac5d9f34b221e5599664f06ea137102132c828f5eb1605736ae838ab8c90f5c2dc5f128e0701c61ee1fc8893149105f8884687d87431e4a1dad7d10a7575a90c577cc8584179afe971ab95bc81717405ab87bc55208e4cc90dd4094e46fb99614eb8d2cfd15bfc31e07eac0ce19143722851b6f548da02b84c6effd3510d27d95c0a816bed35e144391bf970dc8e4418c0a5de5ef9b2e46e78fe1295ef8421195f03ab984e3e71f129ee6450d0d0093bed2fbc66027ce22d067b599f16ce15f14a02b26700ae5c3f2953957d13b46a9a3dac82d81fb9f18e38ff2389ef66ef282732e49ce0ccf66af2cf30acda786e3d50c116f3208f6e96302af78f8bbcc7f792b6c5d8c6fd20891090e1620047c01f8b55e247146497f90ff37546618b5f8afca9048bf4ee2043b2e600ef9d72ef497763bbfdfe78d9c298f652ae9ca111a6325a5004a04ab7f1d209788b10df85b79345050744affb355fedbeeea9a35973de962d2b7f20ed2a468910e140079b0e14a14d654ed47da2163f95db68c408e90af37bc78bc62e9161545b37e4a63586b655e554de06be03c19372ad2db0a4db5adf07cf204a1472b13845dcea9fc9703768ab5e5aa0ec7342aad06b6064f24daa674119658ad4c3a9bbdea73e26644b60e9124cc1b49203b35460c89cf1cdcb9aad56773af08579a85056814b632fced68379fd23764cddee8b6894da9f87db6801d72002b11654e3e26b0dd113d103a63d3479d5e6e335681befc0eb7b6bbc469f6dbf216f32be6fe8115ea7342df9f7dcae17876dd42ee2df064fde49363656a664e9a938807f244b2803f224d583896bcd16b2ac8a78722b311bd0c9a7a5dd81fd930a4bd0022ede64e4ab165b3a1f219019e69f9e45e25e3f5eb38a9e56355d889ef95daa62cc4562b5221e281f3c8e5587c13a5877fae37e60882cd245bcbdb213ef1844c259e7b6a4c3a6d4d2afb9fbfdb8e593c7b8325ce184096054d30027c3f55f495b00592f6c44010e082bd83acf1711c55a5ed3dfe18946ca4a4b0de47896461f0ee6b5d586e31dd0236fc5148d9dd7207cdf3abcfa50f3675344665142ffcc7e8d4cc54d0a558312f4b69aa8606b8f9a2194041d3098c2b344734731594870bdf8b9e850787cc22d6104856c0838e491720b7c3dd6153c804c48ba96a957602a4ad67a0727dd7a6849fb3fad00d3f977366f13595ccf72109b106834a526ee197f03ee0e768f16a0705debe8927f449e1eba25c2d631587c1b74309211780823b46270282ef756a79fe6e16bb95567c12c44274604307a5ededff44b3b6ee71e8a522e9711fd6b9e8eece457bad6e774d5efc111082b380400b72a8c56c5e0fc2726575228fb82d77322087067c45ea6a05459c785a1f3d00b362b6ae0612c1c8f54e5fdb5b1fdee29c755c7c7bb27ef9fe7051b464903fe97f5025b10410bad87ae8189c3ab8f67397e68278782073aff6c6fc9c01b884301306af892d54da9a967ccb2d9dec66f345003160c0ce38d03dddf1db02f33785597b5a573272b1aea25b0257b10cf519fd601bc97a19a442f8e8f89a999fed2a66df404280b41f09e875fb1ed9cc539bbbe9e345831bfb1d910410cadfb92489efca3928c513cb4e1c2ccc6739aaa35b5734f611924fe288ff74be6908575fbddc47fe5a0b10eceacee532cc726b141bf17a55219cc6af53d9ee3bd736660a9f861cfde171c714c9d2ed0439c30ea68abf17ff6849c284455fc17046e3fb649178e7a86c380bd97fc175daae8da6be6b57aedc9573df63792abfdcd5524b84c9925ee67772ee71ee35324b3a01b62722d0ef922ddaaebd039168557479df583a09750e13560e527f88b66477d64ea1e57dced7be3aa89e24e921eda55c0f4d787d28987fe7dc17d721b06a52cda7a4cd4020f9fb32bb137524933034c6a75053f66dcf907a5aa57a808c4f6e564234d66fc239c941295130a8f5883c96a749fec2938d15edba764f4b9afcdef7550a8d1f88206aed9c844c6bae2f6d56a2134300e109e5e44adcdd2de4b0abee8eca3bfe68e0cfd84aceaff7dfb3d10483ae59411e7a2e707c9658d41b33889889424ffa60defab18f5201b00c2690e58ea8e5bb5fb38fc7e968bed8cede49f9b135119d59126cd867cac8577751afa76b5d47f0f4c72f2fcd58f223dddba71cb39c7def746297de6e1f4956dbd8f4466635d87e391239325e046e28a0b83363817eecf8025c61a2159e56f909224cf2cf98681d14c06a37b0356c02b231735fdc68a4978c8a4cc36e3dbee842a87fbc840ec7048b6760828544a15d0a076d3862fed454619306ab78b347e95e638e5ac4d8870e7ee81f82c476042218c8b8d21679cac7a8c2e382e79e719152fcdfed1827834055f38819e04794e1b4a48556d43a51a3ee6c9be2e52bb1bd2bca34de09e612b9be721f66287cc37b8ace669ab2be24f09c98fd756a311005906c229345c51aaee77139906fb5f7874a80db766913b1c9fa810efae7ca9c0d7b7e0ba68d682605ec77590b016cdf1e2276535262c2db672e5697fc4d92907cab198c49c1831b24ff8f6b6d88449586fb19ed5485ae463c607c2610cbe28601a5005da69014bc3207a977050153b07defbfeb7316ebe3c15a54c360f9188523c1336b4536fd5088daf47139e3f523161f651bdeb3cc02ab320ec9107ca043587ecffb2a6e70a1d8d3e2953dcc49f6ae775b84dde9531ac9189c81cf2c814d103abcdd8c2f55a228ca5556ea0ba1d0206acaaaa4cdda7e2ff1be742661d6a91c9f4c9dd8fa6d6a4daf58af185fbf17e739f15af7969d338de1baa4ad14724e48292d9456c64cac078398de832a522efc9c31b149479dbb2c1208a9d54afa83187dd4f2c66fb98200949a071930607abd0815a7fe3bc73c859b227bdbdd5aa8dccfc45d3e714685ad9874938b66033c0545c52e729b1117db5dd1e235ec7088ddd8139d6390514188a18d4cd1d56b807a4c2a5e389f3f8d9a5bfe60b776fc820b18e6e1bab32229f179ea7109f7532db20b4f647caefa494aebee806ee5be7482addecceae1ea20cdd86481ebd518927c3b0ad70db4a909d9f79fc13061abe4fba1f294205ade2c11dd6baa6e9ff65bef28439589c334e9cbebbbcd683a9f7aae9803c12cec3c09703d6a91c0563f53238e74f9daf864ec14538f796ee24254978de5e14279926c4a397dc432a79c5c8d1e08471ea836ea502f473e26e20b4d7be0593bd554213b14ef2d4477bfafc0ba25224ed6a26789e9fb6e787b08677f9e74ebbdabfa0b36f2262108fc4b3aa1f8b0c92bfa01f3020e4d089abc937d376acbf935eb830d22eb0f43969fb3ea165bd50e9a511c4c910694d3304dc7c37b2421d6435453a421706ff91d30638dbba4a7d3fbab8e7fafc2dc4cfa00b3927ba7d8b3f28ec618aad22d9dfa15ebe516f6c81527dd26a16c783b504ffb6821fe481396aa2fa7a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h58c2c2b5a549a9e1238cf547318f46e9f5153175e0673f8fe7df1d3471d3f29da18865865a004126db99d010bdd54265760f1f89bdb6a0b186523cf9351d78d7a0fe003bf11414248fd7d90a6ee0812abe914015fed13a7f4f351714c427aba1671714c3f24a113364557ab7627554e1a628d7192ef5b522746f7bcccf29e01f1c5a67b2296ca03cff01c06f61194c017fe140b0e8fc625ecf990e267fe9a2b870d2b4ff6602961997459b4ff6a0380b81545a1d99e84ce3caba6b7730e31e631b4edf5e552d47006fbfd6247114196838bcd334aca497fb51b35cd0a447b3569fa9f1573509e1d1f7c8eed8cd635668cec58d856d41f960e257d8acd8f9f1eaa1bc05fc628601d17999d29ee6eb1b4ffb908cb15dcbba429aa367fc645db8c8db9100b120cab0721a9dda6476d71d03a5b84f2b476073be8a736596c3d461be445f36f32f8faed0f8d1e489460a661486356b828ec66c60c86297cb10e15e32eacfc1a82ec6b67146b36424feba2d6e526bd1ebcb9fe29a93014f95c75a4ae1ddf69214695d9776b95c60f10dd016095c1a3f2c9d729ae1be98953ba4739b8acab1d1dd5c97c47f7a9155c64e60a4c17bd3ba1d01ac4c6741bac476696cbc7e6a6ff9105b6ac6debabb86bc1ec0b5569590ae734949bfc730e78169b58f444a8db482c3f5a82c4deb3b971bcf9ca523dfb6849627e2898c517b092d13a62982b889224269429db2631030442f5e74ef183feb86e6cd773c421dac20b90328a59c7b12dff725c2e5e698b97f9ab65e799fe71efde57c76b9968c129840e7f8035950c10ab8e9cee56995aff393883f199843ce372e45b79443ae7e3b8bdce897c7a2d73a3b7ea3b20367e6893431e8cf1ba6252195d048dbcdd7cc7afbb3febd8243683f34a5260bfa1dabeb0e2e9e6dec8add0350e8d44b531709b5a1d7f760fe4b319fadf61daad3581de101d9609b79789ff4f41d8be04f81d963799b58cf6fe5a811e9dcbd1e5915d6e9412cd8540f195207da230331fc2e18249fbd39efbf0d160ce3b2664d5d86c7703203e06987e4510cf8e3a1a1978df0aeb7bd0047f286be61fb2a851105d81761e8304f9e7741d15b2a584112e2b5b7faf28f6a3006aa10ef40322c662f33b924e9a8926b015d20863dc94c03b1124c0a725178be131f4dd46c8af82ec71548d0330b2c94cdedfa7bf41aba4b8776958669620c2b17e0cf3c81679ca2d870a23aa9deaa1d4b4f51c3b4fa3c93440f614b73a1fec55d5771861b36f3db13dccc47e11f41a58e8639ad72e86beaa9bc911534dadbf70b77a1e49b370e3138cab595d1181088c32d0af8d3429de16e0266886285348831b92c2277636569300dc19555ac36d103048a0231bc734a0d5e4bc04699e9eef37e0c2032fb0bc4485a78a5adc1d98e4f9435b68d572939164a3cc4f7858229d93d49209542d54e512fbf3bc358b5492e130c3487931edab648d71b8320231bdc22730ea9bb8f67dceb065ce39733988392c31a882c68260b577d9be44ee4beefa4b988d105fe08dc03a1e508a03990ef65bcfdf30ff84a76d7f0a8dcd88ad98755e1a91dece4d0712ee13fdac263c8180f57efa9187d0fbe4777c9937283f890806c8a4d964151c2b656c5d96c1d959f870c6041d0824944e5c3437686b46136b97a2b7cdf051a8c442805fdd17ad79f6b354fb93abf9f936c3ebc46a9e5dea4797c3d349a78bdd07ca706bde36eea5e7f78790b1dfece363f5d2b58b299a1eab0211357633151f5eeca2dbdef45d9a750bcc317edaf2fbd0542424918e190c33eec809edaa2747bd85b9f6619733e476ee3ecee2295268c97d74677027eed04fe364693724e536ffbe477ad5594fa302edea38dbe54890560dbf54ef8ae37de5371581e91681215d7cba87ce20101cbe1cabe18b3046780776c59b1b8b18db119a503866fd27a921aa73e63a1e987ca8868ff269b06a8d1762802e90455f5eeb713993396679810706f134dc589bc4267337cb8ac50bb816d876b0fd6ad70f7399cdbaea2f27ebf07ca43f963bcdfcebc73ae378614e3130caf2a99216cfb011c19cad0d6316b48e7395b3ea42c11921673f9a3ef23c7b7146d4c6a1e9ef6df8e118becf08a44ffa9cba528050efc97a592dda321e416f0a11656719e7fb3a4b8c2e9b2b51307117d181aeb64a9b7af582b146ddfc3aa783cfb55f22be97e1cb58efa03b98120378f2d2bea4a1df9c7a83180a5b00292e5091d7d0b3bbc1cbd00678e179c78da90fee77e0abb6b431e45ad71d5e412bcdaa3b00cfc0b4a4344c30670199ba846ac853ab2f1aa364f856ed33b6d18133bcb3baf0b2bbbfed682703af701ae6cbd3c0be9cbfdc03a97f2e222edf706ca8bdfdb14f01bc89a259d23d2568920ac8d502d292863780fb60bc283d1026257c4da22de48b43957d13d25993997bce6cc7f38ab93ecb62f1bc78d27abd31a3b9819b0ef4e23c057517830ba187a90fa8c60d87708c71cea6e5b51620f8f8ed9d64128abc0593fa6e3e16520b992ceeb612caf5ef248270458a595e613d47e556714f38340f61698d463ce6654f12d577244094d1be083e3a156298b407ca33f3d19582288b9dd8170b96d2b2b937feab28cea8aa9aa8b0f7dbb3062246da7c79f86a671cfa5c0727955d9a53f250fb583d92ab0fc850f264bb7efe6b0a9cfc71eeed0ed1a1e42a36df776c4e4b8804e87e92065ef0c8105aea4d9e22fd04e34e4d73612301619c01179dd4d48dbef43a12b285489f132e6f7b080de6e5f5f9ef061b2cb8b665aa134c57ce30a71106ffb5cdf88d1efc95e31ba14004d2e384c792c7f574f84936ae37863467e3623cde6c4906909664e572108e6390fbc3fc6a6ba0c5fbd571b56718dbf4e92287b780d768c447a3a5bd503fd36b9f9a4cdbab30ed811f3cab23d20520148865b4df5ef4fde97cec3e9b7345c2f7ac90d68d0aca51b7b7a80116c275239817b8a5fab8ccc1cccece3d6190f6fa34f9802fe3a6595dce3059f02519fd32e72a2e6739f92b5c3a728d8a79e1b434cfa9becb244825ff51b939f9bf651c85c6e374366871b27a88b3744c15714c04a4003fd99cb586e294f8ce27616f5781ec4ede22b6214a885f80c7c639f7827ad5dc082f10a17512f91c0c0be528edaeff14bde0d87cc60a28992207eb50fc7605b6501f6198856ec24703ca3183adfa5b2d61395ba69c41c85a523496bda1582c703fbd89c7274e88714ae0d4184c7d830f7716a0af4c2c0d0d858a58d4458b2c6a7a4606932daaaf58d574fb645536120da7ff3fca3018f8a04f798ef1c7c7201510c56f6318e87a411a415c9d259fdcf60b868d51a8822243b06e23091b7caea5918a7b69ee8e221137cf843ce98926056c7b615c1335eb7addb9c075e55e8a13fa6a38934f1fed1597eaac8e74d270a34709bc29bd0525da74eedce0b6b25d9bee18849df8a26b3f99fc87cc19189405422785a4d876227c7b1fd6a75aa8a40d1ed2e5af0b1dce371110dbd8d45e67c95ca7eb464c9e0420a1af8a1ce7f2c1e8634adcd468adfa1b9e45ec14311eeced01530d9c2b0e2148966f2e6fa5b6bd9fa094a116b3d137d488d4ded3c2d03ec85947a97b9bbbd0b6448d944c4067a5bf6fea978ff44456a27cd6257bb30eee95e9f3a3ed35e14d7d1ef9462530fd17014d7c351e3a61b9a5edf0825a72e09032c5902e5f0427ee491cd0891f5302ad7c4502e0f8aca410a59620e8e7d862179d40675db7a6a0286dbc2911eefa4a50058e03f8f2f9a8b95de633d6d24875b60083ec53ca78210a376a6f818d7832f1005501dd1a8ea7447fb09f02764a140ca3cf427d6cf54c764730a894310bffde0cb8ed8adbf735484be3b68dbe1e3e22c1a65a186f153449ddc801b653fca25b6e39c2468fbd63a488a97e23014d24453a9c558b9f3564112a037b3980f3721c151e6852e110643d7347c0ea16e4fc6b448a1fcd5176c5c6773f9ee54ed75f6dfa11cba3c0841d071df9c7a5e7f9ace241d3ae5e8801d98bb6124e7246437e3448f95f688406c6e3da75ebcba9f6840f6bd88d1eaa58c46983e931552d87949cb5bc0878205522d76a614d266093bd79c0215dd9fed58343d64fff10eae5e59a10548deacf99e1a0e76dfca1d04a5d358e3a0ada599ef496496ba04f3e89a23dc3b79e4d21bc42c96bbc9fad27d5b0efab6b81853a31a4b08a4d8ffc4a1916c57c87107994e0ba8ee22fc113b5e324aa40ea1dbf7c4c1ccebf1a4cea7aae2937d113c3d57fecbfb17305ba059f6ac8bfcf91b040de5695e663e1289b35e115a430176e3fbe012bab90db09f27eb41fe3f2ae1388c09dacd91c5cc3bdab1be0bf25804a5167910b7b06093e14ba6862acc3801e2df642d0eceabdcdbcc9c62c97ce3fcb2fc75e77ef2e461dfeef576caaa728be7eb8818584fef0455542dd2b805e2f007bf7d90eee11326603954eab30dc5e7ab166baa1112b2f15959b5e1340e0ce4a68fc7bd64af9a9a2d1381c83d030ef2ec78fb9f23e22ca6e783aa1d2c3bb989e5bbe6cbf63edbc987dc27c50d29407921c690caeb9b707d775fc73721f42cb05e273255fd623cfb5b939850bbd5b3abb652c51c755926ca1eca3f9a3aa2a9bb28bf6f09930696a32c8d10c0fce2bab37034266dc4db7279d6a0e8fd5d14558316ec8dcae602c588d6397f698cd3f87c435b957ac09f4beb78558f580fea2326e939ce652f41c25f24dc923e2dbfcb66fd358a097bf68dfecd60cbeab2e136f31eba6142398f66f1253cdfca6626d8c39ecae5b0a349958fd984cd21690b26cb463244a41c87a487d46885a5fc1481549190409a2755bacd424a2b97bbbceda7eccd229832f46b17557ee0e1f9ea5ea9546814f49f610db220268e69748f9682051bae4b5c15aa54a36ad542fd395c8fc695df071619e4cee39ce4854475694354d2b653a53f37bbd8bc3435239bd48686163d0fef25bebb306a919e787e1d59995ac006f3490e460e76eae007369c5fc9a6707c553421d58cdbdba40a0260570a7da1930b08c64cfd7e7b5fd7dff7f492ee13847165df743be74907f430b1c81e9b60f1b735680e6dd486146ece32a1fa58c444ba1b23c3b6cf5b383ecb676d968472d9e2d1912fdef59a1be24cebb7cf2ea236c675a74735b3c4618e5c068472011174ff5cdebb1f05d0524a904cdb4b659722b95f83cbe23d94d5f57ea7219c358cb7f421c31241d731168c2d752af71a3bb58ca131b1c145110f571794d5b37238d9366ce7d1d35aef812c9f5bf012b6e7845c248f3ad22775ceb04d57eb778e5f04ce68257786a1a50c87bb87f4d6ef09e71afeba374c0d7eb21c848e77c1398b883f400fac83dc93326db2c0e3e4d3ae64844de8337a86df1e2616b65ef820fb11e58c0c07272e71f18fde66b90ba812373aa02ac816dfbea88e37595da93afa215ff8c6e8ba4426510f9654f95f27bde9d54ee457934cc2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc5321b21119b1e501b6262317eb1a2977683b28b4557ad36fbb2df098a41c0f561fdd8d246b2924eee4729ac5c225a2fe6f77ad551d092cba427d45b034bc69d8b8f5857239b6d3a26a80ad49ca5194acef3bef658597538796fa0e7eb1d10f9220ecdbb20221d73bff9920e21f48a9c0d8fc2d293d9d70c383118fa50fcdf8f9d35553e61161703362acb916dad6eaf04a58b38a318acffef5fa1f68dee9a60c22cb56833b6f0c93276d50a63d1cc4a53c71367b1e76aa89e5b00b1c73593fc836fd3695228cf2e218d0911d46acce71db4033b0552efdd047cf3818464645d1f57514a95fd3da802a0584b52a3568e9db33ad36c0514eccf57df6a7cebe6d7bbd819f2cd5237f9249f0a93dc57a057a360170301a386022876f2f84b91bd84aafbb8a51b43a7503905488f2cc8569c6afa6e793161d0a4f8ec8c0f06ed1e79bcc7b917c8e9eda25ae0bf46d037efe22a65294987852d9d6ed1e7b3a7a280d8b3057bdbd8c01de744dba6a719828b5901409d0debb628178d8742389d0cc48e2979cc23191b077d5ce0e5f9b693d1ef318cd1ab03b622e728a04404973b1ed61d8841960b4ac6c358fde38cd309850cf972788f83d66a04b37dab2e25a6f6b70ff10eddd7ce1565ba2b1c1a47b5b4433bb0bbd7b77f8163686dab1a83d60e472d138d7395d37e2836029839321b7c86da6cd96f89e85fe61b0c2961b53d94b2eda2a037aea51f7db556c808a772456a3daa282a08c7f3c73b15e8ecede16b845b8727f996af3e2e90371ec5f6a0496ea7913c2190a86b3c8ed68010c554eaa1fc90e5c5910a4492be31d1d6422238f7db974ffe2a59020306bc5a82c67b2033029b9157191be1bc3a4bf25e8721e47b8ea376b312e6340cecd9d1a4ba83b6662a89c3519a6bdbe85a6b08defad138c23ae47faa16d6c1f0dcc6d10f3fba1869860159b996aaf560a4d8c7cb799ee7021b556a51fc8c0187f8eb7cf134dc82fce54ea932a2722153bf86db3f62fcb085688078f679d13238268baa810d0db57f993b90f4ca14bf52a4f3beceea2c3f430263541c24b74a01ef53f4305c8df4e42ec2944a4e45edc8ef0c01906e4c0d597427e939d4b7815e21cbac85f93ee100ef0ee8ff75e669fcdb6024f878aff3d360720ef58c602a5375d3c609fab5ae51f2af3f049758c6db37112c315f35b956e87d30104300272f647a12f6f8e35fccca2e14b18453471b74c4652e53bf6148f5d3a606e89d9d450e4f2a47500a268a31f824833132772ce0042d94c1badfd60e7996c018386d3aea305a47e82ece907796a07ba120431900e586fa2f8d86ad4db867faf5f839e163e4022541c18a68014e634ec09a6b2855467a08a48eebd8c1f4a52de2c66560a1ca26376136a30f3ea4bf4cbbb0b1a874029d6ebc5730be2da5d9118a40aa96340a4b29746a9a96cd42bcb5d9bdfcc59919cd69c6553dafe6f7330687867268d575beb9c08ff92d2c670d48aff32d6dfa276a13d290fba4987d26ebff07f5f06c035464d50e08010cc3c76d1f0028c602b9228972401fd9039e66d056d9feaea6f092c7808233e13125f419d4e123e0d69e12fac83673fd8d46181fc1ba2c24ab83ab4ebf6b300c82fa8a8a4d603ce41a54277d9b785753e2d0cac64b0911d711da14214ee7685ee517186eff1845e1fde0e08c4c4af9aaa64197d66e1be35ec4d12f84e63067f3ae30bc89bdbc6dfa3ba7319a91d35bdc1bc0a75756ff06c42186b19c9a45095efcf6e92d7a212c0d8fc50563d3ecf3f5dd994b31b987245b559cd5dea875bf92101ceb69f854f571fac954f0f34029d16ef1893710a9a079255afb161593787c1eb03a6ac0c76de08aba7cfe54013ef8ee1edeed0e3a70bf1937e00b63dec55de0c2b590fc4b1c5a25c316805723c97d1439042a5ececd4ccf9f23445db484735b7c95c873dd343bd26b63648c12472ab12630ea16b64b5d061d0d89ccc1875fe98c9f51673c3044c55f58f278b075d67d050afe0d7ef911c758e53ea7ca911122af5e0e1d038c901036e296a562283b2d480ec48017eaedbb50553b60d52fb849c99b5ad35f8869a4bb1cac8d4e32ecdfb39cfbddbf87c178e9d672f7023df712e01b06f4dac23e624f882d6063816ab099b914a5909e1a52ac5db373645f47ddb5e41a674f910948dac9551b8597217d8774328f9a006bbb29d6a245d968a78426c457fc06613d7a2d7334720031471fd3612ba68552292ff6fbd4391cd0a409874c89f7893a71ec887bad2386a1cec59271cb36f50559b92ec0929e8a04b578e393f9233de98ddb558ce3008a0b12ce9068753b4f26383d75871ac5d76dc744a38a1b35636b458f0a51f3f993a58f383166fd75d43931cd201bd3b42ad63c2afa3e78369fffaf715a8b21e5bd2f1f4967e64d4ec28522131b9765b490c11e69c531bdf101da0ccfe1d4511ac826e0a123b5831b08a0db21914ef698077d3af73ffa3f89345115438116ec75ee3ff4011bd9327657194fcfd5a36632e622d276ef8f1ca9568d4378cf60467d09341f521173c21e1f84fcedc227d0d8456122cd662efdb76e5edc48011833af1ffd30d1a1bccc0c139af674cab4df865064e3d841058cf51e257b53d04c9b1548f57b1a12f1bffe25afbdf6cbce0ea77e77e2f804fd79c3970c3248735fb2e2b945dfb0521f46e5e265226cfbf6d803395cec3ec675a18677e4ab90e31ba533e1e55799084d4afc6437cd619221be45e239c97d039404e055cb7e9113b715aa57e379dff0c274af214d7f1413178e6d0812af128246d3e4099d12e02b075dd21bd3ad20223a074ae69ce9c8acdcab02f19d9958e3d0375941ecc5ac9feaaedec8880c2e8e9a28ebb2f77875a16b704f3500f44545502c759603d0b3541a8f5dbd1567c1f8624bc8d72ae3f1b7cfc330a470138e9e9d51494ddae5a2476af50d406c45175348f57e29492e822e91775187c7c277c08e253a6a4625c1bc858165656c7164d00282f629dd8ac3013de9dfb0a3f4ff0e2f94d9f9f72010cd3b6eea429697131e60d62847cdf72f4e3f4eafb082efc91a1e82c0e8bcfd0380f85b23ff99bc7f92b7111db81778b434464569bd2f0e967083ed7a85274e88a5aeb8ee7fa88fd3c6bb76da087e56e7ae224e77b06797fd81623a308c567caaf096b4fff5540ff6b74fb8fba948c97549c6f4d1e9fffc499b29376a9fb831bb022c9f4804b0e410f6fecf0077a60e09a753d35d9e69645b35a3f10361b1f4b399b95d6dae906f82224c599cb1e43779a2033024906134ca81a83398867b8ce59216d6b2f6685e9128d58ffa74b7469f8a7e0bc19a1d75501ffe8d38233f4aefb6a3d0017c982789196ad731e6ba2ca9a415e1651ee479c8c7cc2eee8eb454751d2b437044db9d406605ea29280b8e915256d29c4546cc9e513119fade6b0c73cbde68ef69c167c6b96f2158ddbb1e2da4ebf40f45283199b6650ff78cca1808f03d06cbe02349c377ed11ea042f1da8551cdf0132b9f5b36a3998226c4e21dc177c6446bd755d4e1e69fcd382f21ad27e5fd3b126d40eaf33b7206968959feaf18dd8f6ca9c41c4ec3bedece44c13063941a22a1ad20b19f36f641106921fe6ac7b66eab25ebcf925d25ee825e2eabfe848498a96e7115dc91af533b3f69264e75a2c1c1232ffcb3b32e35be695d395747f63c278058d8c4a5169b65f9432e5d5e53561da054893142b06d14dbdb2ea77e09f0a5d974200b3290dc217d6daca0cbc247af2bb95b455a08ced368a8e8eac5294fcb1a55bb8db4610cf978d3126916dbb855d7e6afdc128508daacaf5e74864e0d6ff9372387d333ea60bea4210ea68390f9b8d2778e06f186abd1f283e085d1a4b3ff5ce6eefad8459bc362df678c1a774b1cec6059d8e64c9dff5f3bd253df3f190ee22adb5b5f2974b4b7ff26ca0a7d54fbb30b33ec23d10b6a7fd5024646b315755c8720f386f298f7e694b00c4e4a79aaad8491cad0dce404f87186ed8cdf2930c0d515158c64b13429258df6ea538cfae84ab6141f0aceca55247f26a700f3fddb63f22fbbb48d42d904b088555af4fbaf26244ef884fa52e00927aa68f969d942d2716b033496efe4c60835ca24d95dc16a2bd778c909554d6aee5c16461a52b41618ce907299252a9e20ab88b8afccff57ebc6bf921bd72f53ab1d7a62bef574865d78e9813121845f126ced435c4a1c639707613ba1fe8c6d83ead2db295ec6ee6be90f825d6a4d2fd2b15f609571e131780fbd4e473f87c0f098c0ca934b13aafffe74b9831e64cdf38809c00136f06ba3efbe0c52ff7ef490edf3deab3f6103146bbcca71844af17921599c256eacd21b88d380ace886b870cd3f660320a8b09282f5bfb1378b3a1367908e64a15195e62710fb100a0d0cf329507393d6e3a91eacaaa9cfd763f3e2c8aa41668d61e4ee9a91e7ca36d2c1042c86098ff14d0e3f0a644db3fed25a02b1181bcc6cb6d519ddfec3cdcdd87b81a939d12be3cb26167898a2c8dc9573432e3ca6ed4d9b6087e2b16cf5b3586ab1d5bc0cdaea16cbe5f819bcd36b76ca0293814269d485999506ef8922a6d6b71faae00c5c1cb41ba06c8c240d1dc09949beb168a4c3e1ef1ac6f12bbd59b999263ef7a36c8ac397a346dbc6ae4c24f2ed22c8334d0c8814f0f365fdf50fcb63eab53927f95420c90901ba899cca239b5f5746ff0a4ae4134c1760e2a0b28f114ec324a7fe34400f5dcdb13b235f7149246bd6b71348c6c06a748308225ff0d5242f4eb50a2b368f24026dcaeda8ff8e26aa538e80234c95cd86a976ea0f4301337511c7e1943c6c854e76d43689f3992df2d63a67229db296384cc455397874c5607e83eba7ad5f3f5d5972b7f1d845278b591ab2e36832b1d1e959888d18705e304a071d874cc98440f2e3772e62655025bc9f6d41812f43fcba2ab77b5669cb3c68ff77cbb4be7bebbb8ccb2ec4838aa85ea62445604ec20a0815dfeede05a011aac080ec76a195c1af776f0d0e6d9ba646921c1e0d079ee2fec3475ab74ad9abe4cb4657ae6208cbb3172bed45277d6ec74b8adca0f79c2d7df352c64974d27ffd9137702939209f9a5f2a5a0ba0ee1e7fa4044b3fff9683734ce06f52573e5a4731d440cbb873fb04f11784ca331aac8bea4e17d2999893e2522efd8f8ce1520117203d96eea57350ba06409aaa46fbc80cf38890454fd29b70f0b474e47b9d74df3f03234cb0a2305688b5745bf04cb42130a543d725951ddc0bb817beea5eb1ff69a5a09adcd75486775abb4c010a7315f07ede80de7d7170355813a7cdef5de389938ee012cd6e8d375f366fe500a87ebe39fad8f07669615d6da388e76aa1d0b1eee78b441db3dfbc7f06bb805f429e1d997d5ab7bfe1b26388bafdf9935303009922749830ac9bb66ae7f07429c77c4046556ca72385210a1d1c333edef796575cbaa54eee8d512958e7f745ee6be91104185;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3be981372ea1850d5605ba6218d4d88179b5483d26e5b825a888526f00010e57ddeaf8fbb03795c74ab739f14a84ef25e20161a576c3861692326bd8575f35871dd0c9658debd7b4ae283351e8557ae0cb14df448cd2bbd195fd7721eb335934b0f3bd303e63f90485b80e5718fb18a0151c2f0963123a6a47b7d6e23a3c81130f44b8f7d74bf092106f0d45e9e37e308c8a54da3b031f5b9a1d8f3525ac3f7d65b907ec693cbf07610006ecb3de1093b3ae6db0b74ed9a5620df60911465509be3bb221b80ac5a1a5db25fbdd33f1e3363239f9cfbee770a2ff82b0db533c149dc005e7f4f6f2dbb4fb0c22c9dfcdcc6f3cb8a8e526994dd999634050b6c2a414ff5e01d4506a9f01e9c4a53e2d7c39665a3319ab12147e954722b4135c8bea07268516194eafa516999ccdba98cf3adfdb478a8640de012fd92dc08e78092e012f712a093c93e01a4c51d284790299ee76c611b0779424a8113275deb053c1a606da47dcfa07ff512dd4d6538059ed4f262ba943ede6013fb2834fd1c480a6e52fa73a5089c18bf035fa5554e667129e3bfbbe83010d53420f6c97390be681f3c4cec4cd03b7e65269f02c22486150eabf23f97e15a5ebd4196223d5a30c80f0a4195f2914f57f1d5fcc4f1d07913b6b45879e8487b67dd881e80a37ffd319c93ae3d1d5d8aeff6ced91e78514e9c5767c6910f7f8f10ba5634137c9407f0eb91eb674ebacfad6cd0e4b7467eac2a4bf60bb345b1b43c8d6016c0ef27ee67243333a206434ba7c48b9f8e8550af7df17e00f69d6c4523df339cb5206c54e04dda5d5218d37920b8880529c30adb818ae63f1cefb8f5a764024ae61aebdcd9b6d355b91c613ccef31bb50e8fabc17a86e60d8283bb35d84eb6c19ade671776124a69548d1a340e87efb1800f6e499842f8554abd7f78fb8d5e37dfaa4fdb9a91028f7365f8ada5063fa7ffff5773121478ccc23fb53d08414a4a3e1679a582748fa8079bf1cfc29da26c77b717051326559488b6716f92b1d4755f5f52be2d78a7874044ac2105e38ef3ac8398dab287ab7078958c56f6ad40c071bf4e1e69d2b9311446711d73151a34c051ae593a85b42dc05796e1ddb631a0416a02a7bef7401ff96b6a40c5a864aab1da27affb5ca8c65e753dbc3420d53a377256ad5ab6324ee8ed19e9f9672032c7af72045edf5d6fb148010a050f9148dcc7275bc37966662b8cad81fbcafebeb8973a4e16f456cb55c959f35acb00b13767495aae49fc154c8b10f47a95b7bc14a29d69374a350b473aa7fd145054589218f39f3a06e3c8a5c067cd3229c19b7803d6f8a578ca534206ee0aee0598dd337150b8425d51c31d6c806ceb1829210e7b105183493be004e0c0eb18fcdc8b9f062f31a571563f817b51a9e650c90b44bd915732408d83001a24806ddb9b9ad3183f9d80fc8766525fa1d2c1a5d5ea7aa62e662c803d34945aad2f99b80f6bcb637d9edcb0a4428905e2250538dca91bf91b5455b9c8afb796f20bcc897928dc95654ff7f836c834c08f883527c5f107f792290a206c022a1ea7aec2133d880257aba82542619b6bb3406989586efa4540b1a958154e5fcd108bf3fe8c3397194ad477fc6f4d7ec9b24e892bdb035bf479bb9c9aceaa523a41b1edbca437574a3b19f15eb1eb23da8c941c60ca17ba70af2ad9b9f50c4d72b5ea8678401476a05a67040265479cc18719d63c81c56c350f01a795d97d1da0d051ce67dcf80e34414d45d512eb8a3bd7a71a723fc457b1fd788c99665b1d5a9307552362ea3b620993a7c312354b3840a5a528156421c5af4efedf4b9ba96ba3d30de978973bb48273a4999af79edc2429dc16d8e0bb45efa601369287b541a8190fcf3d66c834044b2eee03cf7df8d3acd3be19da0a58d332846fc7739bf27fb763728328ab9e9a296fb24c5789fdd15925a7be2cae27f19310d845101b17271eb9fbdb6366ce15b74d313f74952138e124b10cef381648b090f015b8a7fbb4b7940b1a88459530978533f780fac792818325fe200350bdcc777c5ce6d2c2f9e92c8dc7fc7b57167e3896ebd88adccc13249d7796719cbf39777277160bf01f99e02601b25b97e438822190f6e55af2ef0b3a31ec596fbb75fd6f841b88dcb3d43b4929f74afa82fbb905cdf5e01827d5cde688bdf19c11d19881c9fe1342b82620a503de2fd2a52a9703e8d44530c951a5b2d00601f7257e7571ee54838a99aebd5d6526cb0831c27028fd2075a9e1979f19e8674d889f9d2bfd493a069e7f49d22f798b9061640cf27356ed790b3226e2e9d9e0ccd96655dd26a0499c6f9b3b435da4ee3c59c7b5a6e7c1fc62a5a5f7bb68f8fded6d2f639865e43ad6eccc911c8028999f6278e6298124369e345ebd838782f3d6e9ae7bef30a88aae3eac3b1b8e57cd19c60e623d01f8661124bb7b2b13b6978be68624faad084adc305070b6498a4e59e61a2f2d3d7c4f9f5b7d7756927ba3af20dd0467eee728726c85615195152ce63b3bfa4120326e93bb658be3761fad44ee3620a513aeb59755cb5c09aa5d19f02b067bc32675d851cc7b8fd087801d5159a76afdd872a82c98b68891dde2464d7c5bae062974c6412283e5b0675dc2012a309dd6b5aedb467f468f216c641bf43aa8517b8e3a7b085183585e8549d2d741d79aab7a457bc0b91c615d18dc2f4484dd0e8f9bcd105dad237737565363dca432e2bede38593020d0ee5aa1fa5bb37659d1881852a5c84dd051fb0029cf73484c0087c7f85f2960d7b0241b4b0f60625f4dc6403c7d23832553be8b131e1874c247081d7166e9b316af6fa09d8c501bbfb0ace109d9b8d6e3cf285f7cdd59aa1f79ad3a869f6bf824aa5af712c86270b263bf1ef317728385da3ad420bf93e4587daa8252e8fc442a4d199d79320bd7d8ea521ef4aff0673fc1b5c16ea33a3dadd0770c62304454392634b1c9a599fed10d3fbf25162dff657b5fdf1fd119b2b4182ca58ea977a8228d899752d960c98b993b11f1725ff5838f097593f6bf55eb3edfbb5cca8a5d00f1a64478d16e8a957c67f7f1aa2e53c9ebe44d9acc335a9977b4fe9b6ad4b5a54c9e57e9a92d04c5ba74915cf451ebb8f16203cf95b1a7f98aa029271ac434370a574dffafdb2152be093fd7ab0cb29f8b84b8e7442125918ec84df42bba646648890765ad34c9a1415259799623dea514503cd998032a8b3bb00c33461e507168aab7e077b7bc11b1087f836f128b9ff4cc3e373a9542c548df2826cf58c808848e167c0690b85de43a5b6abca0bf5bd5f90d18c0f90205ed7ccd8f210e1b67de0c99f6e187a89e9826bd7adc6c8f60098101a9adc09cb279c672a2ce2741e46a8a8f800f16464647b57b24538fb8f4883a8495f2fed3ea2424423752797a2fbe3c59ef259051493946d99d2fbdaf2f91c08d75a32ac22bd30a118d3203e8c7fe09b48a9b942a7dd4819e0d99544d073a1724c33174790ad4d623e4580df9228e1a56fa2abb67ed976d3c5abb00c690a2c137840267d00e8b46f42fb0cb55d95d9809604a56d0a62c684abfe8321a759fb2af7d37295fd73f08deab769a0b4ea59bd5e55afc5dfeacbaefb4a2559d60def84d5a1e94f94db42e11771bf1ea92e94534c5576cce18df2013467bdbbb9cce24355f6b624bdb345b22e8b5938e902e45a8e9297d8f5906016248f1228b4ae5c0de74ae9e0bd4f237dc330e0e10cebc70fa2d75767e298cb0ac83a290c3e60daa0fc1c41e6034d1575a6da80f8e3b53b73916dc1f403d755b1cdb2870fc501a6e51e722d93e13c58369a939b323033af0b4f7214cac8df918c4462ab3da5cbe5335c2f39170cf783220073cc55a7ff77831ec1279bdc02e51041994b4a4d4ffcf25b2a4f8e99db189341a2bdf8c026e1d7ca8925a809eb0f758757282893ffd32cff3614b1068744d05daed4759b0454ab272ca9a74174b72ccb3fac81c645a8e98fc5b617b9b77d8e0f2167619f67af90f60befc22e8aedeccced54a04ebf50c3abcbb7d2e7c1710cf04f1fc08295d52c1d57b5f656ee3d7fe03d794f360edc2f30d3723a30ac95f0ebff5fe3486c4f9a2e19aa635443ba0c75bd145b9350b5a67c9881019332963882e21d542898ed72c6cdebcc60a59bd4f58e3ba8ba679ff5bc981db2f7fffc6863bb00067e7110ccbcec17fb40de6233253faf2a8ed1c2bd4680beb8652056c80580a435d3d62c4f7d59f608629b0bbd224aca43e8af9227549ee15fe046a9933162aac551dc67c4251f0ca89d95638afa41a04b70640ca87f16460c2a949592aad958bd0188c1bd3e902174d431fcb6f90ec7df9cc9a6909e33b7f877f4dca6ff5ac571e1123efb61f97dc9b081c04704658f71ec9385aae8c04463e63703dc560c9513cd4c8d1eb1cce693afa5e0b48fdf322aeb7db3541269713e91ab91e4ca38cce191b84a2a410263e7e193867fc51b5d574529fbcb2549e041a38b55d0599d37ecd3a6f683ad7b6d3ef0f1d2783bcb1a0d1771f681abfdb4b7c1e661ccbcdc096b402e7440d9239188e7e4dd217957632e3b7925e6d29322291643532adbf7a5079b6b8496e1955af8d713c257821c5bb4b2586c9adf02e8d21a53194e6b8246383d24ce6f8fcbfd8c8cedcc989511081437c103d45f65dc4a08691e57f2c2931b6a2011e27e25c6bb7e8bc2aa798eb8eb91b0e344ea444376ea3d951ce3225ad82cb03501eb69812821e9fd98d02e28c64c726ba6558f87b4ed4b0d4898c9f957626b877f07b645b1bfa611bf16382f4559b4614f0896a5a8057484bb6c7799859f1cd7e8da93eacd6a2b0fb12e04aeb007d06b60eecd4654f1543fe2d139f18f2f64dcd04a59c8f4f9d41d356ca9d9c3a5429f334721f7140e5be5ef7645645528f27cd0f1c370aaa6e2f1f3ad8f42c3796b9c57a8a26642bb0cc5cdd203203ae2c0e725f5b930e9b7314bbf7181dbd00c531f9ee32877db7b13a1a80c733f24974df882e2808a24b83057db7fcedf78626b9e9b076c6fc4541577e4021c939829dd044ee52bb370434c041d38e68da73c40dc741d70ef0e7a6057fc1253c3bd0c36bb7a0c70033fce51d44593e0b9d06a4f81b31cb722d10179d757f50435f3db01f2e50eefe7a0339f310da4222fa1d5a7c324b12123f5b51f39994b0e53d11671711b12f080c406b57bb6ca2c12c1ab2cf6798e2272ff0273e1ded2c312a456a7b9657e93b08dd4895f7d38e02ccf9ad6fdfaa0f41a1a4a3d012f571a0f7547c270e21e904f81d3e3f57c540a169d0fca407e0feb04cd70a8f2ceb9e7b21a811a714160ab03221f544dd5dfaf2fc79573820eff30fb80e243a4952bdd4fffb01da038a13c4fdefc042007538882be76cc9084636f32e16944f31ebf5b021665ba8030c459a69570d976c2743ff3b2095c2752f9e25d63b42397f7921beae1f549da67cb9242001185c98e2ed8c358301ac31c000d76b3723e184d9a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hfac224c5f1318c79a26d1bbb9b743d361cb7defc2126b0b34de3abfdc26a9f022ee5d93ddf3119070c28b28ccc4d9d72b3fb554f2f6210c115d89bbff33b07c1961f6f53814f444c4ece5fad79a89e4ed6a277dec35bf6e5bf857e30dcd5f4dd936bacb91bbaeecc0cf87474447b91dc6314747b361088b9f5cce94db34a050feedf0163d25713075a80f3fe0a979dd57dae230a23b6cdc275b20fef2eb52dc95c1cfda744cc87478b6ad112705de56ab8e0a154e78ce06ca28deb197726db2e014648b40225d51e2347c9badad883bdf5f4b5f25216053795461542f13d2572ef2f3efa48470e008ce70cac76c19503f3af204802d39fc36ccb60c5e27de469f6a065719d9027e47f9f7b1fd70024f845799bccd02a934a69e264f7c0035934989cb56e18362f43070c8936a31e1d21a9361b68840a258de2046a17a996cea1a475625c637fd82ad54da21f541d5b3a4edb25a04f06f28b59e472fa8e6c87a1ccced46ada729d223c6f25edf1a2873d7f801528b485d8e405b0c1801d399c095528e4317a9e354c754b8ee7ca6fe0f3426b5694087a95ac39442126402ce9887e929756dcc2950c83c79fd55fe72e6c51b3ebe45c791bbe3b1720af47857fb5794f9202411269ae863187efb90eacfb392cd7853354a22397e0ee812a418531bfe7c2a62c3e129492ee3199e83a03927681b22acc5743cbd0cf526a742d717cc0d85ddff6cf91d4824aca3fbd83ae5bd8181698f61a6d76fb20fbe72dabf7ae5190cbfb555f5db79345ea7ea632eb0675e135628b18cc38a9ccb5dafb78e4cae11c44f32c8968f91ce551d8e7295aa86758449c02e3f605369bcad7f85e9d4b86140f83ec13b636f4871d57c2e5c583f221c26ac54932084e2b9e3dcc7f8f9c2654a1d049f64ed96bbaff6c615740560b4a4ba9ac62108a575d9be6519c7c6204050e87149d2e287447cd1f5788242eb544d75ab1dc8d151c950a5a59854eaf50ccad605551f2a638a41283ddac0283ce07e47eef74797b6d198c2cf9b679e967d0b883673f2b745f66f114fbaaa287f05a051e761c61a7b8517e6bd3b555c47daedecee5795e74e121b5337f0c9628c1f10d4659acbf7eaa0f1d8f4bf59025bb8c2c24938fe8f64e1e16cf860a89eefe922d0e7396cd2491987fc7a3b7ea0bf0c2e3850fdf7d85a5427e8ab4e15e43a6a461ab89d9231f6cbaa79c6f378b022164e445b51e777f311b94f0a1d5101db5d2c5e4a612b7fbfcb56803f7df6fa611ba71e10fc55ba939ee9e139bdf1baeb1c050365c4bade11d7a48036f0c387eb37df2004c604df088ad45b769434d9ad610d06aa8a9f4b3c8710328633c5bf138ea3969174400bfcb344add1f10464a784aa3ce64237373a6d22fdb9b6a26b1095f20bf61ac8d50a7e20ec96ce35e075289cca028648b9882a67a37a0f23b86939704f0216254c0568af9d16ec1d15e3a7580a7729093e183536406f3818f25054740d7a4a09d5cc440819dff628b6716a77d44d3354897ac8cc14b560c382a96a0c5cc200f16a137748f10f5b7f5a38d6e860dab69a10e4affbf89e97331e5a0b5cbb54d21e4516c61f7a1dfbdd28aa22a7a6fc921ffdb2fc40039eec5473137e0ca5cd22846dcf77481d2dab36b7dd0187e254293825c21801b668d1a19bd56ea366f6495ddd1b92ad1373a4d95b73a72240fd1949b2c743f91fcb3f5068ff10f519de562bd9dbc245fff6bc966fd5bd8b2c27cf3672378a7c959befe43905a3e788536d0fcd8ed2b7dfcf48d064f6f216fe2ea4c33e3eb19a0fec6766df14ce64cc6d66fcf5122e6a6e8f238771018121d92e66de7b34187c4e55de1aa8d058ab75ad3bd0de6b5c9d6fe0bcfaceb5ac4e2b2591297af1cf21628913544b2cdb3be2eeff4e1159c49dd9f566de6b2d266edf1b80522b792218b59a4894e0ce96a844abb1906cbc451eb6e355259c324af596039e46c91ad2850872ed435bfab42499ea80824d93b038b852fbd5b77a23488008412ce0dff40905c5bad052f662d764c887975d20c1c82d25052363b747a6bfaabea869ae0e8d9e44c6e61d3d2c4d01a280e3e6f552f7cb2bbd88cd5fec559bff6cba5ecc782dd0fd4028e9a61b22cea527bb3655f7186840074e3273f36e36a6be82317eafe872d8d5a5301dd2d2a6066fc3372360d2f06d1ec82653787e04d869c1bb97c7c4a4411216a2aa9808990fdf5fc3e6dc6ebc7cf3f1ca8c492fcc2ae7ec689be7f319341914569ba04bd705fa9a22b9ba5d0988fcc2fc241197c1e312e4f06821dd69923fab663cf8a7716e488e5004aa54ffa69ee4b6005dfb3eee26a31a2c1b7d9165f1597247198815785730d5e767d7a1afce9ea5b400ee63233224d47356d001e4aed4dc830043cda67af93bb5615a79267d68fef3633725079668cacd1f5a23b077bd6a239a70e3c4bf28015b6889f06c52701ca7338f4118fb4daae17edef9986c7468e8bbea3016dbffc8e115fe30a186d1f924b00cf249f459995299d260a401508cfe6fac32e0e12cb1af65ceacb57f14d61c8126e49b4271df7b998e6c674aadb4338e638999aa54b8899024c3f905d840d563e92703a410808c65ea7d279eddde08f9b90d8cefc268066516e96aab102d60bbccf087028c71a32fdf9cd504b0cc4a2e6e6238af83b1ccfeaca9a06c5efc680bd9a63c255dc90801eb36f3f5d219110d1005e97cd8ce9460b0651de30300aa743b22d5fa656981fa8872065a46a533abb603125bc97d912863d1d6dbaef7d064f4649d56366fe7ea9270cdc8fd72eb4aa2cafe87011bd2797b0c02bcdce2ba01c48b354bf86fc27fa1f64b75cb5ada3e2d4405ded57ae21aa1d5ee2f9954bcce1f4cfb5ee755feee419f1e2a85ad4fce350a9b9d998036468ea170fccf888191c089c0fea69c4fb6578da24f6a36e43515d64b01a0bec436f37b5f5bfb58690e8d2057ff1d12eec8e6fea156f502c39eb3f6c639415176f9326db85be5d74202d22d141e5749b8f07c5917381a9c6a7daad7e508f560d8eae05b50f65883045cec90f3998da0abe1ac4853645f157228f26e064bc2a8acb7e5bc74270bb8be706f5058e20a42bb3dcb5399f2a9e1928be5ead45ed0568f19eb988511586351005122c19cd267af553087639e0f236904240a75c9ffdfc307252ef4d1e54835d7a1c0c0033dcad521aed62ea00bc6e4ff1b36daad2156c9ed4eef8d741598dddafec870f8c631b0239cf322eea0fc91b41e7fb5535db771ec9f0aed17512a9c41ebe344556975e062f5889c81984a60a60c0691fdf93e4ecd8eda3e9443afcad9251b24efa941d85d9ee823e416eed0d0383cf986054dc0e48c37374f795f5e67161f1aca3b973639471b6e3130d1975bacb0678ee719bd36b105bacd327859bc49bc510630ec7bf89c4fc92b3e44d55336080c8a793cd01170c216904cc2545d0e75ba86e4a2ef2e12f1e841fa57a306cb8e13facfd0e2adcde63cb0d85b1fd0bf547cc7c9cba22fdbefc65027f184f921b1177cf5dd4dbed4e05f8acc161cff53d25c05876df3628fe1000f023327d8328abafb86ed07abdf1849bc73b7da8dd5bb09eab33e434c0108f32a7238fe86ea90f1899c87edd7ff0c953fb6a56bb44dff5fc495c477370ef7d7beebfd183a1033a7674d8999eb7cb15b55fb0cd6c37795d6aa8caf5022c42c49743ffa4be69d44bb779017a402c665c57fcc925668c5a63a9347731cad415f5b59169c80188a743d04eda244a22a52379de796f51116f813b1dac762909cb84a16d838c2d66ab5a19c2a88f79c2978bbd0d1b2fdf79f90b368589b5ce6a3b00c945a2789f8e4a0b86bfe722f422a3ed79267d8ede43b625d0a165f803aeb819db2e34dbb6929b636e6df79bece966d4c18cda230f551b7e40019f77816ca6da088998ebea0464bae5afad81d9a3d5426954ff7aabfa295cdbac2a5e90633e7ca8420e0d7eba97adb08b21842da9f07113716abdae35750dc1f37023295424df2fe46101b7f30255c69397bb762dd5c30d5f6d0cfef951ca9f8c71afcbd84a5bd0d120feb103d6a926948b9ff5c8d8aa021cef627869b49cc7e86787a7f3c5700477c55bd996211baf401d4ea78a79e0509bd9c862609ace795616420b4172624adbf755cb9bf1e256c911999741f511623f85ce4bc9b22dd874e3e6cf4da0f74417aa147ec53f02856e04cfe2430e21471cd155319dd8d513ac57efbd3fcf2b0589e9124fece02fec43f34ba16046b7b3041075527fba635cc632e4926d2caaf5f1769dd96e4a53f5b0b37387735467015c67f37bdfb8cf8dd256ed43b47da5864f8fbd820c7aa85597b31bec8f2db82c9116058cda7fd280fe6b2bd33e50460a89a0da09aad0400c502b22176a3c0b59d4590cc2bb9ede5d7240bb49e32c74104d80b66f7812dda8a26e823fe92ed85589a14314d757707aa195de659078113e734ccc0ff7a7aea11a4af71a3dfa9d43dd4c7aae025da6fd57f4a8010c05af2f27038ccf68ed9d8e82ff6ef5714831d96fe58c46aa4f0e162edb1b5af470138001a859ec8319e558bdb8c5625ce0bb45230b1be91e0a76044b637aa9888fbbdd2dbdd01c61beaf41037929d69996fad8235808a40fd01e2fce4ad9883e08910ada111f7d2252c95e8e624b3d9459b0318555cd6f3328651299deb7b6fbec29c9edde96c41735de57155176bec58483252eee3122aa6936f87f38aa274117e7635081edb865f920b93df2b86244b19b55b1afd800cdc1fe365b8277ea9fb93c22f04019e8ddc00ed1b1e7c1fb67acaafddc83bbab2a82fe82821cd9874e70575213cb9c653f3861cba8f0e270e5942792a9fad2616583854307b0459f05142bd33ea31c356d95c858ae33380e44f17a7a9e3da0802f0848467b0496dcff4ea8b018cdaaa623e775c098f55d072d7e65e72af65177561e91711018de2c6aeac895e8795ccf975c2f19c83d65e5828d2822c7f2b17a39073afe7888458b34ac2cce4f49b913562a9ae0f95568ec1fbab4e2f68a6e7fd4bfca2525c35a122fa51215a2f41096e7a88657d82d4b379fe14fe00c6ada207e8e460183b8a6062a3590e6404c4af209d44d8410322d293b2d14b04d35b7421035931d24262036931b3f4945537da637ba842d5e75a79249a2a467eda91b177a90dc5b4c978a25d9404f6760143256b35829bd586789aaf8bff68d1e3c0e22d28c196e30fb9d4c54f48ffaf25cb74a25d536e8c602989813c9ba421743b288e5c896c9ec21552e974dd482b6eb78c40c7323db29c9ffeb161289d095cd7c5360e9be14e74f0308241860c9e250bbf8b858b332feadda3fd9fb56c4c1b4baf3e983ae8907b06f4067193ea646290181445e19602ecd936c6717ec2c94d23e3a6effb19892f92873b668f56b090d4f3a531761b09c48fe09225ed20b6d5cc486e8b9662a6ba309140dbac52d8b66f853dd92354789e667304991c52b25f92b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he34cb2f8a9fdf6d194d55d0de835397f908e6cb5067dd5ce028710eff2ddd6723f9a2c1e725ab42e1c20da08ac3bc8c8b3c8f9d2548f4745aaaf3a7a0a01745863c45b79e236da5ac7da12a4b7f415471d120ac562469c42e1b0b79f5ba938c38ff5f66593db4a29af49cf46a627342dba08699fd43c00ca1b7254f0f05dbfb2f58bf5b07b622c25f7e47b53848ef0fc5a7a6067292190058276ffd9d28156175db93fb2dac73e400f960562bff3df1d662d98ab66a20124dda881724c8dd4a3a5b28a5dc052e259384fb0089d52861aa81f6fdbfe757292cf1aa02c2f70cef0f0a7cf0f8f766b0da38cfd1aad5ba18aca6fb8694db8928ada4403024a662bf88a067c4d00677591fad8151dbb3709cd56056e679124bcbd39638c37aaa8e2371d489fc777ba88f6eb4aaa03fe9ecc889aa331b16b29af6f0493338d7370a6f2ce6c21757915e076068385a76e395bb3e82377572cc329435389a0686598bfa434492eb72570601da1b47f0c49366c30dbef3de1d06b764dc6bc0b6962c4a04e18753bed4ffcf7a44d32daa4fda5bdbf29f5338b5985640aa0316a4b4f50c02545478a3b6431945d0b7a05be8642fc1e2bd19e9c6d74112b1c31e539cb54b2da75f4887ba482a989434ac35084af7ee27f97fd70617c2a4a0f62d51252e61a3f2b86d81135e62569a400ae2ea9836cddabec4860193e3a6cab5be9d47a1a3cb5864060692b78341f45cba1f5f9866f450eede6d16967417b25d47ab8ed19d83e2ec3496acd9b84b1728357732602f759c2d32074f0764db21c7cc44ff1e2d863d1bcabd9bce2156eef9a6686bb1837c55030d1f801ac689b540446a864047fd53e870f28f06241cd73047164ea7f43ff9923b5ea668261b798a5beeb47d00c82e86445ba454cc8ec8a0863d24a7bc89e2cd19ac0b0b19c605fb2cb9c78bc50e401d1b4d5276dfdee4a6c279130bb0f787884bcbc0fba728c6a889de09697c3ae0e4a1596cef53e5e3c64ff462c4e984eba06039bdac950aa675c8f357e4b55e98af5dfaf2e682504df18a7ac31c60226a8b8a863938d0e5fbd3381712607fe9a3ae9be4d405d6eabb57076f1debf947031f50f3fb3c8697adae65dcc7f660050c0d8effbfeefb687f4824bfdc497950b1b8b30161409792a589e58ea70993ee30a73164120efe352612950aaf78ae2cbba257a79b310b0b8c5d35730534d5f03f167464d63cdac0e0297656e45ca84ceaa4c66df0159edd5f41eac4f171c1f1af00dd275aeda95965348b3e4104cbebcc6cc1f5d31f0ddf32c832f56bc37fb33a842ae4f172244e63facb3642c492d1ae81d8eb9fe69fe7ef7abf711d184d2717a0f597652ae73b9ec68b8ca4297907ed74bd3ffaa7bfb98cc02be07d11def0d275ddeeef8448b7a4a25fe16618ab2f0b1a159ed6ab5da4ab10af193435214c913e21905eec9e551425e4cead9b85e52e289cc986f343d206a3fc130ac37f79d0f2c270ffd28bf699da58b8c4225b7e512630f3ae59ab755ca8f6176a664a9aaddc456e24fa3f10d947654c586cdc650e6cb78093999af1a548b0123e056e374cc27432de578168c873b018d50e49636eea51e09de0fdb94a89d71ce33ca538aca2f798afd38cd4974de54f27b4e64141d356f0d5197f1362b748f2e0db43918f8cc4db3e8325042522fb1eb6ea0a81ad4660b26c37dacfb600d3c9b40d06b964590f4f3d7d324cf90ed7ca1fd95199cf0860a949845d390c447442615e20043efa83b2b5e8364f9937893bd98692a3639083e3c2689c607ebd33ef70b4e7a4c5686a7acbb06d04952279554b753b15cc51f85df7497a0668b3b088df8d63f7979d0d4700434a8b145077ea521dad4d84cb02317b346f6c0b0f9f18c0cf93932477519617f8f9553a6d13d4d74822df1f705b38340bcd7af7faf58ff4f8832ce6199b428b349250b5898cca4e766ea9a4739bdac482d209384f5b42ece6b24158274e3ef1e76eaa1fbe671646d59fe8c6d3cf8a9644b955e70ebbe697f5bae6c801d35364bff412a5cc6a36372f572062e03768cb2fca5d904f4b44c5f76bd4ce86886f3f688479b7337052245a33593c2aa40af29ae0d7fe3fe5407680f6b3b7754cfb918e8fda158956fb29d960c367f5a998b03949d37efe6456db5b87aed60f994a6644e23e1557eefab09660f75c9152cee7a9f0f117b3ed44396155e060f7c1309cf1d47a6c1b61e2df75c80b6a31d262ceb5683eb6aa5bec15dbacea765409d7032f03eb427cefa5f1ce71bc4f50b2c89b922d11f91f74fbeb1f20a45bcb0eaa0bf451a9fd2f87a261f4d177fb86804a474e308fff1915e7fb768e47e7986f2564f6a8bc21b74a907e4701433b4e57d136e90955fd8276be28207e61ea3c155f4299782b6a7a1ed912d81b087a48dc9fbe7a51545c0d1435f88ad523cd34c5261cf8cef7a0408f059319e32f3c549d2d71667fb02d224ff1c0086858bada4ee3e0a0ce22f3eee7dfb23d4daf71e832b8e6921a1e012d566eb8be544ae2700237be7ea208c6dfcf5ffa49f3afe535f11858ef8857e4b5fec6999baa8dc06d290d29dc819a0c0db0c958161c7f536c420c679e2512c203505bc04d156f3e8526c741c4c75e450c6ffef4bb1eef9ab9afa541b065c05a3b1e05a35b15cf3df2b559a2f745c2f0c4d85911994cededa13cbbba773370272173058c616545882ee405e92df1dab0ccc93ec38b4e4535c255236be72909c1359709172a3ef895cb1cef254b700c88e799807e6f49f20023e3d7dc1b549e76b364e7e6e20da24a84d4500396ed59f9b3c4929183c6e240a3bf1dc1bc44586cd524fc48c565142f0de4ca6fa016d94c72b2de1f19f929425c320627e671ce63bbfcf16956928cb80b075764c8fe7f497230993aea404bc2744e27d6b9396d675d6f6e4f0de34ac9138ecfa1d9b83139ab2870bd5f10d701b343b24220082ae3b92ebeacc115a16ce69de422b7a569641ebe174d92d2f9a9ed4ceb7788fc66df637098eba0a420cf1ece9a405e98ef5a9fc23daabaf477a0f90cd0583f7afebb9aefefe5fd59740ee84c14275ae9d65c62a1076ef3e130985fed6b241c769da88e376b074c0f1b81989be958ea22efe3a54bc5726d96f578c586c968d81f5228e19c1722417bbb3ac3414e038d657366538de9499be1d65221bdab9d40ebf550df0c7bb7ff9970233ded03ed6c83eddaaad698bf743f1bd3bf8dfe3b8966889a2996808c1ce0074d6fd05f1ef2487f4551686cc2094bc40ed2af2d5068c4c4fb2449282a9a7235fa8e289c8a644472a21aab063e3d8335469a906a3a61572fa4e275a7d74a75688208bd6a8fa4aade84cb3b9467f0fb4f8330dc80ee2c12d4d6bd6ac180b04dce343ee3ec4facfa450e0eb48bd716242619dfaceb3b0196b20b42e939679c77d944cc86246de9650cadf99512f7834abbb656d64b397fca8e4615b2d7f2ed85317d5b9144c7547193af1e3532b4ca7742998b3e7a7ceddc5191caf58833e878d3bcdf4f4ee48a972c58d486d5a068cf3e0c0709a811e4ac55222e8ee2e6e15837624d833bb91319e97f9dcd50df20f09f0ccc60b964213df11f5bbdf7e20755dbb8ef0d0484073a4b461b229848ec5c5a6f028715f43c4fd40eeac6fd46e84efb553ba785ace1e88e0eb7c28a750b492acaf77203f6d5a2a5a134f636392aeece59311eacb7a521d1a5ad501e78f80fd21f5b3497e0f3a5e813f1fc1e2df7d98bffccaea943619ac6fee3e2e75e000a9a7276260e63ddedf0c0acf3682820f183415d6b30bda3aeb40e149994d05ac660239b9bcaa480a31e0906d05c5b1cd04b3ee35f27e8f28ba16ddba471785b663eb06eff5f02a4a76a9adb709b72b2ac95d64ecea2a3f60093b2a753c7bbfa0bfcedf46f22a4da4013850e6b6420a9594f8040bf4cd5b1d1d3e0746feac10ab854fc797c0926d05adf72aac1cd017f39d40d582457f4a191099c3865074f4c2cd7966138df31b24b97c57b7743d54b843bd4dc9791ff57bccd657b49b901aa2e0a291a59e5c58d8b7b977a44d2cf2966546a5f3a8e9c7a0f3be459d514d5478deeb3205975f6a02d565c7ecbbc224892538cfde4030220a2073c6cd6ad86a82457b9c1ce893653baa5707aab915adac50d605d477a338ea243eca3b39a64554cc34f951d9e286c10c9600e9a8b33aa55d5dc3b94a8bacca91cc27f304a0d67acfb6e821152b62871d4fca3520431c728f49d5f84fa25c4d4696eede4dcb3d3876eebd72207ad77a6dee5713f202f83fe45f4818bfa30798d69f27f036ac6aebbf18b13bf4c287a2d9a85c287f705334c8441be5224c3cdfa8cc24d1fad1aff0e9779bddcb4e10ab66cf2db4f6ebaa0ca737c8ea2e3938647ee44026efe112f32d7fb6baaca3fab74a4cea6b779e594d9b5eb3f7b2d5156c46971771cfd7bcdc6bca3942b6774008b233735db5d2244ada13fd2873e56e6133f01ba01187d24c923b4c34d81b01cb2067f07434d2ac8647d3c5b421bc888434312d5d606bde2a82ccad249f72734ff38b51071d9466ac1b452ef3406e74885ceaa1c6b868b32cd219f69dbb303f46c29b4fd18065e06bdb2b04f1ad828e30b8b21b45cab94f6dc161ff7ec6c7ae262d57cacf7553d82fb7cd50f42774f5de7814febe33b7898acc257ec4b0859cc2308bb1da72d83c81f120a300d19993d0d0901da3f5034dbe8849c4f6286bd250b2d6a691a997a1156ae8c14f52f58e1c1f5278191343254ba5f66dbbad9f8cf709410dde515fbc8ffffce3693c3ed2d5a64a7755676590265fa24c98fb751796902cd9c29dd8b8741b78a9642b6a3323b07e1af30bdd95251a3a7573b2d544540a1ec7cee0ee33faf82d04eaade8768dbf8b0a807b7abc7491ebfb64696674dabacfc6e8422a81d49d71c75992ec8c5d069569e1dd67fa852502f0321d1be2e4dbb1c03bdb8ac3fcbfea9532a966140259e9e158fba0e939cc6b1d4a29a67aecbb9d2a244d9b918a9ac3ee2e72bbc15c129ae83ee5a254d98b2a16288458a0b4ca1cd6b2d815c7ec9a0a90b234428c6d0e56cdfdf618a0b1c4e705a4a8a015d01adfe8569d924e109eb86232d58d5cc469c8b4533bebb59faf97ee24e381651f7d3b9387023542d5ab8e8fc158b53aba9553acd4388a51388e79a1a810a42b3be8d17d4ffa7631661341516dfb0640740400d22c21724d361496c4042a78ef7979eccddcedbd21bad170eb4410313272be2766bda5c94e717f78f38b454dd16179289b81c64eab3aa06e7fa8bf085249f6eafaa0dd485ba25fec048b4a3cf184de684b4a43956c18068319d7b6ec30f38ed07196ef7650beb48e34cfd548c8c6ed1bd47bd8023310579c3c06986ac288827c4b4b577574c3112ad47a6574b57c762e8f1269fae7138f3a08f6b823fd252917416489e75415c16a12bf98af90444766efc1947a461672c3c4d4232fd3b045a3148428e8743bc445;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h7d851792dc590c576d78ba46fede6fec14a961d2dcb8022535d2c7de1f9098428f51e0d055e60861386dc38a8d9a5436be8838402e358d599d8985b15d9a04c09b4e267e3bfc431587ddbca7b3c092be3d2e3d203a5c3053e2198b640f5774f0ba02f79e9c124e80b1b75641230634dd2952c515f191ed2783a6d0ca893c3cc1f2ba88ffd65294a805937272f74489f6b5b378936d084de4291daca62fe646a97baeec0e127abe65256f073670b836de8bfc9816c0fc8d7e67ee74311c516e105d19cd4c989cf4105de55e959e0406b25b20c404cba4dd21de9a881bf5020e0fe3439714dd2c768b67622774fb792213e90fcf8c914dde5540d003c7bb3d19bee85e504e17b5a23e6bc552e2f423deafa7d85a274839c2163953821df1f3c07804b94f2bbba9f87b58a0ee0bc861b297d4f5aa855370525085c170dfd7f13b14ce5f36e6ec800ee48c33eb926368fbbc01a6d4aa13ea888dc4d2d8e92b54cfced2cc37e1430671ab12fc846766b1648a00fc6edd51285ba9d4798a38dc501b2249e61bbd2be4e3ac08543e2cfe09136707281a8f661ffc541f78b53b2155c19fa4428daa8eedb15ffc36d11a4b18a486b38c2349bc86ff6c41ac63dca43d79c33023a30af10e80f925aba2db992f22be646212888f008cadc985e81f25b26131d0a87f903096df6b9892c7e329a7eeb4679523ec876b92d840f26ecadcef3d0f729cad89ccb4d702f2563ff9753d6b75b4c69046ce880843de4d09dbbd00b843ba75b683fa0d01548501e31740b7c0aa03e1b37bdf1a35dc289f52a07e66b5b1ecf271833334cb44e820bb2bbcabe8ad3a3915b1caca64c34c8b26fb748b6287435a66dc06fbbab80b7912039cd374a884d0e628cc45484fd7d4c7246047fe4093b4695dc4e4b64cec16d856c4344fbf398813d63fabad690a5fdf0f604252f69cd30a366e39fe03e0da64a9268ff83e1ecd56eca12025543bf30ab78a726643fab23d429e59e3f3c3f076f8abc388a3b604224a731222478f0ddbad4ffdc8fef576d6efdcfe25626caca23635f9cb4e388dade4f9296f5945d5d4bd5757986ed36270e9330c460252d682148a23d32e320ec21226d977078c535410003921e40284037d99b1bc5a4036208cb024129e34233c2bb220b2d31031ad17b469096e9a0f7a9e6c161e1bd2248be9920c91d4413baddbf58d19c88387353e00c1375c218bcc89c571f3963482b7112f92e9024249bd924cc441cf61dd7bc365ab5b5b4e533f501fbfa7b8332aeda41de6dbf3ab6cbf14242e4143aaa8ed2f382bc30b931a8664648970491ca715d4703f8f4915d78a267d093545629272557aca9b44384afc408cc94eb51f06ca3ce58d99a1d7e22b22abc07cdcff74b954985f54cb77cddf20a7249745e22a83f69eb28907a174171eb7be39a6584055a1f03446e668017b1d27ec79250ebba28bebe90f1b0f662016acd0bb6aebfc5062043d55538c0df8c4cc065416112e174da9db462b06b41c8d8f1311c0faadbab2bcb8a2bdc16b676dbde56e16aeb1bcfd2cbfd2dd22ac58cbd9ca73b05b0835a83e96b578425b7d7ce02bdc823d523969f57bb49fed04bc4e2759fa1e133ece807fca972da8e99f7a607c668adf1d4057a2b2acef0788b09015bf98eee0a3982f483bcd78d244c9194ec72ecd55ea838315188b83d40a5c2ff259935ef6ab8abecbc7ef717b9ed6f1dfa7084fbadf47ca6585d441b0b0c90c21aa0e96f168d3d29ffc23a93188503abad4ae76c735f4aab1e5d0926ea94145ed708179b14481d717ae6701628e98f2764ea1066f821a52573d6ddcc13ba3e846b6a6fe361927995f7275957f897b6c5dd16d7613442aa3bb58fc3149896183480b4eb97e2004e62055aef1e05bee7ffdf1e17cb301208db1e819b100b3900e03f570d8b2d8c0cb13762b4ac2fa5cec8a7892820dc5f9fc584bfa1f4ddec0d66fa5d84e07fdc4a0e6a5d48dda0210925a158d643f37bbd5b562c67144ffcb0e8b4f0e5871a70a83a7a36c1617ccb81567982c9963e32a393f5f924c9a432dba463746a50e7aaa9747fbd2f71f04196f9cec7ca3b56206e2649344775e6ff6545fc4686c46c6a37160cf607c77d43a19ebfb97eaae8f5a83a80e2d1fbd65cd2401cd500c7f0f62dd7543d2ed4cbf604d302537229cef64618bbeabbe06cd5b3476d3edefdb82a15795192fcde26f0330693a22ca099fd626e675302cc78107387e46c1b3810e2569f9c2b39be5e967bd264578a4e142b5f18e9e2597b2d3ab10817af628d56558d3b65a64df3371d0c05e1986e287f0a4ab13c275d0298ef9b4acaa2470f5baecd4f6f9488da5d8953c897d7d94f559253001b84398bbaa80db6939ef5b413b4e54ef7d0ece9cac38fd6e60b77715804ece5f2930eb9dbd0f31b8053b754814773d6b33fb71c573f9d27fbf30b745497f14626ef6c00c01d2c26c0c38e234fe1bf5060844a6b25c0998dba139557cf8804be29a7c671edf89f38fdad42ebf58d01eca1ca94bbd9bf084124b752784e22bcd1f0ccf387ce136791b59d9c4f583817ce63f7528a730cc1c1097f77426bce41829123fa8d74c026d8a09833af0dc538a4666cea935a372057601f4629e6181dbb1074d9268161e3a5542d085903e6863b05fa34a176302b1fd5f68d0e0c08af91719ddfbca13e456c3d4e2145022ec6c6d4aec76c26ede40f01e236e631ee83a6876391dbf39c01e6865dd5206dc1d6bb4ae4a59304afca0c6301bb6eb82d2292fbabe369d7472b816484f0c4fffeb8f4b95ff973cd8f52496bf806eff1edf17599b1c6d5fc5cfa6af189bb7a81d5676ccddf0dae71901803d30e5bf3f1ad2ca794fc2b1f575f8ef23519bc68483a7d5138c41241515b1261f0cf445a94ceef6ba0eff81c9cb5cc87e054179f7f06dd33cc6c3c6425a4ad97ee29bedfe1fce24b57cc7a1f3d00f2b1dc21608767a8c6ddbab992499f574fd9a96e6ba96ed5f15beeda8126b2c803bad13762ddf42e978e6524c45e8ef30b0b98c833e735b349d617bca927cc790d16061a3b6573d115f70626200133e053a9a27c8c8b896e32a16ee985be97ab92dcf54bc820ecded86b49e7e97d5c6e12201fb20a58e6de09f9452e955325c384f3166a5c0140ffc4a9c87f782125b517f0f07b876136aea7db7dcc2dc4d05762a16eafe26a671dfc6a4326abbed946f85760e9361c4bd7a9af44ce1fffe74e9dee860fe8ad5ba39cd8271110aa04ee85c888d240dd81d0c7af9c2a7a7d0ea68851178f19530983594669a120aefe72f4fc3d0a20970011d3c728967823606a0f0ec80a8a8356d11069706905613853b4f5936e07700ff4fda9588196f16e564820dfad118d8569344041ffe3277a16c7c48dc19a1ee6771329d2a0e7af151ba044f2d7665143baf06691c0203fa7bc095450e8584e0f740048c288b5d421de7c05f1ba896b4066df870595dc7a55b040e730adb814a1c53c8222113043f4522cc1c94083fb0d43c4e135f55a48c01f41c38cd8c12df40a17f551e5c27af2a4e0a21570ed7ee4299354379914978adf13ccf580de9c2c42a7218853209f27f3480ae2286337e441b34978eed2e649becd459909b8fa06d7907c8208066ef6233640ac711ff91d4065573c4c21a4f1afdc9c1116e1cee34ed564700b387aab87380eabe21c7b7121a815300c432bd5c3a23f30cd1404e8c774566295adf8928ba9ba8d238cbe286d60d7714fba6ae673f2f06f7f37c1774521c7bf20a08a9faef0091e25cb311824ad907a79d8b955491e8a0141ad8c4338fad018c41c03f1a4a10000564f93b1115b2c6c4fc3acbcbf46c278490bb86d90e3334fee71fdab989b0c899e97860c0f8f23e14aaa215fe093d8d547962e3a77cbad1c62d2cdddefcd6b189ff89678eb5196a535b95a0888c49efcf9c36462e65bdbecff05112878395f624681a76f8c31533c22e41e8c6186b5735eb09eb4ac98f0682d218354b060c7562d56459290da1791cbb26c019259eeda43712580c74d128ac1a3b0efc4dc862ac2c4c23c0d3f88ff3f0c0e74cbfb4128b7876516ae32f24c8f32af51685ecabd1d83a050b7632eedc0e0dc29e103f9747e808ed0b4b9f219d107ab45962cc58fa1dc23c4bd482b6ac32ab80a5820a1e1a43bd1e743d9ea9cee17d7a7b23e0056fd48ca548bfe193c63b8cd90e5c1c43e957a89d3185da78b919f58bd718d57bce24cef9896a3a7c894bbe2e0b0eadfc94036ac1f342cf9f67df4a5d5f9859938fe21f7516f753aad020be546405e3f3f7ed0367f4606071fd14f972cff6c8a2cfd61f7b0b8f67e3caff2ad8375b13b4a36ad5889b68bbbbdc98176ed0e18e5a9a0d2f3c7b7086c32da3750e1529e1f03a1fcb0479bd0964b6296faf4f60b8090a08a5120ca686302687d8d0057de5aa61671a7d2a2fd2abb8bf11abc53020e31489ee417d0e90785d076209e17553395251bcd5e5ef1795fc4f85191cfaf124e1fad7793ff63205f5b3d2d3c4f2f2b4e01ccfd7c5f34347fa1e7ba869f4a5ab56f2c18a0ccc2f9c2b802e2bcf43e7f5bb92e0fa8c9b36c00a0ef95efc779f4c83a426fa622f3184326d03ff39062e38091af85809f1fbe7202d5a18ef446772a9c0fdac52bf9c164556f996824ae259922c8eed59c49a6d6f20e6f595a2dc1a3caa1aedb5fe1a4ae134b537c01f5b4a62498945494f68b3208fb9ee15fb5fa34e7e9697788f7e0cca4af4de06241c7a78eccdbe295cc567d2bcede100596b131bc256a5d278fc461562fbc508527d6dce1f0a9c0f17bd0f0cba00ceb2930ea11a916f7bab8e14c5ec36f4feb9b017f1fd9bf515dae49377e05ebf28e9a9fdc912c4f04a11077c870b07c0287502ff94d41de4a70d5a1e731e5f5b28d6693e96eeee353e187dbf9ab6f971d200bebd69f7b3d50c5d861bdb48268e169362802ae46b0909b067d2e5722466aba11ef4e271fdd231d6e78edfafe40373bf56a5fc0a9dcdcc7c38268f84645efb61ca2f7cc034009a81a7fa82719238c932d3f2b8bfd68ce4aa20aca7b8ab96f2fa55dd88d12f6782f368bae76f17c18265380340fd9a8c2fbc954dc0f239be0dd27b81fe1abd4a47535caf950d68524bb5d529242f508aae46c9e42bb880eb0d57eb99c60c0bd2307aaf546cdf822ee9c17f6d34a4170ccc1b5cbf57912a1b7a5f4343ba624389f3d230983522801cc5c6e0f2849044b3b33f48128e2c87f56131006119fc7ed602d2afa4bdf21c0c500cffed3f48db7830a6cd13e4f3b495e2e085fe7cf7c83d9aa84ece3f9756998c5ae7247cf3b8a1709522ef54441f73651e840a6929660102406dcfefbecad00c37a61e8bc4f779cd24dbc0d9ae4f6735f729dac7df55a016c0f8ec2d7f0fdb91f264d8cf044860ae4b1b86bfdb7c6130079156da94eb958c04d6b17293aa0f759176fd0442df2e2de0e13c9043ffeda7f23e42bb07aaecd9dd5d2bdbbd4100;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hd69e104cdc7705ec41f52e1e3224e0574d27715c515b5764bdaee47497c4b62c9be92a2ab1540d30811f5cbb74cb819c420cf2635c0c3b46d528a1e3125d8ce735ae9329f873fdb3c14509d084971e6557e1e7d31facf98c81134552fb19f42eea06261079a3527bff98ccbc14855f0fb199682240786533f9b0003345f63af8d8bb178a76aca2ea3bc73dadd4b1d80feb6233f02b5bd7262b97bd93c1f5a50a8575aa7f261bd9bcefa2fbc488ff5a335ced4a402c8f7bc4c77471d982cec028d875993e99f7c6fd403426a80ee6b57d2aa0a362a1af6b1c674b1695001dacae156032acf09724c718f25b2018309bc0b190b602495c7042b59d791378725a26c4fccdb5e1cb7b1176a32908b6a19f23e9d0e0152b24f1c7f35c67260d53bc9cdbd47e967427502e2d85374e8c4cb3025dee9323fb506fceed7b3d6bd412e6f883e1e6ab5a0d3d24dc5371139bbb7eb31747f2ae1403abd9a277264ab9faf7af89a286bcd2bcb5bd68d49e64eee92dcb1175314b5bb42159b9f62ea09570f7f692a77a1bcbd7949a4487aad36b1dae71cf8056cff9d3ec588ade576e7bd51976ded94e49d250101ea3c0decc8b2bc3963fb09772a18dfdfb46761ceb7a30ca9ba23086f7dc32e3f38c862fd668181735b0dd8d1d6765ba1f45759bfa27c579adf98e499bb9763a0fb512aef67b1cf4bbc825b8b1db25a4c90bf620823b6b7763c5185734d5a4465257278c3d1d5f195985972a0326e81d912882a3aed80c079ea59bf8bb73e269547e6d16fb1be11fd9c1d563cb0dc4bde82fbf6e41ebd380037a253244dc2c15ccf1aaa5706fad007e7bee50a61049877aa22724bfd865cff3a6a082e640530eaa769fc576c2888f1e7323c9ad7423b59b19718e2ac5b529cfb51154c624032be5a7d43f778b114676ebd8b262be45c4a4e8d5bf0a181f3ae0b5e1dd07f6cea68c5a581bbb95ae6fa54b26d2f91bc5328fa96ea8206bf26c5247f0dd1d4afe3474ea4a96858211c47200bc607a141fd361a9e8405ea292bcbea10c13e6579f9c23cb9daecb853de818b8d091a81172e1b4c6f5f1da7eb0e8c2ec32c832e14d2f5cebb7071652d058416d347f77c9d7bc10983be9f0c42695acc3e082c1630a25c8065d412c2c56d89fa8d395bedef6db38685f5e43ee89fdb45b6b98428f79f92f563eaf061ffbffd43d20a2cf74047105955e8d907350999304e93a24ab601b572defdadd7db1d7d610d3b96099e86cfade0c9b075dd138c74892d88216fd2e7b4abf0d4db1aec8f76eeb05b882c23011f1bf31ffaddfa3b2b8f14a837d54fb853f02fd702bdc55c5f2e5dd8e3b5b6a7fb12dc489b4d3b17b1f3dc5835184afc4b5a632ca1c249a905f55a8aadb7c15cbac31ac23b08646f4d53f5690d7b84172ed49fe7d236fc978fbae48efe35643bd230601a36c380dce26e26a6a2ae246411bce56f832551aa2449931ad094c6006a63a11d6da0dbd734392c0e8b1a43ebb178036c23aabfbb6ee4543f48e1d6c2003124b32443c0f72c0d648d6685470c99f173480d323fade49474d4bf376a83b0929ca454e758bb41adc35ba100b00b34bd852247ec1722a75300ec79b2e7af84563779db5d0d49c4dff4bfd0d9a0fee63f914832025d79c440bc4d78ac90f59a19804ef6c6fdaa95afa2f5d1b0eac3b304271bc5ac0f3be213c87f449e3b57e187593ac48ab40adef5cd2f9daf5ec64af49da3fc7d0d384ab52a0e4e67e2b342fdc9111aa3345b6ad686aefce5d7139c42d463fd79d628c6a1d47c72d60368c2f01b5249906ff37c26eae767c5107703ea17dff5c1b7c7fb1bab7ed86b92915a11a8d68be1b22beadf1740c72adcf62e1b1ffcf79aea9a6c38a8da0bdce38170e076afc1cadb74621daa4c945acf43776e4aabcd4820911e722d799b6bab622a237737cae122b4ecdf1c89c3bb15f2981164021bcb9a31657da51b9c444dce61006e29690c3b4e0a0192ec014d399fc5f1e379376cb9fe81f3f4f20fd5f437ca464f67ce459d5851475a6712a42c520ea08cc69185a85f86d6f9d62ef225457db23cd6310fd868f777a14652c17aa297064a909b3f5388068471fbeafe2bd60736b12a57e36f4da234831ce00678d0c35a3b3de95d529080f690b179bc296a38c0fe1247ae4511fcb937c328efbe354f69a7bfc5c3e7e6c2625ee845a0310f8fbaed4ff8516a0b4ee89aa537657609b4c95a29525e95887f369de99c5028db606c6c56b82025a9d42971d3bcdd2bfec3c58962617474a7d9782c461cca65ca380f5b2bd6cd51e44363e5b5c70bbb58815d99bdbd75bd6e08eae9cff7c9267268a23b115742d017df91dc3a9745045e5681f0b73341ebd047eeed760edea23d7e57ffe6a237d6a5c3f871daaa5af08482eca5978d7df4aad49db391d4b248d606269cdf16533f61185553dab719802659a58b7fec38a037b3cd78b754062fef88f00b7375cefe27b187d95eda9897b237e002b1a92ecb3feadecad11ab74d4727ba83946fc3e5dbbfe44bb51b020ec060dfaf9e241ba95b11a364dabfd4ae23ef52c89db053c8eae4f1a0c90f418108965b63f4169a1c5c9c6e7989cd46fe658c0668b46b18303aa448f5ac6b01b5fe64d49cc4014d0cf8b2f44fe6fe58246a4507bc2908bdcb11194d9f22a0ac8c6e7ad32a4c378dc87dc6b6245be744aa635103d14c128e53a50bffb3098512d150e4a78e6cc524ddb323efd5c64476205f559dcad73f27000467346c621f4243c2b21e54c43b65e10618c5618db076bcf1672a8f8351477febaa36396ee10d9e40cc2888cdd9fd7f3de9ba725b31ac8def94a6c05f4f417104436d66734cfc0ae70d3193d5595587acf7a5ac863dc7e4c38e2a0c4959d4f762d25977a04c24eb1874f8fc76f1940ac33356965de3a81fe20d1a3ff6269e3db28c11a4719f4ed6bb88dd6b074f726715560b64a1986a20774e76c045b77acaf4f7c4f56b2523f3ffb9e5553043bf338d8c17217c41d4fca62fe9645ca98be36c76691ebe4800456144bfffacb0be7673759724559cd939f28f24cccdc0142427f7a40abce6e2c5b7948a266bd572913f852cda58ce0feb977b1c7bdc1f29cc9c25aee783d6767db9163163464683824926fa8ebe4fe4465a07b204e723db7f7afe6f3180e2704c66ba228272bca2d61b0dab24b1551cc89f5feb19e3d732dc106fd0a93c1e74b37299c1fac52d22865c80b601119cb8acd745748f9426603b74f5b92d51ac83d99687162b4215516d246657099792cf1705d4f583e802d83db1307c45b893962a4f6bb2488d6fc5d3ef31e13a79c71a34cbb2ecaab7f33e74f690989d8e7e8ba1dda8ef62a310aba91bde394d76e12b44501947fca49118475f685c0653a600aea3b5d9ca9f2dc976f66a6fc6aedb63f519069ea5b2fe9cdb7268e2fbd1f8d715a5a52f793ccf1878ebc6820a93143b6a188d24c8a6ae3ab14d7e7664d0941e09a5eccedf3779f3add001935523b8e61d71c4f32b9988de35217663950fac6afcdbda5bec2e02dd10e55d11b11cea45e3d0817974dad3edf29e12f61d97c2e58eabd97f4a525f7a38824c12c06cb818715eb57860a547a3d21abbe8f6510811567fd08b39973b42685676098f8c47758b44303365cc28462caee5ea8f005b0286d7d7cbd92a44ab55437fe490a7f5d3133136b4e67cf40dd0f029471d088beda04259fdd76018583fc519ecac4cbd553de9d6b1f87ec6c21bee673a4f444e1b52cfa4bb48f989917c1dbdd15445e108bea00e99d075af8bb2e57dc1bd2328d77a45a3574bb4adfef542ee498a35323758ea3d761162ee91ce41a6a3586cdead1f0f94d5b6cc5ebee776695b443c209024b39d3d4677b0b4cdfedb0c7b35d0f0afad590d27923134b03e66721f51222596305f163d8116a66cad1e1dc46dd1a419943e9669198bc41d92f988e055815e237b3bd16fae66263904c4cba20130312011dee41856782ceb22af7ef8b231c7b057e78bc417700d1dccb4505fb64118976e9878602591534de1fd7aedd4a30c20442dc1f0f7c22754b9927f29a245026d80969f5c25e0f9440cbac5d692efbc362d0323ecfdcce4efe6575a9e6fa1886ff824a89a3e0c6d81350f00c6d4d08dbf862162db23d7e3b711aabf996b18b549430c2085f065aefb5fa6e3a8943667caec95c5d6cf5795f2956abd413cfa2083589f1ee4ead23805430093fe942acfd65517b26c492e49fd9f662f1dc86df5ba768b0a945fc6739a724112acad706aaf757630fe42f2b101da2200c9dbb867497e2e85c1691bbf8e570e25b74d2e4f0512bbfa85324c790f00543fe36ae5b71e8cb6c61b95e283c290879631ab02fa4c93d5d73a27600ea9ece6f05a7b5302f3c1c87b4c15aa15d5ed19d852aeb6b48136b3d564a244dce533048e2127a25a0d29ca9799593155cf61c73e82972c3a5718b6c83d28ee3949a739a32acf5a7ac72cf08d50e1d68f5c7e6ccd4a074c2192d536a2f5f36c4a3fe33954482d6cb45ac6a12be9ac2f3f6d6346f932b0f72027a9762043eefd63d97284346ed70e092b9ea6f8507e75732db8a689c28aa35aecd540982b747d47369756213772c0a8c1a8e0ef8b72d950a113073bb0eb2d366d3f120d46c7962b961680c36cecf8c52eca2990d2992aae5bb044f0e6b2641eb14c7f14f8b3d4477ea9e75c89191587057ceac5eabaddb5cc4d8243267f30b3a10d1801d1a3c44e1920f1bbd08a4c28ee73080f28f038a381e5d6f1dc7c6152256dd523a7642dec850c1dbe4153d8b424edf3958a64ee3ca1b273c3663626ff0c0433fdc58b71ddf6bcad005bd7978cf4d47bfdd0eacae55cf6fff674a523b987930110f386b175867b132ad688e4d4d530f503c112104ba411ca223c898ef1ba4a034e4fe9ee6a7fdc1142dcbecaf89bc60948e0d6bc74e54091f30c5d02a33dad1af141ff2abb9818930cf73e53ce9c6e413f5ed9b9006cd22c0b560673db5640bb07c1a19a2e3094cfd7f1674575a6798029420a315c0a3e76c1de925c80cce88880b6487537b85cfa1231ad62bf196e0c913793721b9544a7ca700e79dafe466e7d7a000f7cb17484d44944b9d5b422e88a641f577d98a0f53b37b5b0baf9cc8758a272b3c78e8cf5a39b585ac59abecf6860f9f6154305f4801747b1063999e5bb0808a06f57350010d39db51c0d2908ae07ab7782d9ca742588d4a82867fb9a8ca741e3315b8d1661c41971ed3c59e09f4ca509f85cad00d96ca21f20796674c83173c2953da3098d02e622b96a78768d774fc8cc3957ce9e8c2fcb86dc0b682bf186910b60d013497849342e60e15e1b2e7ed6f2a24065fa101810a8caeee9d411ef0c8ae197234f809b0efed925ec21c6efb197e0d5fe80c852ed01649390e73b4850ecb7cba86ed7171c3a2666f0b73991df7c5a1dae63dbf829515e642646276b47136889bc005d79b4688bf5514790f5d0c24351a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha1fa1c6528e4c8f204b4c161fdf34b660ab4cd25887e5c1ce20ca8bbb537cc8c3420444b94a0ba4282718353697ca67d848a7096a164cea06ed1840b2ea4394b08614e133526f1b7db7a9b7e94b216ad542b241812f764b74cdba0a8da06a51b84ed72f2ca0ff1ebfd84b8e14b205bd0a81d020b67a775a69cd6dc5eaf811523a5846d0e2053a95e2cf35bb0134488ffa104c21cbc25482ae78922dce5d6f02348b19438a2832cbd5831c0a5586ab5ab148d3bb3cb87592d9302c26ecf96933c49373ed88f0bbc28036f24dacd43927c888d05346fdf2281ee271139a6cc9af613186394e02387b12597c94428433705382e5be41f354870ce7e9ddb73a2c28e239e1f1a92a02a3336f5e02b75f404d6affbaf1b400c5219fdde00015c287fdab3491c114c57c6055a59fe8a8ffadc15d9066cbd73860ee1f749d39758552197f33726aa23e375b5816602cab5856255ebaf9ec61a888a4114098ca952034aa912a2d2461048721797f10ac96518d318768b85b25291763f9ebeb1d0f85a8e40fefcd36f4203254f70782e32ec96b71c19f455b428811285e18e6cdfe203b5fb83ea11e95c929bd51152b3f01f9697653d27740cb5bae831bacba4b085fd347b6b523e9b3c8ab9b93a203dcf8cf7023486f17b63224edd9663dc773e6bd2b925ff4ec672c09c719c3659c44a44a443ef769b51d1dfe76d9634a8dd2a6be8e8976786feb2ef3db970ae419848406437f254450bcb3e5da15eb51e244ac538a7bbc8cccf6b0753ed2615e4ae81cbe9c2a07d82bba9e9425134bb06997794b8e3e78203047d64f299f811cec59b2d6b801040774a44256ff7f40ea9790b189bd8d1384235c8a702b75fb7575e3bd90b0908baf1796fc253b09579f39f43365f83f70bbaba55a3658c220c5d20a3761b3db2a29aeac99b58b8d168fd2cc72d5114bfb5addfd32c60d599f090292e5cc4fb828380b2738d8a243ce78930dcd8f6d3f6e441377edd775762b4dc64e6ade1d82f65184c14b8d1e726dd33d4e9095ca53337b60b8fd8ff360970e29edd017c0dab40683084663279ea83948de9dd8d370a3bed824481c692316603827bea3bf02baef5942b3894524d18fa359f5e5843346c0deb9de1b13d3dbc9bc50ce132ea5ff2a59d77ff63b37ab34b4375463123e0764403a068518e88ec771c07e923dc45b0cae05e833519f63aee71aaa49077b83d0bf0d9c0cd33d0ebed72a4664cb17742453081b5659cd622c4962a50b432b71fa7dab23d0f988b54179dbc385e8b5025f734c7b02b0f6d81280895e3d8c498b78498362d639f8460eeced3bfb0eb23a087843ef27b3e963b96ae9a6e6ce7eba4209b55691ae35f3c9aa3731517314c492b4f5acea53e7943b067b422e69be6f243a8a70c2cd3cd1ee94f1f27c3477a23c01f1dc608e70bf4e0e1b14b41615b2d9462ebf5a8dc666cf36e7582ddc99f84c596a64f16c16c6608e75c9073f0587392a54cae609afa808b9496b19e0c543243f30c0469288e709b79cc50b8ac7d8d9471887cf49dedfa9972cedcffd8df89fa0bb498cecfaa75062ba9437e4b732ec394ff583fe0b54d644839c9af6d00fe065cd477c560244440a770cd8638cd2218f9a97acc15c8921b58ae8f4c42224bb3356bf5b22db40fb968d86def8569603d7b858f6742b26918eff6ddae34cb425fbcda84e490009679b70d3f45487c4c2362d390e01857d8a0e6fbe14ae7293281cac728bc77931fa97f715390fb75f67ebe9d6535f8e848b2c3c1be40f059a97a06c8f7d0d2a38665dcf685e5fdccaec80c4eb7191e1a90c5055d3631889a26091baf21bc08a825d8e85ed1e7308722eb7149369798cbc26156fdfc191939570fdd27c0080b556a798f73f64298fddf2b5bf09948da406f083e3f6eeb63b07692ffe4c5e589fea758528291f404faecac99bfcf4a757e7bb0ddb2f9bbf60cc212d83170b4a5ebed349789a8120d711c83b5ad75ea75c7d9794968181c3b42b15aced2118927f869999f0a9bcbf9edde7d789ca71435a165dd3157b48b75717a2e93ae289b2aa0290c4231480c2dc00e1ab591f7cdf6510ac1dc81ac6eaa62fdff0b9cfb87defb54ce39b30096e0f6c3b170c74a806d624eedd2baf6ca7fd6add2c1a80aefded1b85c01d95f167546b4d45b511eb621e6ce05041b0ca4a54e3e7775690e4f7e5babc24fc150fe5811a85aa592797896a203621968c4e0b0ae7d4bc3e455d5f9dad40f01407ed6d2794491cd8ca93f07d326956048bd7399e77af4d3bfb743c2d9f485c9d494abba9bce2f2f48cc1872e885a75f6e0eb612c4bcf7814f562dab33d10031291e2f87789f6274e6b4b8a238ddfd8d36e6ed6a3b43263c81880df363d0aef62fb014de02e610e1f50fd92df04ab675b50bccad0cdb317eccbcba3c98e0bcc4449e3165794b6fa86c0c10429689cff364ae3f0f3a7819b20ed19528ca9d510a872912d046b610fe75119a8e0cdd6e5e3fba74d94832cbe0cbf3dad2377097e05fdfee205b1ba661abb732ca1aaaba170c2788f3d7d68103c53353aceeb225e990b05fa5c1a3ba16d1bd0d74b85258d746fc20c5b9cea6a3d442999387f999a9097959668712d7900ba725c78704796ebcd3d5df231e96dabd518cb0366c3a25d4c1190ffd46363038256a635e6a33576fd5bdb058c4804de27c780f2ad46acaa3f2412d06c84ca00a46f022e9331183038fc422eed84b203c199c45ae572397e88b93fbe9dcf1ae1404208d29e59e7ba087cc970b82653843b3ba9adf99fb7ef6ab142943511fb45d885cb06139847bfae82f5a21c0129beb37a35256ca0d23316980567216d0f91f7c48245b0eb6a38c48519f8e1af52ae244fcc34364fe6c9908bb29bd4ff5742c50b6d253accf150fb1d4465fac35cedf69d5df733b198d4cb3dbd9d32ecfe399f7fdd16a96df5145807896d01ade4de32ef31b68406d860f1b5ea1ff7945efd62a135911cb3894acd0677af4a459338841aee5acf6528fcbcfef635d9000f5dfcc922d0a55482f1a3b77379a53bedf22e0bc4af3b6b0d32d717b44c12502b09958c8e4177b95f0cdcc3162f7bd7e41658c32cf98cae782bcf7b383a81e7b8fe4593bc195b6363f0785f0447c4c23bff701e42a646a58cd340272353d055e802bc1911d7dc5772d9fe9da827bc58bc9e6d20d377914d146c63a257c3ff95d4dd364e01cbb243a82e0d97d9ff64c724cc4a1eb62acb1a13b12f4ab9b3f6c69702bcc40eee344a0fc83e1c29827b08d6d1510a245bf21ae28a346c44a4aa0ef37413968cc78d35dd7163e6125ddc963f5b40fa286aee6860ee372207be968eabb8a04a44bd419418a74dbb5e2fb54887efc1c8e8803281249e5821ab281cb1b9a5e6b3d8446bfe2d3120f4450d6dc94a9aa55067fc38f5dcc3a6f411044c1fecfb9bad5228b4de446b8835f50629fe1a3eaf257f652745f20f10ad3a454ea6e0f31c803601a69365543017c6d3022a892cb1e1cb05b34176eef8782784bc5833e030fc16e27e695a23c05fa84b233f54bd4713d9615fa1af955fb9ece6d3dfe989561f718f3d15cd5ed970eddd95ccc1efa6557158b1f5c6aaa818ed2671e25ae55a6687a692e7bb8be0890ecad1f81561b8c25de2bf3f652903f3d95dbecfcf026a97362dcef450172752aa9c517a24f6aa37eff1161ea056e22a2f2357de46bc3001ba54c3ee81a5a9106c1738702f4c53cbf0397928c3de61ef9e871bd21d9cbce0974f81179536904bd4fa9d396e72652d6a649eb5cb1a6414167ba9cc76b71d0bc548da79fc66f290cc8354691e4575b8cc765130616194c65b9f96f434a89d091bfcc15d7e21e3c21139d88daae808a28b0e763ba7561c99cd6fe1ded2ed13452de1ae9c1a559355d28aaaba59ada180d40ab749224f701dbe6a3c00b782acc1d43df1ed9c6d411b58cdc7103e364d5ead8bc6ea8671babb3b8d43f5c30900499776b4905358d13d5489ed99f2bb6c156eac8d8908a3e1eb1d5f16db6bd4b6ae69b6eb34ef330e248905990932e78df4e3c864761092dd15f46c82b22a70c362603def2cf1403c2574e6915e695d5ccc60186ef4c947d441974ccda594c2e079408910656e24f0f9397b4b2d39fffdc72cb3ce01620f7de012d1905faf34936dbdab704350fa49d81e8c3a5d7b4c53b7bde86016acac5b3ef6fefac637385bb53b7724ce08e2f3387bb776feb28bf34de26dfa1f9e949ca3794207a6065eecec35134d51973c913cdc6f8ab9840617c6bbf5a722f3021b635ec1a76ffee02781611eadcf76f6d7ae4413fbb2767ae06458aaac9aefb1a33efc77264fdd2713ce0be5db5c6cbf675fde2ea1dc9fa7a6a2390dcdf1d99b9e37c73264c0638069545fad8b7be8c66f4ba078eb0bb216541bf2e060f9b8a125664f0a06d184f4b1acba1d8706617920c1dde04f5961d63186f7a92344bb9b7fce4f3656033cc71d92be48164603beb89c124dde6657c7578fd96e950c12e7c04624220001880eee857af2477deb03247528401599e8f57e8a9b53dc5c203240b8aa775ce352f843ed1cd9c026408a3db94fc2c683b472ceb6664ed1626325bed9b3e18319938f7f575d078f61d6ed6baf1c70cdb36c46d9ac03efe56f2c849b8a1127891946f46576f7ee38bc365133660035cbc5bb12f3342e1baf00301f6c721a7d37c079dbb67245f22af1c056880fa66e208827ea721f47a192763fd3b0c173a8a85900743d415e239f70b6dedcac58e43cef8b4b6d3000f5a6cf776df5c743340f3e15623ed8d0a76b4a8f7179bde45bd926a462a459db43c3c2acaf7b6b9b2f0c8e979ea7b66fc4bf5023a81cef7502194e8d9c4d6f218de0879f73b7764a54ea14b8243d82c260b706f392f317d819bf49284ee79fc7cc74804746a79ac3cea137d5cd77a15dd359d169530e3c8cf85d8dc2f96a8ee4e90c47ee215c2b7931de1f1f4b99deacafb89d0fce5772139efaeb9debf57ae8b945dea5a6f401f3d351bc08e93cdb237e7e2d39150a085ca946944e0df060015ab98c6163379635b4412d58e5961c18ecfb29382812adc19860b6a1a3f90481ed107da9cff77530a6d13f2b3a4956d2fe25fa968e22ddf3b69ce20070194d2df8993f6dfdd5509a2c90aac95eac6f3696126b255c8098305a5446e716d755f319018e6506bdd28bed14f7b9f328ea389e14064e86275d2ea3f115c3f2b7320ffd76cb2f02009592da8c0860cc39e787d37a844d059ec095780b228f4de8fc2df1b1569f769ef44edc9609d47659c0ab3f2b99c24f749aa737874be3a3337e73aff6ceb04139df32b61c62f0b54fae75dc8a65ad0b0676acb1b7e43376bc9974f9074a64140f8a0744f65887bc184e5a25b3dc8965b5ba84e73d943e9068b56c02e7e7224d197653eb7db77cee23e4ba38fa208a7f367caa90d1e1471111886a80e0921bd9a8c6e8c6112c725cbd94cce502e2dad3a88661f59;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h81cbaafb59d8d4d462af162c95ca6d2385281f2c500e83428260becbbc4efac1f66dd09ae246704b35145077cedabeffb89732ceac931e1eac4e7bddad9846de8479f69b198b3754b160573e1cb994ad2370f83cc3376e8f65ef1fd31bafb4de47413d929a01ae77d008460feaef0fff2bfa7d1424e7cda7d090390fcc536e1f42ee5c84676f447b999bfa31cf86939c8f558b54d8d3f6d63ee8b73552c9cdb78fe5a9596bbd5392972feb5ee6a8f9a67b43ecd3f872995cfff8ecc468c43be9329a3a16856400b29b763f944a9574a850797036f8a5739821b3ff5112bacc5e750313584f29c75d7f3b62b017597a3fc2ad1826e2b10c54a579dfc665e1489254508d104248840ba26ab8c34c26dfdfe7106680b0dc73007cd69e3d5ac9cec78ca71da50afbc8d10c34113e853df53f826a18e5a97e1a720fd6337b4da88f1d67287a03868667ca2f3049a8712faff805dce1d6ced427c22c048f601b6eede1c93e8fbef473469274641e9e0fbc13f9d463149c7b110c0af0a73163a9fddb102d8567e19eefb1af9a1337e99786bb6d75b5b15285a9374a7488e75deaf3db2c874217867d7118348918e175d3bef1d10b55da50a53541deab9bc4e75b9de8e50b741800545040cd5fbabad5783dfd7f8fc15af371c181cbd0483542aba0a173b7536bf43435c919699bb62e475d0a31e0197e444c18288a5ddb35afd8d917a4f070c00f385b86f78acb2bdd278d4a45eaef9181b88806a5242a068b51361cb320b2417602afb898a355510f38bb1900143629bea7486fef17644206a4ad308f4f3a9a747a1d0bd850777463f9312245a9f82c18b7a0f080e47f9f92a9f0615736a81426cb8af54e1d750a6f11cb294c4f5e7a32b5c87de7dbbe512bb8189c2f01142dcd7c517c436d526d5ee9c98b19d2077f3452b424fd14d2aa3b285bea5d083df936614322b09412b4f728b1e13af99c4ac65d57d17936886a5e73d6bab0df36e707a55d87e96d2c5285d0c3881fd941171d791c64f74a8ec4885013027aa737400c3f63669c183dd36fef20e2b6cb046b20b35258ff6305004b7d6d766cb885dc7354e4c1dd494271af2bb34a68a66675136cc77a5b3146cbca8af48336bf74c7fb959afa923a11020f3f9abd1aec8f500f1b7b55d905bd4dd40155caf9dadee7b9b5c74ccff1d76f8c171eb565a008c9f531c2cd20430a58ef1d4a9fa0b8dd9bea64fca4876a970b7ca7cf77168305e6a56f43250d8881f882eab3b3c254e47d7f113e3a00a5fe55dd62f99b225665dc97262829d028c461ba77533d7206e6d2f8af4088a53f4d72bdd578d55bc568f2c0cfe6b55f32aa9fb9ccaae097cc233e9769d38841852cb553da124eddbc25abe1a8dd78151f7047a55d9a3c13dc73c2006d6943b6e54666431f4d449f5570012ccbe14f9b4e9985b2b9adb4e8d3c3fc37871a4fe0afb87c4bdb034ae1bc37c2dd6017ad0455b0469aa1b820bbb4298d6e1998765e2329fe9be34c536348337844addc46cff6bb3826e4aa40cc5f51e93adb335fd3049ecb547e6ea9d83e61b3c8bbad8213b19127a6d0a6d7f81df21f43191e329389e5f2a06d572a5429821d46b03523e6d1e00ee767368d4e6f57cf32659cccbed89a1c528bd0081b7ca51335c2475c495dc1328f465194f50c5fa1cf77181a0b5318f19c23dc80e270690e9abaae80dca9ee5bd29922f9b811d85534cbe23977a6d599d25dff74c916bd0a409fa11b749791626bd2447b3cba83bc4a38a0ea814d6c7382b7dce17505bd1289d7d8c983c95a9f2a55d65e4ff11c8a42e699c96cb200696f1c3a5586b13584b6c21677d8d43dd8881b07cf8ed3d6209dfeb422eef3c625898b3a1c3fced41ebd9cbd817004510c7504d16b1175a5111fdac3b8a166bc9f78daaffd02c7b34ce423ce54468d30d20c9b55eeb5e2f14961c9c4f59561bbf92d12ca1bffe2c7b49aa68babf9d7cf7f697d0b346256a56fe3561e658825bec960181ee64f44c578750e5e5f227e188dc48ccd877e74d74b989f31ed5ddbe56d3fdb56feb635e10fa15e84e82cef174b8f04664a31970b32f1612cee7e03e56bc0ce0e58eb5b9a47a7e426eba32fd537ba86f7b489dd9ab6205b1ffa53a64f173c30ff1e15a64d2a21155b0855ea799523d51d13d973b31e70df9171b6c935bb460fc77c9103a164b3bc76a7a6e7c83dee05d238c7e37f82fee990c8befae1150fd1eab72185fe7e050a6cb75c5891d5c253c14228a5779c832b4e550989fe44690ba4353a7fb9e4cf23435c40d0e5642cb782d9b06136ec4337986079c9c7395c19356540dfabc9d537ac9f707d1da199db36cc6e7a46845f8ad078515daa9e7684670aceb9251e0f6c45f4026afcef55fb498c6e77b716462957ed8f050cc6f6388ffaac32951e5e983bfefaeb22ea0317ab9cf5c1ffe8e56874a7b2c81063e9ad1b5cf31ff2d56211ba8fe5e08a2de8bd77962c9181506d452b5fd9607ee5c04865b68cab22b1b7af99b6876db204a22bc72cb495efd500818164d3b03761c12fb21427409627a50a9a0b56da11f07fd99ae8414f02e59b9d5d71a4ab039f53a11e21c69b9833422b2059bf15a096ce5b4cd80482b5f760287423af0c51073f4028388a3ea1b21875f8cd226fc446ba75fb08e4cbb7f476a4156fa4e3059809882818517dfe77484be6ed4c634774ce7955d004ce1b4bdbc534c6932668522aad6edfa3098adb05465b74e25f3e48973c163769bae0b27b91926ae9759900571da0d1c67a328788da8e362aec9d77ca5da42d43b68d8c4ccd0892c2212cab2bf9e363f55e07946bf13abde0c83e14c5732153d83887e8868662d8935bbacde9bde8c5e66e570e3d949bea5c4491256c803fde263d2180a4ec6b6ba295d997e1e64011085ce8a9c55eeff4a8c834d2b5cc95ca352bdd02e80e4f67621b15d851c751960ab2c8733f615a706689077733caf8f2822c7d0bc603bfd792e4edda90cb40d0cda8f37943c2ee7d211da4b3bbeaa566ccaa7b483c804bcbade4d547ef01029491301a8761d77d7c5cff2328b957b287723cc1c40e812bc17d03f973d8e0fa0c260ef343ffea5db706cb590a551d0de8748a8bc4d2b576f81b76215eda4fff89aaa8375ba7b1affd7352167df1618e7212d309e8072d92c079e5cf68e63e245c05e536a0ab33e3f56869d817dedda6bf0b83aedc9ffeb36498c43b46831327e54a569d2ed10a79ba6ab24b154eec1ab08593a5542756e1a2fd60868c9a1c92f76ee53de3d1f5001e6b0e32448e432cc4bf4d39ac28753ce4fe6970b9715ce5414b7cecd1dec0110e81931f506f624fda01dd27a03aa39f911ff9caecfb90f4cee6a150ab36319b3b9fa7d2cb3f774a8b918d3ad19b2ec00d5f0737e7b91db494148f3997976d6eb335141c64b2370f2e4a3eedf67496d90bb106d4fcd34a7b34b8d33de5b558dc8c4ff896cc4bfa2ed429468abc8a4265559095268f3598f3ac72fd562bcc5bcc1bb38aa14c9f82b4a387d4768ac488f626871d229afc1bb2fbed2dd483f44576491149dc981cc7c94868cefa06ac01a527c06dea7d4f409abf18552726918fb5dd1b89197187f9efb9c39e77962112fd75a57d3a2128e3a2fdd1b70042ee83bfbf7431d21629bb22fa552065321731c8782fe46a4c286de04bb986c0e002cff87c65897ffe9125f47341aed13b54daddd58909648dddf2fb2c97189645a84133b22247137c7ff2948d960bacf5009c4bc8c96bd4726fb2f439e5b8ef54741427d0c2d75bc980147b7779ec26586c7a534477df55c4d92e677d6b9403670f5487fb72cd62aa0a62a79c094c30c67d800bb7ba2d93901a75ba0c61d6636ea64eddf7262ed8668aa4184442461b210df348a74262d400f49fb451b44ded8324b31960cd47afa32747a8064ae8bbe0f0fba665f3524f06213f8ca86f16154f48f088cb2055693e69bb97b608c53622c436fd6b5cfba28d838919745ee5272d73cd243ad90bd7763384c15344cb17e906b4a843dd36f71de843e31c9798e124ae74fe052cc2cfd93278166a94ca5e2449055e9d37d5c858645da7ce1b210527c230b69946430709113d855ebdc67a05dfa6c5e87aeda613c44339d50f0394a82f6027abbb6755da6c3040bd6a8866223aa56023577f0a0ba25ccb9675aba0f3b677fa4304db1a3bf7b4ae767042dd58da5971ba693b8fb70817a5de3e73785dd3e9d84ddaddd48edd2356eb63759dffac75706ce84edc336c233586b18a94f470dd73ad7ca6fab7cebb5595261f14fb023382b05d213ca606abad9d4f5a6fdd941dbf8ebb546ce9216dec6f4d67148b789bc393d90aea00b7e04d4cb7c13ea21310eb6a1b4a4a799aecbc8ee277858f5cd43be77f54a713aeda5c5361777a30cce69b8b99709f2bf1ec0d1541df0f5249984a89e26eb58243b32fa95526f08fcc6610f32e613977b689dcb032851070f1326f17e02460a8f83ba1d009817235398809135d37643ded493a266f2202b8be8e7320b2a180a90786b871877fa8db85aa1ded6e6a3ef3293808d39a985bf361dd4fa0376bf916ad0b5706d0388db2e9379301a8a771420b6d15a94f395206828347d1889ee5276518de8bc932409812db75d4cdb48adb5eb83e3edc8c325101976815b6e8352ef1a90c1eb7357260f44a14833f435be7d5c9862704c3ac153970c9ded6eb5118044aac2126316fbf6044bfc540b4804efb7b9b176590ad4937e2a2fa4af874174bb3354d8f14e85965e6c59493f84f15d6ea04dc1aa49e71b94baeaace3206654fc281d4e12a76448cfced5ed842658bf3994630437bb241dcc922f77a1802c2c756d0c62e6a8f30e7871d7585fb4660eed0bce590a250769e67acd163466d2a2d26483a65fc1d2ff41bc2d34076445079c4216c07bf9015d356a3776717b2884a298b1fa120095becf98354e771be4e1a07b0c2926d95b4e7e2c16f80c721eda8f9ac4e817d7bedc977cedc05d1b19c360b78254a61de919d86c07792744a8a2937dbaca05a823e9c7eb83c2c58b842310c70c5c900d9a4dcc184fe5af6ca7632a2e18eb9c12d1ce6740bb1116feddbc55130b198ef1962ac8bdd5da21544c64299c57f6ff71cdd5b9d03331d6a5d25acc07250f1d33da390ccde216b4eec37875a09f49a7292962a08e5e936aaff8fc7135a0c5b1ff0f7fd4968019d21315103ae6f3662632a8c043f8792498bd3e2d0cc28eda733724d3c5778f43711b3caa4a17e05ca5eae915609d16a959fd0b69b9f989011fee949b4b80c263621caaf870b0378b1aed88ea15edf27b33fd504deef41a66b4a797a8cbaa5c455eacf06b698df023dd6c7deebd7c166611ad18b0fff9b9a9c0afeb2eca364bb0aacdc85bc3c7c78edce465ca550688370181cc1e661ff3e98e93c66a178af40378bdc4ce60af6e1fbead659a568d05dcf0e7515c65eb36d91406218ae60b1fbd0ea41052078a2b9f9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h4c40cd1db23ae911b3154b1dc677bdf8e80d61e859609717410dc59cb9152fc508249d45c0f4ea4033071b34c45397737ffdef83ccd2c7441c63fcb3964c918fbca36ca880e9d7fbaa0a3a7afcad8024c1de8c22d8df893415f359e11a7508b4672215971738a84ec28a4bdc86a62501e7739f0ffad35001827d2ac25c1ae381b5ebf3cece6faa53296c98e7025826c4957f70eae515c0a777348b2db3dc37ef1d41179d736d26f2c228a76bb39d3ae990a27c599f8797797d5df0b7099017a3bd51dffbf6506b667f0be545bef6ea5559aaff531cbeadaf8a0730101624f7aba16acf30f7672c7c1c832ef9ec8ebf4adcbeb82aa38a55cf7741407dcceb58d20be07b70779337fc78633fc71d4465089587400800a5922fa44b0c9107091b828fa8500d9a34135ed74d3a31e3d6b2dd4b27fc551924ae761cfac7bb62816238c2527bc479fbc008f3f14be572bdf30134ccca9c36fa22b5c8d989f9910f3451b5c2cdee86374e4240ff9a2b25fdb47e6aac241a8e52ac4c8f9b419ba95e04eb5b713dc34a185af449115925627603cc97d86a55ff7b564fdb5af61701366573b204c675c463b1eade53447708d511b1060415ca4795a4c70bd38e61234c8c359d5a4dbe98c2a408bfc5fb9ed033f08bac91b477ccb24134218f779fe8e4b3991f2985a7e2ca7e09145e5c5ffb04195be530d2c4ab092312c3ad05506d3b31328f40b40114a65364602ea5436b06102899189f1b4528085e9f9592d640a063682c7db3cfb1a99d6b3074631e21cce5afbc4488de6c775c80f783decd8cf6267ab88fb2ae0633c002bb9579c83ecca2af5e7517375cee84ffb8d0c0c0aac5eeee84e1c32b3ee6ff2c42beda0ab9e312d46b036c7c2162ade663bc5d3bce7177afba276f010a1e82c2d2ec320e3418186bfbec69e0a64048d2f42d8fb73f736aeebc1739cd7a643ca28e1465a240c16bb1545e4bb827d5c76c1f8dcfe5b4f615e9c28f3975754cd843e263a32fec7db3c444c432339b9cd9f082a416689358d7de7d46da4d38bd0e11102690830f7fa0f164aee01b2eda505a2e1d35d089a751902254f88c34358d14278b9516f8651820ea98d0ad59e5cf02751a15cd8e9ae105bc341a148110dff9ed30b83e72c7c0591a82b04f3a94824a890d407f3a5bb105bdf1685f34ca0ce7514caa56a40e5b746b78ce9bd8e4950853b88a9cea4c2200eca59c2b2fefda56581ed312434274828280de7a871ff90bfc56e3877be6b0282eaee158da1d08aa102a5867ba4c090542f605a5618a184cbd53bf534467630e6b680c6a02f8ce141eff05365fd654655851a044f0b491f78d4946a7f92ebdfa77a2e46572aab781443d982151a46630e3ff00a9c038cc8361047a37abfc7c1a2c3d4cc0bc906248388eb50207989429387a08bdd0f3cae14e2a6773cf0bfc439a85636b5e29d9ccd74518f3b204036dd4bdfa850cce6396599a3d25efe5b513bb03707037692cc5ad134dc4ba0bd9a8b0db3ac2afa2a56a785145004f2612541fad9c586ab465e132d87783d9189cc92574312f79202f9058c402d12fbdbceba84e6389f425999473fe7f26aef82fa7bd2c5dd4515c46839f21d12a5d772d64537158eb86eb86bc3ac3640abb949b88b6acb29f7e1b9bc04cf0687d250939869491af4d4f41567679489b83bbf3e23ed80aad43a13dac07966c588e3c5eeba1a19477b1904111621edd06bd212b95da9f47f18561f5b506f93458d9a910b96b5888e9c48bdfe16ce461b346641fd880e302c8444d9c4e1744480687f72114832a698852c75dc80bf2a4668e7f504364827d77c312ac3e4e664258d20065e2f7fc739066c9dc4b565863f7727d71c411d20899f6514e572fcf8c0ed16f5f1139b2be14afa0c9d3a25fd4e9c42a2c5e4e8ade94afc1329accd584a8e7ae44df5068ed3fc5c933621f5c97546df8796060cab9916f3c8cafa8cd69d0539e9af24a8124c5079f10c1e802240231aea81cc0d07e98da4a14fe70ed624cd03e7571097e3227edd071dd96555859e9720330ee847b50f739fd78a71f3ee97786a1e1b37527d25080e42e79d8311b257327a97c8dc06740b56a13b10609a62e99c75c6045e1a680699c05d7209f436a69d1855e98cb0b3f00cd38d032dee913adbc7a77b05fe7502a3fd20bd3b9cb1f74676a2b0f4fde03aeffff055191dbfe4e4ce450b87ab3c031bda94d27c9668f97cbeeb39f475ca04055d67690c9985df3fc98541eb1666b141f16f6e3d19043e7b389aea8a96b977ad65405b151a5ce3249952e4770ea234f59f50a8ec721eda037135c8c02c67fec6367430592658cb8cb951718a41fa43bda0796fb42c7585c21e28be9d62f8b414c82b4d732c0dfb45e7618ea1b4ab2b41f15d298f1a2afebb6fa63130ee4260511bc7b47fa6e7bfa547b0b878d17fdb258a5aa718fc6d7fe996b6dce29536e4d8d2a4522500e2204df888c2277a59de1d6ab3abcf034346fd0593fde8ca00e9e4c98f75a79cd607024addb67b13829189fb4d49d37db1834efd65cbc53391e9baa2d45cd0ef4292ecfebd9f0ccb65b2a5d3eafcb52010181867697cc5a1c1dde933ca6049c4bba7c48fdd4d610ee11548c63c42881626273e9b0449bf478567e4a047384ee81a4beba9f5f44b35f069789800eefc5103f150a7fb30e613e7d6e95be3a7e824665405587c360dd19886419cc47f64267b70b29be9877d9371e4d3abc34f9343673a9ba1f9f7d0bd713d2519fb06f67c24b54b7e945f75f39fc4afde3b07bf6363a1ed9692436b2e6c0fd4977412bf035540275d85a47c02fde467a331c4ba3059138b85dceb739980f7673fec7ff635ef2f8946049e84a1bf0b9f7c2a11ce4e723e67cad64ee6e90733593834fe70e13dcc3e54101536adc738508515395d067bce166b1d4b3f5240c0b89241d52f0f19125cba7240226825b998739925734029ad1f5633afeb6ac58966ed77dd81e3480265d7fa3ac872ec1e665c6772a2a53544d61f3a02337c6c62fc97e0db448bfb0bb7e65443d94c9d0bb64f0a472458326abe1dc6b57116245bcd90b45e0182290f3706e169268952da6a6cf544d04c85e628ad3dad508ea54931d3102d3ef14162f8776a7fe959784dae7e69f9bf0f52d73df07c717fdbc3b8acde6924663891eded76a58d488e9f445f44cd83998771aa80bcb58b47d66a85a08c79e94541b48ed6411a27d1339bdf52655eceb3f5df01923883e87504e230b0624cca636b5b0580fa087e6ec1ab6f96cef195188cda136af0fce6ff7e96142e924bbae2f90bb2871852df73137ebaa6625da4b86e8928eb54ba3811f0c439384b592e6a92caac8cc9919baf0a9fd1d816a3972f1c3e1bf8fc0878f9f3c1f30eb2d3777176b260e73796b97fd24a4c28a389ae96762bc56d156ecbeb90c41aef1108ed63e770e637d087333de6c445c193cf7c6ce9e701c788749182f8a3a2aeefd38009d2e1a0deda9e611d8c0521488b39e25cd14dbff50b4f1560bb70debaf64956db922b9960fede957cb410cfc6af8f08548aec1f94a3c7878050cc973c9c32dd38042d7b6ade02272cf1ddb0e25419a38c4465545b22b5fe7fbb5d0b89107ce647c397f12256168970e7f48c9466032de9f55369d82e7539b90b0300ed248e1c75f636655c295d42bb5c400f7844dc4a598d8be9a14ffa72eb2c568935e3af6d940bd728a0c2caf330b10e794e652d446a67299ed84f4bc2fc40bca8cd6f272be92af1147b329a6e54da797fe78d554b3b60388758289a16cdb2525c0997d98d6699f0b3db60a1740cfcc86ee9a3c2cf03b647956704369945fba7060f504b551e0faef38bb5c56717f0778dcebe9ed67f52acb423de8c415b024a60c0951b111c34d535733f4045ba6cdb63eb46ee7e94714f23543d21a674bd677a348f614b39d7b1cc84b6f5560cb9ce40191980b8b3d24f81fb76a6d6e8d4a75354bdb1791fa6f9867fc307eec29f351bcdbec0c7291603cecf1831d38569890a9248713a01bed2e6750cca16dc57242830d3681841ed331f80f994eaa903e796abd1a35731d5873e4c3aaaa07cbe7a5dddac7249f081cf801e13919ca57880b20c4728ec263bce74dc56ca9c45109502c770785ced2959b1ca3b161105c4cd6e554af8b7a194e166d885e46360f23ddd02523c52fbb763e1b672d7e52cda447ece0e82ceaeac30e43300c041e314431a50efe7e374e9cda40d80953f5dd40e6ccf8a9c5769b65776343de429c63f76005a7e20816fd62d3e1b7ab1101a9693ba79c41d0f743388a901958bddcb1a6a5876712822b17538b9b6c4cabd50ae72d7f7b6dc0989a83c7b8dae0c1973655b59e5ee68d995449e306884251b5030ef11cc5a1bd85c0f8f262fd9465a3d28c0626a4009bc6f384b9c5aae69fb7d1e4cda8f905a155d1d31b2b3d93fe600d79baf03a89b3d61d898b6586c8e17c18e713bd640cc2c9fc34b0f992a97f535473fb0ae7c6d6da6a964f3819ed2e940305db451e53dbd46f958a35d2a11b5f67951aec7702278e5f91becffc65f70c3c6b9e795bde75513a3ad1d70a2069a27c4ddcfddf810a0c5be6f43207fea6a9a601b425efe54ee8e1b66c01ad6263ae03b29f9c341d302565d6ab3c44942c14d300970feab660ad87843a9dea538befc33f127d3caaddf05e55d8769cd2f634811dd05955bb13b21884040f5442a81af2abdeaea3ebc182515fb109f4e3fc6b75f54f58f370cd4da8a721e500af501bf17dee0e815df01eb222a467a2ea41053ef28064b1173a2c0e5169caa2c9de016835c563a7eb16d8cf14257279bd0137a5efab23f173f9d8efce329a741d30baf209a327883dc6ab4aed27d2502d73ae7e230de8215496d96032c732ae5df6bb120b99a3b65eca5e3f254b62145878d45edd84582c91f65d2f85de87689123f19cc331bf5bd4270a62e8c77b6575e9909b47fb3bb3525c5f068ae428a1251f824ce2e9d5e2b52419ebb31899b2d84e0eff1ac4f8a079a43ac4bb78e3d1c9aa7bed5c34f9a29be713efaa82334799ab754d9e847c969f4b79119729daaa738ef5bbacdd6122af2d9ca7a1f4fa15807a5ef28551fbc7a1fb0378284a9632ea574a59d86f4b88aaf1cc0752df32d23c2aaf1fbc0bebff473b427dded5bfab588bba5b04f8721f7e69566bd7482b0ef93cbd2cb231539d02a36aa8df121be99c772c297e63af934783286577fae055e8472c099bb48da25db316eea4b5d024f151aff49d9c5383baa4306c06801b45972bec8c1b7f62dc13709ae0aad8d150abfb34fa29dc0b5087991d9e39dd0896c3b362a4637fd5d8f5506b233e96f8fb267682bf98c8dccffe2eec873c2739e592805793b7659b240cd020e9e211d69b19af50ec3a5876317caace257f595b6ab400e013571ade21e0a02d370aad51bcf8eb062d70e5d61236b0b27d21266e71e785392a499ffe296243d47c861c02d2685b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h8323547d51587f7a83892c8dcdfbb7206b5072362abfd4c3f6b9235b1c1432ed22a947a0cdf97005a199d5bd44478f2185c6f3adcf9288dee061d0ade9210340dddc54aaa31002ef273ab4607ca6c1f2a1be76392c426e63dd0cd61b00e0b8809ab5328badf2ffaf12f321611713d64e1bc597a462c73b1dd41b6df3fb10b7a1c2dd5923997250ffbfeac207a7574598f8837ab7634285d7976213aaf93588cef06f0e7dbadcdf190baaa5f0acf53ae2ad9724991b22dc2cbae7ba5da0a1f697e03197c349ad945fe4a61f09d39c76d0fa6d58a2d3abb387b10414112323553fdb6609a3b54ca3f56f28bd26cee2b622e6804f6e7f740cea8fb7839247e2a732bb85d21535b3dc545616e44926951901ff74fbc7979f686aa7726801b2d0a1cbec45bbd3198bf399e930838fb2c02843107b2cfb309c47ab221cb7ba49b996b8271641cd4bb3d9011809eaf3a811fd6208888ea2eb0a31335cfaec7acea743b84adb82955014aa48f43e42014c57cd7848b3a426954ebe482c77de7393e3bf70d0e5e67dc42cc49afcd1c7deadea3c2f9b08b999957957ba987f71e5cf8bc47d06bee23ce97c1e1e7ab60f7218153c43e603bab4cb7a932fa1760059c581cd723b9d07f8cccddf3982763bc9de9b4086e5f87d69f656d096cd605eaccd6c5b42f03077a879bcf877ca792c823f2e9e282be4c57e8360d54e577b377e03a6866ad6050299d9b1728fd9d4cb043462c0d17a13b05d9f5fc6b1dadec00722f41d7e0d3718b948e43b9b9429ed7e8727d7bbcff3bd5a9f0b0a19a4afb389965557accc74ba1ebcc2226d0cc00ea3274d678f37ddd2d662f25bc6e2c8c64312f3b7a2a8673cac6701a42ea957753f6c3fa0fa16277b5cf309d362c5436a75cb6906753929c1113c8045ac41ab6fc3a1ad1af97235e2c2842565439724231f5f171270ae892f1961fc28bbf860e42eb0380d9126f81e093c137ac8c8c84bd77d7e0414f6b77c0782e94801fe2657d3bb0d375ddbc7cf6c5e64c18ec8e0b10c71e52db719d1747d3f4c5fbedf91fa904e4a49646e9f9329e99ec88ce50a10bfbb8d357280120904b485e5ffe10af2a27975f22a917ee76f0b53cd434dd34eec04b47fc89249190797e3e1e15856c976d426beabf69d762c48723b000d57d30a84c6bacd0526edf0d1ea1277acbd5e5c0791c427f8a0a080b6ca1ce11bc882b8ee8a3ccf77142e43996008cdb331d9a3d9587d5037a7366dfb8b927dac714be1239cbce8d572a9da8b2c3ccc78ef75790882b0b9ac1655edee3e9c932fbefa6cae219f8a621e51a22302e938f41cb5bd2411a50a96156171e23314e28d39d0f9f966147114f827bc27ccacd29bdd436265a065aa7400c8d10f9e253852d154b1643ceb5ab18c541065cefa881518f9efeceedb59ec6ddfe0bd6e8dc29c394764b69ad37e3800cf64554f227e5f30f2ceb7eb6bf73ff47c3b3c13761429249f0e8699b09daebcf7f6b70460fc2dba55912d6fde02163445b8afce668d0101941cbbf8edee45c13bca1d7cf8e02b033955d752a330e00d01dca5d7cb33108a6f267d8d12f53bc04f7cb357fdf58e4f3b64f1ac756973935dc135eada77ccd81a399cea17fa1dd0dca4c629f67c98e3b2e85ff74a273f2fec3cf71323b92672d597c6857e3736a4e36990cce636d063be88a3cd687eca601102650245410597d5f8ddd27fb4af1f4d6347be07fd8d53bf1c69bc3ef62ebe401535acb8b5265a97581966e8aefc9594535135b8fbcdd8b23a860281a2588e575c1cc176c0e7bfec0aeefc4cb9b431fd05461d7562e65612d6091a4f49e4ef07a870f2d258e3b5ca215ababff4c703fd1e019002a9f33e2cc44cabc3c83af519c216702a52f3a300fb3cbfe2247d1e6c2eaff7be07e1ca7b894a133ca1ff78ccf3aa08cc29f3e21073fc4384ae8c9830540b3ed506efcb0f121efc97e5e69b080ecb2d6a62a0ec7e0ac3f96eef78181664329c0c7621497962e68f5976aa6751af352b01ac6af7203ac748acb6902202d781ee810abd63d6e9873b018b2130ddc5126bde932f1a0bdb7bb9a42308cc33c82d1daabf79b85634e9a5bfc8b5ecec1edfff59634faf850242b0a33994f3e0804015007fef4189a5236c575f71c7718bcda35c12058f541a0b98ba077b46a1f6b0bb3635955c2b94cccba5fc8d5a46bcca885d694bbf12fcfbad250e654777748d77899630cffb464399948fae407b707842730c0eab1f946f35a51718dee52884e4df6dcf27a3187a2cbd9287103b8812dc8ac3b2e2d39eda0c36c30c746d4eaafa2c5612ef0e9e45ed7247c8ee69cac18cfebc616ec7596fb4894cfa388f4da336a4f94629d29821292469b1ec5644b3f56b7ad7bfc9951b819900b497702e2e5b09d23778ef69f4ba48382ba4163d12169abc3c0ae728389c8bd051edc49e5c735b646966c58a3dbdcab4e9c3b90b0ca4170f14f734730697197ffa169b5da59b244fa9a2ba66277ce395c9ec2337129864bab5c17fc445c9e712cbb4c067fe79e28c51129659a02b714ac66fc7d674e481d9b65e4e0e5101ea19e35ef0650f48d52c95563d213b424ae885bccc20fa009707dd4ec910f85945995aac08e3a6627dc7b8c232570ca37bde0226811068b796dca89538f1358eda9953de251d45a98aec0d1c687fb7cdf44578baf27484678be248bbd6a198f42098d387ac658e275fac2252a7d5ae68db261d146d60d90ed478e9c40449c1f8549f95c1654cfe4904fbc2aa08f633bee3fc925d77246fa9b4079658e1b6d3303996219172fe514cf4de766ab21e35418c80a99849c0302b34ecda04bd74c398e86704b7e453f706c60a7c2927bfd9e1f275abaa7eab28dde476b20bb35ea4f41140d7da841e98a4944f5cdde44ec57e01fc3af7ba3057bb31b0a47e1a3009ca54146bca58c34fb220b7849df206c5b7d05e61dd1aa1024ee6fc7d57613b84bd20142182fe6147cb38f75d5fd350dfdb17d9dc4c85f4a766c58b288f32e66167dbe3dc66b4516f52beb260a21aa9125e4fa053719b07a2d715d25abfc6655c2d33275ed5288553d22adcdc57e12c0359df66752fc471ebe10f5a89c7222a3341115de9db472d58707ac942c9c3e926578a1200fe753f63190f51951ea7392a852f7f72a57b23f6c6f16ca682bbf741c6e08d802c5a36be6f093eff085ecf0a10ffae2b540cdfc52fa48d4aeb2cac28df485a2e0813d293fd32e0d26f2415906ddba093164d0657bc5b85355c8c59b83033c205e10f4aa95be0d93edcaaf4491e4928945ceff87ae589da5b16f682b707b1a8f1dd512ef142e8cfae0a6d2df90441d37321c6baedef912d5c73e2d3cce95026b0bf810bc66d6d9f454050548b1525221726ea5b684251721889772ae59e3fa5d8b7a02c12a461e9bd3a52cace12d50a7b76cd7e83ee0053c69e0294bcc2203753ce6781f35c6f0dc7aa37bec0e50ed366b7db8472d62037d2f440d8c03965ded3a7b09c500161e89993c6eb1eacc0e02e88e02a19cda39579d5cf5ddd000d93e0dbdfa4fe8f4838c7907ad2a701efc81aa561259d32d635bb4af65d05c6630be26ed0796c4e103bf597fe4ca985ec4cf9fc58982b6eae2a24f5ee814e44ab84a37f714d78a15b7d49c368415734de5636f5267ff28811b8c475b6dd5306c25af8145007407774be2fb6302362233d280b3f8a161c6b4741206e939da42d2a533ea2d795b39572680023a8f051bb611042c80b97c04ee7c87e6f179de7702b96271ed0e98b2f4cef32989fe19acf9c77644c6e57a212a1da4f39913aa06ed4c4f303d08323c7aa9056cc9f32effcaf8eaf79b7d885c3c02008d14a1e7f29fac5647c88c29733804c966c7b2e4b7c199082860ebe43effe990ba2d3a534ef92a2839baffd8b869ec3c5fc5520f48f763cfea4117873131540f01695ca58a277e3902e565b244c93df566ddd35b94785e1867e91a3a3735291517d4c9dce6e04f4038d42eded8866077313277e4802f3830e53cff0b353a83b117bf8dc61c3926840ac940fcddc38725f953d734bd284716522eede6a9b9ea91317d676f9c0d3f3338f4a16c5ef4b0634e8310169ca8d1117cb3a1c0378edfcb11f927ff43539e110d53905636999a755c860b3469106c3bdfcb2b0414790afccdbccf28c8ff571a72924a9d451f86efec6ff432c202566c3ec4c882edbd4cfdc936a012c8ed99d822248738c6e96f9f1ce8387736b99d2770833e96d1deb6901e6c777c35a6e2d9184f10006b4efae95198fa224a84f48a8b41a685408c8f8aec12cef936ea78cbcca37f32c1a27b28768b61c27e4b2bd9015847562d055aae535f927a34922a92615c609c7b68469120d8ec751963707198db6ca559865c717ae3361b4ccf2c9ac1c898868fea2c205b17ea7f7149fef6425465704444354e4333e1d720b7dd60d8ddf2ff3b89e4687d104749363f7fd3baf8db0199821a048652bc97a90c66d7d1d6160366a50eb8a5accb19385d206194090be788ff87f54b760dc3e2ba530b0f67fa60c7dd026531d6b83ec0fcb7a29ffe6d530f420ea380df56a547fe9d3abe7e73b28d108276a9ba8a080e089ff39d46925c78eabbf27ffc3f6441d1bb409c5bf4933ff085454381c384b2480cf6913e2de1d8edfd714744a0d1b4be2ab0a34eb6c79df85b83a3d4e43ff540f1152352c61897552e41092872d7a29606e0c23211eb8d2bc60f787f0a6fc3a2785bb476b70b122963c2f87e917ac9950ee19ea2b50b94c5d9ed27a4a3b0a12289a361ef400e8d614e3c31ef1557daf2f09570d030d87e3f511d6891f4e583095b7e64d70ee58738e750f326ed7afc5cd95c7bb14b13ddfa826de45f31ca5e6ed10a1acd91b62e5aa71b2eb8104ee75f7d842448ffbbb239aceac9df07c07730356126c3ad9961fb8b1c5e572b0c9aacfc520c9869afdf6cc629bfbffdf7e1bc7a4afbe997ec003e461e7191b3e8169ce07efd8612f26161c4bc662e345a93a065b3ca8b8b71e15f72089a2f91b6b750810eb3dd6149f89fc5377405479e69866e0b3b6eecc53d2f112e078933c6ba2e147e83f6fedf2303580fc5995c265c7137356889df2b44372fd59f20252bda285594c23dc505a92aae40ff3bd0f50585262a4b55749cf68bbd55a01d979fac82783ac4db819ffa5b14911406dac4a171df1e8468b25ac47eafca025555d380a6a402f863cf27c817c10a13a1152ceb5d6299f111f2e6af3831a176e65e292a334a808459e2e467ccecfd0af9ec794c047a1e23497570602b144c40638d1ebb0234ae68b07b0eb37a4d6875ebb3bc0af75cbd978757200ba5cec800989b9a0d5171a424aae7e8e13863765b10ffc28c72e901e74a10767b1edc74ed14d9f32a72b79c2fae0b7f602750f2752af6cfb2128e2f1a6c3f43bd7fd5acf89e620254696de0609e1411e27bc13a7bee9ac1c403eafc202d5a15f254a24d877e734066b0ebc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h59edb9136f5081baee3a0875e038fbfa7c3f9d983d3c57a4ee24d83f13532d9c330363c8b26fd95fe5c45391260d7dfd85e441605eff53340749a43e889e6d36fe67522bdba529cf8c700b61bb1aaad0bd1a44818d8442f4cf69639ed4254d4ab093dc7f365da6b513369351938084bbcdfccd96cc599221e40f74d202d68e10287d7c74c9a335916ad8164731f0c510ccb793f4ce5f83bbd1e2e6cf98e19aeb6441a00d559c555d6fc3ee34d0990dc3602720bded5354f3b0cfdb6afc7a3949ace685009f0b5891ef57ca07158b02eec095c9fcfd8045d34225189b1cc1c0c9d705ebd40e9dbea185bc2dd246cd5c127f05760cdcdc694a41faafe7f7363a09a90922103f17de117691fb7df0555b0170ac9840a4c9c132fe5fcc210bcffb97bcbd138cdfa21161a13b791957e9b5baf73a12f7ded8ffe40d3600d97aec2bc7719742a32401cebb02782cfc80bc2bffff9d46d268ecb631ba707b5b4817954bedbac3fb100e2d595e77eee8b2f014654bc6a31c9307d5503240d5ecd1f8a398663510ba95f5ef741579669890c56871075580ac4ec453003ae48fe104560edf131039684ca440c9679e20a640c28eb6d3de2de28afe2b5c887e253fa0183a9e8f5c6528bc1f88f4e68c6d5d4caa9860b346646b4e0c72799bb9fa891316e25108f4b2720804a623ce27d4a0a069670758c8d2beedb48d1ffbe36f8781e4a5132cbcb6f770880d59d8fcbe9264d56de85588126f66f0a7b55129f223b29f51844f0fee3c36ecbe21dcd0ae561c220dd52a890df706e56d0f6518ce0a109c77f52e2c205fdb0e039fde2eddae785c7e9b686262f4f2016eb4912b37a4f0d6a8d6186915db8f96a862f10667dc341e26663dd082ad606d0f20b2c88a63f87568fd1cc1d0caf916b71277b6f36a56f46f1ce74eb4f88f541c8254360cf7e1804c42fa010640a319c41ae67eca7c6d6feab29654b4b29bb93ceb1844593b8bfe4aa5ce99ed391264db7c0cebf55f0658b89e687d384f895a0d5182bec4ee991119ad3b430c4640c95af6b1bbbb5b43055e94fa4e415d3df3cfc022edd40f64faa473bd4ff197cd98f84337542bfd680d43856e9f348681cb87fa8a93605d12dda8dedd4832bc71478bb5f8e1859ee43848a6430c8b2f09748233ceaaa581c4ece603a430847c185596f49efa2319e1bc2f2191bded1087957063b2c79dd82d1a410349987ffac1f4fa1466f0ca86edd7ced46df284b9172eb1e49d5cb909112cdf8811a400cdebf0fb4d6e6cd5ad48a7e3c345863cdae8c89e2f5553e154c512322aaf3d9a8fe7b258d4b8719c9d4d30293a82bd53ee24c7d728fbc9644aff1414c789fd58e215958df4def34554cb1719127e4e9a9a43a424aa860b4005056bda8d732a1bc0a25ebe6a2244286b0e748b17d2faf29f31e2cc60afdefa2dac2633e1d4c39bb643cae6c7d58b2b80eac598909010d5e3d3638aa906d39828a3ff69501fc63a1afccc2401948221d630e8cdd4de4dea6d66b069bf43a1cab35de42ee4fc3dd64612eaf419ee17345a67701205a02fed53f952a9e6235f84266d5f3daf752793219600384dea9b7193786b001c088f636083a49683aa840ca50cbbe35c173c542425bdc62eee2c1ebd0a5d2ac082699732ed26606c81d40b2b6e84ae74d76cf6e3fdf213f6b83ebd6918c54dac543880856e9c07c5349afa2003895b0f9da7eb6b0b952c45697f98cb799bda7c876495765f1a66329390a1b04db13f3c34c4abf7a6cf3046974587ba15a714dba726c1d39cf7d42fefa6a16debc9f0f0a4141e800190c014eaec5ff6045346d7ac5b3ba05b10499e258659d0ace6a1abc91f553a5ddbb84607448297208ce280f9f7a8360cbeae732179116d15951732ecb74e5e1e5767ad8f2967acec1fc42533a0ad77838b45043796ee8889e1a8312465f668df8312f450c185be3a82162ef5820ee2556a01c624c5e50ee15a0d42e95378739e1558aa9ebe95d354bf361d18466344a29ae6b4fba1650e97ca5e1fe4ff12d2172720a86108fa5f40d2e9255c23508c6588c8e60f2e6c2d339ac95c210071280768c9b38e2046a1e2e2a6fcd53c167b02be04b77a862fbcb39ab4cf0f37f0ad7d087758abe2d593bd7dcb7497493f0619b33f46e478d3c9c049bfbd49bbda4c8b2c3568d721ea5ec667193e1f477ceb3e039d99a020a4ad97047cb457a77f4d907c25fc9a6d98d5ef2440582787a605e32e522548d0ef041c595665c4f333cd24e928fe815130147a6a0fb728c064beeb2773238b82712f74d439234acbc3a8d9681da943590f105f3a12f5572223a7b368d8e011d0a6611aa278161e86abafe85a9833daf6310bebbd80d3b2424fc6d2c7e092a096f74d09aa25c716abf2529473c00f77d2649ccb14950c46e5a2e007bcb6623a2679d7423c4b0244669e05edccd14f4f6c8482572c2b63f081f177c4f783b4e9bc8210c67e228567ae7ae49ec0c353c14e7d316caf1fad3ff3a151161b829cd8f2b7972227d9fbddec3904e9229507db951ea472c72ec94363b71134a9ca2e39401df7f884ea8a0df2153e2000dc470016b5aea24f2514c687863bb95ad67d147104b88a5406057c65fd5d790ce0b02aa28b1b62ce0dbf902d0dd73930af4de75e3d7c58e5ee2be7298a6c67523256e77416a561aa807069084eaa2b0edc79467b842d084a46390ad79ece34afe6966a68a61aa281bf90a4c56c34c6c47c59b44149b6ee860f0311b3d7d295a33dea675118d7ea2be3b886a2ca826ff5005e4b7502ed837bce1a7e09424ef86f1b2ce2055e490aa058569e6e02ae8236c91c6988f80be78fc3eddfb5945c87567e9432a6c6e950e6dc94e28e0303ca24100e972faf042be97d73e1928f4c992c785c1319a855cbc674e1a28ab8105f775707ebbc018af9e473de3ca17711dffd3849e6b9c54f08ed6039fbadef1ff55c57a6d485fd500abf3c5788eace9ffbe21c7f72352b13557a5fe97d9546f859996eafdcbdbeb450b2173f587ef52137225ad57ae064b49af5117f3d5468821f1b5f56ce32b42c609e187846e9af53d407399a3255903e403aed15b924570bd39336b8999b0b82876db569e991eda35f437ea0e6ff7a85eb4d0bb10babf83e4c6cfbf7fe259072ce1e8edae44ad81fe21f31d25e0ad9e4b126bc79816693850d9c71bb8e013590c5ce00590b9ae7e2a394ee9c28bf82a374fdf14cb67b788d4787363823cec6677d3dc4906316d07b2be951df61e551fb60cce5e3df9a4a2fc6e35a7ce0c4387c00aa220ce63f4020663070269a7a800ea8fa7eb723a2ee917f66a1aaf36a019ff10c82ddc18de82a2b62d4d9ec48c37d084e4c2c8a724411babfa464d407e53ccb863579b64f8c9ef29d8e29032033019f7cc658afde1fe1db3d744e62a704544a6c6c3c4b08161a47a6ffbd2e9f62d024d9eaaa23934d686d9d637a3eaadd077cadb6e19dd96eee3541d40ff02b7428bb9e534e94fc2cba711158f46f36342e7765414f4bbe4fd7f61493db3ba29181fd2026a9a0fdd069f663b284c0994eb4cedb80596bd6756d11ff148dd0beaba312d96a9319c50bcf4de7d31117d564952a93047d17499a0d8e1542eaf3c7e6d369936ac550b6c2135da7a31b795e96a4e4d9fa87894f18469bec097264bb98beabe604693fe0211b3e4cfbc97079ff11bedcae3081aab54582a0a6bb37e13f8a75e3ad1585b57962d83ac717e7908bbdbf47ce2440b7eba59a217e26ed4f462f1afdcefecfd7d429aaf7bc5a6f61e35a7baed63887e7de6e812e8c8baf25c4330d511c970542d0f5bc673c35aa5a989c33b87c5a78b1672713c3225e5f22e103cc44787c50d6999897b21cdd5be1c28e8abf8037fc73e8f76ce0fbd36748cbc7c5d98b98ecd136571c13817c4b90c4e0792da924ac174f017c6d5762fc07b01f10123dac030d3b7002d509cedc5fb0464a05ff39fb1dabfc45755b62eeeac5203a8c4569560cc89a3b78a43bf640d6da102e16564641d310c865a6455e118a3e7a07e14c45c4ee4af9ec04e2ebd7f4a3062f0f70ead3b44be3aad9d2dd127f27db0f29066ede9cae65562d04e89ac8acba146888c83d92d80489b0186054456ca2c47c353b510466879d94c4046856675b3b3cf59a6642c077d50457b58a5ead516a81af68192c91fd605d2c1184f0d4ccfa402e05598e16ab9c9f1f0c2b67cf83ee38597e8c451aeb3f557c0fd27f592cfabf78cca6f1f473a1c985d5b5b3085ab00fedd11bff8ea241a680bf252bb55357949bc312a16a9f55370a41150220301e81ca33779e729a74b95628e25c4fc7e9cada0e6c47cadd2e3122b593fcd4bfe6cc60564d07ba27c16d8a7644428115f463ba6f6deafc7f98e9884f38413053c7010e838264c1c45c4261f5fb5d9245e536429f0f2a984bb71243797a9145f9cfcc4e89879915f64894a0dc97cb7c6d7d2f6fadd7f616746da601c25113b419fcb5456863b86289d7563baf60c16d8fe10e9c20a7817e74336912bcf0da20b9b303f3f22c3aa2764c53657f7ef481e19d7daf9b9b97a3654854cd8e38d81dcf6f22a986cc4ad7a6cac51165b7171acd6b613898578572b36e205fdbdab2b88fc1d97a9ed0f7547e5cd9501f6c4f4be31bdf09e51b2aae9c87f7e5f12ac3a6c8463041bf8520971ddd0f4af7d05c36b092b08702fe09528096056ade52bbe558e020e15bda7ae4060420953dd9c12be2e7931f313a054772d29475d620d79cbd6c8135095245e714ab951bc7a6377f9d59f1fd724ea8e2bf3f6cb804846fa8e692b816912cf8670254839a14ad29202db452f0bcda4361ec5804424c57d523a016d626e5ec98c1e161bb4fa98d4e807b65b369c32ad8c2deac9a6a5d5d52bc13ac655ce69f57ec0f8575f85885d4fe3bf2434ed88a401b2206c7126b9699169c7f290b26ac526deaf7ce608ae50269b9b6ef807398299590c088241acf88bd99a96d612a5a9a8907587af9e7f773b664d4ea9440568bb7872acee18b8238ce27e5369e97c825cd4552e41e22b10415d3996088ce4f0a3ed8ced3bcd99155853a81411f3368e75d93b4509efa9b5f57c806fe8b0f43c598831c4122ea515a06bb61aa5f41c93364b8052eb59990de27a0d91f52b60f82f729794a95739008018df55ce206725f2577dddf34998de7181dca1c94b672cef225908a59d02ab8c15d4ad12653e8d5670e65a91a08294aff967f19749eb870d413864a48ca6fcb0b7932aaa6f387d3f4110e0ac2fdeacb43ed947affa3f795aa29b4e788a36d167ee3664ac1b7f6cd8aad999c588d07c4812943056c6aac395d354a5270dc22404670ce7728607873b66ecd4a2253c84c30978971cf7c0337db536e698f945af7a6e9a07ec51b8b2c5393ce66be4e5c7967fb8537e6efc41fabfba78a8ec5b8b2985aaa6552d861d55d82c7190beccb1cabb2856bb60002638f533bab600f83b555f893379e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h4bdb8eae1ecd26da000db276c7cf56cb999ea6aaed1b70288a169ed0774353e3d256482e87b14acb451628edca9dfdd04f6f3894d871d2bb9a4e19698fd904a175cf0bc50cb63fdefe0a270fb490f30ac294cfc9b3385f72529494ea0071ec524fc387d9679f8d26288b7fa389d0e1827f8a2f9284a538538558dc55128192ce76a43175c7bc5ac571aed59234f9cd444a0cfceaa7a7462c204b8ad893120dc0ff8faec73e37f62e19212ab4425a27553a699417c054206cb1e4b9b18538c8aac5a8979a7b305b0b0689491ee32f001147493b498305638a437c15b55d4a481cf064f95ec01f4ec9c5c9c0917fb7395488b648b739f15ed3a437c97f608e3b2d371c18c26e9a484b8766b35d705056848b8342eafe17fa3e6f3a7c84abc7039b1099783b305d3340e06741b0de94baabac485ea1fd39a7d2254b9321c34efc419051aa31f1df1d8625664cf4848c6142ba669d57a6730e7b3fb41fe2da8c6c81c40fc1e934e6b4d82b558bfb7ece6c94d5d25eec57a0c4c0281a7d8764bc8ec9ec3e64a7c65a0f24c97b69aa82964d2bf8282d10238cf3c99d0d2b8e2fab7df5fecfe827cb2c79da2307e246c7b5a1a0cd0b5e323948c23e49705575605eedf1f55f5b8caed1f30a8ad320b79182f2f9f990ae31a5e2e064961222cbfc7421ae3f0bfce9cca9ac902e316dfad68347cb4b38a91599e9cb5dceb09a4e49452adb1b26c6dfedddfb4923c8c4d1204007e7cc0e78c5b2399658ecd8b57b0696c6a9f28f7e9344a18431ee84615f51ba19d84ecccd5449d0d81308de87c1aab9ff03169e13fae61c20e6a26126214d2f888db459926bbffc794cded23786346536f08c08fb3ac489c375450db9ce22cb69fb4b029538bf6a328e4240e929cc09c3ef533609c1115bc2d27319b7c60b9d4d3b5c20ec7a585c6c375b092de78e2d2e77a0141028dc2396b7b3aad321ec3da554ba8b8d8024c24403aba685c72843187eeeba64aef1421ae986134b54545bfcb38e8b62ccaacdf94cba2263b17d90770e492ecc3715fe3f0abd8243f561080e7055b5a37929c09a1bc884f04aaf78f14ec1ffce709dbc9bc4fe11c953528ff8c6c2eb5f9acb8146a06a40f21dd5577a81dfb6d4d013ec324dede22a2719cd774f6ba74aa08adbf4e7fb5a4e671f15107d10f51d46adc6d7b977516ef9d3f18031bc478261196248e988b2891b41c1cd810482c665171a93375a14f12b22082ee2c3578b370a87929e76baf2297496a153b119aa4da494fa328b9263595f4144963a56869f66306591f51f238d933500ea0575ba0a0a04178ed603c8c303cad0a94d042f33ee077e6934bfc6865358625d04f8b5c04c3627b16662e1f6a22a8daa5915685c09bbc856faaedde8e81bcdebdc5cd1cc4a969875c21578f9c496b3bf64e285c1721185e8f7f02c911c3bb34d9deceee1f78612aa7b33f2d363ef465aec571f68927ff0f31c9a2cd41884ae5952b28fe46c24ef166f690ebf1755243e3a6b904025c38b132d6502a42cfc4b3721afc04b6a762ba8d406bff343ca0c439929fc6adff4c2cbc5770576d31e3713a35617da789bfa479b4dfc4a183b5404868ce0a5fa7f3ee072d11291f0ad267d6da12a18fec98fd8c899c02d9155f32dbf73fe5c471b55929d15318856927b68d861c1ed93796bbd9dee6a7c91ba6edd59a13038201d8af71e8c7a571ae8c129e029b8136caede1d19e82f2c02bbf01da465a649cb919a6cf016bdf284c7e71e1c88200810d4f656007ae5ae601ed000568523c08557487aa5c3f0b63a3d8370eac6fba9eab9680fcf9b4581ec29e125001837becdae56960778ee4b30cb80bbea98efb62ff58e1d56b34f1b1d5559335b9d2c11c708e34e5233ca775bd4facfa6af3760665ad1b44657631a3a4e21805117f94d2842128c23599a6384f48c432ad033480efbc2cf109279b12af75f70bf3c6eff66ad5713243a4a6134aef9fcf60ba8d4d22a02a71fab36da9d3f8ed42284df79c243a835de5ccfa3dc34f11a023577b13288a1f8fa6b55312c6fa372057262a65b8d175fb852baed8d7c4a08b0c5658d8e88fd70b5096c2b45ea8f4d06ab774de6d3cc8770d3cb2ecbc0e5b43dd41b36fab352b8028cad2dfe07a18653bf5e03840e7a07661a018517f02432a497e5d7e58e25025afed7f0c69c917b6f9a0a46a77806dd8ce5645e2c083ec2c0992cdb556863a65c2828ab8b074703f4435552cd25b4e5d0296ecfc081faad5d1238f9058a6f9ffcd04ae4df7fa6fcd2d6d8b50b45178e9e1c365ec253ca7140f3d6f0dfcaa051416b17ab33e6af2e117d89ec5db5df12d15986cfcc5de86e26dafe9884afcba7fdccfd631e1eeaf0cc86b99dccbabeec2f6ef8589d19e9e69f329409cc88678b2aba9de28d713585fe2cf060a64b95d8a6469dd9ea08a99cf3154cc44deb82094efb7e4f8ab98e7b1b72e1ba821de641715595ba5bfda675630f9be84d6d72c54428f50fa3194062e3dddfd8fc08513e9f7b5c82d56b4d3430d555c83f55626ecc58a5efe4589868d6117069a5a65f47d04d5bee81aa0e79f4f01bd6d0947402c4b8560fe82a4531ec2fd8a9bf07598c3054f9504081fea3372773e04d1d9ea44b075514f807866ea093388bb0a31e25eea51eefd8c214c7521d1edb6e0c3c0e376b3116223827ac2edeb1e4e773e9f1391b5fe04bb0a2f44f6cb79d2cf239c1e95842935ba93251961240f16af9307d4a7235e8ced13a3b682321f7641aaf93831b0a36942da99b45e34042da77b628772b88b34349c0cbd0f544491bba12cffd6054bc53aa22320333a784724b78b746cc855fe962a7eceabdac6e5190ffdaa3cecc5a49a91264526ebef847f85be2a2c89170d2d2a506801a318911b2532ec7437cb0f1d4671bf7dd81d4990e40d59e8b734de93ef8bb65547bb41bd4726bfc0b09dc60ba7e8a6009c61e4e3a9dfc827b57c674be871b6ccaf0f1b0f2227f2218ee5b3c03b5573d4d95c8733c80f46114488b2f60d0ff770dd2a2a520e7154ef71e5a0e5927c19ef62869ffbefb5f6ef86d81221f456c61ebbfd4543dad2df5213855f2c72329a471a35e5db705355089e2546e0172f559c06a15e0bddf6c91df6022796f30f22dbc75c1f0bd23a1e1e46c0fdcd3183bf6f3af1186fdefa3cc440bcf899283d4232f7860f1b4a167efa018fb2cdbf3241f790fd42f9d40b0a21e8590b45a9de73c23097331a6487368c573a6d2d8459f97b950f1bde6e3a25f65b7b9b4fafd55b6acd2353479f8a5324444f6864c3f59bf6873dbc1d0ea8df08271d5dc62981df5d33791f29543426b7fc57aa3cfe0ff2f4449a5c518aaafbe725591dc758296d7e8aca336e8fdb9ec1dd0ba97993f6ada834f7243e9de442c844174fa4dd157ca90ef14f368f66066563ac9b79940eb87ee34edf064a7ef4a8decd19eddf17d174d2404aa212feb858585e2ab218aba6a46ff3bfc6514f9149a1c7bc1f9a76134986b21368c835842558b448e88c40c2fc5bab66573ed8c38c20fd45f7db40b066158ea071b09f3505661e6cb1d8b0742ae6f0161b1c3ff97e99555eb9d227cc89e4b14a1451f4fae184f665b0e80fce10857967604eaf8c4c4a2eb5e8e07a1290fc30cb77d4073034819a50a6c1c7c2fe6238911cdb4286f68c67e0ff5b81acbc37330fbb1d27c2f636da8719d620f91a70ad450663eb21d5c3b54e76347687583fdfb0d3abf6525a5f33942ac59a74ef7475cf688180e4ca336c6140cd29b943b4cbc3fdd3f0d870ef5efd0c2e2a1faa562e6c836a00a6024706ac800ab9eff25e45233c626f4a89972098fd0a7fc70e8c83821f610567047b6bba3ad62e189b9d9c3a157f3f785bf0265270f74b842a89ee257180b7529426bea7693a13b7b355342bdddb53687fa00a5722cdbd7083ab3007cae538a53a86c8c7531598da4a01922480e6d89d38e5c78f8e25114a776368c9c5b5c5ca0373921e611d0d4f43a75945e1ad8cccc7cbda9d5394e068974decfb2b57daf3ffb3b3c3b292104ce3b407c84d52866f1affe690e5e680b0bca1a675002e1934c438ca7274125f6b9b52b0a236db3003cbf9ded8ac0a0c6b977cd809847be14e0fd74c109162943ab0dac8d1328f2cf8dcbc421f1990464a2eaf1d653ec3a44c4ae91f20985b024e6f25beebb89989efcbedb636638d5d03596596270b1e4a37cb51eb7df24a1502164093a8658361b6c75d1fb89799b574e13bd5b99f76ee3c19f9ce1ac1602b40bf4103afdb589d179ea0727512d19f931018286fe40cb952eb891a275f2a18e5ea54b9ebcacb9e24525f840a510308383ef1ee4564b6886b1f06d459ade4f44c45044756ef4e1709db28b30a8841d5fbf7406b8135c89d6bf3bf449327411e2431e72198b425273592bb41d7786d5d3cc60de43e845b196236e22ad07f04d8b9e62b3a33bfdaf5e53a6a9534afcc2e0fcbab646a74b590fbd945f4a71eae4249a790a107b6cad6e4bab048529ea56aeeff5978f89b1b5e0ada3a39026f8163a83eab91dbedf0083ddab904f682acadd7931b3c084f2e1fbc809505457cf45bbde9038afbe437ecc7538ac4ea68e7753dbc2c95fb0b64b860594dc285595d665a8e3a4b373e5443004604b3b7a1c76dd0f8a4bca7240b42874a484d24fdd46d87f1e60f585512051db976864e3b3f9313cc1f1fe7f731f0aded90ce1b2d98e511e36652ba2d4f7f4de45d76a4a244fd9b5b014512f8ce955e509d82942651f81195034c33c645072d0726a83c9268da3b151fb214b690def27b24b9a99b6904cb8e58b455469a252010884cfdd40b41a7708ba8bdbf04972c0a10307846c966b8c477601daf99339ae2770a750dd7f0635ecd6dc4bf60628b7fa2c2179532e9b99eaa5a1eae81ab4589642f5dea2bec871327e4a305dedb5c6f0ccd758102e47ea906a71f434eaac8c665b066d7f609c6ad1d7dbcbdd674f6a6ddba3a48de3d47d5fd3712c30b1d1d2d4dab6d266c3a8167beed43e9e9714bd6cb7edd72588ddb53839f2be51afbe4914ad9d357308ac8d43f62bee2db525c83698a429d215dd4870a67332fcc10723493f282e5af4155dfc89fa840c629b9a9b3936f4bc2c47837d902c124455defacaa25f12c4ca0cd85784153eb73f979a2f32a5996d13a0e17a44b54fd76740e92098ed28c09a001f88bd8ec97945b433681c0cc30b288bf31c5da1690ece2dd8395d81053a3fd23cb9fa67a1e6c8310aa3bbd3688c414c5dc0b1234b914422d83d699fe489a5cba344832ddba874ea87a565189e4a5a07c1edacf80fdc20be577be69bed4706d08043f2576ba269173f5fed76c94da55b7ad0b5058dd8e05ba292028e96f4885d381ad1890a9431d756857213b2f31d5d0a9140741ef9266357923fbe0c66e5fc13477cc3c273ee17836f5bc86c35482abe349ca1e0db69f2adafa12b5b7eeed6ce0cd40559c66e6fb9f96f58adc3b1d0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hc71edb6823c965af98a024859926cd9964a3fe6e8d75eb89e0020fec2a338ac5582b2bb0e840cb561c24e8eae674ff92da170ac368588034dedf67a4a212cbb6abcaf96dfdd1ee86fd81fdd59333a87c7e00ef1a95c4d9050085c08608be83231cee0ac736a7cac165fb6081b4b539865a3505acbdf9d56dd3a7cbbf9af25a7584fb96135ff7357a705a4c21c10d984d86f95cc640da3297e05af7feac27a39ff281602599e0962d3b0a2ccfdedfaf0b2ce17230791bebb88b68bc51218c6627e33440508246d45acc869f758bf8b1522f5f92d4d46aded1c5ecd7fb0753aa41bba1851e03d586d7615b59f0445e7db145cce384e94e757751634a32fd3d07fd428e58c0efa28c209fcd052011b3443942c50014b8cb17180988957a21133dd5113977d0f2eb3bf57720865fff69f50024a0cbf4fb7d2d9f9cf4f542ded8095d83bc32ab196ca18ba30b8d66e302c38366557b0dc1d7a4bf9ff525fa2429ae83f6f563b463c329d8935b1903e9ad62675468ffa733f977bfeba6e359db3ddd423e43baf11841e8bc6c5ea9f7094829888b3d89b2a155ad36cd5d268f5c459d8f9c09beb0f76ef78297e46c87f0fbc02183213c1a134f4f7acab3d3fbd47fb011ae55caf9ddaff8ce63f30ca1f0455cf67824f711724226dac7842920fec330a6b77602d6833912110b84b5fb0e543afb3a93f01727331f986223423f4b2055db278553a2ed03166eb87748d6f20797437c01f3969698da13bdb7a7eaa75df301337bd8906d7ac8b232e48b67b21838995319bf007826a7ea7d44ae7965b2fda9f262665c231ca34a1f742739f128fcd6c74b09baf5d83e894833738b07a32fbc783bcef6b99bd2c0e4884adf35e95889ee03cccc201b6661476f850e56da90fed77fbba92d18e32911e0e29abf8da9e39272c0af45d9fdfc231c6521b91b7573732332ccce66a4ffd47bd3c42c076803941071e883132911a0cd84871bd6da7dd1f666153f82e789c0925023f6e4ff4c77ecd2b34e5dafe5722a1c084797380b9e91c355e0703e5f1f038b9ae036ad35b0be99e089522fad7fac03083f14454d372b70144ca360dd1d2421ffb8df212a290815c01d4a1d9c84abaad7736388c16f3e58a7c24e00e27ab8796d626c0c02329f76883b90e07311c4ae458bbcc1086388a4ca465deac0afa12807376844af370fc1d0684a535659555f1edde449c8a3e2269d851ad03a317955bb6413de4f872d930421fe4e984f88c87bd77d99f1ab2d747626326df3d808ea08a84aa8c8d42e35420ba040b819c54722d2caac3cd75922b89af03532fcc6a90f3c7753c3caa37379ae8191dd3d2cf0658161270823bfea9747ae6bff2c26e76c71f989cfb40f79ab0fe6d7d67a179ab05b01eb57965e894d4cef310d7618c63b71bf9367cda5ab63911d5d336fe835ded1d9e4f574675e81245906d8a1fc360e3acc424d025cb5ee6e493fc8586bd89604c3876880e68c8169474c79eb840757980fa341685d995f3ef09f6ab34bd7ef8ab0c577cdd4b96b478274837a3857975c36ecddb6ca55594fa5628d49860d5ee24281eda7aa56134d4d3478d561c23559e10ddb1ae79f1a6086832e5d78b5acf025eaa631297dca59a7d30c0d5dece506e3c6c625975873cbf8bc080579f30d8ae2e284c3183a60b852f36801661355de9114d56a2582343bb3d7a8ee2743e7677ce3503c304633c5dbf175cd37b37c7f27551b2ecea6ffe4ad41b3fd48268527311e9369eaa29f8a1e4ec4cd07b24a52dab11a6f04a28bd8453631e6b7462e61281c95bc87eacd6120a66109cd1370ee335815e55c169eebdc291a15ae945cdd61275926f4c0969953b8142fa1028fd0453e1adc6a674709326d7645ea3ad2d45ff2f973971124567fa2986cdde90f366abcd40346e7eaace1e8a8304bc61ccfb4c3a3146e9b6b19c42f19b9704fa4628e4997118dc0e83d9567e8daf5daa6810b9943a50d425128fc133aaee67aeed4c6113e0a2c8ef2451ccd7404b9f638011d63bcb59fa15004376d68c5b47f6f1de082c04146b9f8dd79e6da74d31bf513291c8a4f1bc7087092b1c87da8ae7fcb4c476a8f2ec488c50e5a3459cc1514fac8aac3276f9680b37cb7c2151003f9be983b698a54e4a165af24538b5ebc74bb609fdab9749b39ed0cf4ecb9fe22878a27ac219c9132bb434b450a6ef6bf12c03cde31396e3fbd92916f411dcfab4e6b919bfb62b203a2abca8eba606c39c39adc0313de2eead7e1c5f67abbf7f6a71071df5f031e4ee1d1f45be64cec52f64be44fdd81bd31ba20785e24991283940a07d863317c25a92a610a2b3284051ea2c32b9e6f0f83098d5c9f98aa244e2e7443376f99aeb0278b3b323f5809875ada15142b31bdbe2d96d2ec7eebb1839f7e5ce83b1b0186d68a0403ee46f5486f103652f8aa272105a57861553a2eb6fe118b324b27d305759fea4b8a60e450202171ca6f27de589d260c46914fd6ebb3618fcc5e088bd52b5eddc84cc8feff0a7327f07fff91002a50c83a83869dc47daa478bbcd95bc512fcc829a5bc325e87cf99be07e39a6a0e543187f9cddbb199e852eba34a1cbd7a39af1a251f1b8ce921b019e5d8cd4c52e920d94fab2115b1f5f32b5af27632ff5870bb7243a1e1c0ecbf4d9b33b06263febd477f4ce0f0b726e5e417b12e2316fe1fdbb287dca5171c1609e8fb270d5e0d60c92e28e1a14133212ba6e1c02e068c2f7349aef4efdd4a7d2d04bf8281db1f805b73e43efa1ca97cbfea175b6fdcafa6ebb578b43e10de8a3c9bab93af817ab1114c96dddd301b008ae24bd8b6c67dae8dc4d9358f1198f4c0e2bdf3a1ca75aa5acc4f1605d06c509c5377bdcc24f0467589b8d531f2923ab98cf2fc7fc969c2ba6ba932f7fcc7d750ab728daf8ecd8317a4c553cb3fa3fc8d19b741894ae6dd1944ecaef44d7c1f8f0d13597b91f3258b8a535c407cfc15ffeb3ee91a9ae382e076c0b3e25e21339013425c68b4f8c5f2c68cc772733fc8666e90ea277593f533ac66f05d2d4d0f7b843a5925d0e9fc96702e12e73f13147b6e85456d5a859f77dc8eb1d09ab542bfa24ce25d50d73fd5c90e6b16065efce7c44b57ca3514d67376f754bc8d9dd85b7ee628036773a9460d7465074ad5aec018184628ce9aae890f8d7166e2c88effaa7729e0a7e8b89b5599e09565cb2e595498684394faaf958970aff17edd35dcfe0bc858ee54f004d103f7b1492dedec88ea611b5f65be2f583a755f68dea16d891f183416b8a82e5b240704700b90e5f745ec93d8f664f8127986a1c92aaef2489b16d0dbaf4f54ffd1169f2757080a5f6ac82d5dcbc192eabd0be0f25e2a1b0bc03e2e3d1346463b4562e576548a56cfc145bc81eb9ddbd4148f4b725b92733f0bd185922e5909132d1b1afd9b0d2bffe18ed7ec6333a501df7b2e8094aa7dbb0693e7ff8dda60fa43d0adb7436cf4a159d6c366b298099b09628d3e65c983eaa9cbffff00f8600551a7a10a945804fc4c5dbaad2e3b90670f35554a9b4d72d1c7a4570f54355cda532ccba4e47ff8455782045c19b754c3ea00e9432f9e6f4a8707e8e756a7a1b47d19b17ab69be8e934e75d8d3284bb957a3f6d17af2ddb435ccd7ffdb235f8afef9cbf8519e3f311e912e6804e4219860ef31e30f83c78d9a264331dbb7634fe92d73a576ecdbf15c1fa8691e7795b1775ea527eb0b2997f40a1951ac1cca0619ec40ee2c4cfc13c9e61bb303abc530adf88f161fa823394b2aa33eb650e6580fb67ca70343ea186e94d02929943acb1276b03fc1c143d787c6066ee99cd8ea4fa6c7fea3661bcb30e475e80b0d0d3751a09caabc05d4335c34d8e096257a58bf8c590b0c9a4d640fa4129adcbdfcb3c9a00239f8d74f8fda47da514e543ae0ac5b506c52e39a2c2e02c96fc995393607ebdca46f4fdfd0b7ea333c425a53682fde598cd25242a652b58876f1db2e607561223bf153ead4030279c442405f61b3d6ac0df7308a99bbbdd5c33842f4873378e49fdc7a78f2d84a216e01903b3e0f8682215f8e96b4b1deb64b0c7f9fae403967f2cbe8521d820fdbbbc42519fa4eb1544378ee25e5846be46b43198006fd242cbedbee1a141434f97912d9cf7c74862cef5ac8bca75515bbcf80c5a861e08165d45dac5350ec12342bd0ecb2a72e1eb6c34741a5af931aad3505842d92df02004f1b4d173c21fbddcf1d90b6035f52f3251d3fe80e6005af2ab2f0ce5a1378f07583a469ad9b03c490b3a2725ccb697d48cafc3190f2ac83fb9cb70c4e9df3fab60fb03dbcc27351905410f8ad840970817bae4894397d915f83991e9517c17e3723e18ad26fc7ba6d706560d33829a187465d1221abdacc8ce238ad4e9de7ff13f007ba5914aba443a6298d4d31619a6e679aec5d7b4804552bdde10102a5864c84ee7edb0cac0837ba7fce6f9d581d3f15e8fd29573460f129d9753d3582f2aaca1b482fdafa38bfa8b49bfbfa014f320e1d1812216c382af62949f9d745d23e64a1d5ede9ad03de976bc08df35b64c02786d922e80fc4ed46c5d6b4412545d88990f2a81b86db77d67dd71af4d9ae4389e44a952250498a1d23ff8121139f9c4dd0265183274b6174c8747dd36de3d637016d61fc4dad16a058747ab2f5f395203cfe054e59568d22c701771b426082d0930f4dc9e2b1aa7ec3cffb001146a1c86f81dfe84763bc03dcdb9532db37582bf20a0ea7a21c071fab44b03d3845a1d947b03ffe5c50130241ea8c5edd0581d565619a6ae09bef46f5d97ed5af6428dfe80efe38a78bb6fee0c5d5de1558e05fdcfeb407a98f6d283c35491720dc2e0cd3acbfec072cb37da37c44d887cfb4d93e396c55a21ef772dc561f5e408e9b1b35c70ef2a8ddf621706fe99903d63ad4866e0f19ddff5334b26e558838adfb3bbb160227bf6e83be427a3ad0db96d89490d4a3d7cc9f7511d6028bfef6fb0667c41e8d4eef0adecddfeebd30d60424f056f9952454e4b967dc86d3489cd938da4d8ab4618501e720b4db26929750f7721175f2e79c02cc5562f10e7c35a3d4f66de76cc3d3c417960c4b082d87663dec2cb7bce87224f1bf91c51be4e8b18791c7e2fdcf229757863b8743c5847f83c9a15beab46cbd63188efc656fb73b664fd0445b2d4b96ae531ae6ab967753e7a0f439e88965eb9f20c7d800047e0244cfb453ee50c0698dad6378cfcc4857a49abe08baabc2f7f4bac05139eb937ea7e4c094a23507cb03095cbd9ecf19c517a573ef498a7ed4563c6650882b4b54f10fa12b155fd3d6f0ac0db395566cb9fe12d90bfd9016521dbefb23b74b0e322a080f04e4b8e6c5f130232ddf6230090e083ffe938771f7d1c6aa75eba52bb0f0dbca34f740c68e1d032366f8636ea3a887598b6e543158d0256ef13af94d6f212d6c58c78c19e0548b3f4c62408bca398a8108282126892f323171afc0b8343615a0b4b61;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h1f588b9400a4087d45b3dc6ff5a6d630cd6c2d25caeea598b5a499613a3585b7ef369ceb2462826807abef664b54f8242caa8ff53ab18a5574f9c347685eebbb5550ac82f01749a21bab9ff82b4701c79fc9a6caccec1b5b9f788a7521c7aac1418d69f18e7a4eeafc60b222755c162a3044b565683c6888ad43083a898d5c4c17f30b207c3cfb7f802552a586deec0119edb672836ea941dc55149509c31b056a3aff143796d8e246e1909d4794eba0aca63ad5d4c787c4756ef5d3daf66b436d2ba88060896760faf33c05dbcdde2256aa2856adfc0c0e33d670607fb9fa4b7c0dfaf82b2b76f437c1bd2d12f7276d64b66fa2b4048edbb4d0ce7ce20b2210c81d12d09f29363ba038e26450deacd05ae172612404a289ad3df75e08a9b3fa9942d45fa366b9b3845631996eda89cb67278e1750cb00ecb2d05faa4d510af8a530ad32c16d3a62045ac6f3f018910e7f45657dee30928a8c439dacd4933f30b814d7a0a46c8656eeb07449e51740db69afb87ef1e91420578abfde9b0dec3ec8d39aadd040164fdf944ed7208b382d5edad0e1b044929413595d94588dae9088d3a5a8af1efba696d476b5c0f762ef02bb14e17eea84ad3cbafb18bf6e9856fdd680327dadd3563715c862ad4a99fe487444bb49b4781c54d6ee0194c3037aadef065220ca631bab66f5764839162e3dcffff72dc1d6ad40ab437d5aa2c6484081a2b15b9bc96a66510a39d048a81490f255ca8bfb1ce2eb4bf2e52f812ef9b4a56e3419ceb68f0c6727e2d7661f92a8ecf94eb2a7c08eff679084003bbe4f099d2f25934ad4a3c9156c430ef3aa36dea6d84553a2f9de43e1649df7d58756e4c4b8d5777b1a3e498e1479e429125c856ad738b270f5c168ea9a29fd12a23ba15e37daca182802abf6d46a2473d7832abd9558f9a30d877bde135f1e91c76cfa69713a31a12aeb6e497d5b7d5d2d20c36eba0098a60f52950caa82be090f92b2fd64ab18f644b3653ee8f23b4832c1c01912d9c84816349da9fda84b0ca513a53ffd2ba35dd7878bf311f8a14003f259b638218584300fb5367f0be3b6b52ba4607d11a2b683cd3df3cb915e2f7db5a634a5b43772e3327f3f1c06c4b7e5ba35f63b2f04abf71a12ece03b77cff31286cc17443a206c5d557792021f83f5239236450d9d9b0c7a487e7382608664f706516e28814268586b414d75685ce5c326999354096b278bd485adeca9080d367f8eef173a7df99754d4940619db409bd08b80c3c68bdac350100c472c7a9571286767cc1597af577e5f90686f8dd864d187c134fd7cb1af7268f36cd689468a3bbfdc74eb5f7f6595edbdd5b53db6c646a7596f72414a675049b5cb5d30054d0df8caab5b1388f749c6a36cc1791380c2e668bfb73cb5605ff540e6285e0a67d20daed3e8d6df151a08bcaa00c9ccdd4150a193e18f02dc67644b4579474a8f9111cc5e0b24980a0077cbb471a5819f54fa8e7d74e72e9781e2618a18b1ae3584bf3ea69dd8c5a0ff1ff1542a478d7349cb6f12b8f10b6db4f3becb411f1e8804820099e14516be6e9a70a24ab0f6157c7842ec330f52ee647c5992a5d7a4da19882ce69b6b0fa9cbff75c9cc3084ae42511f6c463c5f20d36e9f81800b900458ec01099e1da71938a73e024b9e5a865f04fb05cf42d0fdcdb45e0408c45fd7bf516342c8279e2f3feb3087522172e990f585d17f8b7bad634b78810c51348e8fca01ce2e5e42c9df1a88255f867c63d209471290b07915c3603a594d9bd15b115cd80ffc5f1c7b11992a5f86f54eb7a7a8d7c196d2af6701ae93e9cd76022a4f18b0da0a097ad492dbbd33fcbd8f82d4c2994f846096c81a7ee712f22f7c741658503fa11e7564be9e174d8f33d68ea26b951052198726ad7303dd264680d98981159341d9375d86eb26ceb3b1d3ff884805fd67cc1fb01bc7d95eb7cf9117480e0a79c4811b5c1988e3f2f563e98dc1833b9494e86ba555595c6f4d0ed8fe7f3657a1cf9ba9721d13353b1560054bd19e6efda6847418ab7a06315199de809db42ac801fd7a6c9100a5d458905c89f253b24b1c2b4c69cfd9e301f4cd9d58768add49402b49981340277ef6f1aff8e62f52d46add6a41f19a4b85f9629aaa03bcc15815b044f0b4d4c3f9ca6ad2ad2340cf8fd28ba3e212f2edd5f539675c43a8acee1a5e0f854585a3fc2ccf60b27174417ffccd3420800e13f13e620c67733ede91ee2802e3ac61db2e74b0c98cae287f1bd215a2bfb6f1ba570f3d27721edbf6ea0f024b9c70efbb2f63893984c76494a7b5ecc49fc1f479019b757ab61718b65ceb4980effaceee92e33339774e4ee4bf81bde201b2977164239f7fb7648b6479e9f62a3c519bb4c622fd49f3075f4f3167acdbcf4e3d93112f456d5e429a914e79f1088f58623565a62a995cca4e1fe59b68349b0bcbfef1a214037d11633c9d27fee674f82fd0e0f3ce82825183e9778b8fd486e8c4801cdbe23b43fb2fa68bc051b4bf333cc780e7cb64477d520dae26482822627f4d113579d57f934e5a168a4163f075ae47fcf31ff0bcbdcb1e850cc077739ac1a49743b25669857962cdc15d281ebe715519836c8219ef5506d8632bc13aa42d8a379affc8faaa9ad51d237eeabef6d02fff71becac09ce28358e52a24192f85b180369e1b738b35b3c45b5236cd5ea4cf2d4df83464692b07684d5ff28829401f9116f2f2c4424a8c7b8bf658f428edf4c75df68bc528083d53b1c98b979d76ca72d7d6ad73c7bf4e7c493bb06b94678efafb6245107e7f2398dd1c78b4177acece3c496d8abe68d04c0ca3f449c1e3ed18caf8099c603b54384eb564e7d5d0c2fef852e5ecb637c07173d285967ead8889048cff64ca931b3fb6f38c12b4f11999206ffacf99cf60892bcf9c9c491b8a390e56b70e60e225e563798f9ec0cf660ece253ecb2684fdead4f16170ed02175cba8ba4b6bdd369b5a604cbfe33599aef56a436fc92ddb9c98a6d6c5ea48ff1d843f44cb1adeaa4bc3d84571e2392922d385a58d54d02636b0446ff61a5a51ebc9874957d86ee997931b4deb9d8af205fbb421dfef6884b6aad0c9a2050da039dbfa57937dd1fcadfd854b047842f2be84e512de83e76a4aa1d7d81fed09c59f19f1ca060793a5c143ccd7488416287f4b4f784eb1bab4478dabcf69f8b8cb58b1f76047333f9beba41bf2484ed7bbb8ed175acc30c6d0f0deaa4509ac6f754a9f16130f3c7aad7c6094b4e1cba1fecf55efa145c3af541ca97f1cee66f24d4570419fed56da5a4d04df8d35c39a6f210c741913211d71b0b7e25698c32d783c2b11fad2b6c085c0889a75abb583cc8db0c8e61e6c0249132c30a69b1fc18fc57b199051e66d541a1081f8f1e171a2c36a02da26ba4e7db5ac70772bb5267bceba40797d4ce7b5c2609105e5ed6e790441fa8c56ec7f1a672759016b1e363ae93b5985bdf1a92ee7d0161c88eb40a2be919ffbe52acaa142ef86cf16d5dbd46a636c880695262de9a6e5b07e75dd47c39f05bfee4b4f09bd06f3bf52dd7d2346ce7259bd5a724f11f58601977cf9c0c5983284ce7b1b70f13c8d8cab80f49312b377309f3c9a9388ec343fc0099edd96d7e53b8582d7689106c4b1288c538920b8763530f85dbefbf08f5ab9b2059bb3df717ae617ec9d93229ff0bc651647e3fc68de4b450f7057b50bd2f704f8884dc5dcd549e99033960e2cd51fc8c27f2144bc08af68aea5eb53ec0bb560130bbe03f89395f90ddaa1d18e7c40a9d833272a87ab2867c4bfa769cad4e944f7f4575cce540b3b80dbb9740deed479aa344f81fd487dc9dab538c0efcf9717b9156ba9f666f1144cd6bf6c62f09453fa7a4f8ac5a38a7a31c66c035fd0b05b7bff4f6c331b2af76efb8b15d96519cb114cfa5a9e51cab6bd03a9eee2e8bcc274753d1f544863c974b7db643858c50698a929c8344c40af6198f9fd72470ac6f2d368fdb7f5d110486459f1807c00b0e361326b2c5a0923880798b8636f19f54ca997c9b2f27f5d507682283a969a6e19871987ba2a4a6ff73fedb8c6a41d22b78b0d932f419c89e12f870625557b1135fef39b2882277b6628d9a8ae5feec59fefa8ef34a145a12aa5090956078743d945a6e649afeb9198058ef0bf54f64866b922a542b7760ea15582b31246635265ef8cf2c2a028306cd5706c39eebd3ea1349655f1bedf688aa446b7d798f5c8a9c2b068262fac0b40fe242b7fee59ef7e8fb9a3bc48cba7afc55b36795b87865e4f89543a7781f5e5db425efdb0d35af9444489212aca66f33452fcb04a32f5055186a962996599aeedd8fdcdfcb8d9c9070fe2b9659b526d3ece77d596663078bdb6234cd360c05095e6d5fdd79e8cf164163c633af3515d1586306a39f9c6651802aaeb3d88179f2b0ee51e5faf260cac2b715839f0db2e1dbb08e0b76e7ab41f6a4e4dc7a892a70f9b47f71638f6c4e3d03947662ebb4c15ff7baac66dca2ec5fdf7728ed195879a3baecc929714d2ac557c54b6cb290b21d8fe40f1e5cc13e0685195b9d4880d073a0055ec9b72e189c127fbc338034b383a8724b1443d2367411caa5ce897a066a6575b47f26f6c0519fecb03354efc010f3ba0ca74a4f9c32f5060d9aabfd4a0863887e56ea36b46d0787598c15e9fde5ab88351231e623871b4e18fff7012c7ef9daf05b0262cf8548fc04b688718e8ecfa7fdaafe835fb1b783d8a477d6ca3c0210193d587f341f29d12fafc9628e4254409b52200adac770a737535ede68dfc1e8302b4a5d5605b6df78bd10e0ce2daa14434ae9a6980ae673ecc848123a1edada2681e47ddb463fa8bd700f15facf00e22583269490654e995768d2b49b373f81621f285e9e5d33cbd676015350b372faf32ca16e6713e72da644cd1610b449b5cfa2e531f54d140d76505b393e9f58bcdb884aefeac0b5269ebfd9431a6df8ff331cf526801c764d4f3b0425c8a3c46b448a4960bdc38e08c84439a29f6acebb51bafbdc05a9e6b20e25807e3c90bf6f477911ba3c456bb7eb89983116d9d993d67f5814d0eaf809fd0f5a8400bd33daf327b26db5ed1829b86fe838765b2d94249e4508df5d3ea528a0dfc91bb8041e2152b819b6e0f17415cf5d50c1b6890451a9ecfe9c965527d967a425bed37b5af0d0f8a34d2f7868315b816c3d3451e38d883b96055fe742447c076afccf62a9d992f3d82aed280fc85c12aaba0adfb9cd82cd99be7a3f08afed5961966ec721055f792d9722723ca7f59c3ef5248a920edff326550ac4349f884429daf4b8dbe3a622019a889a5d510c5ebda82f4f71435b00f570a8e4950d0cc76b67dbc42598654966bc44a14fa5b46e470d289f058984a8229efbf5adc7856d48c0d5c267764e7f568c3afe91c737da8827b26dee98b856cdd02fb5f0568daf9d7c8592b94652ee8a229e0e6938f63eb0d2e99e1918966db4c60d436d0a63e0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hefe9b8a51114350d5a72b0b6eddef0509ced5f2d7bd404b1a2f8b342ece643a855ca6e12384187c7c02419564cd6019c7d31a2df4cd51e4504a88d635fdf9901971da050a92df7d956589d1359874fd76bdcc1d2335b3c552d0be0c16651cdd08529eee09b61f075c69a63b23ea67c700e1638ca2410c9b44adceca281b550c177df6b609900914302f9ef09c9252085979560dded10306b9b819050a043d3b82a517e43897f0a98d76469513dfbc1f2d4368807ede7eea4850d2a0329796f25d0b65aabb9008fa3246abcf49aa8074b5d27aa52785ae9eb53b56ab2c11d05aefd7f18a469596d7786c84949e3c63970741a275e932d67614398bbfa3b7669f0a06b79810e5172da768b0011513855e07f5fb2a575f715991edcedfb8fbfad720c7ba4999c7125769ed960154a3f6b57ec9d8b3b91e7f2dfbcc3650b2a57e5469473283e13397d6dbbddd689e925a45a3b03f6a9f25d933a18a934246c944bddc8af12d8d38741076a9c0d2dd74aae3ba1383a9cab939911d974c663fd23ac38db25eb87e8024b0a91664a18c285642a3a9a81a529c23249a194d661465089b15011456d416cf215caac3b1739d37df41d2ae3b7b1126847ac80dfa6de4f4b64ff3f6c86b644a0f4b15f38c4e980fca7ab3db0f39f130cd9bda92ff76a27db0d29ad5908dae710000a9e823ab3ac1f2b70509c4647e400e913194806ffa4957e3bd1629a3f798c6788df222b82b45b77cc9dd3c0e5e09e6f73d9b0f75eaa5e6b939c485b0795e7ce754b95a849d649156d4b0dad4cf6bda26834f23f9ffdb39e95f9ad9d2932a2e76e9af7b168fbeaf7003fc80414f617af07ac95f141505bb5e390a2e31c861ab1f2be64b1c72cc3e86326c37bda55e35e56074d246a4a0b4c7af43a78d5e0d18e61d848fd35fcbb092881ec9174fba0bc0a12aa7f37ada4ce2da3f412be8e13d95721776702ec36f37fe4af07c36c225dea02a5ad4ffd786b96ddc94dea469dbb7ef066a167e03e1cf43929bd57e69b81c27835ed09f7b9646ecade654699fedd01975ab8cb26d7b0b8d491f69e642ffb9938b0690699c602e48f59d684cb2d6fbbe64e4b0fa2cb14761ce25d0f952fe96b7093c76f179dc1d8c5d377dbc291d7c2ded7a4711b3b5d09fe7ad90f7648159ebc03d012565485a848764e9d74d644e206416925b2907b72fc92359beb5db1caab500da6d3465aea1c90f0432e1697df920b93824ff33f62aaf6999e1601ae09e1a5dc68a3b05379c77ee0e85d855bbecd7a43f5684a272048e3069893f624e0196f8680b9dcefd917870e255bb30ff413132d2d2a0454ff55e40f166d97f99711fc8fbb0e1370ad67517dab1056c9b88c5f77597ac817ee8cb213112142bda7b5eb081492f15044024cb6161d8a1364491b7661f0f7ed6cd2633c2054834bd57a7fe0de86f8aa133df1932a9c9fc6544b28dfbfc9c1584efdb3f818ad64539cf3a58397b01308cfeb6dff121487c3f4a0a8875f5f7750ffa468eb6b6801f9c0daed38b608a24d3b2a8f983c57447a53659337b718a1c19ca35873c7c73c438a3d305f15e8b45bce163d47b22ec27f8afd53f48b4c5dc111e98e0fb46eeb838603dbcd2faaac4a42b5ff7a96ba1be128fca2d10188026eb19ec60de2c423d1265d8558fa7e8feddf3495a10cc60025835c7c2c4764d6f8bdb52320f42ad01abaf5a49a43a589273ad5fb15e102b9bc1377cd67d548447ebf383218ccc810802619e7e106c7098325fc7c1f339136cfeb0702804812f77df1ac7a9e5afa268bccdf9c8a1f10a278f8d3a41bd2bf71337780baf6055528ab29744e70d76fbd9e9e08a58fbd63ab3ceb45beaf222abbebd5ea27bb8a43ad994806f065e28a7d6ad51aa95431a0d1651cbd7da55a432f9af99639a7e6913daff1fc196811f9a56838d620afff45dd9cbc64edcfe562c7efaaca056b1ce9d3ecad97537ab8fe525ab47868648c38d280137bdd9caea3a7e88b827c5907a8ab78aaa0cc4559c651f0f784a4cec589348bf614780ea951c9348aa9a90d63fba1c344e336385156f40f1a35069cd935fa18f144d12080722c0d202bb88855c24ba27d1b908f99ee86b744a3a646a50de538982c33efcdba23db3ba1e62dcb9a04b98aa7799e46957e4606158d54b39d1a7386852f1b8e861ce937040523786393ea3173446bd8a9168a244b414b6b288c71ed1aeb7023ec0dfb0a0454ceb22eab9dbe50f9cbc6039d539859e1588b29589fc1f1e31a6ca6dabd5fe6fa3508e719d2493a705fbe9550c37425e51ef97c0e632b5cb57ba347e510dc43a5a70aacacd2ffa9f98c1a7f507ec4860a462a47a11641cb7d27fcd4c67102ada4a3b03e8e414f4830c17b74e32fa6134581ffefb2cf5e315c8daf4d1ff90b80543620c10811b73514471c7032a7d9c323be0df7787234e8cb65c051a6ef7ecea24293542ae16e798f6bfa115fb58f1d686083f1777d6f62352bf7536cb80a0e2eb4f553d735a6deaa1f5b554ff8f804047becc1191307238ca4f58847f12a027fc088ea3ea25bf2b79a3910b7e1e058c62523167e89244239768f38693ba37db9dd89a04ac204efbda156c6f327dff9e3e3295f22049f7611ab727dc2a6c6ebfc7c3a0bd083bc811a7d9721b61fe4b460f5f1308447af5ee11c93569893459c37a647b21ae5140fabf66894a889681c4112b77a29b66bf87a75355c8716082e50117b2565af6b5334713e0d7b6e57482f7ab0f30643f50a5121a226d6df3c46ffc0f73b4d9a4c7172545af8dea57f85cd7da80547f6706f7c58eace129074eaf287fa10c5941b98b2fdbe08976035e02afb16abf9dde2de47d8991777186bf5c43c60acc62374216a9883ee9eca8b02c551c3ac240a44c7911b7276d93fa93b45acdc7e29a75e75c88e6aa0753c68ca0b3b9dfbb36f998c17ee83a329dc7192d00480196e4b44ca3c9ba0635de8988b13dc87d703d605f410aa7e9fb67b2e3f5de0e17a3804bf4a96adc626a05d58499306ef0bb21d499518c0ed6a1abb5ea9a164e4cc388c45ac8c683c001d7ed660334497d6b9e426a264978bdd8c55805f941f27e64e0f3f735231cf6ae4f46eaa253807399795f2a7cc517f8e8a71ed60d538b4f02b2a4b3732afc22674e9a71b222f061a33f728b364afceeb90318255796b8dc9dadccadda96dec8e3c87133e10270e05538952bdd4c79acd32b5a643752c4d1be96fc1a78416e3014e881676d633d299688ec8d086b017231f72057a140cef76652bc6930a2fd1019b8dbf1a6296e87a67610554cbbb0e3db48f2e806d462a71e726da3f5e4c151a50eba5c15fd0daf9635608add0ea48e863df6878f68016d686fbdefd005a6de8a40eee5fda1de545bad7b1bb4e406ed5a8ac5f9519806db61e9ccc7d931d6510c55b0b627545c620416a792f8933c523dd4087e72e8c72373eaff9c4381bb6e05f20bbbcf7c8312847910b3c842caa67c9aaa0ffd90a4dde58f3778c4a9979d71f5a05f4291c2fd2a2a3f212b32fbf1f8a808b49381d9d981e5a8bde9cfa0c1102dccca226d9684debfcd8f41ba6fb6ff1a15f6a010d21984bb4d9b7eb5747f6d2663a66304f46371f221f448d14a100a7328940a4e5169fe9168bf12a04196d3ee736d2e2e7014cfb25e2c344fade83cf34a6fddbe39b058e4933c5ec3ae6e09fd1639f0036ea46d0f8ba0923191dd434f8fc7fec78758141cb57bc95bb6d0c82afe5706652d4084d23d802888a5592b1b3a2008d847a7b598691b7e5e1bb7a0501fa99ea0de30a9fd33c1f0af6f43715b57c8ac8c19394069197776c22d9e93cad7471554bdbaaeeb9edb2f2562eabb4ed10a73b3041deb094c77ef3b7db24acfd2234b718d30480efe68f2feb8e087da52f1f7005b5e1766b1afbdbae00aee988a9c5ecbdf20c5fcfa2f9f4e3d1a2319cd83baaf09352a5705db130f2bd41fb5f32f8a96c3e1cfd9b11115e3c1d37785482ffd3442c8053041a38998610a0b56280dac844ed213addbc03b93567810e0c22a95390cddc5439c119dae1cf4699862d3001806e7221efff5af6198dd08c6fe5fa75e0e3d7ae2875b9a6e047a86a20c1c2a6aba00697d231ca26267818f66f3f422166adc3cb0242110704a88f393b30124b6e8ebdacb9a8f46b4b575e1cce621111bf5c4016734eb6e8a9251abc806a731fa7e6fa64461351788b925e46f57a9249d08abc1917ab6de8fe9b9244765537d711314c1a398886b8890b1df76fe276ef641d13c7d9637226f7d1844b22aaf2afe2fdecf6eb6173310aa3bd3abc70565b7691445816389d00e8b77b461972ad55fffbf3239e80340cc9c762f36e7376b093ca87295230a270451b00478d7c241ad35cda7495a6c4877e5b4963ba760412650d51fb994fd637041aeaa0e1a86743f3c72ab3364c246819a8fb027bf1220884376ce74ef4e65651f0571c62e5ceceb4042699d1e3aa2eb384eaa6d189aea1744be2cfbd62cc18601d90831609d835d56c76072cab231b3f66e78d5cb5ba829b3e872eac2954b9fdaa8a6a54caf1a87283453e9e9e6b8f329988069b82bce5801c226f01f14f262eaa2e174d46447ec921fdb6881b7c12433f2175c9f87c6d7f6b98153ae7071d49f9cff590377d7e7b37bf24a068270ed2c1e65e3a41f747c489ce0ca07c5c74ab480c9418fd8585a36234d45da972098483a248db220f1d623062569c380a1d72c21e1c11de818a01129c960a2b0292baad53d872b2424e2f1174efef7a7ee80204f26b41f9893b95b1053ec1d7b3402a4c0f1a28ad2f73d7bce54d895166d507ab3182b46489e2b792eff679c6ae7f2dedd2f2193b253bcfb45ea01639f435c7cd392cb906cc73cb4aca986aaa72e8bdf91e9b52755903f520713379dcb515d0ddc78aa59e9db34c161df0ea6c63db48ee20f10be5edd0f22334908c9f5ec26e672480a57b72d66c579c50807858ca0c743bccdce94590557cf650df1323e0edcee5c0f9b9de700e9fa3c9591052a99a82f42b54125bfba010e200530d7e951ea02608400ef6b159954693d5fc0cd2f8c315254fe9268e521cfa4af4f99e82dda6d8a72db51e12068e2b481eb54f7f9b146de16e99b8777b57cfb8db0be35e8f5a4002cf8961f05d6d39121134a397908354b7b3aa048d0aa8702d6bf28b63eaced020d0a6fec11affef46b932b068d6a67793192321b6f7db49639c520bae0c218d5786ff46e280c97523280132724abcacf5f7899c91857bafbff9c018f1a972e101b46242fe7b9b7df772e1135e956ee0f4c69c15c14f9a5210cec5ba81fbed7dc172c139c0b48d44a2f08b48e3b143e8c80bc051155ec86e87655d6cdf21dc316021a526fdc0389001e7ac1eed939b5caa9518028cd3c00e623a523bea8a28bd0f8fe99a239384b907e745eae74881724290f5cc7f34a50858fd29b6b2911bed88d0221e67f7d8b75fc020965534aea1ea1838c11bd3b14db42e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'ha48bcf7bcd8d9d4a3cb2534e75803e58c6e7734da823152e952bc8f380d4b0be609b0a6181e77eb76035c3c8422867f19876c8b0fc0a8f1dbe887577390d765bcd814a037b6be826c5d19d7abc4176167d139a6173ea32eb85bd980c99f295ad6949747840f380c76fe4bae22dcda3d117f35cc643bab45d8988cbfce5a6d379ae9f8b5e5c4f6ec42d2ed64ed58bb9185cf8c2d31244317cb78190c962ae303bdf575d388c81743006a306e79dddfdb4125f1bc605223914eb0e8d028db5fc660aed1a3ba325b0795e1ddb9480a4feb4b6ef6769e7eee53b2fc13e306612aeb83492fb470f3aec5240330d5d8b69a2af879474c1f447e2db8b711c679350ca582631cf312c445a410fd0924485d720709c3d311cecaf898f061b1424238d23cff11466914958afbd9cfe736971ce4e7b6d578aef581a9b8c7692bf8a250bdb4582b65eb11f47bde27a2fa0a31913899cb7327135f2cbdfa7bc1210acbc97597bf67773313f357e6d76116202a5427315c5c3e3ac7e8daeea6b16d99825c88816446a7105ef2b28c6ef8e57ad7a521076a6704ebeff301524739c9fb449dc00a3913e7d97ee1f711ac6c5c040241dc43ab4d93b8a940ba524840be8bb9342da92db3077434f8140a41d8eee7caa1294c84d4fd73f2e428c73045c133ff25062d21b22e38824c3a70979a25caf6af9049c74df75ea613ba192f69a840a89df8177784b250ed1e0439c9616efc718efd689bba213ff5f1fd19aec72392aaac331896f23c81e01ff7e7043dc8ba27e36ae3f861ed6770bdaa2c538e805cc77d8650fd33bd69a57e8182a355a604bfccaf6eacfea2c412ff81d5576f63bab4fddcc98e2f0207e0c17570c54284c54416477795ea351f7e6d68cd9b348295d29df06a4ae82f28b8c3576d14191a3392963f164b21138bd0563f68f197777df602fd6638b3ecdbda4c793cfec0527953f83d374d400439916ff9a16a6bfd0cb2d925de47fd128cf56e69b5bfc361797e61446635ff49a94c96415bdf49f19d7b9ffd9f7efdf717db4d2f0148b47207f09869cfcc8ec6cea31cc3630419b98d2b1818fd0705d13d35a2b1c26854a3447e46c14723f494923ccaf7c50d46425581d89776153f461194432fde89266b4e7152688d649ff415dc447970940e1f75308180bac32329a5fe50dfdb23a968fa527d196f839a0e3813073aa15f84a4fdd30b3e6d4bbb778d10c5158d237853a78af21b79f01a0ad32849d7381c8ccaa4e57e2216feca7e30f6784acaa9170059adbe4a8c01648d096e76ce92b15a85e5997cb02e6b8190222322974417b920202c976900a7a0680ce51a5326cfabe4436f6a94f18b6d9a3bca980c80672a4d80888442bb09ef6732ed269d97b896c41aea55f7340fe7965bd48cd20749f87bf934ccec0c5f8d33d78963031a3cbefd9afd0172ed48a37e14f353faef4750d3220fbfb8b593e593a8f15258bf6fef6b8b1bc437ec3d04d6f3db9875d8a0dfd078807ed9f6d8c2cb46872d73f55b254b22f5e8d0f3cf5b22433e2ee12d3d50aac027bc1f46b2bc6fd63a10413e2b1df1a0b8781622ddfd7829e15bb55d9cd88d8ab2bfc94f32587666adce723d5ff4140967bc2bf3e86884cef8e077936f5f68147121fc41eaf5a6d6bca2edfb47a055f8ea9451806f1c53ef8e3cfa9b6a3bdde166fcdd7c5d1b046d6eee3b4fe81b01c16a690167bcbba3c059e3d81ef4ffe013d99bd038a69c715627873ae472a04fda5c89c038415a0e52e191f183bea9ae1abe5beed781fb93c0f09ddcb0bfc3bae229debeba9393263371b4ae37d63159645695a40def52e1a44df89fad7fceccb0a1ad091b43a2be7f25969dc386ee6f9a45136171b8173a2dfbef15f801279e79091bfa7bd38b90d32885b082df43a851d0dfca4433f60172ccd27a115af3554ac4e41ea3833c494b0a4420c405e165e36bf92669f6c0ee1e9f24fcefcd42529f3334d5f5a1ad28ecaa7314086e2214c3e66c10346aa2d8d06a4a189f11fe827f1e4c2d0317032071b1ace507ada4a56e4c35c1fa08a54d697df50eb8da5e63b104b55b559cc6a0d9bdc48977e7883e19a4720954c0ebdd37c56c9aa1e14ec09524b4a48e731852de1f57c82e1f01348a588f275016792cfbfb25271fd162193414913fbf02a1e0183e1f74093f2fc6c475c191e00ebbae07fa6a28eac653d702102b184f77b137a334c9ffe8ec1c0fcc879711476f15acf6cbd21ddfdfeecc14f37367eea3d7f64fbe24a54a7f0c9bd094d6a11f670918579e2021925d37676bb208e22377a88f6b32a9e7244df10cad4d5c2699f2494ef665818801d15f0d46742a949b039eb954eb6226bf2f1f8808e06c71d4db632ea93e9fb5ac5990158f062a9213ba1229954dc17c08a6272934ab414f52355ea39d30293f011d10c84b4c499741331bcdf2d12ff12e3322897fb2a3d2fd703da8b064d9fc226d61eb8f2cc6754d125e811786b1aade65dc98e125a0fb63d2ba7d509e3cd518e2f213e47e83991da5f5b2f533d493e1323bd1640bf58022965fbeaf8fb259c7d50fb3b78e710a25fbda64563f36483176d3bd77bc07f9369ac71eacd079387960f96fd568ddb20ca65584a1e3047d47ac4be2d24d3b32e09ecfb12e717101eed4432b395f665baba2fe9f33e17073db9cd87f09c92127dcfeb34625f4267df9a5c2a34483d255ee5d61be5754adfed6fca754807c687ed5f61b35681190f913bc412bd2f1ead15f6257e93f5dfa7abafcafeadbeeda5f53dd5ce9d1ffa8544c44517740268bc56466c36e99158e25f6665709d691b1e831d58430413425de79a8aa167e2f13cda73c97fedd7faa5e55660693f546bd1283abd50a169de5a6d185d93971b916e40fa6b843fb637f160598cbfa9d40d30362f096c1fcaf45e1970f6f8e1085dba1d2a3ba590d66c51043dc2ea16088a3c1720c52fdd5aa3516404a3c89ae226187cbb84271723f790a782f8826a47cb4e37e3fa8cfb0ad109c55cec903ccc2592fd3d76d6cb393b60399b5e47d505c159e1615b70bc677faf79f7095d3b8e3eb4d3692a1517c103469cf92bbef9c1e45285d4ea3048e44fc4e4447449b384c02f808a0e40208e6e272d5dfa09e5da040a92788f77d0b0f64070d923ddc26b09696832a2454d333d2843d370175eccf5c193ef68ec538a11c82fd75d9402dc8e5b72ea67288b4d5617f4491c2bc4e3f1c62509d996978a408bed206081b38dd9f5435a540f7401daa49e3c1dc71c5c129c02050baab2ba6608d4bf0128069e6dd9594c4e648b48969f601c13a57cc3f37f46a746929330a70306f61d38f281463a93e844f7e2d61b2593abfd8512a4e04d4390d26455aed5d91b57ecfaf2720d75b3c651478596b632aeb069747737805d2d9d8e9bf1b450cb0cf46069d636364454c9c43e2879c8a4cf22517c13e3943d9410a1c33db1892a9c2eccc2566146f1e93cb49ecabe1af7153140ed11c3f91c81bd7a7ee0397aae195f4d8873af6749ea014ed12f7c5e5cffa01dfe7c69cc9b7bf51b362248f7a4069f3e45fecacc0c20b174a4fe3835b2557eba2ad74eaf92eb48c042dd3a9904073482ab6059d7e8167e2f22c7050caeeb74d84f536709df8e138140fa343cb139e58c1857c1ba678da0413467b1cf6a0a208d46563c20a1876cdeae08c89a19705e692600bc35d27d49a5667ac5a8ff54d9dce85357692d28b6a213d5117f0b40c7ba10954ac2cf23c4cf6e23af65a518a53eda7e44da49909c2a35a819adbe5aaffd431b5437f772cb37f0f13907575e3467e0ca29a9f5c0d15e7b8c5a9d021eaecbb0fa06d5956da873a90e45bb640422bf4001a5afc72825512d7245a4338a0732a978544eef5ce038432bd9b216de9bd65ddc90c08438a948deb8ff6e9812fa36a5e7826702b5177d1550e7d53b93efe92df73dfe2b82404576958c55545748fa7bfe14a99ae494dd657d98c799bd133f0206b97c669fadaee39d0d2d6a9873ce0ad937b9fa439aa37f1e4e02f397c9fd9823a76f9aacf817deec018f29ff3d44198ddd47351471ea4bb28706a1b85e1c78c2ab4294b1f2439064d7b68d6d53d4999d355df94bf05dc79dccfc12168d8fc9af06dd601416f8cc615473343ada86347c2fa87fd479048226c15f5741c1efd310aef48fe5b8c2fdcee854e360dbe4086769a63ca9ea87bbb85b6840b0d239a4d3d91b44207987b0e0a8fb457d9caafb37d2d49dffe0021749d64577bcf91344bfb02dc7b1dc6651e90052f2c6423d1b514ae1ec83abd2dba92d1db7e2e734b8720a813d9ba450c0f8c6a46fe4ae5421d88eeb0227e1627d21187ca78bca5ed9ad556a0a1b1fc810f75273fee4bc9404db8ed369b3b679ee2bcc87c5f90d9337ae1f82cb14e585e935aa5e8a0c60c08c23f4bceb26e10460b5103deefec92fff7d5bf2e41def4e067653f4accd6e2669bf29c140c172cadd022c6aed67f9a7496e800b36b3b1a5b94874f698a5968a8ad546f77726e0f02428f67d41d5bc9cf0dcbd364dba69c51ddf2ce0d413928c65cdbb2119a69f59d9e02231cc778b535d6ac83af72938de5ae56b2bde3ef99db659edf778232ffcf5975b0318411bcdb1ae4cafa4b5a881ad3f2478dd1b2ae0e0fd818aa7bbac492d5b502d148152b66c3fca45fdcdc379dcaec3d18f650d6f1806630c560c918e6a3c199fc24672b6a593480ab8d47e759deaf0257bef018a7f3ebc10e0082fe85c734854232b52669af105bb8fca6d543e6249486778e0c1653fbbbae0ff192176ccc778f96adae836c0e0cd3ab5f1c2abbf5e6361a8a3b1115b877b8b524683682b7c85b4e7d7d3946d2dd59a1e121e42248bd776e12ae521bea851e835368cdeecdbbb31195d98662b7a009074578b63ca81abedf77384bff8fb592d1b88caf5d504e1a30499751e2fbd5dec523acbf800d4da8ff4a8dd9d5fe22f380d378098cb990d4c8b768259b81c678c176b93d5fecc7c0b0004253d46eb607c2b796ca6ccb5b161206f1355a277fc7f830b8e9ff9de09394d862fa198bce7dd01fda5b4b23a6f460e4bc4925c95e65dd3591a1d65503153d4d3e666f31eecd915fda78d1e76dce0f5241cafab5f2f6bd51cf468656c88f2647b8fbda79682d9d9788ec08f7d759df45c1904951fc3efb31a7a919b3697febbb3ca8a7a68e5d475395113dd7ef3d282348a6cfcd7ccd63f3bc502480ae6296d33da4859630a812d05409e9e34da344a268df6eee6a08594b5191bfb7aed4b581ddfa20195f052aff6b28e653ed178bcee35fd1c622dff64b4752eeea95dfe0d777f52192e234f9024f99431f826024aeaaa0dd83e9819839bcf394498a6e0aee04cfad30fc020c60c7f6585d4192908e22b895376bf9b95306495cb0a785552ba22cf11851f575fd30f504ec09000d27fb2214803857a3a4ef027052d4c3a64c67a74ab1fe6c982c074332f7282781b6e7e550839e66f6f80;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h1ba6393410aa1e3e1f693f93a9e85ff73b18f89e94c4066bda7855cb275df1902ef859d50179e8a5be95cad0b4b9e9336eade06d39cf9b7b302efa48def39f9026cc3acacfb17c88cbea90d943d3d3c72cb995d408fdc864070b989a52c2a97ec4f01bfff5a8048c3bd1c7a01780e28293cbae0a4c4ecdedd60405b2631a32f1434821ca87b7ca1cfe01296d37fd7586a5db788e782723581ca4ced2fa8935710b8b388503db793dd14053328cc3fc8cd287b618ac92d37c1910e9dc9f38a72f3020cd94de7cd15b98fe789de6da223a1497c21805b34acb0efb082f555f863baea85e49ebf81669f477b77b2735adb4ea65eb937965080f0752b9a0ef7da04553a51b1908b9fb20380d4a3914f32c30980ac670ff46afcb4a0bf356714d71ac8054956bc376d4d355ccbcc4efbc04dc435b52160ce9433f1e9e60b829f6b8f314082b704c2078d33ad978207d4d67c78340829605a8fc5473f4f700d7c5754988f8a1085c8ff50b7e4b9635e17b881a67e93f073dbb07e92fb9edd2766c1ebd37494b092e34a1d160e76393a69de498e5b6558a1a88ba56da842795f1a614ea0ba6fa618bc3ecc03ee536ccf1ee0afe54e54f33aadcf3683902288c1ced7540b1b406ac98832ecca1a5f1332dfc5a0c318fd49f85ee3c3b3944b4db94d8ba2da473cec757b8910c22752d8941373587b1f02ed79f10fb930ba61f19d83274b87c9c14988f33212fc75d271f5c64c9187def7a05f0f86d4cca19c48e54f1afb6307a3d9832094f824edd5a7cd3122535389eb8180b537c8a1b87cfc8032f75574d006f518c194684004ac79c3030030db647ce63317c46ff30a2863803369d4b788475c914737f6418522f991006707d72b93a8e112dae965726091ebba9c395a4cb44d998ac613535f33c7768f861c863e449afa22c583b47db2d54d65654fc2e47e7337309d0cdbca5df55f02df8034090078bcb95a07ca7156dc5e2719e57cac2efa05902dc18e0a6e8044fbc9585f2cb6b89d7b36366dcbbb77c4689e7ea337e985e03c3c4fc40327ee43ba5aeff3b54970bf48b9ca8a378ab135e1092058e38ce0b3d1abf9bfaa502676e51be672b22dee8ed37674b410c5d3356cde93737974dc0185ac860447ce0a4275ab528e4161a809722f8f132def00987a24c935e35db1c051fac3e866d13ae6b00271f0e2fa68a9c2bc7cc7276bc1a4c1f5555c32a54d9e4f4f1e717d009b476b97af0912100fa9f929a0bae2cfa8bf059b951214731daf1d88696b0586f4a281643a3e1b9ef929e338322d958e4b4737f21a8d74e1d4308740831aa0aed97fa2b7006b9d947ef80f489ebfb5cd3441c3843356e4356757782b34c48e936090609c6f984eea4cbb7f592747c97e4b43b83a8a0b3424633e98899218253a6ad3dab8913767f944e98e402100c337c41f911e177d646211f4e3b52b5d06875c4254ae144c9b8dac8795a0b0777182e42c246c833d217a1d5abe26d696a46073067a1d4abbab9e6717ea36d15993a7758139ef02faf1c87c21425b1bfc8837a40b1f8daa9c965f4dbb5fc30286b331ab59773af39ec77d06da413a5119194cfbdc150e35fe3d1f63c27a0a6b330e84943059459222d3dad14b5080fcc953b873ac154edaaeb51da76140f1982b793f73f62a82ef35a5e9c81555524003097044a60ab1a29da9ba291c5caeff576ab045ac20d6f855e0696fd417ff76421303e5bce78caa1189f9e14fb419b434041cac83c82e7f91b5b6d3c5a2b2761c2e1f18ed66d1a4f145661bb86f3fc1c747b0d219f284b8636012c8c6912955722bae3bb4da459a5fc183503a57643ba53240091846d6a40cc7cfb62f65e6b94da29ffeb5d098a2c09c4b7983d26100d3342c0c95fffbe6611118ebfe10a7f5919cd828b58fc05648c8ef7e27ee9f0039102cce3946703355b4105ffb0371ad795d3969d09aa915f1e98ce651e92db7b3321d18b1d23848a29d69a7fd9ce9118cf7666bbb8661f9a411e7a21c7e4a8d02c15059242d6896e274f05956d293118972b68dd910933fdd5c8221db114879ba2e6d21c4ac1a6bd82ba5adcf6defc3c2dd77319a8fcd50742365857c7ffec8d514e953da73dfe8853908f44400498fd70cd4b1c5b1951891204a9187ac33f3a03e728a5a9b18dc4953830ddd943b37847d66337d250f2b41eaeee97517d01c060c07bf00a48d535da8c1e3de271e8f4b7def29bc2c41aab306d3de8b2f747ccd560baf9dab053e6bfaa56b73086ea19a1d340f04a1056ec92daeeb976693308c1a1bfc75529c9a6acd47ecfe4df09d6f0e7aa4b0f5779dead7b4651b1e51ee05c401dc606c9ee22719736f0c76d4d2f5a4d905d2374cadf31cecda6a12eaac6a0bfa84c00a3526b2fcbc241634a5c2cc153e9e496596175ed426a19c2badc0b8d156cd39d173dad8842d03a187414cb47a1afaf8fb67f9b842b33c488d927a11ba32ab424c9ef90fc96c8f1d78c2e23e31331b02f5473d92eda1d8db555e93d6be69d78dac1069d15141aefd447ae77ea7fdf77529cc1c057412ff6cc584c5f0606adc2a501b53e744e75e305dddc0edcf828b22611e93f72af60dbe5cd25e43360d53ed00b0bfafa01fdfed76d5729937525fed4cef22805859f07f0b06efe48cf11f240f45ee78455132a7eaa1e9393a374c950ed943ec7ed32cfe11f7cb7d15e956b5a3887a2e1c31fa111acf091fcc4bf3cad2aa6bef523ce016182cefbb2d2d500acb98d000eb76e0e9b31c3b8489d2c6a420b29148652ce0894cf4c757199e8cea2e661c8390fb268d806721cf3368859c42cdbacf507fec3faf7b88ae38a1408158fd04acabc77db95b69bbfce5add05bced525dc03d67c0d0bc5b0ee1146d4dacfbab431889385171866ad3e54e6427d93a30a4e4ce87d2c636b99fe9c95feab7f2d34ea67bd3c789233f38944fc09dd3392e529148bc6e019aa5a37a7b140c3239ff7184f310754e60d245b93513b54a1a42feb24b524b7712eed0f80691f697be97a26bbdd0e64230446119adef18048073b678f05b01ac5c1f4c177cfb3e06ee7782fb5ae16d5c6561b74ea9196999134f8de119fa2a1ee2371af22e17decc440deb80ec168f65a39002d6155a8587f7c8101af0335fabcdd5590c92a3c5db00586d4cd3c785b396656999b9d982e153c566ecf71b5d6b7bacd4c5d380531060a50fbc2f58ae7b439fbcefb7d860974bda02650e3f645ed316f853bfb5086a8637752246615f529c18a7fbf94e81cce1c01658b8157f41538bac877d32dcb19fb9bda48a79d0c88d5a9e7cbfb8bb8f96795fe06df2d0aa025dfe93515bd10958c2355d2bbf486632559164cb6c524e290f2c175d36454a3c45ffd57b4d283038fe8b97f78daeda43f4333d2fce79cbf91622c06d108796d099cb9b7a1531c64becc3ab931a5da70b0727f868e0c059ae2135d8dd3188a0b244db9d27c3cd0c7a169b76eafaeacb866acd55b8d53c0bd430aa96666f842f55edd3eaad05409eca30c5057f728fbf2375872acbaf6c7051214ac2bd8e28e61371e4823f6fb995307f03fae43def7af3c768ff43855efc645af03d95d7bfb486f77ecb08d26e5f4a9ec5dd18517d8224b15c2d0dbb95515adfa31053fde503f8efc8bfc02b1e349deed2d9aa8696add3080fe3e9a3254cd990323841ea7185e5a8fbe0188655795ba64ad8cce31c6ffaa486a8b1a7444f051bf43226be984dd765a117885b87e2c6956b62a56a0045fb0252ed0eef04db962b86f9632cf18864bec4a200db91f8fdf83ba6e74826d2d4c2de8ee506c14fc050c1d6dc440a1572e9c674b65c4597d98026781a62ab60a188c02a9bc827303fd71470fa9637391ca2a005a298b4d77d1ac11b6bfe10656df03e5563a1f6042865ce5c6c2b82803d808ce9d061d59ef0d355ee7662ef34dfb044be3f429bd3bacd62ea034172962466539da2544964de1d3f54a479ead1a113627e9270aed0edd9164ca3ee01611addf8ed47b2cc5fbacf39f942d24f8af609b343bfab19d6a5f25998ca7e24cb4f289e40b8105bb74ca67cea12c0a450aeffb135e15c378829b6e093a7a7e812c55a4d13ca4625439f5a3837a2a35acc72ce7ed5d23b5f8f20b47c423df55593e2b4d73bf7e07a0feeeacf7b930fbe2189653623cdab533d1241f7d773a1111da34fc86e87d35689d821aa7473454d6b31a2dbf476a61c189c8ee687e30351b96f406df39ec1439dc86b0a350dbe5a04a77feb12a137054b70a9043cdde6cd737bfe6a9daab2c2a3a9be8bb5586e881694339c637efd64e80b6f75389a2effbc07ffd7b9b4c50c05d2cdb435d16c56fe9191ce2b77fd03b0e71740d189966207b78fa7e87b86cd6f7b0202b98c833323a09b673ad69674565d9e871241300c0cb228c14390750c612e674f29d417a30578d8762d956a9b5f8d6b0164e9e0f426c879b417429bc9121f31f77ce11c41eadee6bee9e1e739ac57cccc095f155e86fc3e5dcadf65a8b7b9679fd6c5858d3f82aa0cbd5d1ece40e0370479de68166d2b49adcbf2c809b4297a9fb2249e9c182a4f690c4cf580cd40954d69e79747b99369164483bfadf97e62d00dd4e96541a1afee7be8c55b1d228b9d336d16b1a5c2b06c03487a3b869aea2a15bb80919e2164a76ba394388f19db0f5b76db7a5b7da20f3becf3909972078111df48196ae9b46c5b843666da0e92c5757c217b94f0f3a1755ea11b8381e0cda43e965f6c47a34116119f3a2c1a39b9f1edb970d0c4c2fd99e2cca722cf396b8dd6836b2c4381297422d4d166856f37fc569ebab3274becd31769a1a06113cfc4de850e458d2467aa6a0d5d238726b134d67065bdb7d02eb135ddef3715e23992308f1843b1ff3dd820666fa5dcf630a04781fc5557480520a505ebaf7d1c929a6995744a05de13161e8a8c63a533819502da31b91a693bb9b0aa91e52012af6df46e8a99b6aa75d622b44d8dad556817f8069b83b01e1f97caa0be431f8b4bbdcdf6e8c503d89d118e1cb5d646ffde66f875815505d7446b1cc2feb7760299f0d781cf2f2f4465dace58da88fd4d7a21b578384f062684ba83f7de3ac4530f13036974007e137f27e8e5ef92c0885bcf5f3987bf956060aa6293fec5182237f8f08e702c783dd2a3d9bbb98ce56c0a08c11701f60cfac6d3faa343ccc198a5e19783b72a31fb5931300c6eb1cb4870ec492e0fa6fc537717b95901149ec4bd9f7bf61ac5745b483ae46ba8ba8b634d68925f9149d0dc8c8ee7e97f02ba4ad717375df3aad329ef59a305029ea21107317bf0fad6c8e990230fad4fd2f4e4b6fccc5ecd4f239727775fa4f6f5e54c94b4a2460fff593733ed5aa8e05681a51235db49245672338b978c55fdb57eb845c87bd4f4877d3b74f0086169d8cbf33275e74b1db25ebb7317233930460d4b3c97666e73708be7afd5d2fc253f58ceba39ae56912cb14f664048a7370dcb58dd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he88f68eb32c13d49fe32c7a22ce782e87b371348f5af821a702e7f2b79571fcbf8dbf338009e4fc4e70baaacaadba127c1ebe762fd41befabda9ccb0bf01fbdc3949c7fcb327384d56968aca66844d07c54cd1eebe9b55e5dc885b94c2be1ab32237114f3487702aaf91f67ec3e8586c9bcf062e8d1355b77106e6a0c90d6c392ab9ed102844a4ecc003836017209e063fac095bad87813bd91dd141d36223b9678fad6d7dd5318c1a4ef3d9061513f14da739580194e5dfb2352dd38c2689d8b8bb225be2a114ca217fda7b15379a41e5def840162c85c7782aae2b5d41c83daa94a5220a4703a469e0c7de8321da5dd748873f3d10a9b9035a43f9ccebbe61d37ce2a130468745263dade2738c7c2e3478b526a4ebae253ef423944957e20c451a38a67b9c9b10fff14cd8e553747e65502391c65960986042e395da0716f0603d8f1ccc672ed5dcc729c02fa5ccd7df61368b0ed5e6614290ec75e015876291815ddd22dc9edc640609c9d212daaaf51c5d6a9b18952d3852ccc77ed3e32c76a92fd872f9c5ab2482d51092cd02dc9b4d9b49f6bd31e8e93dd27605c50afcbdc3c166c1acccfcdc1d778ad325290854256ac6e255a97ba0179b7924bb8fe1e5a0e8e83c02651ccde2078d2fff86101ab5db4416f22f5a08c70f41226cf3ba3fefbc1f4e75740fd5dc6b2c4717b1e0c410d224434351bd744cd01a94ac98dc614b60da0c64f74b4d9b7733a895546d95d08c48f30739c8afdab227c53b206859f4d581ff131f27a1be6a1748c9a096616c9f1fbc745cd78d20c050468c32e41732a9210abef4dc0e33265e1b87af6dd413fd2db65addb9b696839d88e6db97ea5e382da7f081fb4013d67bded39e7936180e226af8b816d085b92db2ac82072974e82d22b201c9b8933d7b15cbe5bacae84f73548aa9fd5746fac812338587df8e52413513cca639854db9bb91442854f55d1aa56d0ca4428193c19c3ee892af5971ff7429d6dcc037094067d1b8afc1898f1d626c3e8a0267bf4ea658ff9d52de6c675fd34e9636dbaba01c63800726e2227fad17d756505fbae2b24d7e972ebebb62dbe40493bca4b4301763bb2cb1d1a888722f30ef08765c6b3a123bdc3066869b44d55a0e95a7c409741a17801c8a02fd1797113c8f3f52800125300502c5d50003efc76b758a4f22ee8b5ee0842f014e37afad5dbf956f8f87998d948213e634c6874f854c0c904ca9ead578c57358cecc8ee924b224db9c4b72138514bdd45b4b9d1674ca855e77152fc14384afd09bf9a688f6350214f4202924c657f3f28570ab13389ed0511b24dc34ef412c15893ab2444fce556714e5778f38667791a12790c1de83623585a5bebb33b1e012702e743808f14995f17f4d5904fd6f6e39f4341a3be63f2fa2a604c66fb7b076750f3bb07d5cca72f2e3ecd8a384d15b78c751e42330d98e81e88982a76dc0aac029c84cccdd5d7e1317ef62dff6e34604970f159faeb3331579107afe1d3cdd687b4bc5567e7239e492f1cfffb6cacb953fc4426d61cf805d8ec2a707466b2809a3e0341ca18ac4abf0322656c82fd8883043adac563ac4557ebd3c015b41a79c0949665f4ee41f86a0c7172ad38effe769492d58b6db7b6668f8dd26472adc488623de0d9ba5fb55b860b130bf61fe98154720d4d25ae5915b7c92a879a493724351b6f6a50fde1dd777326841e62426338253ae63388b52e679d467324402fcc0bae6a69ce0c962882a7e2980e92d21dab68e8d3c43b1010eafec76a03afcf15259fd3a24b1ddf8d14eef7dcdfe41b92c0058f47ad02976428d8ec16157f33cf108b4bc322bb1e4b52247dc0f0b09c36df43dc267956183c8fa5438dff6c3a6d65e1c68a72aa2160d671d73d7c4bd96ef9885456847f7adad131bc1e4471ca9d4748a28784a9c95890b3ce12ce566be251fe4c7e8e7e1a2ce8838fe081d8012809d022383851ed2974619aa331d574fcd849dbc4ec549546e1609e79ef317c10a55bb3941eb03c93a78dc5fd03dc6d3b78a100fc03b6e7ca584e3aca6587fec022f4fea411192d2a188c4f6d6d125fe87f039f4aa3b28552b6d7002c5fbbf12ec2c0e935ea8867fed6eb7828b2f1992fe8fb4feaba50f3e1262d3ab0fd924e90299e0b75d57a22f8a0b6973d0cfd548595b49d562d3058a30b482007439c3e7a9b427e2e5107761bf74a79036489dc66aa04ec70e02ea8600a14b562724941775950cc72a6e767e3adbee0db092752e1b0a644e47bac30e69f01fd64ab6e0898d8a304d55d3cdde0fdabe5dede3bfa3561faf9e5220bd17ec3f33ee7bf21aa3aa958bb9e5a4027692c73774749cf67d91e206bced6e23708f81105540b7e7c5213e5fc6c5cbf5c464d7f757bb91d4e60b2130fc3572b3826bbb08a43ca789d8094dee9cba97a2fad0abcc49b41083f47fdd12b9e8215bd730794e6a466dcadf0c3fbc6e24fe4770ddfecde1a9be340af24c5d505f5d7437d032192b4aa75c204fe8d4c3d6640a7c587025f108bc3efaf23e4a5d25f1c9bcc4149e8183e49431860779bb151b6247abfe86b374fbc0613415603d465596c84d61f5f3b952faa4ad0b920042f8fc951b4d30c667672a1cf17c1f9803326a6b8649670fd414d5a726066dcf393dd4a6dfda9ca605356a7d8e6e0f150dd3be2ddd6462686ed3761911bddbbfc826a5be309ba75f1ca315bf49181250f43dff1abde69df65025a3cdff2902efefbcb3f69c3449f8030b0160166c7a797f123d9d09c8077a1e04c375c28526de69d863a2cf51e0cd3b61a883419f5a38a13ababa0db234b06e4b8f720bf0f427e19cd5f65d2803cd345199ca687007b14a90c90a19fb556d1bcbe888547da1a9dd456d7658c6657ce51a0d16ee99a2c4335ef646f77264aa077babb7a863c97085a96a5f3784e48b1ba7e57238fddbe2a4c97c8d27847b5bd6a9cbece34a0d60dd9adf9d5341735017c11f947d2ffad50887d617d00dc734d42621d1db5229434ea56c409ee2208003430885c29da2ad0d446ac58f409d6581d179f3fb7c57e06e0ff04e1615828b1997d062f11283d8b6afe471e927626202096e72f2465338f80c27d719bb1529b11b8cb837016fd0eb6ea7546fa2ec10435797f90b106fa18a81f8c08fc1dec5c366ef0a1bf1a99f50d777d145955cd5750b1c30005a54d484475f76613a7babe69be63f381b6042bcd8ee7c6efa69a8f555ca418d11114282a6a9fa592247019ce730e40566a08d660bf8ba562c372e1ad606a7407525d4eca7b92fd3c24067e70798c7dddf35312892305884cd895c42643f73d726e7d8335c99d75130dc9eb7f5bf8aa66bcef083dce798efdc526cc2fda5ee6031e92adcea49475647d6181901c9f639b29a1820c1e19af9f8b48d873f81a352411d72171555405118d2c9f8c3e6fa796822e517d132f432ee7ff6793c14f98d9aeaa46c397fcbeda208f5d3013d2f670ef3158e6347f006272fa560d91bce73c538eb78c1e82b81a2ae7aa20161122feca799c6ec936250909fb67643c69303cb8985b24d10636c6d28b767134f1424ffb3a4f34992f28d337b24ff2ebee77bf5ca2e33574fd6ebfc7f9ac4e2ec20b448edf5d47f4e94fece7a74e718ce84339f78751e51ade53ba8a9a16aefa60d0d1b1586b302646c7b30fdd514a944474e7f3c21ebc6a9f9f1ba3999536780d1894a70fd6a52569333113cff61cb593f077ff5eab44d89310a88f158b3f91fc328709d016f01184a33589fa068c7679955132dd3639b650b82469006fb0064a36e2b468bf6da9b3c7bb22225121ff90a2b4e30e95847daefcdabc238dca1aeda5f4a2c976fa15cbca709c02e7fd4bd862f7521056358c752cafd1160a3391471b09710670db7880eb05472b4cece440d127abf47b83436303d7b4770608b8268e247901c12c9005a559d7c94609a0384acdc4ab24f831d3ad5b62a38c7963726fb9034056dea29b23335a53e1f979dfa9688ddc117591629281946c6619c0dcedf78c684332883bf9f17d24241413b0a513795820cbeac88606d503b13201830d25e570b99aaf27bc885963dfc9d12b8cfd52c78ffb9d02b4f23136978b8c7b6baf48ed8958790da10d3c56cf6ee07283fc44f4f7afd58cbd2201410fbce013afbda8ae424c51c730033cc19911d2817916676aad5dfad1011f3cd8da5c082ecf6df7d1a9c6309b5d7c03355d2db036fb1e03bd096429a26d433694a69a539371d45c5225be1d51dc9acbc105691ab8f902e376086a38c133697cdd4a92edef8280deaa32025397e61f81f5f902a638b8326a57bb442f6a945fb8d16e47452a2789717235b15dce5b7be540f58e9f2d67386b72bb3f80e1f6606d880ffbc5a4d8ed966799e694e6615e644d3daece21da4c4e43cd69dc083fd683ee0fc0f181b591afb67eef86c779d4d4cda6089292742ef14d6f7de64ed7f669a613f81ec8b83899d05f691dbe5b471e4a5b21aa4ed92ab8e70ef679bb11373db488f4ca2b639ef5b2dd843d760d74183ea7386f066c14d92dcbc7323272c325aefb78a2e1935216a4f40fb68bf78386c8be269bc9a4848d8e2d87f6a5247940c06f4e134bd7fc675433062ba9c49d53edb249ca479ae3fd218db24c0d6eeb7c23dbd581d5096b97662ba641938cd9c138d96449bd0377074de6f9aab4173ad7261dda7bdd23acf75f1ff56e04e2d9a86c3223245b8ba4e444070df1192801687380aec4ae1a89ed04af078bd4246885edd69b466da21f748f3f6cba7805e917957401dab30e17cb9066e72b71ca34d0838dbda217677167cddceae161bf4d18f02c7f164b960c88d7af9dbee900cd75409233fbb116434b500bc9d5422485ecdc7a774e0ed1f2a766d949685ceccda2214ebb5c9353b97adbf1ef419330a90d902bf40a167e399d21ca01f62a67d771e1c0501630860256237cc0ebe99524aa50761bd0c9b686094aefbe1a452b13d53c57c8e899ae6e395669e6254e3a37265b4613f591f339db0f9147d36d00c6348771deea7c5bfcb37af7b34de22472fc9bc3203c678559ab90dd539a69013f24e5581da69110bc580393ff21f867389ff43baa110b64bc15239734ce640489f1725a13a517535d49ddced8e59645e4c22e52904b015cd09e032352bbc9125c3cbb3a2b569820260f1dbb536c870f702e3a63c5ffb91e0c5c05bcf03014a7575d3ea3cb056324840f790ac94ec3002688559a40a2caf371f9ed1cda9074a336bac63b2dcab1ea729e2f81f6a5fb4e56df4869a2dc6c51a3582d1e15420755bcec011a6911ee1269df4a534c2d8d8cca96c62eb664050e2a263ff974598bd4050a9da2f165bc5b75fe92b438406c4564cf472dfb5674a276bc3cfb23655522297136a92ae83e0591c6439444a200f2492b2992a932487c20538fc33be73aacfc505d92a5500de2eb2f239f47feb4c955d68e7dc849288e1e691d15764f9559594b84f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h7d8cd2c30e1fb6b6dd2be90cf86d2d4a84a0e7b9da0a38049412cede10f81af561ebdcf36b4d40a985bb10b1aaa8c2ab58c9583f4313d938f69ac4296b67e621069a5aff7e7ec0941b62068ae27c0cb68cbc814e3e66190bf6fe3ab64e06d08a3f09e7c9f9e9dfc13d026e2615c5049e3fa8b94188c09260b986f193d04781616def403efb32ad1e4a3af08681cc113b78b73505a43d01a2ec72753df0671ee2c5101c3da7da93607854cbb5134e0009f3eb8b22d97b9902c938f3e81cff45393ede75fd524ccf03f7f871f052e5656e0a95725fdd86facaa363a530680ebb9297849832f076d4a439da819cc11e874c4db53fa6db07107b55f9df08295b8494c223b06ea93dad54d706589221715d5502b1cb5422ea26ed0c470e11908e4cb7fb1ffad74dc6ab8eaaf1e5b65df71ff464253e92e7699080dc0dacc5e0a7e66a2477b39ea954fa2892f299986b1e7b6989bf22532bd2fb4494b44f63b7e7b1c772f84d1a4e727d532206c52ff66304c78744ec39c87bb2146d424b62692991d3184ed60429f9ccd5befbc1ab308f91566f29b49aeb310646d2543d0eea57531666310718a33c709164348e618673b026a927f58cba7808143338d8ad0a518b3175d3ec6fa26e37831bf6d776c935a243e3add57000f2834db4a5e929151b5f27622bfb0b2c94dc6254cb642acb9f7cc9b803d0dcb6b15b17cd785e7e4b105dcf12b582f3a1984f3d2ac2f6456d9b3f9356279a6c4cfe362226a1e0e7ea0fe30a2a1796817f1896969828abb04a4ede17333d30cd6abe333943a2bd8be53a4f33a149eb6353817537e55e71de8f4d2c10eafa444719254356ac34269cafb21a4afd08e916044a14bbf5ee0c33be502c58f51f7a29660eee56e78b16995f1ab2305b42f2566bf235ac26555a9a77157871c6c68f4ec10851fe5fd57283468037d6e2c3a512f45705f75de53007042410c659c37bde7925035b6c65970ca1c5366abc680f6f2776b7373360dd7474ec33c3db2567ddff99a592b1b39cf51066f5dd1c704f94061d959dd1e52ab423e47d958c1f3b838ef28c7b774934d3737d0b3aaa1d1bb8965c3ccbe43a27c8b3d6e60df581f6de283b0319f8f52c43498208bdffc9de2a8ce90050c1c123d9a4c0974fb46c714e65c93a4199becc8920b57d848b9ca8772c1bb58f19e0b75f78f37a341eba19892964074e3965aa1ce615986cac4d2180dd386ea008f6098c5a7492a2c5687792446ed82d3a843abd03f11a1903a103b0aec7cefb39599fe7335a1125fdff6c54bceeee7205eef6869a9b123d9a1ad885a1b3e06fe802f3b23a607f7c4e26efed0ea47e3bb1a5ec356b112157ada8e25342a0adeb914d9d30e5c0ff907208682e49966c1e8d9b4777f0df5d330d14e0826687a2513581aa5d401ba44da384b19ed466f94c4782667b8944914a2cc844bd41999513a4f4547952d039de7c0b725974be76fc9870110fc307ec3028420ab29743f0ab206b3eb29db21f80d6515a80fb5985d43c05894a2e760ccf026cc095f5738a2dcd2a94f85456d11cdcdcdf0c8b7fc893939f6624b2be157dc95f2011858c68623e5506c759ad160b9ffcddb25888d0896e15891797c4231db35d716d9f4d07a5ae116e4743e546abfe161234696eb24cf792820b33df397d28f4497ddb963bfe95e7cb6dcfa938bd1fe38240830d581c1f96c32d60ae32b7bee14e3874d8d49a1613f7b5d096e94e1d8f7b1943f628cafd6ed2d99928ca965cc44ff15575ce05089694b10a71ee75ea53c532d4f1b2848b6f5e3ff36d115cdff394996de6402a88210b5bf2682761557343e2c9cf83afd89ed79c6bda5705bb463e4b3393a8e0d9510558a6337765f49e65bb5888072f862fb3b32b1c8783af466b214c337de74743c44fb9753c61acd8c9ea7f7162fb9c2d9368f108fe41cd6a94b1748efe5893775a637bf94b4319a2c13abbf48412e6e200ca1ce5d9bb6770cce3076381c065757762a86fd4caeb7afbc67eddf0468b7b2a6b69056b2ff8183e3bf3827cb289dce5dac502766f725a9b62109a2c2b136abf5946bb7e2aaacdfe4d64adba3726b3170c754a8bee8276d47ab2fcca566a930dad4867f61db5e2145e727f8e67de29f353ea1c3e7f7a70c2aec307fb9986465702d21671783cdd0cf073ef7da92ec0f5a29b62c3e3f0ac7b56b2cc7d3a76f44fb326440564a9a88adb33410974d45c2e363c4eaeaa240e99900e27db166fb8c411bb31a437e88384f34d957b88fef45a9b1b91ed2b911851c53aab2a0f43f95c1eb2ea3407a8ebf93116bcdf5a144262ba4334bc902e2aa138cd65198ec00fc40f7dc88fbce6f80c62a0917780b013b7ac9bf64679b02a7c7d3f209acb01c55f90ffc26b0613061d2ce1ba73e89613c2851bbbcb774038903cf1e2c4ee36da640266b17034fec8ba8818b127eadd717a6eade9a7a13f21e9c7047186f66dabf3d39b8b5640a407a0cace9e4c0521a622559aa2870ba2c896115cab394cefa2e6e928b8ab6daeb3a0ade7b8b2f0f502eee99ecad88ce213f73abcad700dc6bf1e8c1f1fa3c579e8c04ed15a7bc62a74cbf1de1dde6c8804059355f5bf83df7b9660fc01ed174de47de41346d461c00cb9066446eda9c2824a4e5c48da2aee375a9f0e7da4dd11bac300a902a7984a5644612bf955e2b5423ab43deab7b6d350d21665ba8c43bb98f934760f3696fcf6dbffefd5fcda5f57bac3d9f159185ce2a96b6671563850f3f3f9524bda0e1c9cfdfd236e0a88749fcce17f6ef49a48532cff91ce1c40e03770bc238a4262b82ed156f58d553c969ec7ab9b315ecf678c24e4b1d88841f22e32c67930c2373b7fe4c24d72448af79fff1246056fcd661125b6e3bb4c1e6ceb5b789bea4a6963ff5be52c2a5cd35d8b3579422a7171eef7cfad312c89a1e9a66b7b72f41d120bc4b791c9b5b66f93fe51b2303ea33b63f6f049bd32b79f7d5f8d803adacecc723cb3ca6c73df0bead45f938fbe52d7a200224e9495952052bed9400df7e46a73322b575bb26f3bb3632d11e03e97f2865981c30efc040d7e948baf6e55cebf5fa396e765dcb4f4949abb2c240fe6d742421d78658171ed72eca52bcebf67d3b35726d5f4b00b053d6e0ee3b4713e4b7fe3a221ac46165a69f78ecf19ce4452adcee0ba9ca4da3c306757092b981ecf27d10cc45d630006a5193c20f470a7a94c8e9d53ed7f0a82a39389d5967be0d21c1a66d4855f006c3a7ec80ad861d2ea2e0290f7bdcafe9f10d5a5e6927667acc81c2916e28b8ce16421c8e466b9f7cae9168f38b2d86de33b771db04795b863b8d7d9b554a8cec4a2f2bf3b9d7e658a6d7acdd1714e45e01e31f38232bd52b1131291f840c637c58aed77bbf749259cfae6760c17309e72204bd799e43bee9adfc87b39555ada5024350534134957f4a55f206dcbd192a94779e3312154661582dffcc0b612ecd96dd87fec0732d861bd83cc4d321ffffdc52005944736d1911c26389c60d80883c41c84203900bbdf1898046d0cee8ebd9036a795c8194fa721ca3c12c6ffb2e4401a25a875512fddd701df691c8a761ed4e675322adb28bcf78eadd55a9a77c79bb83132ffb7092dca75c97fb1474b1a9cb67f941d5b07257b78e4b2e830c28cc7ea00f3b36fc53c11ba9886236bd028f54cfa7f4a1bc71a6690dadfa0230cc4b39bd8f454875d1656e2c20e6d7ecefef040e78fe08a3785ff29a77f89d0185eb3e6666f666c665edd0723636de2937f1eafe81cc8308ca2ccdf48deaa10f6112cce47e4f59e5071182313b2f5ede4b93cdcba7fea47da4322451a1700f5485b8f44f6b824645a9b7dae4d595a00e1ce4684e720bd19fb4640050703557e6ba54079efcb5685dfa84b52468a7b1cf3b175ca54dd45cbe957c160decaa21c161a76bca4a0e7ba6457c3a00a79e767c3c4d4a81d0c4f13be0346b95859024d44d1ad51f05ac7dfa8d182a91073e21b01c7ec4d19f3b9b15e403afcb16a86eb92a1319fc734ef1bdef9dd35e4a902bd2b71c619ff4beb6fae0a2988e6e514117adc0185b1cad6e0c32a0cef53b421a28d3dabca62d2e982194d57d2abeaea3f20e74c46d095171a8b96e71ddf5117a6a1ebaff1fe1ba96bd74a2d3e89ba54af70e4e50902ca0a90906e40d8b16dc432f63cda0ae5374aeca74dab6238e7039d549f341bdf3f66fddd51c5c287c86e15622a6a14be1f91b8a58cd3ba46076afd83b256239a8fb53e0b47e3134357c308a5c7e7e853bacd5c9bff50456bcb86f53c6a7ed0a2fc1a741de0ef4935cfbe1e0a8b1568f4998c73a770a0aea091199ea4fc14fb1f5e83867f321a059e06feb773d6a0810a416b5fcd84bbdd3f097ac2707a715cf7f358b3f20c25c638cfcc27463c2fd1f1d0481027d71fe450312adc30cdde504e4fcb30b541f11f8a20f8cc33b5397a66579c5a34b2d61e9c29edb0d8db4553b0371b96fb347f6db3bbad0134ea8dfd257c216e5a3961ce570923ed258f24b615ecea983aa761e1a75bf2e5e5f8e98d308ee732851497536389183d9ea5a9b19c2f803a523ac4c7537041a14a7dafcb84c4b544e11b6e45ca0bf3efc71f25c55334984213899d18f7e629681fd98224fbfc432538abe05b1bae06109887922859a824e964443d58885238f54fb477abd8792bb8df3c42767a2aa070ef8ad99166faa8da0eac24c242c02f61b4407168aef15365c01782e7669264081cf09fee43f3ae0c33acdaf2bec050bcb3ab933813a029e8156dc8abe8332c16f25b73d8b99f806faeb436fab81e1d39409d5063b070f395a5bef529a525d5f1913e78cbd091f692b3bdd029cebe2eb8a4c977f9d3f33c9ac67f0aae96150bdf1be6809d867d4c4743b45999ab032c0225cfc01eb03e6e38e20f0e91ff57f7c67cd584ff699605a52c989ffde8fe0f2a496eee2e0f04b3a77ce6d35ba177e58cebb154d9c562edad5c38c6e9ae491fad5a06cacd381ea8d9d2a97f2b9b0e92d850d54b874188a7d3fba76be3f664514f7a8f0388b7973762bcdc5b4f6d4c20c4ea809af516d51154e924706c8714f800ae991b574f560e1786f503ba8f636d4e00732977ed34e38acc5fc4a9789df117183f69f81d3e3aec10aaa83053e05edb8363c900df9a59b9058c594710d5d33cdcebff314cc638b932ae3229e75eca95fe218d45e2ee6805dbd3765db9d09978f709707ea31cad79f3290d4a32f38e6418257f94af6376d79226d34ed98af7ff5e01705e4cb46eb21f86a9f75ff369b9a8537c0ad8b2871bd986fe181e7f702ffc23023ff6f80f1b9adb13a5d57816af99f53e715cafd5cbbbfd3965d2ed9e42e877f9bd05e416a52d27373b923b9aed3bce7283efd81919fe62b936bbbf98b1dd91ce2503764ce8491b253c8dd451866db8654209a6930276bf81a765e3b1414554d2d746a5302be0b5923d2cfb5cca6accaa34e419f37bb9bb1f6c840556f453fd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3e3926ad227a6bdd147a9e2e8fda04ef97ca35289a4c1c1fae93a47008add99d1beb72365b4d3d58621193aea6fca67d9a4b86f3f4aaf81fe9d3edc006ae0aa0bda07d31dee88f0cfb06d01d0ca8fc56407515e9f6287143647c08b252ca4b1fe7b99158ea26dd702f943a6ca19328aefd9dcadaf209ea6608ff31e3978bdd9ce35d9d27d90a330a03018c068e452f3f21eddfe02193ec6c92786c9b59896d68ca5dd67c1cd4ba942c245f2b38b58ce08604fa76c698298c44d3c3875112eedf3203c899f1e036beb97781ef9d553f09ddb9502a04b8c6db87265db9d0ad93bb6d97222cbdcfe21ced8aba2780bae005680f50aa2428b75d036741b87b37af384cfed8a121edb068fe4aef5503135db02c3eb261932b4b86d47a7106d4e045c47cc5da688d31f68a07fe8c597cbdd5507a6186cf4ee10b2d86e28ad518f8607253b50ac75073797f95fe9a2d02e62fce14f26a48872c922caa33aef2212217ce058466569595ec3b5e342cc85f36a9ce6c86b37085f28eb6d5714d9c81ba2a69f50e4412852b6caaaabc6989627e96859703a72f0aa79f20752ca2dcc0260413043b2109793e433393daa53ad36727f9045a64f32b2c3c498c32aac8d2d81ccfb6de4576fb24a70226023ad1d8fe78c241ac91eaf3f1e715e9b7a24294cee1822d0cb88daec4c84ef9ce67e637f820135a1f664f24fee2cb94167014814c14b896c6343626ecfac9bc1bc9d0c466ece8770dad8fce19aa80a70ee3424b984c5bf1511b29990f534d58c0d666a4d20c13458d862f31be3e5a73aeba908ed313a003cf18ca42f1a6efb42b03f7a2eabcbbc87f2ec6159403690b07bd35b9cc3439fa8859412bdc09a8fb26e5a36a5a655b79b5928f8826dd787c7d60cff6c7a0d89634d9c67b0e82c1f7199e76dd21129ed2490d8113abed671b71daf9dd2c3891996369b74ffb2edcd98b472c01822f92a81b79d00b6d8b45f6f44cafa3b590a210696cfaef2528d19721d02bc4fba8ec7530489848ce3a236358c91e8c1457b1fef160c737daef503611d9a735fd13522a16e4bf9b3ac750846b5d41ff77aff70f27655b87f8e0c495ecb7bd314fd31d05bbec2081c360350d2d170844d68aa3fc706f0801d936c6ab707080d64b3dcfae42ecf6c615b44b27d8337ca72673245c09fe27ea24c8d9b705837403e279c2982652d91985fcdec1a8566b651c74ebcdb699f26baa84c3a29987beece313daea3e2dc86c2872ca13ce0429a1ce660bfae2c3d7889de56e6abd524627b4826bf4554509094b010d247442428ca1108950410a3a657820b2fd7dafaed0abc74aab12c3c4e3001a2fd4b16ba76c7fbf92f01e03f9ef4d967120ec8fbe3a8368bd7b221520fe231dc2cb0717a3124c3a4e3cbd9689b4d2c11e6fd1be9d724024ea78d2871708dd504efb741d476d7be798c65385cc348a64e5d3a5d8705006389bbed77ceaf0e3fde355c20f4903357113d136be626498179280e8c6150ff30559c067bcce4de23f813ff9f4ae594c301a332fd4fecdbcca1c3ca3530537b96e22a5a46fad1a9bccb85f0b75cf2f86080e3b041765ea240c4dffe650b00b84b08dc7b40957573e26bac585eee30d918bd3b165fd91952a5bda6f24c0bdc98a40698679687fca7144e831f83246da78ae3f3d470b110445b931db8e74cdcdfaf7e9ad3e8c0a6dec60e379965282490a24a8eecc4df1e46ffe6a1716986c90226cf400cd7db6f71bc99b4b8f4fde2546b1c45c45a534d71055d1c2498f56413e93a2d2cb6468d7c765d421c040d62fd7b1e764eba27d6621791e1fd41616751d7a1d86cfb9270a4c54c70eb90e899721cb7200bd1898db3dc4a020265b3e83e6b1c848d77fe5a82388f5ddbf289c646378a9c3d58f45925c6445b33739cc3c6cac6efaffe3807a5c595ae566df087fa3975df347b127f8ecba466b6936a75f2257deb2c0100e814164e2c3ee479a63db429a028e1f1e235549a377ab88057218a02d5a149559502bda648fa2de891a491c09d72fcd8680aea2fde9a83754960579bd4f478c704dbad1d2ac4c73bf200dc7e84e7f994d43fe2f74a70c52b36a95deecfa1c5663a033da1ee81a3f41cc3b73d88b215c8716f36281527df84c41807d17224a5b8bfb53620a3bc67f9e2095faa6c05d86cbcc044db25e751a1bf64d25d487fc97dcc95622d174f9cb11e1e306239b16069fc40317bb43cc3346eb06a726836c4fac80705f3f9380a94e7eac43b23165bc380e7b5a470639e65b89cfe8f0301718cac502e2f69c8c2bcae2167af8a8584cdb0f0ad7cf7c65e527b5da198e4ae77c5e67f74bc36b242a3277cfc49e80e22f33a86ec2ab1c9783c6ced2e41995c2e1ff6af7d595fce5b18c1f0d7f473b2b3e130ccc5d7e76026b1c475f5f0ef5729a2ab2539d19613266ef3cf9b89f1aa82b4d3041611a677d5239c37c1c60b636d24aac67dc425e726886f2f96251be5eb85e6a49eef90fe65f3ab97cd730eccad39a26b39f30be1b9c033949c14ac368bac77b51d81ec815ea6cfbed214229fe9ad8d2ade245b715ca74a9b6bce88eeaf1334a47d7834bad84436bc815a45f9efec76dc7f9ad0ea11aca210f83632117256302f8ba7801a5025477b76179a7b7c7f836abc4d630b9aaa577517f926b00be00fa5a537a33881e21f99c446316ee31a9d4eaec4cce92b6c4045531fbb3785bbc33c90a17ce5e546f086f970bfc7db14a435405b63705382d22ae3fa1500519eadd7213a052a59f0724b894e29bf721054a2d74cfd0930f9054eb6f55506e06ee7fc6c555c3ab7a36f681cddad4027400ac4685fc0ea4e8f2d9eefdd029e177ca2cfd4981a952b14cd4a65ff763d52f0da6ff5d79c0bf0e0dc8036873148876f9cdf2a191d63b7656f0c227e3af4bcad374d4ef50f0064d9def7d91e2c3bc21df46d98a94516d908b1557990a9c518837952bd9b3a080c6c8ecfa65bd9ae199e9cfb03edc744aedaa22d819375665c18a8cba01d1e62f882861d05930c1e86f870a86d504ee90b209a860673a772991a354131c8b49cc48118cd32c4d17ad5bf94961f60db6b5ecae1604bde8f5474264b738d205581f0f2ab0b3b0d6b433af6eb07b2e1a6d23f83cb305ba8ec83d3d5e5d6b64ae9d514fb8908daae2c68b9e44da6504edfca2b4c65b6fef7dbf08f04d12ca667b48b43c42b7313416f6e72f1eed57587a91adcfcb3f20064ff3913959d2d66edd531779007207f7e063ea6d0816ba2f1f7652bbadfd6d2eb8d3894c2e5caef3a4de024e23a28d6d728198124323568457aad92a2b98820a444402520266cc8678a46c0f5f725082400ffa81d2c482873038ad81bb2f8be413e39a936841fb7e65308d3109229e5de54a391eaa1346c700467a4bfc329306609ec38bd952de598425e5d78eb34c64b7e24e31729ee41738387246dc86d9434d4a1e8712ca21ea1354f0c12c14b79a856a383268a3d6a22987806a5c441337850ea31ee4a1085a61ae957ff094ab4160de37b9a1c61a89ca5e2a8d87fc28827dd0cbbc6d0e18346404725492fc8998fbc671bf8a0dd311fe13a00ce80260e1401220d98c96a9a014a19fbbfa3d9544fe500c4b2deafa52819f518969d9cee9a0e1461a9c1a5c9d0b2de05de3d8afdf3254c232050d5557a698495320c202d9f78a7f3c7500742f2b158a4facc0a9487f116c3bf48b0c21782bd83459a715a44f23fc77b16554a5b6ed57a09e8484cc2f095412387832b4ba1c74ed27cb0c10ac8d565b785b49e2413155f3b8ab81344a89ceb8770307000bdceb718b48339349a7ad4449961400eddbac9d4aa1a79fa2e7b4e0d561194ca739b618beee63a5a42a87ad0d3f896292a5319edc92be2517124b1576e8762768ecaab5336b8571edfc53829e11a0a70bcb59e6610c87a92fdc1bb29247b8a400c90fa773e1983f8ec2acbe84c622f1310f7d95157b3861e3547ed6d32df37571081bcf0057addba8dc67958e9a5a66d2e4f53b38e8e84a1cf41aed9c9e61f24bc3fe9f27d4d7b121d1aa14705b55176accdce4ff76bcaa38b19df60e5a012d77b453926e6ca01282153f3533396a6daa201f0c4e31995c0a92598e5c94b5b15cb036662a4326486175b13d893d8f8f4f72417df2793539a462b261c54c94621dbd4dd60bf7a97c917601492c96172cb394945fae1a213938ca3a2e9e0b6ff886b8701385b31fba1db4490c013ca7a7f4e8af78a263320987287922513eeb8558d11f86f5d3cc514ed5823cf680c2631fd5b2916a96481210a9c8b73fc31dbc818831b188f492afeb6bc66b2c34f1ce5d50498148ccb1fbcc634d963cb54c9c1f8454220bd1a56464cdd800718992b964e68bcd90181083ad0cc9822ccd58efac426eafdfc6a42c6b9fddfe3f0870e3dac20c194e6b8bdafa1db3913dc1bf6607e1aac58b67fb3cfc395eadeae17c3470fa7a8d40f1d790e466590f2fdcd9a1ff2c29173327533ed8e919512a7117654110a5420e7cefb8fdbd1510f8eda2a643e635a8fb988420f2c1f4f44678205403a60edd84b8a4fa2f13afdde86f058efb5133f8f3c1048def33e2a3c1e6761858575875c57555c4aa8ce0195208db30f92a2db1efc8c0b0b727fc70c785ccbfeeec93ebb1efd64fee9945c7dd35f78bdf167f71f1b5c48fff58c7efe2f4d171a670cfd636581664a335e205d7e12d0284b36400181d40e82e6127d3b64f9d5d33841aa85993d473153cd380a476938dbfd273e1527486158c7c3d81b57cdce0042863b73a4cda67891adc43ea0550dd49ed533329142fc139dd41467d31ffd9e54ab1d13fc6a908c0298163f879c853283180b9f69bbda13daff67d6feddc59fe9b76b8ae2f0ce7969a81f1dd25f18e1cf5272ee4de7f2dd06aaafead2253701ae8a278144a3177495ed2fc56282b0aa6ce8f5397fa04478991179660dd67e5b476f272d3b2a3452b57d948d2d59d3c9372445c7d51b16ed543c9b813a53376d51f4183b1548a5965f52504c2d905dd97ca64d93ad531603c8b8735ea4fe9c301147acdb5c2a2abb7e8dfb9d15e4c5181f20e5dbeb55fdc081e8dc0fb681e68e0b66b6f74c42aad7fb0ee1643acfc17a090da15389882aa3360d5507ad2d326f8783c00c269c1154641473e7359a7b658f62d4ab69692598e34be83a76629493fc5199bb72d58c37b4deebe7dad0a66ff1f1aa8b958eb27b66164bb594b79a163fb97e0413d8e83e5d5f112ab843f0da3beb506925b9e2ee48020b45bedf8d55dab67133bb2ed51b54decd090d5f8f17a047bb9818341df85cd429cbf7f125631ec345cae49d03e281d5a1b1079b1ea3c8fb22c83e155391be8e9a0d718f5d86833e9bef401de8694b92beeb7fe783d18ae24e2a158b2221d188a871428f531a1773d12f0306292b582d6a49dbed208a5e4bb391a95beaeb6a1cb8bb5126974e730bc5b05f5bca71f7bebdd7a26da749c3a3b653b17e292d4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h80fa2ea8fe57f1bca409e54e4525d870746f56c64057f063855deddcc6b2e07189103e3a097733631b4972993e666093602a158bd0c9d431dc29e413dd0c8dfedfc21ebdc1fa882a6388c5e02e6d59e05f227cc1d82ccf958d4acb18f79095cc98a17cfc0e76121c6add5f8e07ac6fa679b5d66b5b615f073195b25958718f36ef9884b4958539f527823638f449463df4e6494f92fdff73e41a542df20c90367a9bde8eff7a1dbfd94761b28480a36a18e2a6a846965f11c8c7fbc81d671ae2c720c6ef2046cd4ec5684d7035a16f4a85a4950eb9d66a2dfd3254bcd9383f29c9826fe86f39cd5b029722f1a19c0c8706f33bc78c8b72f740573a6396d839b1529e582ce7ba50f75787190f1ce0609f09ef822e49ff523a71838490f1a61d7170873baa47a155dc48b67f75f6e96add2e4bf14ce097d276a56ce0572fbf0e807ef086887c4626af6cedffb9b138316320e6e7456e3749a778d523ae8a7f75d1ca98230e51c9e15b78f4abbd5de84ed3bc699f916bfb0fdffb4e61b9e0885746693f39351393ff242d6bb5295342808b0f004837473b4fad7707356ae6cd727820844f8e965fa527796974b02647997e7967498f1a9cd4a2f221ae4dd657aab7865292eef94cb7a70cd8f8e308c971c92ec73f3c1306ed79e5e5d754e34004cde86b63958515b9a8e988cf0c23aab93e92af69264b64e13fec97045816bb25883c3a40a7fc27c9b8d91fe76d86c6df18eeb92b6dc23586d891f8c9b8a2d63bcca98c1ad8c0625568f5255f4811a6c175f7f06ce2a8d52ec97d17fa2abb8b57045b62aab6e4ba7bba6240a7cd151a7551bcd109395e3cebfe8115865ba212ea33e07fc5530e6381c8be562471cd2d54035886e070f770a0ee1cfa5d32696bd4c1c01b997498650d959157617d48f39750230ad1a0f4e00e8b1270be30f76bba45c4a3e809a409b075eeb34e790fc85574691f7f814d5b4e8e290de25da0d3248fefadab42806150981f453530192eb5c28d7497f8b06bed72608543fef94043ff3b70206acbd7b11b6a6d376a1d6575e8068bcc409e691b8e0e022d510610624e1bd7c92e540e317eb47cd3e7a0e43e50e59678a1822ba8b6ad43064f9d1d6363e235b590efa0191b5fbce2b3cf1a2189e1f3b4aadbb77ec34d891222c7d17f0d26dcc5b1326b4c9ce05466f424136baf6948068ec85d41355292117fba19c11067af3e8e500066c472a6ee0cb2bfc41f485e46a3bb4c8fe7c16fe2abbed8d5fe9b47cc6ab118cd98c3ad160135ac8dcdacd94047ce0c946d5c809edaa4ddb94e42dc4d5854782d84da4a0963c9c9bd3a3314b716ab2f6d5052926212394d27f6efff80aaa48eb1767046f491cf1c353bbfed513f8438b6734eeeb098f726f32d8b5ac26957078d03f8d9d9d5678403f9deabc94c1d6110ec111b749dcb9598d4f95c06ed7658f17bf648c18abd152ee1815be157d5e25122d90f376f350876ea1e1fc553f5ac38bd9e27dc06e4a1a5917c6523bd1480ca43a966077c486d4074489a662add066df176482d888db4372bd87cc447bc2f45086c21992752ad17544ccde57045d9739e2d25f8edb33a426c912158b12c3341be1dc3e41e845f78283176a58730bd64857fe753eec098b73211dd47dac52e0555afec30972ce1486fa5a36dc4b3e99e3069fe922d36a856ef0d4ef9c502eb04c7cd2edadbce2b16a37f208ccc3e3fae777848998d8ddb626fa2c0a9edd2d13192d2e6a148fe219fa3b48c7365dfb588c8f0a94c99764ec979c00a1d7813146f4d81f1735cb189e728b1b3c8ac0e3585aecbeafcd030744e79d9f86bf286b5fe44eb5d2d4e5503c4b723758ffe4c44881f61bf77bc9abbf90a770de56c5245642be80e0d4d9504733f51f77d54aca8fee23032c343a89978729d3562be8416587035cff34cc2e6b04b51bc750c66995cc21c6c1515bdc96f079e5fa269ef761b233617dd92f31ccd890519e38ae2e11392d94c5317211c588f2279151e9e8a64cdcf88ec09000d6f8b15fe3549b91f6804c77f8b85dc4a5f9d04adb4c179b830553d38367d1eb424e14e78e518cddbecc4cdf31ea2e39daa314633b0da94fa2503d6dd6022c44ae14983bdefe52a209479eaa6a5a38db832f8d5917d58293b01220faf8cae76d3141df63677f94eec8c3b1fbc4145fd1c82e23eda88a4a8e6a81c5deeaaceed3c68f461732c20ca97ed7a0184dc69a1db52525e56bf6e05e7e9a7545154f9afb942f7e754b271886bcf73c5490b37d5629206a32a3513f3fbacabf1c25d8a2ca06425468a1458430e1dbbfa3f3b295e973b85e19a3897cd618342a19c63c9af19fff22285de50b71ea4d7d2d5d769704a2c4f0216ebf7e60bac86d4ed76bc98890c1f7b2aeee429aad8974f70fe2e591d680982a2eb6d2e0f2463681e611ccfdda662e5743a8a77ad41b0ccc8ca740912ba26f9e87b5aabbd587ef8c81dcdecbc5ab0a325f80fefbd33d7df199f333201ad141defe6bd87c6fdf6b67d264883291b08b2b20454ce2e60dcd0ce2407f2415c0430675cb3c394c523f5b71c7e4c6d787559d681837d1be212a058a9b405ee3b31d4846a98ad268931dd50dbc6d5107e8bcd180c8e93c2edcbcb7ed4a5f61af4102eda418abae8813e410cb405c8f5e95588dc60d7471dc15ffdcce55f175677db6f751053e21b8896a2225cc2352845d73ae34e860a1152a4c296d9debacde5e068c8b604a347186bf94533caed2a297ec4ec6b1bbf1bf68584693e3dc2eee671dbdf7bbf7e093d406db13e1c49d7edfb801a284ff5ade573abbd4224e8bc7223c8c1d2b3e834da3e8b5710afb3ca2fc235f69d0969208e44c8c4393dc2c89bfd4ec0c784f6e32cb99504241544c9c8bfa1052f25340061fbe1523d44b642e7af86e1d5f714bc1f48eb403ce8d2e3436b84d3eac08be7ffc7f3ec087d6b1b8c4248b4ec1321946dd183d8af6453eac19f5b1b0d1737952d6393d15e3e23b91c46eee1b0f368887293a94cc0d9335c9b7b581842681f28add5a26bd50b7ca5f0ac2eea2155cee1a7dbc2eee6e8c66e59044802124a17b978d244e1193f2c0658282ad70c5929689a2953f77e9eb7e85b9912f301143a360036911ccb5e8a617ef74e521e73b5ca0518cdcd5185984666522b5f0f1256681ee1846f9edd1dbc6045270649a4ff0e05042b8196576f034f17bc46648c6c0c341ce1b024607d966a1cc501e15a1cda8a47501f88bb1462a9a602e29771d84342196fade3ba6736fc1dce4977c8c4d3ddb664595dcd15137c2523fe6b1efa7c362b0ad7dfa38a3b8dfd21b57a55377d3cc5fd52b7471280217aa42d8a4edd3dccd75771d5d1faca8c73d999d7f42c60e9a5bcee64c3d2b2f79c3cfd73bf12531a8b8ac7916fc1a1e53f9a2bdd6f48412c62f599e8d2175adb4740230350d31db14bab2a1392800463440a0b85e784616f039857223b300ee542b5b2b8f137442ceb6665fe8ae0bf08846fa4ce0b253c1bce1f32f923e8e916dba9d25bd7bc285a4e1fd8c570d5252280b2bf4e9dfd5825671799f1be9916513af90b4298bc5bfba58143c8bab7fa45b64f6ef7775812c81d00ff7ed70b486c3139dc70c588ae4dd5722ba63a5ee13562742c8e49c1e659e898ff913b311645dd6b1d27887b43d1587d68b0f7a5053dbd396d6e0310ed930b7c54e7f0d58ad99d99798c74119231e12b991ef3e8719cb3afc801c22127c32140bbe749aaf0821f37aa71e1689faba69267914795a1bb96cec39dd378b892afdf5d2e86d37e700e89d2cffb8506a492d9fd7fe4772bea7b3a7e92bad46d5c38527ec18be6f916f9f8aa616034cd5d6dbe12498b01dfe5ec2155734ba32f1660cd2e836b8dc3af4e0f0985b970629df857e2a7efefb8dc7876d71e74015d0d303f2874cc76d34dba655ea581ff1a4c8c659e741b7da0b014cd6b7166f1617ea340ffe5df196c7c122eef197d32196f4f0d16a9eed7af1bd7306e7c4205dfbe8a73e349117eabd72edd5554f3cb8986f2bf5950568760975a8ec6c2e13d2b74d8f50c56cc3af8d682b7584adcb265163f3e6dca9ea1b07f7fd07aa50cc5801439062b32282446d195bf5a4469c65855b7b7d02024197dce9d015c3d1cfc3d5b0611b12ea5d75ebe9826651297f52afb9830beb4b4804ed0fe800c09a6c4b2cd2c1d49abe6d40afc774152b972714e4460a7c8a974ff26665c2a5361d3e92ac16531a8e42fca2f8edbdcba335f58fbf3359dee27ffacd21e236fa6973cd83f608427b1f8aa512bf7b055664dffb1208ebd20875b7f654dcc655392e9827193534c7ca88f5a1296e1d507d66762d9b64bbe49f8db7ac1118ee84bbc8f19ec9421fb8907c32813426477990eb909e161d2daeb5e005f0dd30484979bc96ae8353915063fa06c46986b892d05c87d10ab03b1bb9606d61c1628a40bec4665dd9f6d927fbbd8d32ab6aeb4a9d2c16caf239a5fe55f9f138e7102b0c3e08792270af0adba5e99aae128242503c96053350df82b0c5b5471114278928dd538517d67f204dff52dfc052bf57530e2f215ffd36f2205eb8bd60e76e2b0f9cee9aa7c2a721a252e7874a54d54de6bbb0ff0c5821e981a58474a5182ba9264879897f70243176c5ef9a88d4475655590969a94dc4b5c6edffa8d25799bcbf8adb3ca8d9202d324895d5ce91fd19c95f76ea33aa62649b0f6fe14f20e05059e76e346f88846e4a38645a6272e163aad8d0fe68d51bf82c2c0766d1e98abcbf906864b16a646f4f6b6f246b3d393aabd785e2419c8ebb8a1975a0f86f6ba02976f3e79b31c6f9bbf2334eca6c0c77bcc5e5e51d4b664ad611c0572d275cca53ecc2c94bc095918c25a973b2dcfcee6e835775e9158aadf555fea23a419cadf05b6d044a158f4a16d7b99ddac893f406a0e1708a612f562883aac2b2f4affb696a963ad3daa351d9008e8963c38e2cfb4aef79d62fe4069e59df98b21847c99b3c14917351035084028d214011f51e9324f64bc9a363e040e8d39b0e2ccf7758098e7e0c29800cf9990f3adda684e9a793dd9a8c2c25af10cae77d2c101ba11cff657007863f24d38406c7725a5d8e3e55b8c6f319a8bbe2fbd45100b125b3fd32a7d665ce47a81122774c400c8a6f8d62d6dc0cdb2ef8c55ed3fa2bb563ca8f1764a1b40b6ad9a03aebe49856dad8a15be6c06fdb306a053908dd81e0948776f1fef8c71259c658e959cf1d88cf2e908a9075f26bbfd73e93a1d7b9d1b1836048eebb3e851cc5aed29592da8f10a3b34e5ec2cbca5360849cc2e0120ab817277e96b6d001f272c281d459d86d327e7c80b789cb16b2afb03a4d3665b9e2ab8d0ea22ab149415e072e3e8f6c035ce9532e5486baf85fe809d8b0fc6210cf288297978b306cfab4bef4c33b074e7e12c23950a3ec211531501009d95da9b577c022bee490a30e35e1d40a73e61a949cc7edc2c58f2509a794bd281f4b55a3f57;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3e8df3fd8da33b69a492798cabf58b10abff208eb034195387652c3f9234f04a5c6479ff87f98eb6659fe55eefe72290649007b15fcd49e2f2cef2aeada2a099bde625076783df86d71c1ea1adf7b47a5eeff4ad60c065cd86bcc31325f74a5c077c2e1d97f744f292d148eadb012cfbacff64d5442d3adb933376bcc027d23c9d21211a909937f382d13022e3294d62193179a53b1ca02838dac2ba8b9f45c5c83a2460675e053199e401e681266bdccb539c64faaa87a602b85ee2421871b1b77cb242ae64321c0a77c52e877ca429cc4d82ba2602b42a0ac9ffcdecfdfcc95ff50b1b150a881b4de7aaee117709c7bfee6c65a8b0c14e27ac8b163519a5e619f802325cdc3361bb2d6bb70acff6da1d6c6f336da1ffd9ec394a3346cdaf7768706df731a37d809825460d50819c26d2f18fa1c8222961a24b44a5912888d84b9921848ad48e2060a2a22742fb10524595bcc260fe4833c6a7378061be62598efb26c719b0d7c40479308271ca904521a73950aa5c6d15b12cac603ef12c8c669ac989ebee61ee0df0fd99d0b55005bf1bb77f10cb41e93859943d64ecf18e522b4531f66eef0eb5cf1e8e65d2adfd03f931ef879cd7562a99b42a1533267bb080135a9f8e3bf97421c699f248254b89e9c4f13f44c7ddb5527292907f9995e6693341effbd5e24526c2b1cdaae9e24ebecd3eb394c6198328eb68cf712c6c56b3e19da547373d3dcf1a15884425cbdae30f03172a1ae9ee65854ec8ff01fff4fc7d76ac3f75987b41494f80fba198aa98598d50a647347cc87496e872616ca7a7e0fca4b221b9fd34d44c1267206975c170d9a5e2ffe74f197cc849eae944508d9e85a77c4e073c051837bee9f8eaa6beb5214e9eafad45ce8543c544dcceb4a1a6f7ebc30073ba36710c58e62eb5d58370d3c7df0d4cff79699446a92cdcc764b8550de2720b0d175f4fc9db5a4838b8dc3a61b24ac4e75ed912b087f139bfcf60a5e247556dc438ca4ebd61722df6274fac5a21d0605aaed3a2e1ef51c66ee586feaf8118565b3b4a92d1af82c6b0981cab32fa2cb1e84e8730ba66b8e0066718d34eb8ce41eb2e02d1e33c0723a1d228739fdb4bf8b4380445f6b3e1daefacfe2bb535f8b47a21ef495601ac0035ad9881fb13228fbeca42e9c57fdcdb0906780b799ff74912a20dbc59f7e7a447dccc99dbdc78c42aad99097ffd007b2b43f9f95a5a332fbfd5d327df6b1e17f535ef3690052482a3d7476657a350acb4c8ffba27275d7a91cba3d2ea526a385b484f91ec16d28bdf481b0652466e7a86aa097ab3fd201a2aa961b6184002f696b52be1fa1085d0d2e40bdb3112fd47f35a7da4dbf4e4dc3ae57440edc835464db399830592cc64d6297c9db6bd37cc1bc8027a461e09c47914db562c567801415e89252564873952b52d1550fbebc6b7fff0cf4530035e6294dc9e25bbea4d2c53323068d1e3fa3a116cfac9d2fbcbfa447072602406571d9f158b8427724c8e59174d78e005a81dbc737662557b1ddf2754324f6061eeeb70443d84134d2f7c1743a5f8010c839a227cb606a400a8a62064e0a9e18d9e526697bdd3f6502446334e1722995a7ab48ebdaa64ea90d97ad9e6cad85a16e730727f90e1bb74470b960f8e9c20a65d8c9824b721b3f3ef9efaf90b2bb8f8b0aa02d01b84a0d2d3d4e2aa81dc253d68556410eba4b253e65ff1bceb67732a9cae3f886579043fb62af759299d965f1835c056592e4aceadf692bc6df498e3a6a8d4c1002bd251d4b3ff1fd84dfc8104cf9db7d611cd8bd1efb1104a52c0793e3496dfc4f175995b9170f8656a2fd854bdb46926585339cacbc2f80142527abd970c2ba4e17264f44bccf54a114ae4b2d960322f8e2693388f20a1100acf5f14851335b0979aabeb14e53c08474154a997817812824edc54d21558b3ae257ec888a9f53730565ce12acfc965215f4eaf7f41328c14c029a6f89a9a6fcae00e6c762de2ba2a7c4a2997666b0c9869b47ac6310f4a622d1dbf89d4345467f50289af314c534e144b0d8d522fd82bcaaf9491c3dbc73267863ca5931a89e8640dec257a4d13035bbf224ecf05060d0cc21a5bfdbe31b65e573424875b69b4b7d4ad3aa92293b2d661b4d99b7cef1cbc68ee7cfb605fde149ac13e9b3ab095e1286ce2a36b78d89a4e915fa3fdc40c18c4186856837f08cec6f0ffe31b97cd383f2a2a1b75281836fb5e07e1131cae5f7b17135c0ce8b336854e91852ceba8d98c9d7a51b9ed22e8240187d143e1ce552e2c1f7941600ded437bd1979166c4a1fc1bd6afea1501d2579d182bab530145c42e3471a339637338b7f7d740d4c312e9153bac5b21805622529320c44bf747db4448cc140b433c0ae1f707f8b7e8637d1b695b49546658d578174ffe3ccea562dd372456fde9cb2dc41903c94926100e2b10a5182fd4b9d539bf7932114e1e2d7a1825b093fdc7512a9cbe6fba5c731ab606ba076fc786609952f766591e50dac14ce9fe5ab339c90d28f417615b8f3cd197eba563a8743f978faba3c7d53c0919ef5260eed0bdbab1cecddf097d71ca78c162d0d9d7e5ac73f7ebb4170739d6322765b68809831088e2bd225e3ee05405b8bb6678b27377e915dcfd6ae8cac482e48e930c6b18081fe9dca76a92b562ab12eb706334830d34c923be6ea065bf54911d5dd89f6748a7f4468f00b9d2cb262fcc286edd389973d2b83b8d5e3512e2faed73b42225b0bc3aab9dd45e5a5ba44a14667d133d565dcf355b5214e185edd8373fc181b1afe70f35e2dbeffef64f6e9ec84e20f8c92a3223e12175ab50cdd8b95fca77eea39b7d438d3bb8ed7994652bdf18def24d1beb4b5e9cd3181afe1f3c487899815de93e19cde0083ce9f1f78abc529bbd20529e5d74c3190b87c07a1ded8de7483c0aa93f6fa1df32fca448e1268815d208efec0e1144e916508420158ee4eea1838324e532b803074cab15ddc013df1030132f459758926a6498e631e08668ac3a8ea2e9450cbd1605978f501572d1acd1e88019b9547d5f539e47584b97003ac63cd10e31faf8fe353bfbd368b81af1c6a2d09150dfd5293fc7e1ad331755a1297b08afe9802d9ea0506eaf859626fb604a46fe65006e8b08b5279316a7706e2977e708130e3c153eb58cbc3ce5255e58bb04acaea4e0a3cf12d1344f0cb47f8e7d58695c05ba15e6f2ef64456fcf6d8c7c5967b574fb8744841e7de8422ee249da259b7b28aa0546c9e23170ca32a11070499568ee357598b8a0afda59595968a6c10c7a2afe7647a3593c352ee53e98b638c46126b5a8321039e565bf35fe0f5f89138af382938083bba78a8ef27d40d91d07c0250dddb0160afb7607cf9babd8ff7ca2cad5abede292e0d730229e6062b3e1aac2f0e3d441cea83d157788d6630c3a6b1269180e3f297c5dee4f81aa9130f2d2c9281081ba3ecd7dc4f6a55e96ce397a1bd67ff5bfff0d6870743f63431832150153df3147ae3154d3412ed8bc8d7380cba08c1b7c2a14cae429eb125d9436949008b283ab6b665d7c229fbfb484b96326d2d6536f38acc9bcc6637c350ba8df2ce48b5ac831e3e6682de12a7ed8b8a63c002baec6c35eefe486f24145a0e02bd294bbab5199667b2e81b528d2d8085cebc3f2ad12142d229f4f8c02d435810021acf3aa6ac7ab1464b3911787f5c37a81f29ad505c136cd601b165b7a0a6aa9916eef6c9eff7a1e425e0755c411458e381b05964de51ccedefab2ff4ed1d9f2199c7d66f82596e448b81a18f845723a16d2d9ee57ca422613eceff2eafb671ddc586bd9ba1d873f5764e852c57cd61b23b7a4536c15c2cfc45485785a96dc198b796631529d7cda959556549fe8dfb25e0b8323b2d3832b91c5861e25d38640e947c1f4b7bd447cef53426f6287272cea46e02472ca68fa6066e2aa84b52e542555b658835d6671a9701d4b3e1fe378fad5dca080594183c9b665073b9a49c41877f3852f43a0d2fd17ca60c152d6b9b81de923b47cac0d27f73f5b78a259b34ce7caa02a036fb279f0267fda7b925baf77333cab3047c845b527a087320938d6e625db0c84105db300c3ea056b2c58129ec7180a2abcf2c17cafbcea6dc01a232f43660719a62aefb570df207c3cfe599ad9f3660b08219484b53ea6782e0f6c9c9b52ba32b9a912de574bd84b4283447b4057c31e045b3ae3a83c7636d8a1dcaa10d57bfe09ff014fce1a6ff779c63e6cec742407d66bcdc28121ad1ebe172abac74676b8f13e91e3e72be9b4f37119900cdbe27ec47293e9d143680ded5109f32b367bec88bcd9550c9900e7594685cc1c3fb71c88464d938363e70c0d59ad20a0cc27bce661a5eed6f4e83e3a84ad57c0971eca95d346a08de225e357326c111f168e9dd2f3f949bcff2df35fb608df747ef0a8e4e8e6156c14a880dfa28cd87bcb519b387b7e875e93e814b4d182239a9b73500936130c0984be7a3c88cb91e3a136cdfb45af37a2a3b3eb532f151963b2aa79be62782593afbc98828a77bcf766dbb767c2dfbcd6737af8780b52e598c9333b47d4d2dd6397871810965819295e3ca0179ce253eeab60afff5a34a4befc220b77c26615f7fbbd51953e149d79d05c31856289325157db49d25c584fa96380052b74a3b48171985573f159fdc41a995230169b42a3fd931b298e898f77469d6a9534b12720bd30cfd29c39f7b509fdab4ed9d836ccfb83c475253565a859640f8da338da8782436ddf185b52c3dde18249f2a93ed8e0208e0310bc59dd939b6fb5fd532ad49f1c4e454a6b31430f31bdb012ab3e0654a784924027ada2d1bbe4a97dc5e678a057bebb4d65f7e2afc74ce3b092d480822e18db095dc17092ddd537e6fa7ba27f160ef759156b4bf6e321310c2b379e9c5ee1aff120020b9dac7eff623b8f0bc7dafe07d5f10cd55060afab722028626583dbc4bd93da53e43c9c323047d08ac413ea845f40cdfe27e7763ba4002581a310e78695634ed6ed55064bde9323e12ed99589526e52694e49626799daf311129becaa7c07a7736e4330ce4c2c7c64790be20ef240c64a3b31a9997741e2f97f336f593486028542189caa1b77bef5168ac04fab678cd6265a4b42d176588ac93291bee2a460cdf6ae44ebccfd522e36edce12e26081ddc08597c46b050d4f8f8e775657f4318015467510ed703457b3228347c083638a535292b5f1f1c4a7a828bad538a6358722302587811af5a10919eac339b42e02937650d9ea04c146b2c509145f604a7fa5e69963a608187f7db4c004be1729e4c681279433ab8c4a2ff041c59009f884856bae6c6e7c81cdca27c9d7738e26dac85d585b16513b34aad4d24e9b3e401a5a6727ab86aecfd5c75f40c9ac6af40c158d6acfbfc4c8bda447a55c8695aaa84425996584c19c40a324bba13137c5ed1bf0b262ba692a31bcaedc4ad0584c653168a9189e07c70b82aa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hef31a845875a83ab0f2ee1b3fa19443231188139008b34f4e4dc256d7e6dcf23c4423931233da9b867a83cb7f8cc319748fce41d89ddc7aaaddcfa2cf2588dc57664d058d318fecd27385eaf0b55bbc00b258778153a6a08ac8bdcb645b621adc415ecf440bae685982ea366d8e51ae9836ae9365d3a1faf393c80ed16c733c45598e30bc4996c40767ceb62ae5cf3e795d6f2fc945717b61666c7a5852d96cef49f2e6ad83f3e40a0a341ecd191e31d9541fd7432cb3f3ee78c8ab63120b8f9d7cedcecd12223286110b37350cabaef3b213449182df2afc278e60cf73ffb1b9beebe28369d1a1b9a3e8576f2221d4298a38a223f89cb9e467b74028339669b6a6e6fb2447751d83913122379840801760343518fc9d96e59aae6927487165e7ee13914999aae7e8547e251b358ff3fdda259a4db321c72668c9cee6a169d8fc563f4e6407c713a2b12af17ba14ed7befb57e2cce4e2d6a8fc1d3b988f8a833524a7fa8c53356b62a184765623dc5fc0edbcf642443e6c2eeab009e24110c15591eac5c5204506b35fcb4a986b3e5408e237ed55d36b51baf1053d9d7357492c31a84a33b48e7eb22848b3e38b073b4786f2060c4146533c060b7a576b1640eef753ec747a789c3b586f647cc15ab86c630a428ccabfef60996feabb0a3eec26535a447a373f05754ca8564930fecef8171474816f2d273c566bf2e451250671ca744834a463ea798bfb94e246606db4f7351e0cc101051676e10212810a157e32b5ba1495e094df56af0e87f2d343d85180fad34cfca2d3849bf897fdd2d9147f1e1d900814ea6a52c39c01aaed4688349ee101e58856a45f05fa3c7c906bdb8041d1145d278f1cde9eaee753a0d1f77aa234874eaee3b0f0150c000bc1d85442800898687474b56ddde761cc2528203022e72e0e9c8029c8ba176d15784ef017cad9a6920d525235750745c65fe3381a7ef58f366cbadf48770480363ed6a3645a3a04f2c89ce24afd7947ab6e78d1e2f8a630e588147ad0743918ec77b1d462cec8c37a3000cf6b6d6b053f8064576dda3bde9496807d1326e9baa87a16bb3da869ee2bbdb6bbad5a26d220a5163011f979ca5858ec893e6aca047eeb2b145c7c019f1c53f6ec280308f3444025d2988baef3d2874aef86c51e4bd1342819dcc7f16f86031477d6c119fefff3eaf4605b02406f45ff2a8992f07746bd5f5690cbce4d44bc29482003e2effdf609f6ccfd94eba64f8de71b0e6b763e4e3f46a13b918a1de7cb98b3da255878fe7f947af09a9eefb5d2b67b201eca5e024bc63b19a6685c5ea7d814d9a87e96dcf0004cdc28eb9a57c2eeb60e6d45804ae6ce1d4711a5e3dd72efff74f7b1e30d260239f82cc5dafba1e3bf3afe8e2c5f14fcbb1ea673c839eed998495fbbd5a44900cda44bd8933ff1d497dc206def9223714d421171df6623236ee23fa98fcb000a760328683711fd59fbb1d68fdae3248f23b9210c8058660ab17a1a344320a9bea4a1685b8b848b6923837a304d5c27570d9ba3c10f7e35d9ebe9542eb76f0c1c998cf15497ac2a58165078b21870f9e96c56d2b71c4ef0e56279257238385b9acc82bfe71575b12ac85d471e91f9e96df60768c7d4efcdd5bebeaf496555214263c2e24a942e4e1e646a793aa28016caba334612ce237f318fb4bed73f8bb4f65da682a1d2747032f5f334dd1ccd089ae6947b877fdc142ad4e2327435cb8bd1bab91c54201b785a2997aca21ccb972399566ac69558d1cdb27f0075ab4666eaf97aa9c029502fcb26115b6a5468514cde87166fbf465b10f29f2e356980cf4f826b094587cb49a9ef7e85a78f72706188a092d15e5492a7b0d48702383d72a51496b8860f0c9c6a99a1a10bd6c24c05d9d0407b47c622759aa377aaaffdfe090c54f7800210993aa29d7cb518e39154b2692227941f8e6e4611155116ce3a62e323550a19772608ebec495974cefee4be79ea9d1c60314ac3d453f6992a48f48053ef3594d2fd6e2a9e33e24395d91875a0270ed28d9e99222231c747d511939ab23d13953946081462e27519c720057013ae910e507922b04c9208167483bce65afd724d5059623b6854f53e43f54a1ad041b9dced51e3095d742a8746905b724ff503efc62aeb0add408f72c499ee8be6accaad9ec8f6e9e535b5f9ec8184353f9d4c7faf4a63481193fa3aca7d1bc2d3d7e99d3c2f8be247bc34a342f09ef9d0b3c168b424fdcca5d66833f18a4ccb01019debe3cedaa9493d4dbffbcf3555ea0862bad9b043b91fbf8716621e5645ed703c3088fb13631f3a5af62010a2108ae358b3f1d4d496d309dfc973fd6f56ef2e9298f8d9e675c20510758c0695148a8b8554b6cb8ac1676127c77fa3317b0eda5af9e21ab0c46b35f7b896bffbf87f3d711dfa1dd4ed7b16c463716f9ddf237fcb06a770561c70403a74cac49924091b855ea838a2597b12175e773debc61841e64f60ea391057fadd79d410d7054079c6b6455afb83ce61a4081772f1b8d60acfce9c7d3f6fb69a36c78b06e54418498ab786eb6d048a3f29b97db00e8cc0261af6d8647e722b837026ebb26be2d7c1cf837b3425e60f64064fed72c816905f5977b245884db4f0e6c295bd564956a261993df61c6c5ec88c9b7e585cdb0b6278f5e18b82cacf60b792632cb45c417889f8cf7e793a193c7089e46a77a2631739c2bef14cad32ca907c0df34745d994e7b975a91697e2f4fc0265e71ebdad31f796645859fae78148ef70959cac657abc278264927a66d046c883164c0368f010df94da7c9b58df7597409506c9cc4372097767de66d90030ccc3582c8757fc6f064e94702829cffdeb9dc155c8ec6eb4092266c245bd08b171591c03bce748d1483c4c01630c4f7c09137657cacd4bba61643cbf2578bbcd1713c0924eae2b76ece0e12fe52333bfda945c38926ada05c1bcad9be1613f4ab92ceff2a449fac766e69ce48933b1f03bb774eed9338a1b71e981b1dfa405806678819e2d94f48dad6e4de4efb3d4ab1b5fd25660a6a86ce1a296a00f4afdab12c91768990adec1881d6dd077bebf8ebb77dbb2c9287d067e851307796b2c795d331ad17d64b3a81d939f32928fe859249625a9a41554caef7ff70eef7a4f1c44e9004bf287098d1cd408d8a090884ee13bfe75067e211fe17496267469d8e33b098d647cfd975402fbcae26d12ed7f852549254811753a96735c155dbf181b761abb8eb31c2a7bc10f6d8520f72fe229951eb18aa6db01dcb057351c5e5b55b53101cdb0674e72467093711e7d742ec33caf659ded5690bd2da23e3022ac7fffc8543289b5ce3c272265538a492fda6539fc70a7a7a3f5711b767c7383a1239a91b33d1aef118b8ed11b1f0d6c6df6e92947b76184e36a59ff83cbe548d65a0294fabb9dd4a7574797294414db8ace9a3c7404af2d31838ab742b2dc44f70772266c73be530b0db55307d646f749b202d993805605017e884407a2555fc1ecc4de8a7f355f32a647379c6f226496082c879d7765d29ae5825eaa5702ca0524ac2f157269e063322879f0753551b856e6a4c8516d28dc39d2b9d2c36dfdf1d28d3f07dcca9f0f8e40fddaa392bdc5b16ed35b7ae486e1b68f80f8cb99c11c024ceb54e08a140e993c1cf9b3f99ff75c6b368e7b82a348ce79ee42ef7023d291ffa955ac41de664895b41be8d5a7728a75855911ca6e540c7d967de693563988914e970c37543ff9d7e61e7a6a09292116852927573b45095d55f0cf1d30bdf9225829c76875a06a60f75086966e0d50c6603640aab405743675191e37eb0cba480883403193db49ca954d7cda277ce681133a1689b38f758ca6b054cbcdf8a337aa10f64ecbd665af161101260154f60f0415200715936a5e0618c36b028757b48e6fbc6e183b1399f42f3f2fd1959bb386b3029097c6977f25e9d21eb6c86e51a32ee2195eef098c3920ec7bee359659730e57675a2eec94cfc53af8f927683206e3afa58930219002334ee512a2ed998e4c91dcaf5fd8f35f82e6cbea84cf316d04419d7611a86d2c493d3e1cafdc28e9a6fc176d0fc4967535720cfacf84fdcefa96c9555625a7853d56f5e6a8af132b78c3bb3b153400ee39b8a8342d7d15276cd5d67121e7ed3834f291e03c37ef8df09cddc1a98580539632e909e78f4d79849da924a980a69453c3544417dcf24a38800f4ac0334336da9b24f8227938f1f61cf7191c6c926fc131189fecec7f55c29bd465db754967905db344f50ccf3e774fc5e73556a64379595458dc36b4403482c880b5fcf9e04153311ec4bd648a58e49957ff53c0d7cc186b47eee4d5651199e249182434bdb37ee81cb7110dceca6fdd1514cd1df5cfc215daa3288dec45855cbb03733399f3d6512e1699f75c325c854a4538331476c7bedd7b2af61e049f73530d6429c0d963f24553a4cf6912ddf4d7abf5b47035a0fa61c06b6fcfa9989394b4dbcb808f9e538d349bb9cdf9dfa27d2b31ab7ab1e23062838c744626a5c98cfac687ef54a7d59535c4cae8e9221122ff0432ec167ca86ab5b08da65d7223e335269218a1c0a8b2ebb44e69516132c11144aeca9cc532eef27e2d7cf4ca7993535ba21bba22fb74e771029bde0c21d27d589ec0be352743d25e0d72e467dc489386c9ff1f4a60af96de07c9b7303f38712411d102f82f54a956264e70f20d32ba62ee776d4951f804106af6cb02895593b0e947815f4e889d3d50c6e3558581d159ab010c883fc0d4d6b2d8081658eb2fc2e3a13f85b372cab93d7cc3a3cb8f121cc87c098e0a8f8ce130cc52c40f8591be3b92f4a786b578e069bd3e927576d162e2d3a9fce9c2d9fd81df6740694a7f24f8c207738cd2d0beb31a1d880504ae9933288a84c5fc3b8182004096d6c66a1e77e6462626fc849efe1d5fdf2c5f2e7736eefd4e6b3dd9777ec69247325cce55d1272afa05ca65a594dbd0c00b42efe698482d5be1c52bedcd345c0f71964b16bfc738e765299e1c5a78fd8a90d096b40865b486fea38cfab1eb8dac7f6319cf970f5a4f9b11a77e15c0ec0194b1c93196f6bc2b5acd9b976ae99fa73266aa7db09c7ee75b47464c0c433b0422db06b28cfa440b0344dd85c760a37045d28386eaf772b00ee4af90647c7ff138f15099c9313626a5c9d0524d78266f41c1a50397a4555e9cdcdf34f07fa4f3e11566a1e5fb61ab13bf6cca4a69cac8c7286ffe089ebf3bfc2da7b22a57de4da988f4396bac532cd1c1ebe861630155b57174f3a7d945a8ad5bcfd02b55b36bd28067ad2d4d700020b0c57eaf47a29508503d04fd660205e9e68d5c0eb4433187f948b0bbcafb942bb7bc71144d45e0cb277b3a81c37e8ff0d5f5d3bd7faee590ec0813fb60efde3c101d998db8b3075b03c1ffb0b81bea8a5ab3abe0d2265e1f6405422eb28610d89e5da04153cdff925b6c306b83f8525d76672e57c9334;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5e3318233b31413c45464fec8eb1258a69fb3d5ed7b21a5e8d12b53bf83dc06131458cc74aa7a4db0695499a214c9932ea55727601f1d01941b28f16ff8e3d4adcbcaeb34f5ab920e23eacad726264eedb965582a8aec933aff3d2e5e974af3cb199839fc8372b29e107387783e0ada87b41d54b1428bf96b34f4bf55577c6952e6cac7d9c1046b1bf7f455843c88bb9733b4cc1189c6eaeab48ee114814d3e20716cf28df434d95b8eb45e33373210591dbddd55ab12be209865fc95c21e8b9064da54332a8fd9dd2c551fb7c808a12614e21e38dbf50c3c6fde4093e50f9d9493d45551bc6a0041f080e32ddc5a063b7e1c78fea8c3bce5cabe08c0651a919e4dd4d0c60d9318e047d23cde1e9f158b0795ca127377d5e56572b8202569e35afc207b014e643f30ea4833b1bd8f39711c889850474d1f6bcc5bee35cb964958c48f930a4d6b51cf08d3bfdf81340d329dff6f6dd8fcee5567f5f03f6da72425abbac8fed3f724d621624fa90454d09783653bd2c49e3d8ac4a87da26dfed96bb73e3093609582fea752d2b6472eeb8ec38da6e38103a4f70862e94db456f004f2a15ef6a898b03c7d672ee7abdf99696fcd7edc040a10edbfff64901b92ee814f9cb8112a66fe57569a9db4cda7ddfc9c69e5f7ff734a6e9195088de74fd2ec45d557e2cb29f96367798c9e141026176604429a926e9eabb14aab8bfad795c5a5f27c8ae6fbb1e81ee2963039fdd0bbe7908ee47ad3f8576ceb7408c16bb6835536382f335831bde2acd08515559de0f7b4e0381c5e879488db07b6fc0d52490b1dcc03c324025c2a66e9228ffe4c51281b0bba3a50080ff88c7a4a354dd7e9bf5ea3ce66dd5b74a7b30aafc3efab983acc2d5e4a3be5108264a72a09d9fb95d241f27faa8c1be4edd486291f63928a2ab130f703d42ed46c0dd23365af2305bc0f7bda5317c0f664dfa881ddb8e35d7927be2e039f8505d517beba7e59108869c4d0526f4fe339e3ec1d310b77721f60f258c1652de710bc9c5d5629a88e4e2997bb56aae97e4652755ac378b3c10bfe16e98e46d0fd727a441a9c6beb08d919385028ba8d9678f21d6afc031a4a539767fa28809decd6a9ac6f3e2f08e8f799240a3047022f296bc43a9009bf2927bfb9536de9376346292de579747b15be7bc72fd0ba0cbcf2850e264cf5ccf5685673693bf42ea97fd19ccc1070293fe0ebf0e4a41538921559408ce6f16ec44a793260690c232cf85d059fd913f00457c41203b58c1ccf4c337d25408a8b60525b56249181cfd0577dd751bd32ce7830f53c3d05e5ec15960eae9040d409853742e18d38b29fdbe651d67abae1e6aa5f809c8cb58ae9ead9371a1879092a9c2854e2e0ffb5ba73a03c4bf231a6410ed31f942deedd4c7bd3c96832ea4fe1c516fda9a82dd68d53b2e04f0fccdd3eb72d5f14abc7a5a36b53934e726839b7c252f480fa59ac5844d5a6fe90fe0f1e2f75445cef06aefcf30b35ed0d60a042ef10392af1520cbbc0a57512b03630d21981e670e0e740abc9fb9f3b6807097143c06bd480d59901aa257183ec28dc9d34f496ff75b3761054e93b9d07c4c871f8b8997967f38e064a77f765e3bb4e68f8158ec384d28d03466fc505ff4f71358aa319879d09c95870536fe90eee9881e047e5db2a4d18bb7f6ea48fb6f1cc606d4c446ba7fc861d8bf752041b57594a5f1ccc16f57a383a0f1b30f9c1d1a22fd24ba97ec1e64348e49d9c5436a395092363bf5ac0741102ed2184e985db00b92ccc7b49a03de265f587ed2f6dc7163bffbcfcb5a363d32d90e57f475fd9cd0f68acd589ac4cf80f99f07bfa4bce734c8935ef5d5eb30f8c7cbbb953570b9420cbb6fab0dc4eaf50fb0d02cdc78c36c67202f556841ede9c9c5388cebcf26acd1666855da384820e8ef7c9ac674263564aff03557bef300b73c9cca229e96a74a82bc8266420ecea0d29fcb2cd3987ed3125473e82103141e3aa6c052f797e7ae8924e53ebbdf832c60d064b13c41e2a189b7815dbc977d3d881369536216f163c4a74e25f2e0a74f9db8a22f9b4951aba502cd67945b247a5bca32af3915217bc6371106854a39723d472d3fafab4ca13480dfae18a5a57d3bbba1db49432c663d7f241c7993198b783a59224f78181cac735639bc442b017148818e025dfb88323ae83f9c3f48db1adff961e37847abedc326db921b113d1cbbbda085a111d13c96f0277f9f9384d9b47735ccaea17a072f37e644f7f7539dc78f2769a25ffafbffd93d1e9a203b3f3f70ca90652e19e1d13086346aade99c90b902791c66c2dc410eca4d3cbc86e8740f8ae4fa9431a6edab3c405fbb65134731ba572db0881566e29390455353321ec2309e84ce9c66baccd07a41257b43d1d431de6c970dba838d002bd0c6e81b93f6c1a6199fdca4bf098208e2351969e47aa4f320c70e471dd46e480b1e4019128a6cf4637885a6ce47351d9559daa0f1ddb5c2b4c8023bfb7c526cea968c6a079d89caf6ce67102b45bd517328d8561a366c0236b3d9a140defd49342eb1b26bdcbdb30b5895ae8acf1f32df14cfbab570a7770e78f80fa87b3c6a6bf1183d2a8174dcf44c5d0e9ea2e80104983b8756c9bc9e558ed3d72f18b65575f90f1e4ab9c30d32fa162c4c8710f5ae2afbac59590cfcaf7a27986c818447a20b972ec8762851752bbe3e4e89ea4961a11d972fccf26f8cedca08778d3a15b1d9be2d846d1e8629106238608163f0581e9c4e8b2427da30b1f4c4ff68ec94f970e03ef95dc2046797c3b775e4f609b74624a5a63ff82abd05383dabb5be0f5e63107bcf3b45f4b55db01e638d9617fa7089676d96cf168e89502191641900b1d3f7985391135bdc2d7c1a99c6edb81281462dba7e2191172891336422f15f064bae453d3e0543d53ba6ca825f080a4da557e598dca42085acd0400c03498910c93a0ce93ddaaeb536f4a018df38dd7f565f6a79fa91bee9c39ab61603533f505f94ff40d6fe40142e2cf2cd75287e05873754f1281ab8d1611501a97c9a46a48bcd36b0fa308608ed282b395bb8ef152f18c5b6851b44ba77c491ced0902de89dedeadcfbd8b67a0cee8d69df423a7e9a8b30ba989ccd497726beb01cb11db31d77c5d0b50ab0a06839fd043f569c9c1223e8b475be4ba06bb4f4186d483d1eaeb44acca8989b819584b344235b8b1268c232a566c502e4f4812103942177c497c70f89f47d8006b6de79baac6c805a5ed3742975eb54bb0abfe52df5a1c9f38b2942b534d75a82716a901767069f134739ddd706a0fe3a6947ef9593ea04c3b2e8d4c08342b1645496696dd78c100ff7d184a302404defda7270652108a58eb59763fc9a0f6e9c50cac15d118c16274c2d1515a6f997fc56e71bd37231aa12c4429dfe1a95bbb98ef5e4a28e4fdb379b696397c06c6799de57aa78b1895b2ec2dc63888a1096f9038ecbdddc14a616786622e066b288f6e5f09aaf1b9a160aef39066460fad3f8a0aaba599becdd99b83503915550534870f15e77e570950218b06592ba6a8f692d5f72a56de40fe454bf900dacb6e3a7467b531188e13aeed78fdf3d1e913185f1101a53b4962b5a77a41287590e9edaf52c88f997dd940b8a5840363d364898aa63965c7c142d147d12300530449775f823c588fbf0075349684a64932c710a0f55482f8602e40cbb68d837f49f43e1728e46008f0e721c026d9003b2992012c9d888e04040ea0c95dd66f3ed73f483a1599915f356dd89ed6b9089eb46f369fa69ffdb8b56c87dd644eceaf0174270d3862ef11eda8dd37dae9f5bab2b47ff835b12162c4bd4a699676b9e84195a8e90f93a892ae77caf502bae19281c02f1fbac46963ff401d8c3c1d4d0a86f4d0a7af22ccc8520e0b65f551028e46d83c65b284ec7550a9dee2a5ee0b17a84f4b50ea4855084e62a8d5e53d1114a000a474dbb5d60d43790797da5ea8bb0fd7487ec83bcf8a8f0531a0387870ad07852deea55e5942b0853833a2313f8c82dc178ea328e4e5b1b0bfd7923592b74c00d337bbc1b8809617cf263ce0a5958c03981463aac98843089987af78dcbf0f6f5affaa862ab8f2e7c60d7858bfbdf0970012e010aaa5545003ad0e3a6d092ab62d0bc6a4a38e0dae97c84e1eddb8c0186dc4cde99772f1789bea6bc5fee105d282ae65ebc76ce1d9188719ce4c583205396a2a742a237ac230513b6c173beb78e6cdfc4e8dce3fa36e1c685c0102afc196e445401714e92b6ba17ebcd1f2bc9e180fdf8f11055107aff5d173a58b6b65d342dcd5349bbe7b169ee2e7d9174631ea890277237f98e3dc206c5109c5c5fb98245c4fbef83356c376f45f31f536ed36f11dc2bdf1c13ec7728efcd6c3122d2b3be1e552a9b5e0723bddb7d90f3a8579d4e488525c7a71588a3a5931db5baeed541f0e2558f4711e9fe7cfae405718a0885e0d93471418edebe95620e0bb2a645ae07b817ba0dc150924a9a8f6f842d35edba66ac2da34633839036c8bb1e2f999236afaa78e025544b0e219f54b96d9b0e9afd07946e671bd6cda2c35a8eefc89b2ef36449fb4c41c25c8baa4525719a5f9a3bc224f24264f695ad37b22a70163b365be12f5d540962d4f59a75d92cab16e275a31f6f19126e3bd03ae729f5b9460747e44fbb264f4e2dee8e5fb14aa115b11f21c7524507e3fea48e2b59a5a62d8e6eec3294891404ece3ff60034f3335c28708392b8270c249eba43e7e57572e7ec89106feac9b55cf7ebb61d1c13a2099d764a3afce536688993326c19ec6e391008761afdec90100663d7a5e989d0122f880551b61ac3ed4e28fce711e8287c9b9928a5c9926652b10f9d1e4682c15f1ec917fbce73c8b9ad5699263ee1ad5843af55252b6310f40b8eed79b1adff333230ee38cf50b9846a8fec120663c924ba573dca162c5ca2d6508f7b81a07af5f8cb89d031fa20d8df002829c9d691a495046c58be99f5a956c24440db2afe38778069a4dad5bfeb139b4964d705e4bbcc71946f0c176c851756f0b303e514e4204e173cab138abab95244935475e5bd5407829286ecfec1297c4d433a9b04b02145047579c63595fb8d6acb20076380b0a677f09f2bd30c21bd8f0bc432ed01638e3c676e8b2566269168bdaf4eb61c43d395926ade33bd2748e1d9e65681dd924f77a55764b02cd554020b1137b22b8ce77421fd88d0d3ad42e1f563cd4f1ed7ebc0b385e77352cb2a970586fd3e6c36e1415fecb19daaa2a6491fc04d0bb106879a46be54b03df67a9767f23dcbdced3fff3eb2cab2a42159a9b4e2a8f35ecdcfed9ec1347dc54ff9c706970b653653edaad20cfcf4d72cb5f3f4337b7e1f192b4e588f43025fdb5c3b87a0236f9283f34fa52833987cc5f471cd20f0d4787a5dba156dab62b6b026883e7cb7a7aace983d0432fa2eeed4fcd3bc8bc91facb3360b04562cc3e351046d4a29829c8f68c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h974f6105374407840e017a71357f06517f8c587040410bbe05903c88df4ec882879afa882f0a11061276eda81d8b4be8f58e5be97929444c5f18b672665b3389808c42142826244481774b6bbe783f37999609480420532da23dcb263b38bb757328377cb99502a28727929ba6d0d43011c039a05f6152f96b7c20ccf2502f6969e50ed1c833312f441fb294a8e0a646a4596e1303a47979a75ecf7db0d8693a6ded471746c51465548225fab9bbf9c7301fc34fe0b0813e5b8a3121bb492922512fa6a7b44be7a2bf2c3531256b3ea2755071723d1b85435ece5239d7615838b1fbf5fe6b54a53bc3dbc03f4c41ec39f10cac4b5e3edf820f97e4d4607a09b9a6771ee585d40e0b4f7fbe03c526b7764a64167210fd39cf5c0bdb60d4a59b47c02c1701539e2c0d96c4e7d25f305d2c8cba9f80b6a34e6fe73f39dc19f7ecfd4df93c5593452679d3c641aa2f8c1d05732c04bd0ae98ef20496fa254a056d7f28ee5ed8a28f0adedd1de0978c826f5f53821be2d58762d5879039d0c8b476aa19ba164e0cd89018c4f6d8aa4d884ad12222b560246a058c8d0f8708abb1aad73e3361babbd30b4cfa87242c19a96e282e30fa6b48633eb85e6647d599d889cb84dbeadc49d13b32d051784745cdc1ab548d3cb231f1a60648426beec76337c6d8ac1d54607f163dd0c602909785c6605d18a9b8db7aee748ad6703755d255a24e92f3edeb49baa82495efa4b120d7a707ae08a9f6370b342b3b120ad2388b4b1936fb0b20b5a0607e4fda71d800f4453ec9fee1933a09928e31bc6526b5e8508ae1b7ef4075ef706d1a3f204fa2213af545902be85d20024d0c3e67721b50b8925bb86152692410a7a4571079d47127847c0de156661a2dcfda77e6ef2e984cdebf0703b85ff376ee1b6e116ec225ee905afd5a03a90288d2b8c9fa7af1a1494c39f3b66f8626490035bda021ca227ed104c194acd7bd0ef2b46ad1fd35d6780d639b1787abb354d908928eda6ae6e482467dda0352fc4087f1e335e5737147cdfaadeea7d5255537a60d177de1d64d0958b9b87406828a2bb5da013d59fa757315e28ced058360d690c250db7837add72857c3e7e05614f750bd49b5cfdee5feb4822c002158ece7386f5911b9151c7e306f7af9d3d7d27e940e5586ab08ec6ef196425d0f441d9ee7091a383aa40131dc9535557f360d781bd5553ead910d4a87ee2c72eace5dbbfadec3b08332add703e83a5a241176dc3393354d8fd7a29c997f6afb892cb3bc1ab2502472f76d5c568d6e4d890e04c3887d169aa717c3c958c9f98aee2be619b80749aba99e7026b0d95d947d1fdfebabaa85d251c90e76c33a5a5def73162870f2a068b33761992062c163e5409bf1e04e5c9d83a00b064f7be2783727d8e740d1c93b8f28cd39d04b68559485526e90e79c8aebb32219e7590c8ee353f4bd42a644d2b145f84fa2437ba50c6a8189075ddc537c52f4519e40cf1c0b963c4116a59287b294689686ada728ad940b1d6058f36f84dfd3ec6f00ae152acba1d04ab625268d9ccbb1241a7c4cfae490d88f2779df831dcda9f7cdd7cc6fdc33645bc02ebf0e26b3d27399d54d1415490a5a62909cb0f404d76fbe57eadfc238a9aa4893e0f21d9008a453b35001e67dc13a9720171b3b8760f73cf94b5819860b3747f4a3409a516893194cda322400daa6be7abf7a094b1d997a8a07cae61537eeac3291237ea210289b6b0d7973a1d4268ac54f2fdeacac838efdc5e460a22252e58c2b811e39921f887fb0aa103d4d923d7ff0516db6fcb9e8a28986fb5aa753be5e4cffc28fda8bf041f4637942aff45524ed73218c229c463209612e0068bf9661801b989e339754ca3e565c4472f8d9a60864d9baab892bee8df3c3262ab9a97fac7a954158c3f7075429d5bb868e68a9730a662b26ce97cd4ea285a92a8a63e0aaad7e372f53537e0e75f9ceffceb733087506351dd5491ac2ddb145813a9616a2b559ffb7e79c82f65a7cbbed9c0725d5239c0e513978cd3073aae3d704c2b2aadbc67660570b3b16e78d3408f7e4521a84e6d6c9facd1ad73bb58f785fa745d9c89e059daf261361fd4c224662139b80e070d40ee4844d43d4d21289d8e1941f4db79f9e671a04503bfd525818afc98756611f49e233e26a2054935fe29f85d5b8fc8f6008ab3ef1cc8d42462ed0dc9cd5c32510a6588fe1eee4f2b390bb2474920b8eeddac0a444eaae897ed839c71502ba618df3007aca6b8d9be34384dd8affc156c934e365c099073de7d5e37eec18165a5a12c490c94764f88f1533b02bb0bea91bdc2d4df054a88609afeca1e41ff9766c3ee949f09b6b33a3aa8898fdaf39e824287b22473b818090332a43fa4bdf6997bf628c781c14ad60e4fcca3f030d39bd1a3dce43a83273cb94af529ffdf84d683b812249279e8bc439318e5040414b2f269dd44b60998239eefdaa0d6f174e30235b1f6d3f6a1077ea5f8991c2c7312623739675e05e56dc2530c159cf0826cf8fd43ce9ba07104eef56a4974189b85e5f2f287625733045d880eb14b1e4ca701ff18650a3781643d0005a0229cd3795a3416ec8fa631409845fff580359ccdd90f09a7faed6125683f6d0d72070a5b5b6acac44311d96e2f32c7ed16ab984c8ee340ff78c282060670caa03ee41991c870834e5a12f74d73361a7d81c19bd9f3d5ebd7238cefd949db945ef78a3c96452122f30904328ca7125ce1733342801c6a9d6dfc21ca6a7b1cd0e0f8602b8895cd486dee3191897bfad978833fe5b4d5522fc238239617b02e7b3d96b0b28fa9a4703f7339fe79492f757b0ef3370206f5c393ed31702a743257abd0aed9e1b50975327325ca8b084646659d14d2a0cc07cf6afb0b0928f6778d493c2d748fa2c4d62c8de5212139cff0a5e06f312671de97b15995d9c4e0a1fbf1b41f42ed3d84c065a20f20c62163ee4444b3dbe3a3948e20006dd7f18faa90e5d8a3a3a37a6beef8863a2592225d564acb7a2fde87ea005f53801ead3eecf9e3ffbde020ae395a41b9e744350591b82e998ca5e8faa2eaa45cf9a48b0265830931fa7181272337e47bc20bfa79e225f52b16863c86ecd06d0f4d5595dfc7b88c93208263cb97b306d5ed1cdf6049001eb803a9459c44e3847437f0f6267b8c5684611c69fc5837e64bd819b45985b819dbae1b0c6d9e1cf7267fecb76d48564be1f831f2242300010f9926c5b6bf6d8f0231838947852f4d7815014a3a2773083e341b3fed45a6b2b5107a6abb077261ab2cb044039433f44f0ca43e751729798e711fcaf0f1074369c10742af081a8e9fcc11bfacabb7f44559e753d1b598548dafc9b6b82e96f7b955de41786a63149158dfc1f19712cfde8d7e1d980d5c30fe21478aec710e1a9a679a41306583422053c0c51e456d632c55d1dbfb9ed1b2a4bcdb6f1798db82885e272fd8e00cf9a365193251ed095502984c68de278bd3f90edadf33dc2ec506c249304747f84fe2e0a57c5cc58bd84e6fb1723f47f885b49e133f9241c5802ff3bce148b8b4fb51202ac77b538061f60b2a05295cceedcbf110f695b6a1ca277fa2f8c32c659f274d86920cb7ea9554423f9976b8ad30a49101e2f5968eca819e6fe4f516983da06b5b1203480bbe671fd457adca5cf117f144ebfeb284123b047d3aa0e15c332675c72562202e889c733d3dd7db39948543a49a0bb29cc8b793e64d694ec009d347f0fe43693ba38d2cad3cd1242539128483f9d2d0105316df68a768155af0770ce553b6bf65147999b4e1c598bc01f3c00d90a22f2d6c396a4b2b6faff1d4a5c20e5ce9c3568aa8ce53af0ada9f45738b38e3b32884fbd8aaa9fa89e969bd8eda001e49424ed26cff463e4d8aa1540c0cfe57c141d6d84f19d58f0605aa5f9b47de92c9f9db12c23c1574caf244d9a4fa9e589aeb53dae9f144fb9be717c0310aa461df4167df86a95d3f2cc27f42bc33153c293111cad0b25f484ede6768277f97b6ff50776d96ac1c72840ae5992455a43f471056cd9e33fe7a8f46634678b0ac2b56ecf4062c30a2a61c23c25bf8b5992ea2e3d0ccb0fb1e5ce88da4885ac45a5036ee8f5840988a9d2d934024ec8073a2bbcf9b79109566e61da682f6ae6c052c4e550dbe710a192d0c5d5145002caf03b4a66da8a6b86645e4df23850a488efea001f117196149215d171e578f9b992923c2b1681e0950af01c38898c66f9bdcd0bb353e200bc4abfa189b2888c013875529320e32bff3de93a19a33188ad6ed667a05f946d3757ad232a8e578a17aa877adebd46bbe56c285a90c93376569d45e61fc1c7606aae01c753c03bca04cdd8b76cef3ab0f13932dfcb8ebb212fad737df6e272eb1271ffa6e84128c781cb168510ee8c7abc8908a6afdd4fa328f373f17a55dbd95d3b8b96366502c1411bddbd297560b761057522fc2241d68dc309e3f40d05f01fc1784b9c7ae05c5dffbca1fc52b2b464c5a003d9637c1a4a4a592c036709f176d2f0493b6a291e7969f6e4e0b9098e29b06d92c139c07434b7d29f03807f6dde0167c14e1d4270fca2b47fdc9638c57842ec852390621b23127bc703e3e39b2e0019294321b0d5d9d14ae72b35750bbaad5b92d9afbae04bda5f2aeb93da1ad41b3d2834d34a086f987859121153c67f86e046a91ceaa3aae226322319a4f71bcf78b677101706affd9c0c0e08b2c233bb030be86867758dd7268842c2cd30a5f821ccfbf9b0f0e3718827c249b776bfc1ed8fe25e85d5e93da835f6c28a26cdc52f7c3c86a872c4a74478f0426c28921f7569fdc18ed45d917e601e2e7a4837096d8caa7828bf8d552306abae78af5c145459a150e324fec7b93c2e04cae5f8f5a37e50407d575efb4a00fc2c8b2e8e840d229f6afd07b9741bb3c8fe58c00829a57f6f4720aa7f66f0544c0d764de9165d4195b7eb29d60e23d00d9bb1adb8da3af6c0b173c02d1e8d651693b3e7adfd6e9074a4aca4f1cb0644a5ce47ceb70e536297a16a090033cf196555dabec0fbd10fecd2c7391cd2ec5b1f0bcf6908f1aab43f9b0fa82b9714f0a93786b4da7552665a168f9c1b0b1684d3ff8b7c01f5dc316571cc542f2858214c0e55b99b1fc63f8044323acce625f57d302613b7ae3c197284550a95434af8563c7ec4138a211e143e6a80efc7412057080fd3790f5e1ebd543f94906db1b5063fa788abb8c32661905391669fdc0cff40b0c18433816cce466eea0759ebff8eb4e68634e38b532f42765454d79a89e82c0b36e6272b9b966f8ead39b90de2b257b76824080e045336009a7b8035f6eadc87e5b64dc3df8c668c497f4a005ed60b622e7de21f4f2b0fc2e6a24774f2ef31c0866d89fb360cfd400718252bdfe6d4c562464468a896d4a7a704cd80b8f805e6f8aef50b0a3020a35a0e85d71bbfc44e087e218766beba4bd095b9dfd218c5c974bfefb6a7de146b8a7957;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5d2864e370a128933f24aff52bbbed71ae1e2dae6b469c5daeb4e3784c803965869e4f8ec36c974a952ed3cd28bb1b09a2659c417eb79f33799e7e6037ed2084efc38c4485c5cc7e50079ca783f2e7cc635ebe38a7016d539f5ebf502a8048b6380d3c3219d1735cea49863f3db627603220923558229b8cd5d5734287da3604a026ac6ce4a12ab67c33a052c59c968a41accecdbe3288a126775565ed12f29a2ef9c608bab7537a1199982c1acfbd635c765d9da5f8c1056106f4a0323e4463a5300cb9b1f3352dfd5eaa09045dc97ff1d3c72124f5e865207f880e6a6a1bd787d9f57c22d6ae76a8a4cde1498ebe403293129354bde8d2cee0e047b8a24db0cdeb377892bf3a401868c00fcaaa3b6879a2271b38e57e3a08a98968d6ff3d544d20f74e0ce6ac3349887fba15be749a676e21e71fed3f148c1d3ade24af6bd407b2575f07744d9748b20030ed87008857da44b388687b119893356bec4f1773624f27b9a029d2161b90fe52992e91934c64e5a2346b6953a10319fcfff6fcd9176272df1f675b097bd921749446c3adcc0c35e8a45a7b4d35ca96a22eb29bb0af9a40a9ed412a8fbd2b560e868d88b887c8ac1ce656656bfdc32573750c59fec396454cfd35940714b19755d3af1b18bc5a31175c11894386bd7393fbc6db00630b0d572878b96a7b89cac6a9b967d5e801fd3983969b4e3c397d3733f8ba934ffc38ee13a26e1b68c7382adca1c51c520fa7c809d73e399fcc7c559500485f14f678af3d532d469d879a3979b7133d52e3dbe623e10adbef010c537f26110db04528d3c2645a3233f10f60df24aaee5431af7a0ad4cba6760967a14f2698d4e1a8334a57b336d2680266e70571c0d1dda75ee8e9037579a2d4796738968e2d1c40e7946b988acb187d57752d843156c49d1e9867064b305561c85fde68e00edde225accd7a0283123c9d7fd0f3b45c6b229db5df4cb2d573dcaf07b4649139bd8acffdd8c975791a7c6664926461f698d3ab1085fec9b8680565f2510e556528a8c4c2c8abb0ff79866dc1fef170cc2fc43df479b227913cd207748c6514df97fbd65a1e94ee239fb64188a20a1cca658eaede4beaa55e0a5a7a16ebaba43532e7c1fd80bc3c5adf57e432dc826e6ba2e70f59a0d3b25324b475bc95f3af4595739444113ccf52d1ab6abf4d30c2da97d9613ac1c7429b092777b66fc22581a19f8f385c4efe4a4e53480e17259d5b0ca24a55d93e596bde35738c71ea33c58e16d3027b37bb014b12d426ba556ce3362c48c208c84c16fcbb99453123359ace68e6bee8d35448bfcea008161ca9c7f37ec2f181f5b5fa06480618fc5a5a7b8c74184fc9af16ccec0efea557be84bdda864efcfa00cb85c1a5a45728dd417b94f6ac0ab0ed30266bd84aec4b95cd37a2b6e15f9dc7f34b3793a965e7bea4e29331cf03683cb50a0b0a14dbe076c7835142e7a09bcd1120af1ae709457505816e8dadc496a29b83d76b9611a6f3505a41e1101b7fc526aa03924ecb1a263ad53778b35b4ca10636ebaf25e3f230cd619abb33f501c4804ef10f517482616bc3b01cb84b5ee0407b8b9095b8a2a3c477a816ab6a9a9b5b4b942691d85e3d3b3936aa18ccd071ca778622fe7429d5cd2546822ae000690d606da091ef9dd2f9844a9ace9f1c3b5f904eed6a22d3e6703880a900c9f942f5a9908863f9d73c78c031045205f818ca095adeb0aae5416d9d892370fddb3d864dec24d7f360fcef9c31733debb008ce3da8b800b0c7711cc9aa7804170cbb171b4b569081e26e874aca834a21015a5e402ff4a7bdc1f367c9081e9f0f24e93ad6e417f1649cae0375b6d91fea9de76cbda009f04043310d8b3dd507d346ae823f763dbad47b70f8f16390d497b03fa1019a2b68f0cf3b495724269af5ada226fe2d82c7cb7e5b2c5d726821121746f4decadda8e9aa0b1722dc30408986e9ea80b6fa1339483cf24cf3fe9c340a9c252d9c0e7d242e135b35f2e5048508d38f9ea2c040b5f4a8518e4ad145dbf2dc65dad0fca66f22caedcd130e1ba19d548c7778ace8dd80603698eef8930568cc6c9bff2e816b7267fd2e1bd2d6278bd8253f79906c530c7d04ad0fe50c3128a282fccef09295e2bd8ddc0887163a9b0748fbf4d112e175b7f8d674edb2a8c96fe9306477bb246c92680791bac3089456cc1a18a2696eab27ac84ff8e0744c54e4b7dc9df818d029aa92a0a7f2579a2116f3701a2adc4174d37ded703d5bdb108832f0c3cc03acfb770646e88c75fdf88c6bec874ca5c0b75238cd6021f04572926d71a0c64eefc5d9e050db328a23552c23f8ccd2e48f6cbae2696e76fae43ae77a87ce85b34e8771ce2a1f8c4cb3eb2cdf2078af428d0892644dfe298b589750948d6402a81f7ce8f8a958df7a8c59cc6b14529efbd6a7b6f16d9fe4a468dae1dbeca09dcccb8792ddf3fa6d550691699b6b0354ffbd6dacb75db7aedd0237f34a3a093976e8a5329e8fb2e6c63c64689379902807bccc5182db04b4f7dc47618480dd35acd7e18afb8ce898eb75c3135386a0192ad31167fbdd4d4129e4591c603799801ee209ed43f20866bb13f235ed2c7ff7fdb75609e31abca3db84b561d28014f3d9468ae9bb5682a5b0eb5078236266c449b049b83ee0c2f43ba5fd3dafbbbe77c28b2d797014839d70f1eb837fbb55497ee3e11d20abcd43ec4a4b63ed738f66be45c444fdc39fcdc475ffa8bcfe22a5439aba70b69cbe0966d46fe18883d0ee652cec5ce5a17132d30c8e4085501cbbd379aa4c6ae02dfeee338aa45c1eedb2ec84966217928270745695900ce39a1ba5bce5d774c1be9c4dd997708a69990741886913a884ebfc4846241fb4fbdc98a2f559f8995bd280a4ed7eacffb147c876f6af9df5517ec358cc875eb9dcbdf8a1080e8efe425651eea6da5759acb9e28f620df8340df85ec473ad2edc7f086cbfe986f90d01681b0c47aed813cb0592a407ca95cc3cf57d699925e7836de7b7a18cb53dd3b38e5121e190394aa0a22782aff0f3bea788aaed1df68713f0a63958f81eead83d50adcb5fee44cf83000e89cb0dd6abf2a8805d8d411f7acbf83bb377e18195d9a8258b00d2ad9845bcf26ee06429a55fb5c8c073f0db51158db856296be77f9218c020acd22fd59ebfd5986cc73958ce5ea1e9bed4494a9e8890da77fe183a6e34df6b848d15834fcd5a51d1e1df17f62906c1b243e659fdafa98a009ad3061131eb73015bae5efdfedaf3cc677961c24fbf3ff1fdcbfef375f683d93487e9b68b6901a5ffdcfb92c1b153772dfae5c9788b8e9942d55cdf96b4a72884e02a5212865178335e6c811b227b028c7b6f1364fbfaf44c6fd0541957c39443014501c254a816222fb66fbbaf6cda4488fc372724caee01c3c2690c1f7f43aeea0072f7b34c7f349fa9838230a60370c36b5cb82c3bb32a75628b22262c7e6207e83191bbba30de321d6eb4ffab22f55182fb0db22045b10cce5d9781999f81406bb5bcf6404c7b1f5dccee723420ec007c7bc502044018007a02ba7fb14c13e3e0f55fa9d00c0a11439ec2e3fd0ab08dbbb1a0cda080176291d382b8639368ca2ee8e2638bf4c5fa842b8e082249356bf808eeb18f21f9af7c11a5b491cc020ebdda4e58a8dec099abe570384d8c52c86aa5e7b731bdd16b4323a9905e23fa9e00f610ed10de76121c25e2ee34e85adcf9f3d9704e247fee4cb39b528d5823118ad0ec8485b984dfd318ef6d0d1d6d8000edced03d4cbb1ba934a913efe94bef68dd92d474c23a0c32a8b5fb3e8fcec36349851bfae099e1c513941f3f39cf3e585dd0fb389bdafba214652d2704fac776846d1db827246d7b9e982413a65d8aec12c2708c55c2a09460462a500e157f4d2ee855954539e08cd035690b0bac84f2fbb47580329d684241da122a69b427f37fd28d91c222d01a6360205574f1f0e2826c32c5d6361c7e479d123522b3ba5831ded0d91e247aaf065f4ee811555f9b9a76791f3824699055688f6ba531aec120b6f9058a62f3fcc8c209dc06510eaa1e7bf625fb97a5c0365fd7ed6a3033f38c70311dd4dacc0503928c477e23edc9f7313b425b67b283eed3467cdfcd2abb29f510f4fcf86f7e856dc43b8b85e0077eca39bd6c6ed65657390e1c6e878ab0b74aa72a7c3b2a699f43b8ac2de17b57de2a2a359cd8a17dfa54d943866f74edb767728cf736be72ede60c61f90be73eed610db1a6a7a176ea103ad227f62a815ef092d97fbae70fcfae468b57c1224cdc73958bc315b39b1f4b20b7351097d7fd75ff8e7c9f368989a6126506e16437c09010eb091219e70ed5df5f6400ac899204ebdb6ade5bd97212b0f317c3ad3bbc27b9c4653210be06dcefcd05f9c5680765415d2f0fb104cd822c36af2805bfd055947524df782b73c9854c4904785f514c5e00f4fb7f4bf2344aa0d883a6fad7a908953ba3a321b45ca826bcfab290ade64066f972005f28ce32f80e0ae0f951ad58bd9be8c4c7f89bc112067a9b081ea6b7d9d3d427c0d770df3464b6754bfcfcffac50853308283514cd195eb7fd982942df03f5e52d13e9143a6806432bcb34e953487a3d21f0a030384e4e5298f1e3b3cce9b8e90c99389edffdf0d132b443936f37672e4fed23fc3f70534cd9d74618ba4d8c3912a54a54dd4ca1e6da7a524aa8061dae3a8677b1d1e5c4e8b1efe5b8c5e79228ecffccae55794c8bd6778d67b459f57d9ad87b6753e6f6e3e98b260ff0e9b05cf7ac8e3bfa6cec08bc2f3073760ce31282041375f7a9e6718e8b3c6f4ef4a78f80739fb7b587f4756bad945a61b3aa8b1faaae78e71573d4fd3d9a37af25959962a20d370f2b59990fecd4bb8079d55c065f4a3d78ca78bcd49117bdfb7c62c32689ae80c805cb071abcbf598c5013e0bd1bc7a0ccc2c565b6cc24a9396faa5a3dee2467a2a0a996623553856340f5a5c957a6591c34a6ca568bcfe28219fd15485eff8ea770c6b7f909b5e33fb2f9d1ba94fe7b93e19eba6332baf2ff59434ee04619868a3f4f907f570f91d89c3f8ab5f75784ce2552b55d8b146b0e09aac69336387eabcc41f4f4667a3f038e9c3f365518605e46c9a391cfa0d85c3e78c74c2f002c09f03cccbfaae84cc0b39e67a8159f2da12d708256c7a8462b2a72f9123201de0c5407797132171362c1086b867df5828f9a7852db1423ef434ed30b06605a12dc922257941baebacaee5da179c81aad97d39db2e43ebf22124d3ddbb45b5ded566eb92cbd86118755fa8ed6ade25077f453b7adaaec5b26bfbbb855d4a7400629aa604dc12450fb8889ee212e95f54900257df7151b1ce4f0ae65354d974a3953cc46c18bbf2a0bd93d89f0014faf4d2090b7124aed83e1fe6d410ad900cb83a14dbd3e3212915341aa20a0a14c99bd34d5dc8aa363813f07fc83d14598eff1379f9ebd89a85f99a1ea74a6ddc315af2b805a081f7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h9581c97be81e51c73c2b9754f6506822bc522a9016f2cfe1a1d70e5607d87b9d42536769f376e5a65b1a2820134806dcfb9a03cf7203705b75b5f144e11d4531315f964ca352ceabccb2e99ef679e28ce05172f22174716f10fe9784b093889adaec0d010b8b322976ead81dcbc298c7137879a4a29b24d7f9d4319f17858b2fad53b4db39eb1f9fcb2108def25dd7582b61c2ef7c56a91d7f61b519a5733cf4913431c96777db3edbc81607c040efd7fd42d3b1335a6749e2d69ee0170b936bd527213f6c8745cb3377ffbc7832d4ceaeee70a43541dd7b4495c9fe2dd9a2f750cadda0b08f9d3b7731e1c814154e4692380ee357f296fb0e2c208d4f1b150baed9b6c333ac13c0a4b586f00258cd3caef95e37db5d58f9a7eb867e0257d65b4f856374553813ceedf3081cadc425120ef4c3e92adf68cc1f6f717d1f8d02da6e32454fe6998da5c83670a04663ec761a7635e9fd32545ad59749d651712f5189e5882740781e84134edbadfcdeda78cb2eddde2dca9938b92dc810c5f4c02039b388b2dcc2fc1734568db09142c10fe01fecb8049f4eddf3f1b0f80dd71c8393b9022976d82ee6b32c819019b3dc604e5509825fe0532347c83ed0f68d491e08363282130d7bcbea9eb89c96b0a810808820af3d0dc37dd444072b9f750120a4daa9817b70da0239bdca9354bbe835ed20311e6c731df5bc4c7ef841efc058cc6d1dd2fb4a3cb9b95327b25692d0eef690a80ebb36586f9394decd14095f09ff07b32703119612c05bedc465f10c6a514e7e207de860e0abad35efdf6bd19ca37f8536dacd85057e2a466cecba1143e1c51c5bb382c6fe736fb7f6dbacf4105bfcddf6c8e1c71dca7cf865ba64699d6c1a0fcb518f9d3390a49b0a6c5cad30ed7918f92b0de699ca67988d0bb536f09e4997268983de5ae21d978d2bb3cf6519b01821c01dfd19f4bc3d3e488d7f9f2b15f67a3df60a72cc05b48cd63bb7e5f4bca685cfadd521d3817227a1148a856712dd29b0a689c0248c6612dec8d2945e41bf57747421106ba5e2104fbdb209fc709571c7eff35f4fd09d6c01e30e4abf8f8b1773371c11c841a6339ef1a10a538ede8672df78fc7b801daa49ee3ec0af3d896b8a960e6fa612e58f11877cf3d9b8a6d146f2851612998e00dc436d392a0be3721ac3e97e2c5c2fb3fa1cc930b6d5b580bb26477dc58cee38fee4604cd147e4368ad9a308b6c3935d1a31ce9e4de8689c3cc796a1322bf5da8deceac2692b2009d6287ec718a26db59f76f847550222ba3bc6b2ecbf3c1c6c7ab86650e674b6b21d431bc8541e87173d0a0a44446dc220ee035b193ae8f8116bf7b2c04be1001dd5ff7f5a3b9d7e1e5c0009e0491c850d96f8e89c56633ab44aeaec68b6c1ce814c43007cb48bcb91803c66b5e7008879e22d3d1950069f45c9c145a87b98bebd719208d608770ecb8675808e9e1a2c2958022d40a4b80ed8e18d4df3980e2055eabfeab013bfbb0bf8190c3ecf842c5c5870ae0b84144c9bc98526fb4fe54961c799f6dfa080b0fb4c6f51f1749c0387460aa158109b363d0ac9ee0e49036c5e0bc825678943eb8f15a370773a08b3907bf8b36f36d4fd31b1f743aae200b6292e10213a548ca3688aabd0a8f1d2e49bd86b28ae519eb05a7beaea7b7fd1ea8508e9c207c35da533f359070e5c016c98ba5be0879dbb316f724c787fd3568e4bdee9d28f0002c81f189811134c4322ae70fede5b049b1627d585629be72069ff99d33496ba92f83e141c454091645d923cb048b8a7fc52e8fcad60d701dd533738b5457e98ef181d72d6b51e0cca936e2a5020a25d178341f4f54a8662519337ed261aaf4c2053f54e48e686607882e686be470b126c04d8b4e1a8ea64584e06807e371dfb5cf0907a656898213b1198cc4683994096ae572d71f99ee5375a6bd62f996d3497371de8595b610dc96c209fcf05d66cc8d7239c6e4cf226cf0f6c1609330ce520fa0be92cf3c00fce9026df3346b8bd34727d63a45c8eafda7d703e75ebfc0f864b1a6722d28e001b56d716b431366016380c96a808aee0784ea48b8692e18cf3a001b40aae6ed441449f007c80f2c2fbb889d4abd66c10cdc0c2bb1e92777bb657a2d6b77c29eaccc69a4dafbbb793e3dfa68986b308282c5b4441a5b575ac36f29dfb2613e271ae90520b5c8f7d3ef563bb99191728e8b607653aa47036642e5079faa9ec5a155502524cbd0be69eaebd704e1f9401a0be9a6cf2c996b9172d46a1e1f1fd26313c39ccb3451bd7334eca5b73332c48947ad0716b6f6ecf8e928e48e8546243d4aabaf284eb51a861cbb661435268c64ea43e979177f094daa6c0ac862d34ddfab5010fa114c7d81d72ad354e8d97d8d8e97d03b378a17dd0874a054a26f5318770e99b97c0f8640cce6a52046320014684eb4b4a9c197a447fa6f2162c6367205ba3d87ebf68fb0a9621f7ce3d3d3a1c576de076515ca07669c761ddc3d42954b042156bfb824bcda6be734ee3972b3aac7e8f790e86d77fc699f6ead0ae4d70e745c771c1e693869aa354de6a706b6962b108e5d49378d1d3922f96c85cb2d721ba8cb14edada34067f7c612a639927600d592fda5b9559d59327a0be75a026443cff0139775d9a5fdce666626ab4420bf44d91fe87d2d370b602667f00ab8d6a8593cf18bc69ef78cc1b36341e141ce13f7781697f82e50f4404302d273f3c614cb1f53da6cd7f5c6b5932a56fe82f260721728b14ebdb2438baa7a274fe29e6868a48c5a54098bc4dffd16d23dc4c884dd6c496e633a240d867459ee20dddbce97388cd5c72b40bae956fc519f94a476fdab6e232d300b6dadfa4a967cc55fb1f7dc366f7755da79e03fc4e8a685fd34a127c651a7ae27237ac936ede394ca0dcc02b4fa706d28a9fc4748cdd20fed9ae0828ca9c5df040d35dc1eef00886541de44ca654ad34487b3e4b9a7f39f862ef2343f20775c97e48622fd886f6181d4634a6fce31e9702c64e1f6ee6ac75d53eddd376924b7583c4a1ff0f0ee62063cb63e6f9111f85b2a82e8aac7792888c2ccbd581a613404798701013783f58b07a990b205e6b985c2c747177c62bf2001326abb34f9a9f47ed23c6636f8ae22ab2735fa939c1e799261c7d986a4f911f3c6b40a4832dbe0002c90b26c335a9d72de32859495c05ff73fd98f4465a429952d8a39379b1c678fe52977e87e4a0b464ce0c1b3fdc10b387d93679d2fee3302dbfb2a1d2705c01a243ac347451ec4fc557855f41b508e94692e3432e85f8246529780165cc933bf06593063affe5726c01a549a28ba6c7675e8034e9e071fcba199a9829b112fd4cda69ae4706e8c8a781340d85ef483e726c5871e3401ab7e294e0f4df5b32effe8108bac190e65c6142defd67a396b73385736d8dc8545eaee6001b291020f2ffe2e1f26bba26f6fb224ab181132619841f5b2f69e55a2fe656b19d1deeb93b4e0f455424bd064d6fd68e250f73438640704919447a5b2e2f9a499a52fcd3e7d1fc91b5ee855b60e42d9bfe1ab55febbf0b7b69ba07de7b6b0fa8225fca8ad552df21e54b75cee43fdc2ce57608f3c8afe09c622fce0df05111912ee241cf5ca3b63c5ed77098641a0a0cc02bba9e742b8aa6aad3ad884969de9d922e26e0d4f3f07eef93dd4d58123f3889e09e06a81d91f9889b5fb5df60d3433af35478df8f752135930c72bc641b784e82974ed607320784cfbfa594f2f1aceec3d7b2a4980255e9559fa30fb3eb148f16df380253d55569515cc572b9ce0154b73032a75c3cfeea78e60ed1dee684c1e69df03b24b7026c08a15341ccdb3d2a4d52a00bdf805870ad778f4cd08e2d9b28048adb728e46c1ff5dd03cf39cb6acde55817d124f3826cc08221e263847a7769bb847f96f8ef47d25e933987db334a62b4fe77a15bcac2f6bc3bae9388887150303054bbb5cc345e6d85f056d39617ee86d6ad7b8c256c8aa587af16b758e99d2fd42fc6deb830ff05e346921b760cd29d275e9093693bd59892868503b0de5f61356222ac8a954d2340332c2dafdc2a88e96e82dc9d23479a0d4f0917331963ab5e0937b6269e7299aed15f2aaf0bc6149c65fd708d54c80cec1a50e077360a8300549e45e5023b8bce57a82c11be5202acd6d378bf38673ca3234beca111f20d10b85dad6b44f051db998799668383007a5ebf3f8368d6d11234d020ddfdc8911cb7b95ae842521de97dde7cd702345e11f499dbeaacc22738ec581f3fdf14709b5df9641ad3f2068672337aad5b029a4c0131290a01ac8537a1fb6265bdf81e32cbb0c771779e4ed00be120697029219f8e3e4bbbe8021f43308df415e5e4920e25e6e5c571a0227141bc789868e3ffd099ffdcc9a507d59457677d514480c1241d2d6d64191b54b140b2aefdecc880cb49a285b593442cd0509b38ebd508f9eefff630d91e21d60955c0431f01ce0d352cb27123182ef58d030a3d0241e3a7b5aa5f8d63c307ce25427330c3911b352f01c3c9155d5b0b60ebdb547dafe9dd579e4ddb3a615d6d5037bc982c06952100f23f5272ad53f72262a80b50881fa069b78efeed201d7c4518ecc737b629644f0e1bcf60431ae3739d218565a20491f19f2e5ff4e5cd4d43b452d3d6cfc7b2a4ae058936256acd2a1e034641392c9a6f3323ffa7841836436d9121018a2d33ec3f74514556814d8e538a540d2ccfafc6e8c3d8766bfadf167e064a039f4a5f869fc02d540c29ef6365eeed1cff7fa72c102e383653c851677d0f549ef488309c0619db3d204e80a7b953d0439da55ce0c5ffd6c2d2e671f0f7874162f54bf86448e4dd416bde654b9f428d2d7c015766a2759f4904bf5767e2311cf9b6d10d372edfd989986f4684a61c6f4c09d1a4a0f5bb9be46a2b49ac4d4d42b2140f44ad3797caa3977e2971bce6b6520d157531cd9fcd1450a8ba0aa560810dbba995edf64811f95be30f499435006c166cb24ba16f6f85680820a2d226e8e3222a93cd2e5d1c5b2d10a8723fd35c1880d79ca9fa34a37645f0ca810016cde106aad6ae7685e725f0dce7d6cad5c44d573ce2f8ad657eb8b9227c2a33b85651e449e011d799cd1d33d9f153815a0f8f6c4cd55ecbca7e19a10e6192d54f777417af0e72cab044525b9a8535bb3f14ba1264050dc23bd8e7b0995e40638a673a3a107cff7e133b646f83d201ede53562767bd80d2fca4dee279a2bbaa6cf9cb277e8751d80508659fb0f7a3a09a536d671948365918d9dd10ad7f0caf70022c85f67d4057421f89700bbb651b7ba90aa60b4b3b6b40cdb38db33bd99d289d245c840477d4da731c157b566d2e887634235fe0695bd9fc228993c9555e9b6a0c90c697587c9afcde36491f098b377281928ef03941476e362fb17991af6c6b2403db11c080c81bad7f283059627a963c53c873bd6aa46e6edf018cf933765685be84b17d61a376333aed9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hb139d2f14fe7a34d0bb8b4cfc1ecb312bffceb5fe752bdd446853f12dd6da91ec5ee7deebae245070b358ce69ef3160f3a5d6619fe723fd8ce6a75c3a37c044c629ad72051e39f9d4ac960a8692014c3d305ffdc1430c33d4047703f4a9a7967198ce7c368a5d27e5e3745a481d4f7b29605713374d574eb7b77f45a96ae64eba850605f12f44d250c0aa32f725e832fe1ceedb657711fdf0c3e6ffa847233049cd3403b4ac1ac019076a0262260ae1077b1b44eb249bd71c8fb25c76a770a3f46b8d677f83f4d52af01a9d71ecc222bf494443320e21153371b474c85b8411bcebb840efb32d8b6fb2dfe68bb48111a0b445840015037c2d09502c6e1d02ce78ce5724419f44f1de783073c8b79902b770747a38a686b8f2426b89dad457f9b6efd7b26a7ac4e77808475d9d044c6c1cc5b6225f99dc28212ac1d7c5b6db0b1873b7f76322d2f5fcf8cf37dc66adb49c5eae8f99395c608220ca3cefb0d1e9543e478026312efe39179ceb6617c160a6555f7775d5dd9301fe196ded64f4ac556823f484f02ff4d72e0ee852956b48a01cb3f124efae5c157d0774cb992e386765005d9edb56fe0634ab4a6fe88e19521efb590729322530a5658c1054b681702c8e109438d1cb3c2e1501dba0050187ab2c41a5271be6dbbcc6b85a341f10a2ce6644e42010a11ec4777626f559c1d521bdbddf258b01aca9a0f8ebf0bcb9c8650c28fa09e523e48cc4fac8c3d27e86fd16654edb14c4a555ff4bd8cbd73c1df015e07f2fe322b38fbb588edbf660f1d9a2b7b44b0c1042d0b614b81157603a00d7ca06998b3dfaf935e14b7f67e8bc7e52b29b9385672e3cf47498fb2346d5a8623d5916e8b27111d10ea757d70a60446fd68fd6a890aa06ce2eca3389e26091d1b5d3226d1bf4f8f1ac8f2de5b5ff33618f10a98d9c67f1038efa8552c42f283466259c8810777e723a6eba304ba949232407b6a35d60aa9ad557939e404c30f7f42dd88607cb0d37df407a18e923700e0b9bc75b5029590fb3b253c24a5f5d489ffbb8daac6bd50841ec61aa5ea3b2b8fd8cf676bdc89b04aef6d67e2f4a1fd63c2ac5e30b4b80ed9bb5aaef12ce1b9dd0e8bc2b69f9db6d18e1be93b386a9fa8caacc28329d95e603805d0f5ecf8d7348878388d9cb7bdeb6afb6078733b76e50e5cf8b8b6d6968923981a02fc973ae27be9bdca27d8ff9134cee831be773073ba558a9d3ee9a61748c230159b2e9f36aae9065f59aacc053c21dab81d55620e7938e5190ca9d35691d0262a6990e3f76e4432751b04465ad2260eb8bfbf323be82d0e44a754f3a0df1e89dc7c32e866e562529ec7057b9d18842c49ad7077bfe249a7aff42dff1b4e4c28e132b612d678344bf2fe0562674ed737d88dc9a6adee227c5b78060ca987853f22532588b32b267f67a8777677b48a50038d92b764139ddc5f463614a3a4879ce1f60c0a8768271e101790f223a8e74f3b2911dd0229d3a81bbea9e3161e64801aae5a4f586bbeb2ef265d9780e25345d256c356b3c7ed708cc722080150418778ac669062adb771a54de72e9f8f99c8377120660601819846d469b92772d1754a9d3192b12f58356e4938ba6189c7718aabd430d9d4bd493d8c79e51653ed03548211bc2a94f4ed2eaf5cf536b3f89faea3aed0ee92697287bfa5283e59a984fef6422c15240c0addbc9d0e1e8652e43cde1504a55c5e0d434784703bb0ce85eeebf54ebf04f94a0569822ef3e54d07ccb442ce4ab24cf169d180350bb4e147d88d07327c135b908adfd6811980e3c977daeb9d0c183a8c73ccc400e714e7ed49f9996ad6c0f0ab2ad46106ee1ce43a13ae7c4d7eef5ab6df2b35af1a1b891ec47e18427560c31dc9dc5f4361f9d45c90a47fcb8f05fe47b4aae98acd06fda2d03a447186c74e375a5b4a80018ebb69010d282f346bb14b8afe196f6a831d4d94d04071818fed035d99a55cca3983cb6d6a25dd4d90d0f0382c5210f5aae85fb3a2fb9a7c484c4385556c4b550d8afc0ff7ed0fe341c9c2aa22b9a32ecd2eb8e0ef2630c000edbf92184c3edb957253a2f030eb08fde5635ca677612c5a81ac5a66a95fe0a14a8ab2d4da667986945f38aa094d818504a39f3a36739b37f875e0f6ac6d1b346e0288ff3e65e158a172c25c67faf081a1b0372d5b318cd22510e729104ce863c5b6bb8bed0933a640f269cf48ad5234ae45260e1b519d5f48b9685ca6ac2b7365a7e15ed7ace1c56eb466e21cb61548f86dc120b1f3fdb7289a2376cca6ed964209e6362f446dea03810a227a3360d6cf62cb1a6b4b11e19ede5264dfd73449c212b0fa63fe418e62d841b1fb861f1401f6f52d794bc55aa6847472f9efdc07d59f074da23a73d46033134a9a5bbc53139d593c3287d32921916f2d980d07504fd987a5c6ee765f835ab4372eab863d7df8587593ca098d981ac9228b71af212d0fa597cfad14c6e8181b475adef62a9b1d5302671444f4624682d910239ef138989567b75865c3006349b8d46c3f7a06d199559bff3c8c6daeb62c18174dd7f6beaf74a5fe2cb30a8ca3da05bee86178797def3c8d4ea22381b8df1a3a78761d9d11eabd8a76b93d1178bbf41188aee85eee138c690f16a3630ae459bdaced0ef313fd59fe18ac3269645d35e62fed1411f36f372ccaca208471996d9c824c41d3d7ea86e1a1774825179101410080f9d0c42c433d17d9bc3ab336c22308db43abc946eaca474e387f09445d5c061aa80964fdf92ebdf033967517eb1a048088e81db751ada7df6d0fed1de4d8327a8cad40c3317d7c8b959e48df031f66b5c78c50310c523bd65f547ab6c6986300c5e2e4df3eeb98c2f53efc6a260b0650dd1c58c211a0dbb0634daecb8af9a6061f02e63ea801fa5f55cc2e1feb0a65169f2a18cc7475d3cee669b15e57154f548b91fc75519de4d80fd114464ba1a11601a0e8d08074f8b18041701fbf3357aca8e13c00937102af2d49b4d863cd55a1f14b8a09cbd312c8d49d886487b39b880d113ed46ee18258c53f2d75bda05e603cd6db0fc4969a6f222070dcaa4ed0058f091d28d60e063a2637f44cfd1ec9da5e44588f61258476d754c03975e9182c737d2e31ba36d11d152bb9c7013c5c016dd03b4db6cc65466b2d5be4b19200ab9a3b126a8cd032e6e30365f881c8ad08b03cb270a83723433df91eb68ad287f81df371089abe309f4b600d73932e2a1219d884428c59decfb40046efc2d1004a5784a427f94dc8156cb252a412a4154942ef6c9618276eb78ae8a44af449538aaead049f9da12c5920d0da7528a867f4b965cf46b1f4918803fec6adee4ee4f92622003bda2e50d9e10b189e119228dbd1186498333f0f3cd88cf3b36533d283641a092cbc4dbe9cd7f3dc665ee03776ef6e5daf33db86d85e28c5d13bdbfd07da6e51a9e31811b965cb80b8bf7a0ad4a20faebb5d5f8329a445db5acfc3c8edbbee75d3040df42f7ea7c14af97656f67e853d4a6d4382966681831e79dd58a0ae07bd6cf6ec45fc6b9c695e083661d717e4145750a982f4cae2b43dd244d7d0db353d2eb31265bcd5ee1d2bb2523370d65c610cc9c78a26200ec97f14f91f1f3803e7ec5c78df24426be6336a3e1be3fd3d72ce9f4a82caf2fc22d4a464d7a4451d10689a8894ed26b7aa69e2e40af817b2f19325265598f6977390fc1c35f0cc85395aff452789552e6326ed6799f099bc80ac5d4831aef1e597687d165545794ca6310340e94f834c5f9955ee419943d251230bfe409e0dec2e403c4e4f3a77a28ae4113eb86538084f285e29a97f48891141a5da7aa43dcdfd32e9803d83db6447045e3a5c50f4ee7f651d9ffb7a9d10d6bf81b2209fd23672729b9d914384f4332c7820a0ed70736bd084e78adef11e97a93506d3729c8945bf20151c70385f5a9bde0530ab244eabbbac6a6aea7f7375e9441daa8b76d88b410c25438e7f8aaa3ab8d307dc179c7b0b5d2ced80220c68517309030f8195932ba6baa7cc0f83ded4a2edfe422af0213a1b4a0c702b731bcfa6fd393b3237304a7b56b57aac86c2b4d5a2266c30018412d94e794693f34880ea9e7e11c41edefc4e4625ea3c744ec3ed5e12f9743a75be3ed55334180a2c4ea6f0d7ed705c68443e67338ffa4e9ff40666687458031d4360de438759866847e36b50de9e332e642b147d53cbe6cdadf4c335ee00c425a4c522290c244f3070f932442dbc6050c58daa6104e9a6144f00070ee215a12fab8bfe3fa4c84679e01da26c7fab86cefe0d22f6ea9cff20ae91fe961904b8bfcf72cabdfe1da10895803b4c952d28fc16c7875fed90750d900d4fb113c7ecd6211a32784b82f54bed717a5798e3fe9753a491c482b829f3ae1e6d396abc5799f4e81d4c4ad4ef2cd61493cddb0c0a7d7e7df63f701faf49713c21ba82fee5acb5f4129368eb3dbc3536e68d93b6349cedc2b65165267e8edd5123b8b03d45131435a3f5a913d8657e3d833a717a8e8201808d12e06591270d32cc7ca361b9ec99ca8e58bb3fab384239f1795cb4897611423d06bddaa450c1abb64a45c62710229e5547e7230b60e5a6b84d651cf841633f2ac4e693653d7c6bd13a4e84c4bc6ec58fe5a51b7b68aedf04dac720fee164c38168f50ae4ddd238b673c64c4377a8d0e289327062f617bfd34bce4ba90b174645c7e94f60657c295b3d6a1e213a60f5e12e40569b7a3a297c05351520b42738920aef1c090bc24d51a8c2e9b799241edb43d64641154cf7d012d7e6bf37e27c32c54394a1c3549f5bdb9d62d734f86126f8e96a0c5866265cb2fe593aa66b7844642937a32134af97ae6ec2e6ab78b72a33b9f8ef8fac563755ca03eb407c4309e66ee0ff2bcc10579642d279a9693a53cc645b2bcfb1a7d6bcf6991832aad33a0a456d845e55a2c81f07e00875b34f8aadad4b9d83857e87bbac8f4d185e935ba5015431900548e263f12d2bbc28f84836a9bf385618dfe4976839ae5933c0816396e0885475fe6565ed39a3dda573702ac2d3df37a81730d9f8c21c24c0e1a49129c338e04fc7c3797c4ed255601d1100abfacdd9e7267a9d7bec391c746856a8547e61c038acc77180eddb9d42f7e13c002be9cf487adce0667dfd00170a8c9236720139cb56baa59f23b69c01ab875a79753378f3b34d34371bb450d6001ec5bcd4abe1fd9c9de742f9ce3533a6eedd1440c155580ac96d08e8eb75860492a089c6811b4eb12cc7b47c7512a7973dfcf0fe5518e8235815fce7380e3947d5042c4f71ef5b8db02640c9ae327d65a39ea0620ef717f2ddb7861cfcc8d1c077d578a770725ae32959b0112a7ca670d89366a671937b884db873080949e0e54dda4265e1ddf99bcdb3ea3097d0099aac3e91202cc410cdadbaa9b64bfd8d389ac3a4f8c27706ac13ffbd1ad7999341a153dd266bfa3ddb5c261942977ba10f7ba234e0570d4c09e5e75ff78fb19a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hf8f1b8ddd06a5fe4ee49f8f9751d23ffee6dc78a603686b7ad9d90866a233b9408b871df1f0c167f1967669f5ae9c842b14d7c1d2ee40e9ef55df8f189aa153b15aa76dddd713f06d512ceabe5d44b2df3336c5f8c968169a70b94a608855a7ed7882810c7d80ab18956ea44138cbfe23ff14cee23edb3c99c7993da5654c8d40d7150e5178d8e32816fa65b2d2816c9efd271901e33106849536f49fb6889c74c2b4f188aa8328efd9ff9847e8c7b69271bb034e0eb98b288acec6ea08c9d51d3cd2ebcecfde833e594313e0c2d39bb99dc621b60ce2d3f7bcb7fc887e4ee20f3d0f8f86bb7a6f2d74040cc602fa62c4a22a70434f85ae597c849e9407c81dbe8307566c3a17ff6220082cad583034ee360b85da6a107ae0dda6f614d141df25d605a0d90d0ed1dbf061abea3d33eeb0ebc0c51bbf0e2b104891756f9948bba6486e64e1c56f4a379d287e00ec6fc53ee97dc4457279725de1a399498bd37e700dc068419dfce53618ac16ef437de7171983d13e5ea4ca0f435b1f4866bb1fe752db7c2ab41d7c95d1834393ec74f525dc106af3f48e66f8f1e864d275352e74391ebecde598dbf7d1b6f777148463c66756145c2a3f4b9f508d415a2ab9f9d366a78dc5562c8b1f772ca51ac887a22019f7d38345f6a522cfbfe9d92657309886cfee7f554d217122cc0c87d6975d4a2fa77462b16054d1bab699424a7cf446a7bcf327a16e395bb1b11f3895454bdfb1f71b33b3d828755b676cd6c8ebde3f52640125a9886271cd84565eca37997be90c1978e44b02ea2b2d20a487505989b30564980ca83f8b0b48b576d638f22feca9879de2d0dacd9e4d2b2581ee45ea75f9d0675615a6bf2a9c95786c77e0988eef387ca0b114393156432d53da5b0eaa627fd279cf4ff243f8ecaeeeea3aac6819e35ab2326f3b297cfd3089133970a8ef11ede300ec3aa5ee60951df0bb31ef66ee7dc5b31d000dd3f223a5224a3f04a2a8167badd7f45fc5e7ef974eb48445fef4fc4b45e94ac628a5f10d035c9e6280bc5a0d116619176564c659b9e597764ba117ad952add5507a6347d18a69c8972f3af93f8dee1889d6dee008bfec25c3b0886bf242aaeaae7ebbe57d65984d28643b3de7c0d1ba5688fb07b91daf7af28ff961f91cb02c59807c266173198325a70e8c45f69f2487d0a25ac94be5acb3776f31b923506a3c51b1f764c42a3399fc79b220691426d725a2583443b9b8ac19b96245fe10810ce102aa59d1fa4ee61ca7d032a5a1e182d4b8d0c631d838abd32f6dc99b4549938b3fcf9dd697b6b2d43032b7b6cb1a9072601b7299d116f6b6aa6a9f7dfd2eab0f08f43b1489ad9d3e7a4e3b1cad1e036ea52fd98df6660ab2a472e3c8bb2712b3a161f518c51984d25941b8ca033bc8626b22dc3323aa208ea497ebea404b2ab853548d3caa49b95ff21fc6b9aee003e6c7289933f90cc481c73ff5a8fa83614e925ac4715772490ffbe882db5f2d973d4596d2b5f27225fd8e2b1bed344a0220b1d25162012e9c4dc41db25fde86690c362d6568fa931eb1733d60ac09b1bcf5ff0fb86d8fb88d23606050f4ec6cc9ca28fd73fd61bc46b1e463884ebbf6d4d299bddab5862baf4b99a651aa76f27586279fbb10e6ebc766495c42b6324c3f91a4a814075ad24aa224befa4bd44d5fd9a6bef7b5ec2d2ed93bc6634075e0f593e7fb5eba13972e588abd7fdd133538da9cde396700924927a979b1760816ee18af1c4d10d2324df70cdf150a536551f37da124dcbbe459d797d5da6bb31ead747d1eac8c32b0fc74b19d8488798b846d56aafa67192cd042da6f9c0ff13c4204be03ebf2b00870d101dbf4e70e7fe2a2f3d280dcd0ccc09a5e0ed6acc05f8d8d8a7e462c6de1620b0c407001144f6f49a25295689d1b13093bde7e7916379dad9824a7b3aaeea7a0c6a16179db619298f40d9b8ba878cad2616f98a2ecec933d1f617082166d2e5a60741df5ddeb764592abd6cc8dbd2a282b978b65af522f3444e0cdc2b427823deccb008a63185af16acc78647d719a10d5723a885b5abbaebc70b7019e71d741ce585c45d2d02875750567dbb3172ce6250646f52fa3a63e7d105dbeded599090994c74da65cb7f3b1199c417f4591d842191eccb18c9ff715401e1862e9c584a1774837e5af97805488f7b27bf859e1669f512b5f5ffb02361107f8fe043bf5b8a92b292f8b75362fafb575ce489cd81c34c682012bcef8dd05f61e4e60fb1466daf7307a1c3261ea7ff1615b1c9e084573828e0e81c53db56a24de9ff376df7d007c2ce19df991af468b253245eae388f5a685375e3a4866b5f47440c7ad8dc9d6d3ddb43254496be559f38fafb5223b8524e89ca2861ab8ef4477d85cc093faa95db41ad6728bec2ca628574adc8c45aac27285ba51393c9429806bc4f3eb7ba450cae6030fa1e47a5336d8590e1395343968c0d972f0dd1de8ce2aa557ce1a087a1db38e85aced3ac96a0b1469ca424a046f929abe80009c9f46cc4a83187a81e643af03f9b825c313182da5b20f746a3dbf667fc23de44a94dc09b8202d9d5f755e7f2306bf155d5962437fdc96639af9e2f40dabe95412ff745f5b8ecb026c4533d9fb0c03700e31e6ba0fe77495d6067799a44df9d350c450e47bb560734efae1d99ba565da0dfaab959a053650db2c1801b8778a56d810db6f767ead6d55b564799350e1f8e57a68d38d999459ef055ca4222b9c6a4553bb0b51dd6ad3c25386d27ac6b06114172f20f1f5700298543022217af9382f4463fa5ab2a1084bfb399100b48291cf0581d4564444a0445356a14c750e220a7ecf8c5ca0e4d66af3957dbb8247fcc70ee74afeb5db35173e2403665b9ae6724a0cfdd0678094f87ad1e665ed5551c648ce2bf3a3ea67e388af7cfec32b679e4c81bb9a0b8f7260ed9766da03c539ad155faa07190e58fe5d75f0542ce721bf485df54f02885c86d24f6473b112c28960604b5588da0a1a4ac4dc88bfc20104004b19c629d9ed56c32fb38bca7db72c6c40e08dcb44552ba9e896953be71b6fbc83b530536fdcdd892702a6e2c9425ab8ba7e8df491c664038400bd077e90adf18f12b05d36fad2d8d60ad9b8c1df3670cdbcdabe5c3aae7cad35b83fe2c602f6f1f601611641df871e424ecd6142d6bdf8c27101f9950271e547433ebdb3a240479237d9394b20977d01c79cf4e7efaf21b7f925a179713ca27783fe38c2e3b31578d96e3d3411cf710c388a9912a97c78947ffd6493aab813797a58bba7d959a927a3d0533ad7888102b9ab2b2c54e60402d6e65b787779c553cf7741035a06d6330b8ea9c2f1b866a55e685c43da1b5b013b9760433591eb23acea0c2119edc0a0d614dec149dec4ee464fb6f09700ae342f613c7fd6a7a3f5b7cdb257ad1de7819498b9fc8fd0f0e17649966c1638f87fe4ba80227616584e39da0150d325c325857f713590540ffdd09dfd56d513ff0502ca977e64d284a27b9ff396f5c450724bce67160d0cddfbf6bb11e935c7bda0a8d9a5691786056e326e7faa615a5abd1afc0bfa270ffde87f8bf15690009e133c5b767174aaea3392b18bd6cee68845df8b091a0a7dd654c7e67b11f242374798b7d9d6069e4634120bcc1d658e372e266bdc4c19a022bfedf7e3dfff56f1622b934db8274764f4021be6184655c44a5ab7c471b6218f146799d46723fdb2e8702c1c907d1226126873a1e790008f3a85b96028e30f88737ec6c9c6a59477399a558043151c383bb795c6d88b3c3917149e30d638d75221f203da414cc3adb84c28a894fb868476c68c4f25d475ebede78c96b609d7e66dd5df7f7249d8340fa1362c1f4c6cd67b623c34f25bd3e7a28729c795f2a802fb2f7a00c75d64f5fe16b7c4cd822baae20236a9127a6bb0920120ef7b16dc1e93341e549ec4db1d42e5d153ed572286abd5431b59568b2b6009c3ea6afbe72d985b6321b5ff85ff20bd662e3ed589b1f861ceeda2b1e66a69d54f3a8bc8697488ae6ba0ce16a2dbe220af611178655b492109e4653385e83c1d951d0a1347e091ec3107049e0292b91a10d3c451db6616900bd0729b2e78bafd57b949f48fc3ab131907c83d26b9019c2708029fb86f43fa44cd9fc3073b2e8416f43a68396806e885235e0ace3699023cb1c8bbe6252bf25cf10595e8bf9f559cc2c48977725d0750e93f46f44b4b8b41ff041369ab1321363b1adecde308f47e5b6fefffde9d4e601cd62c03136702f853a4c40867963d5377be5a67197bc1533ab12e744782787aa157c32f574a5a638a90b66f9c5dc64705765eb6cb60238ca8ab3df468745b95f939cddf68e11b7042cd974f65ea10310b95c62b9f18af65a6722f239dcd7b48e0d5af9aa2c6b5598674036d76484a9d4d284a427926b2a600f87d2420c6415431f49842aa44c27aab97702c2cbfcb3cb9cca4ba8b01b9cedb887cc951fcbaee7c7c66e81c683cf9e390e3769979e814f22638b18d575fdbf3105567c5875e44b420688824be091d83f4d2a516db33bc4925cb6b07f64456c8c92e2f5494cb76b3603922e1b1ae5572e7c546af2c192a3a1ea69b44ab5250f0e8e061c0d898bb3e41201cf1f6109a468c589c188e680a8ffe9c316701de9fac817264583c7dab02abe4c271f97c8dabb0f56e74ea338f192ef9176ad2b18bd4d279d5afef7b65fb7598619f3ee34d59b071edc54e4928c43401e70ab40bd3d7fd6201d91afc4c21b79959103698c046950280351cd082804ebfab70175b522b2c7cae3cc8d0f002c6515579146391bda091a69f09828146fbf80f2e90c8e4a7ddf85ab69857f32f088066b765d47a18faac517a52ab7a32b61ae74def50062f1e5bf6f987e19b3674ce3b9f683a41422bdc25c61e556e994d31adc55fd6d07bdf845a7631a37a2ff2a9551849f2528a850ce3bd22845fd95d2ce5c1080d591285453fc08a789fff59ba653559c183a0261ccedcb96507b9ac5c802d393b7c37cca18398dc4f20f18897687c915be787461f0b0c6d500315d3791584a93c3e1f88406f3e3a36af0b8027a5f8b4f85eb44943bd0edf08fcf5c589195f53bcda5f770bdd31da7e2b3703f513baf102ef1592794ccffbee754ca8e3c26df4f9cb1e3a226911c16bb965439c37422d48c0d1159ca2cec494297a47b11331771ef620d48717b26891bf6c0be3d8c84b7f733abfc215b0917b91e1b12fba27cb48da487e841bf12df19a9eb4888092e516a3862fe44b87aeeca94931877321951f3c832cf9c79cc8d4c87bfd8b70946a14baf6b5493a67a3b1c97aa7ebf388c195663d1f638d8e0c3f0b263dc5c00963135862205a07d6241cdb14d30edc9ccd1fe71335919c72255a866652661b6b5e2e031158799cd0e0227d60171c074273f3ecef524bfcaca89a57c41d59bdcd86e23efce7d5cf44c5fa77a1096134cab99bf8eb8bd334e19d88597071b451ad9a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h5696f09d18cb7eaad85c0a40bc8c160a23a61d8840e4d5b383bab3e7d1e7cf4cf12255c4adbc42836ef45e9daef7ab42233ecfe6a25f56d013ca60f8c7e6dfa841ae2d1c0c123210ddce777a353cd059538c5b80f38cbaa079fbff6bddecf3b96f846c75479bd4c52b1569cf28e78554d218fc5da5597def422446c64f7797d418eda4435d3173f26b070ea40dcbc4303cd7a3b41ffcda35a16372bfca4755e0a5bb99df1d6064e80a309f18eb0d473f32f5207f2cafcb2cd1ab9cfb2accd6f6783cef91a738ca19ea21b02a9d2768672f8a070a607e709344955e2a0b2f1bfb8d976fd0b42392b1c2d1014c210ffac1b500a6f571a268d81c8a69ec73f550caf56aa2da87df59bfc23c00856db08c49c64d0b9409afef6e5a60d42fd0210f73755b9ebdf53e9a0e9232213418bbbd10eb270879cfafccead32489a9fca37b96ba30230d19efcb0143ad2c2c9b567f8dcdbc7d93c100e8d57deafdecbcc809a44895e4f5f160e56ac726bba25f04c3030c52acf190cf5a8f62b9f113cf1b7a9ef7dce5446d3cfd40baebc3d8bf6ed77094c2d58e2ddbb357be2f52f8503636319a139e990ad0d700c2841d257bc69d9da983d05ef910fd8bb23ce0b7518adbe8c53dd5e7603e1143ef6a6ae80a2c224104d4eefbff70fd2f2ef5199814b5adc57fd8c409ac6d6bf821226b27ffd7a0b0655352629d84499a3475a4bbe4fc156048fa4bc2581fea00e74950821b1cd6a196dbc5b5baf4b779034c062c5367073c208a049bf964cb9bee638ae67b571b3ff764f70c327150df35b97f6098f0a4a18413913b0ba432eee98cedaa6af29972c744f1e155cc4874eb499c7e164ad4a0f08b2ebcbba619764806e5ab66f8d1fc279d6d0f7ddb1ef8d72fde8bd5aca995d47c4768241a87821b4d4512ead56d820ef31917843c3356dfa6372f6598064be9d3557eaa9938d123b9b62877b3920c15b0b2bcafd45a31e97cb87c5545d6078c74c6f3facf6f9a4289515e9b404a3deac860258af00be8ac5d1eda1f5aaf5d877d71665591fa364dbfbcdaee9ac14bfb45b2a85112cd77a64f81587b8d5f9b9f792040c136bab3958a06f4c623407fe3d4f870e7accbd7dc5a50aa5d0e55b188d5f3654147e7d997afa4f721be7c78661d28d237dc6b37b7a9726479801af14bfa8f45f7aad39134ab502d241c48e552816c6a0f93f17cc35070b25c7f2ea1c61c5b0430008d90d8c60a79436e7c463c9994ba166a7c6f22089a84faa7176ed4bb10104d68e63f682c138b3decd587000281230dcd37db96ed2b6588f0f0de68ae8e5d698ec55391e20bad8bc7b70f7cc5ab15678ff89b582d4b9b436cb36164ab7d5e137cfe963ae054fafdd9d04dc26978af41f613a6ff631fe4f58a2e6400c0ef67a0495481afb95ba543ba26b5a88cf8001bbad4e4bf691cbf310d4933f43a9a98bee6cc3154563fa8a380cfbc781074ddb5391a0e7d6df3872c6793ccbe3da75b9abaeff2e023ecab1f618fae13cf1cf7eba630806a60e0e2b3fc8d7ba5b45db0e4096663b2d8d96c04a9ec9d2b1f50c4ccf89b3f01b3f7fe27abd50bdefdbc33e0c4923f2678d81ae6afd524232ed9d26e1572d18fdd3a5d5dcdbbf3adf38207c7e7adc2ae2b95eee2f2b75133a6f62ef6b07a389f711aa98049bc514cbf605b7df4f76d0ec56dd092050c260413dbae1f156c0cbada6dbe379c2d8b8411a3ac48720e41d086f1d9fffbbc75fd348afb4d64ac89081f1104d3c00261d80dd294feb8bdfa0405b13ddd4490fb4f929d3781aea0783ab7d338b7a47a449bd6da74cc542797f70d9ed3ae87343f6eae58be47be518221cb109d8f9061eb1205fe649b1540e9170fb439b6329dd373c68456cf9c9da9748c0bf1ad638e45535e4ceebfd4b2f0730036d2d6201e08f6bf041e91ecaef74dfd27ac48cb8f492bb8fb382e69dfc85f5c0cf024ca6e2c9bf8df367d9405fb38003bdb8fddc172dacab31a7c305afe9e34118c90c6102cb42ad7e0d4505643214831f9bcf615bf466b142899f100fa27ac8e089816c67d4dbd0dc7c51bba10295385193a94a32ef55593db403700a44b231c79e3bfe7bf84e644f3be6d502ba6658d12a2bd3b04af4263dda298ee4526dcc8f7cc45ccc13b543fb499111198c33fe249b89ec0e7b6c1ebd4343e5bd293266850cdf8c907738d2e6d69fc6c633588294de109f425885775d0464af6acc41ff6a0f80f72cf5cf5fe5652e0b9e48f962034c45b332440e7acd23ea8e58b4477bd82c5d995eb0bb4c2cf85b802c0793edb22a2f4e1bfb1c73f83aac65b0456ac0423fccb0d63f62175064c861a1349b7ed34e132bcccd5c28fc4cd1f006aa54d04953b204e03cc073d9c83afb2abc907d663c347fa4f83dfc184b8e2aeba9ea516cafa2b514c779f21146013e8641734e4f07333a6397e52b8ac34a66facf901ea1448d9e9beb6b5aaf08acf48f708c7ed08ca2e31071af4a67f22e31733bfd8ebb616c70363138ef956a6748e4eba1b488da84cacee9826d53e842b8a73945d66f2760c05759a20d8e3819e49b6eea14abc16ffb8e1c2f88ec5529ed0077f4fb50f292d2eec3657c524455a7c5a5b49dd84b07f7d18349aeee0f4f9985c952dfb795b9307219e0c3dd10c493f1fd0b3fceae6debfe9267c101dfbd4ad29e91d47883a70295504182864e2f70e9bff1a4aacbd268fbff0b9b43d96e65c4872fe53db6b15fd6e4ee724c75ad70dcc2cfe4e305ea09e06290ec4a80a431375cba84bdf89f96fb8a9123ade5d93589bf7b0d5711f79c5207e8c27efc42e7777d1980f351d2c561494caa3c8f1ceadf1b183fa95f3dc0140a6a0f0434b95c11dddb629c97a37ef0e496b7a2306daaf618db7c3602c4555676c005d49aad1336dc8770ab1b872a85f0c37b7758df12e3384a9f445869a83fd44d0e7d4b103615ed70add476642c54e7edde964e193b1ad48fe5f7067eb867b7fe8397194b6608a9d1f7518c68dd6e8b5f2f78ed6e87a8a021ea179187b4f73dde5be8d3f02d8cdb91ceb6ca7ad2d245f3dde9145a37bfde3ab7ad639327345aa14f516d9d4f95f915339ed64ef11677424ab1c0a234ad748c511fe0d38acdacea9f396b7b1f658ba5b754e0352f0fd5219932e93b088ebee199b9e53ad619c034c7f9107957f6d14d5cfb619553296baa375e015b6a8fe4ed2301c3165373d0692ee6341aad035ff27474c30c6dff992e990748f662ef85ae4c212f315ee5318ee72fc30e7379b2b987555408e0cfe9f88d14c1dbb3e6eb70b7a026e71b18f4acca46a05205d5b79d294611b31829d161425364dc4f87c3c3d84240252956f1dc536864b73e98a0e6a3ebc45904e94885ecadb324eaeaba155b7230a5735a46368fe85b0d7fac70a95a824d3d0e9f8476ceaf865e7e87961dd76be7179c65d2286f4d40c24e15af5c997535b41c6fd2d5fc6c22f547b7e40c7cdf3413c2c46ef75730fbedc7458a654e4e0ff4093a4c1fb00ece24c5f4d43e2ac700280bfa9a7ca829705bc6b10ec8344dd797b92582088535bbe176d65f7a817b8e71ad0b0fd5c2f553b787dfc9ad8147bc9e58b4c542a926cf2bbc3a9a75cb1e24f149ccfc1a100b879624b7d8c2290ceb63f17d76e1fba3d6e63a2155ba415e8fdb2f7734bdd5f65762f7f0a179216e744164240f8de107a628453bdd167d9b079deb4be2c94f46ad09cd36d02d5ae1b99b37dd77998aedb6dda6492034cd664e2e16925443e56e6755228bdc67adf00a4157108684da9269b965a1613d64c4a0a05f041c17f93f765107f026b55d3adeb6870db7e27d908a94761d213bf2587dde82e1d4f6e6e1a8bc43b28597e8b1c9e6ed8f1a469d90d23ccff0a644f2eb5fdbcf6b5c26d3e859e3252b0e2545f268a2d2e82d6a5f84b662d0cd6a235fbaa4c366e077057efd0731d52367806bf7eca9dac8da594fb37fa51c5eede49779f858d3777949a1c3ffda6c9d5c20c7fb4c4a34be1026c7a1ecf71534b8736c50b310bb7a5c5979c3523ab0788a7e4e8576f26c0cb7defa2018d86018d520188107188582ba41f7933b011fd9bb8cccda886b216dd13ec4173b7aac0d57c61fa94d6f704abb1fa25d9db3ffb5b6d28e9a47ee161ed05cfc41ee94c21292d9a3b450d94d6a7b409566a2ef46553fe2a8e39859ef58c7187b8b9eeaf44c42d3d27d1a0813063b7d5f4a3297bebafcfd1fcc8feaf5fcdcfc85547bbafa643c29e5e9aba3bf7dedff253a788a0b5a7d4a2cca1458ba560c9297827f8868752f3767543d33acf5fc73aee09cacc6ee3a79b1fa818da928a10a5a832e6bedf6020185b4dae457ddd064ce388623fb1fcfe2dd312d1caebd66a163a91dbbb5ee2dcc906c5d0e7a42460eeefc724ca984c9aded3be3bfc513dfd7f5a8b799b7c5c7cd75cfb385714881fb216eb56ca278923c6f6c10d4a05587b296e605d46433391511fc1467df781dc52babe184bd83531cfa590f1b1b529b00a7ecea69afb23a66bdc1b57d86491b87987890e509530ae8df8a32ea93d018cbb9771866ed1eae01fc90113b74a2e0d4994ea00d54e3b095eb9be3f32673e80b587b18b54948bdaaa55d62b2655e2f2a5d7eef2798d32809d5a8dad4fc776b028c1156a1beefabe01bab11e6c8b2502880ec67ba3e782f4a85e6d62baccfd75116635d4a4c4be9074a705c4e04e5e8a1cd24a212ea54cd5fa50db23cbdf6d1490fb117efec965bdc24d1e6cb5711db55f178fc2fb1c88ba0fcabcf03ee7cdd5cbe27718b88f51f296cae114f1d5bfa1ce34eeb3735eeccfb78c3df652bc6e96e9639d2e0e86ed55f7bc931a505525acc166a001bcdc5cf9a3482b52d37df24064af650a7c626859ba657ec47388ecdb5f6de18d5f475bf26c0ae0895236109b3fa86ed4f8d1ed9861d11898c84e1d5936ccaf7654784f99801183b3e498538b7d6c7f98b9401528016dba51654e3010b23c526e72b895d94fa1f526d33cdb0076bbd9bca56cda88ef01fb4068eb2d30437d1d653d77f7711cb691c2237f7c5813b05d6f4c024d574b73fdbae184afdf599fe02054982455762158da552a6f059e083239c14f361beb4370bc6a508517dd7298b6a2000eb1d1d46370fa8af3cd2597e18d7db32b132d0412049d0444fa52ad939eec89fe1013501312c34e9b56f107d52dad63ae76a036a53581f8341023199d38956975d46975582c9d49e36b0ba1d4f3121a1bafa47c8f289ea2e1d08b92fde681e4b1becdf94a7875bc2a926668504a96f32baa70147afd9ac444634484c59b76d91d335e36e896987b01abd776e6765803e84cbe9707e5cb89c879a42bd5191478c81a00ef22cdd9eb74d5ffe45c6d8c25c6df54577be91584cefe8e1fb810f64646c263b005afb3204c23eda2e3420c9a3738a12886527c376bc5d0177c63f916fc97f81dae25d33ecdcbf150f86f3019c78a5470fbb3c272cc936c7d6219722850621a2d7ef91351eb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hd338205a1d933e5e0f4b6494060c3d6140e7d7a297ea7044730e7306185abcea9db631216c8f212e7b5a2f9d68d9bdd3205c54d48757563bd34840ad849b302b24c7c7ebab73cbd20f36e5d33754856a76c89f37fe8f9af6dc372b9dfb539e3d9c5fd0bf1492156a2be97d812f9a9f5960afbc9c95aedfafa3e283d1fe2fd17e365aeeefc47c063357beeb2aed735851f2829d30c0cd571ba84853d756fbcb3999880ceead68a9753ee0f894aafd02147114d64ffb87f0523c00478f635330dfbbe0f6dc288f923b262a8b66c348668931b562d91ae2377759614f98e5fa68bc757ff7338338d90802da31beb5ba6e6047bdf202266071fb78047724db4b939ee23687e6febb3078743d1773a9fc7f91f7e99fe5c7747e1b49439dc17fe48fc59d24edf5aea123255d025b26fa693fa5c7c2ed6b6f78b33b5ae2b4a64b8eeac287d99a025d900ef0cf739e6ce8b76a44dbdbe9292fe0ee9b296539640a3e3b29d7c9ee7b682623fdcc14e05362cab7f1974d240bbecbe719598ecc63630bc342fcb0d1ad6d226e6c18bb281ec8f56976a8a147b214c892e08b08d1ce731ea38c71a29558cf97d4f3fc72459416f982b66ff7de31bb8851c890b3e92dbd11ba9ee1b970d4651f20202b2bd2032b88a285ab0a977fe42bc785b99914ac51417cb2101653fa15faa94c1a567a3ec6314c1ee8a356cadedc7a36ba6a6fb410d0e0364811e8b37c096305d7d9487153a1c6f79d77b92622b174ebbf1fb07be64da31c337250df607c50bf25ee77205652cdb1f8369527cd4651329f9b42d337ce74b74799c3986acdf01faf0f389432a9a7d617bbd40cca900c1c35e0bee4302394e8d12deaea0601237ebc19916e0c816e13e8c2cbd82c58716d4e715ccc8fdbe7d8e2bc4f7fb2f48b31241f87e9c6720c58d6f2133274472abe6dc667d463ff151700fb03c8b6b59649890c526f81eca777fad5477a8243989d80ead13b96db9de5b57182a618a974440fee50aaa107f4419f99bbeb2eba5da2c60a369683c552d18d697be244e41d740445f9aedd0929e0330715c00f4068c087fb8ed8dbc0b6a0fe075f37bf1c93bbb35d1a1c2262a005c1b7be9912ea20a9be7c04bf6c19c1ed20ca0358f8655c8076989a7f334e816ba3c7c5927a0eda1e36a397fc4396179250da6edb171343273ebf6276d4e3a1812c7a9aa7883e28d5d659da2c134cbf425da4b7c86bec55cad7120fa906cfd1b3c6b245d5e1e01e524b2df5973630bf59643e2308d623cf807630d86c3f661745b9fc8a898ef8670e366a7223d86dc92cd47dd89cd42a5a86c202087ee313c9cc00c5672798ec7049cb9f98b1443e834cad1bb9c9ec535e7b9cd4486630f5b745f22a88df1268a6b79497c65fe1ab264d34621eca832f497061b02b6409933946fd540832d3a1ae08cb34c7abad87d90ea868f753f2008d5e1a3ff4d9a70e702d25bd983dcfe057f6d68750cf39fcc705e99973ac5c567cf083ed816487e5a2c5802223c3e2041a258d340bdaf3134d363331851e48b4253828b5b828d66ea458565ae872054c5a73281d0919769381b4ed8f181d56b438d1efe215db61d494671367d0af6383469d4b3bf40b6c1212db0a7a512a8bf162dd50e20f9c01f538a03ae8811e8c4c44868eb051c38c88e3ee6882f56ed083281f4c1773385a4b969ac746fc09e5d286214c9021b3483d7104d9ae1037d2202d3424f4db00ff5c8fe83e1fe393dae040a1ede742dc83f06bd8c828cd5ed5912cf9b923d1eee795c78ed452e1891cf6ed9dc871427487d4afa7f751d0ea06437aa1ccee05b09e7251689de6a39b7a927ff7e56fbf0ca2cc957c8f86f209656944f6115b82918e343d34ea978f178ec02bf9a06f8217b5054d46493fbe3c55157f42b0d996e5b884a181af50bb7716cb8cd81a2d11cea49627ac153b8a26795561f595177be591cf17d5598d87d4e19bd3b163056f1829a5c3d976ad6c5c6a38e25506c9ac13538a96b89ec35a7458741eeabde34de03e6f1a50efd0c7bc923554ceaa5d3d304cf20575402d20e1dc7e51d119b5fb597f8e26a23a1b051e508561db73ce8c8f2f9da83efceb848042779570b7160210be8c05c9016136ed843f126fd059f36ee64a3446c5830aac898d25be31a0fb9f5bc4519793898c6084742b157237abc0c13141788a0953e1e5fbdd6ee93d7ec9046ff5959e5e19f8b2be08f324c55f41b3b4bd53196013099a155f36af885608d8cb4faf898575fb5914e461a1f3df1b24b8cf25639133b9da2f617fb17725fd55f5185c6895e3d93fe52832b691a1448406442dbd5b03e6c55a1e7218cac75c641b232919878521630b8157c8d779fad83be78f6969b09cdf7231725666fa41a810469e0ac5af060d19000a62ee3ec58c24c51dea348f5a0a750de49329aa07392f5b31b80f2c2e9bbbe186916a59776b1c40353d2cdbf30263b609d4e76f9a51bf6f9c1f5af5d3c75ab2afdb073ed58194596e79bde1e4135e12caf79645f7b35ec052eab2d1541b6766afb7894a565de3cbb00ab5762841e3841504a8d70fc29c37ebec44aab7aaa480ebd833415313aaa11d977e27e662450e23e943879fc36ffeb7153941ab5a8f498dc9716c2e23dba296e5e5bcc20b5bb50887a044b1aba8ebd0bfa33e649245085bdb6e6816a3fb9a32db7202d16f7ae5ea36be174ad07870457c6fadc4eef5cde15c153284ce8957093cca6d00e0736da78a2d1f21ac4734a73f7aca3de634fa401f96842cb563547416d87c5ac319800d3bf753ad598e3b43979d6f68093684df6b413d532fdc6ae5d918ea0203f197f72ae3d7bc6ed97c236013de0f02bd0bbcadad5b49462c275f533c9301027ee0690fc6e45fb0547500a7a7387b4d52365349e614aae3b09ddfc440a71b5f226807924fe67d069fdc11471b84132078de11b6a9b6f266d48383a75cd8dc510635a574e2ef3d386fcfd25c78db5b8bc686587de4930ce6564a6f7e86dfda375480d7060a33ee1dfcc9af56c7f626c7fa4b6431a94940570affeb11e863033463229ba7c53bd959fb4e52c3438dd1d18a48c2fe70113c9bf01640ec7051ba494db994c2401b1b13706a9012f205bc97a23398b7c6c76348037734b3a90f656f3ab80be98d178207789935750215911c93591d6d1e5fd10e0547a74a5af16ec7b71a03fdb8b40a7378fa1212383b1dee73c4bc95c849e55c69bb5a95b0ac9f3a3a7c10edc6cca5d0783cace8e954a2f0fa757b01f984cbf243b3c55f6c9bd4441d1b1fc3b8b0f140399147e0bf754be9d10d2a89927a59012d43daf3144470b1f5e547e78974013c87d807c7bcc10099b5b8221502618b92742f4186fbaa062242c79de7b43c9ca8bb045eb3c9fbfe976e818dd73640bfe8bbfd9ed5606d87cf945179db4d4852c44fc5717a8efb3ad165dbdbc2ae3d5b150ccbfa16f669dd60de797a0d12b95cc74bf402255422bd276c994572fbb5e82e591e33261fee25c352150c0c9d861352a404b9b9c7dde9c344853daf0276766fcfa1b85ec3deca2a84c3b2b5b32b687098f13c05a9434f89945596cffd780baec136b0183d2d4ce78168d308e4a40471f5362ac2784128fd7a04b962668e92f0d1a7f18b7d4cd14d3d310a26474fd2ea9329b09534c29e7f9cbc434fa089db48ff041dd73473d7b6566bfa57516c00191b60684b5e473801841d651a2ee9ccf725650ebb8e9127fc9b58753014eab45f1c97b410728446cf36734f4e7948747733923c5d0f1b923aa5080faec315acd869a546b2d21f4c1c261f82213e6344523d51465b0a0221e2250ae22a23f759a16c9ea7617d902c85160e2e75f91de8753dfb2bd77152616c9a49afc27ba54e27c1b49c28421be7fd4a8d80626c5618fcc7ca843376a65f40cf9d6f3ea00d38e78e1c0a161b5e2c801375621e79ab5c666c95296d825c01cc1085d2d2d8788ed1846876b2cc242194fbbb6c649c82bfaadd78c0b802a9ef1998f326437f9cdf0d9eaaa39af676fd7651ff6b23bd1d38453984db316735e17a3bed6d1d8635e59155e53eb6fb0c3288945fe3ed9afacc4b4b63f991969290334092029fe6dce161a53e7b92b742f6ffc49b734fef2a61964f2584bab3511e04dc2e285f38c05db486da0675ff8e76e0b5db7871ca2325abae1f90db75d5810e7580db152d485dc8fd409e0bfd1be6ca740776a1119440879c5ad1e43350f3b6f24c450217d351829ab87c6e465b170099f954678018fda886eed3505d9f885fffb3019429175af21ee213763bc4096f1758fc7adda6077408b146ccb3f8c9aba240f78c6dc96b450db29fb3b9ffd1090cf62424b729fe0be41efa506e8d80241493eeb41b69a439f83a0612b167db518956080d53f6dcb980aaeee62fe5791942d46104cd6767081eefcfc5d694b868b635d1ee4be8849a9ce1359962f559823ce8fcfadf7294db3439cf7ee81042aa5b413aa7fb3eb369d92bc1967be9b07d9bdb3fe2e3f54284d5e045091560b1285622ded0e53f79aac520e9cd9cff155d976ec83a9d33a663faf3575c254ce03e02d824fedf482f0be10d3686efa19a50464a770456ee38392cbc367a17eae20749e30b0e8c4ca85596d82bf3a8ecb1cda60bb1a6fca207da50f57b3c4e881d3a2cdcd827e99d03cbcab852cff06d0e6e8ffa49b4968310b8c5961c28069625e312a547a3b4cd4b5902ebc73790c4c80607f814ab902ffdc7d84bb17e6aa7fd0a1b49f4cc36123a1195cd1c71b35549ab9f0eb350103cd5d551b34bb1b538775e7abd84dfa2f00897efd80e50d8cf88ae47fbe6a81631478c49a0680c5ce97d4341675b99919ff9229c43400f8f56de125996e7514b3db1023e1ad0fdea4d401474de143f6f1218685978dbe2801df143f13f1d93332c8a8d4d7bee6afc1352318dae9ada5f558b6ec3a65a9662cee6c96b6dbc18d820f91356f602ed99743ff8d67bfc5b229ec1f506a31be32e7183e1763508cb1694a3e0c6bbfd63c0b5e2154f14696c6dcf42985573510fcc78244ce1ce3248872c51da5c4485c14e546379b25e70793ba7d32470af6c3a92fc60197bfcd617fc8c09050c80174e33f469d9adfac132ff0055a0b1d16ba165bf94ccd176316b076f4bc8d4bf28859ec42054cd55f670875bc6641bcc312b68cdc8df027c9289b566d72873fb7ee6cbd3dab3aef65904590f1fb171c6ecc134c66d1910732bcdd9970b84e628756a7889035a2d7067bd6ff87c0c51e58f4405b01db843f07d62b80eb2c6cce24977860029c2b652f44d170842b4606669aaeea478d6598715b4ccfdc427e253efe4a4098694e8343065ee5804fc5340c9b9623d7f9b09a50dd2cc43097073ad25d0766bdaf65316837cb9428d9076a7af977fdffca75d70bd11653fe9e0725a241e116ffb30f6f4d5642cd002414d741f38f8795eaaea78636fd2c5c8327f015d279a5553542077f57ab2875bc82b8100;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h37bbc3a8394ad3d171288cab93482cb0b0c0dfc719a8ac4dfc5b8ca4d0ec1aa96c83df2952a55ea5bc0ef83da3822dfd73ac0bb591402f07cdf984d2e1753cdfaa7b409e7dceb4909b8373aa8eaf764d83bc98ecce79e9654794aa1afe9825b641fdb68447f82d168a87e007ed5f604b9067400603fa438dcdb45aa14d6e049bdabfdcaebe4f18110230a0caae75e4e29ae2283c568463925d2f00a2a5bd5f8e411ccfd5cef43b92a7f8e4f013081baba01308072bfd1d3272b468d1b3d9e98a88d526aa4876b28c1b38d52968f86d12534128abbab31e97ceb52d9884860737c23481b729c17692e555fa9ee537bc4fc217b79e0262cfc309f58b8009aa992651c9ddda95bc741dce0599ed219022755abdd0e8b891366533e0d78ec7d03ceb535b6d418c52444c16131a3c4678634282cadb1152478a7821c4d68532fe1d79e73099a118d6a867832c7f6755c8ebddb721438e57255bd11c27742b5bc2cde37c3a975275542e344c93c9e68954cbca8a0bb72ea81e5fad64343739b265bf96acdcd1311908a20ef03de37c8241c6773f2c1455c2511b63fbed4afcc5949e996138646a9a7b815b99f73944fcbfe53e407a552db129664efd13ff4b8a94334d5ab2dc5d1ca885b5fd917551755b8b1d055b040cb0dd5d685bd2712ee1ba6f055ccb52f82c00e27302f9caa2d011a75aefe395c0621ce1232c6b0dccc2390e9c15f83aa54a7d2fd39f9df885e51e1f9d18f4fbde2adc31f2e79bdc0516662c293a70fe73e7d111b6b5cd5dc391498a36bc3ca1fd769b866cb548ddf27412c4fdc3979301b3a429788eb11024f8b533e7e83c03444c0f52800001177649663cdc384d0b942fef4b9fd1a42e28d45b3a9d3179ffa0228021b30e5463667cde31eb01f180db7fa1d7e6664b4385287b024c1fa31c0d040467d21c76d3cd09ff11188924615aab2e9f9a403451d89800db7be532f59cdf4b8990aa08862f0d2902d8a35f7f7fe6756c65772eab2f6cf72a7f543aacae9864c8fa0340e03cf3ee70100d44d86a23b2b270cdae9ae6d4311a9738b29cd4aa7affb91f32944ad1d8ec6c7b40ccdf322bb050b70275c6ac2d5acf1ee7e896b020a893f3476682b576699921a029e3b013cfdb6401db443d276c286f83de4c8e4796b0351abe0b776b9c2dae3e04d3cf17dbd652db23a4d5d2117e40e83145139a90034a31cea78376370c79f7c044336709d61c029bbfb1d05e6b5bd770ea106320bf9d63273335b59ca6e72d315ddc77543389a4332276db0d06a33891c19e2913495f08fa82495e61a543603e170228ac1da4d428acd8806770dd555641ec62d44466eb6817e2d6dc138ae7158a27a0550faf7053e33e80fdc8cd0dd3d7157954f317b3816c9d024e9d1a13c886798d10617e2d9c5146ea72a545436941f84a0f7771288f856685879fc911a6089d70c404d38db46ce3e65d51213a3727d7f3fa5ef29b5c27740f2ae749d1d52e686a53d90e1e0e5e0625597457cbdc689a91ce5ca590c4f54b87e5fb9b1d4d528355f282ccd386779c32536ff27c5b17eb4caeb04c06d0aba84c703f3d0704505ccd7001f538ef2bfe61ca79e177644d381091115e7e88133d38588d182d7693c2187d17dda3587c3e964dd722d3ed0b2d76df00a10660923fc48e881f25a7af29cd7b7ab25dbd901fe0e9ab4254ecc90502b1cbf4cc6161bf23ddcdc52df2c1b82c62e566ca3ea4d148024118760b30f5196b575e2455b47ee5322a4f4ff9eb0c973286c595934d741876fff633e28d8a75db2753e4a1049e10ca8edd19d024adb3759a5851faaf2ad0e0316186dc391c6d954ebb9b6823639d5f9afc90ae1729e2695ba711c36ba4f92d5be1e665be3f9c3499839430aab361c1beda894ca0dbc119d040c455d8c615a5d339139588162b31eeb67a5b0e9382c82a28ad08a752817a4201558e10b3bf7bd7458eed1814d565940716df474863bce2613a194fcdc625361f7641232f22e3a8d1906f6f6a2307aab52cd87960e1be0f9cafb6fdb3c67820dd87448e077982f65c809f687edf3d9d34d34bddceabe0cbb48cb8f233780d5753695be9099b6003ad243afca4ca02e44a2d432d5e0f438196033ed7c5534f54f2df88329e81b83ac6e61defd20edbe387a06400557f20068f8fa8b67824c03664751a0cc60c533f5171e02b54ea162d51968723e2f59b5382413d069ce478012a64e7e4f4d2244cb54d52e74adaadfa3784bf6623b083b5b8ab172acb7fd32782f5d087b476bc8cecc89dd7480cdea24e6024ac87e79f0825ce3af6ce91bcf054bbcc684777e9898761c6f2f5ddf8ff3fc738ce98a3efdf5a3f6410f6d70569ae17e22d96e04f4bdb65cdf0355077c21312819cc8f5636a03be5b8f3c21812c606feffcbdc4f9fa708c9b61a3a9a7f4845ec4b1b0c2aadbb7a6dd9b262fc6ac79ed5efa552000cf39a24f2f813b8ff6972b04b42aee33e921be4fa0e0ee4508e00e44b5989176b09a8d8de91cf327ea67929757cfe11edae5b0e38b39e285a46eb5fa4661345b010dffaa902e785b90b957d63f9361f49dafc0ad475001248260fc9812e25bc9e00bd3cf2aeec1f0c06235e27e1c6109e15f280a7f241753da361da6033861057231cf75a139bd9f10664e9a8893f0e63417965b12b80f32ef98f097268cac2952c2dcbb00178d7dab52b40130c7a111e0c8e81ebdc29c891daf0af91b532482740dffbc4a172e229ab859b0344e696a87f79f208ecd5d1be7b062411ca33cd60ff8d5dcd57b5476fd534302d76e1400f71d08e693cb3bc806c73068dc1a9af88e3b202e41b050dca78a7470f7c199d84188869ff7d0e9a8ee9a9f8cd1b1ff786e88b6276450aa1772e03474b86c912e48f1778ca60a6e0c2dc72b7d8a69d8c05349fb0ca50f6addd86f900b4db7cf70e7a83ce8a84b7345eb40ff9d3fbc72d6d2ce5a00c3287b3c751b2bdecbda84f9b3968315e36b3bad9ffee5fabdcb3d4f1ec4c38b41f7358d0416f07fbd013e55318ecb74a9cb9d502651434f6503c6a7df2b43b04d7ade1bb3381d5c8806b69ec57310c6a49872ef25a48d8760976a1c1f5356ffc560044d7578bb14ad1f51280d556de60e1f3c4ca9d12e391f82254e10fc66a475cce2d5361c7b691ed541ed8a205b8ea0e9443ad565a66c888b7f717cd89e5bde02f52c35d347dbc7957760b089680d66a463ee61e267152d5a7066f809ec31ab05f8db129221619656cc31bb27565c006ca455eb24207a0162ccef336f9571987b694bd51eacb1ae5ded6c8e1e1fb01c13e92570f35d822fae2f810c92f32f5f235121c8b6314dcee40f5e92aa0613253e00db753560193562ba25241e31debb9da8cb29a5a2916ba5ac4ce89f9387b899d18bec277d8b0a4f1ea582d5e8213b221bd3416d1c1d3cc4e980993e71201dc3282b13b22c1841f751f468e4f9979c9f2ab0f7656b449e908ebb6a03bef0eb4363bd49dedbc5316c841eff1d5576dc229c00f6b2ade33057303933fe3b1d0474c214e69340af8717bd846475c9fc232bc5f629872d97ce39689e7a116b297919ea143f59412c23d89929d60e3a1b469aaa58ae0fb2c317340c36c00ff3050116950c78a7dc8aa9602361b4b25c7ce4e7db2b0c7135e558eb3b518726fef94dd169905d10caa587398238b067aa6f064b89974b4ffa95737d9c4a263c9316e166a226e1f240fa7f64ea0b7bcb07b9135827e3cfe2dd95556ce9fee4bd08fe3bb203f6fe3d0d123289167664774fde700339e798855d19bbd6054f6abc3a5b2f8c5b4f0dbccbc4bf320b70be1ce1387ff3024d4f1c9b1cc0fed78e91d64e8677c0d05388026bdc95a10351f0a48e7637b8d3ceec916b946b14b1c89859c0557813f52a8cc4e955adc8b88652363cbdd2f412f168fa131eb4e823d5010c1d350fe872b46984a59526b737ff9273a5263c88687f3d7eabc19877fb4b834abfafd047f63b87645891a09d48f179b8562546a307cfd04cf739d9b212a9dd05bbb92f290757a28a919bf25eb327f3bd13c2d4cd6c10df84fb0d451b2d47def52cede27ff6a7b1d0875665871398900044d60bbbed4321233b32fad4c567a065ae8cfd0c30880358aebb050160e260cc225185a2a83ee74ec35920ab6fd707bf53ad61a19005c68c0ada26c88371002142bcf6174d4c31d1d1aca9a14d9ca4c504135126e565c3cdf113d70652c291340abe5bf43d6ebf6105620b4e3f8778d39b587b4d7dd7df7229535a09dd06cc62055e26163e36f84bbb1e4340f0b433546a3c9ccd7a0cebcfd9ebecdff89fd8eea4bc1e567a3ddf3cede8af323eed1f25f362a6c21f3928f378ec870179705eccef358027d6a998c22304093df2c15554d39c4355f15e3e61646f1eef7cf682d66d331732c9b92a9e49569a43554fe3a148a921faa5efbac88b148b23e490fcdf7a0054459e8da4d90dd0f6a29514601957f29faf25cffbbd4048a8ad2bceca46975d21833a6b646bd55124cd3c65afc0702c3582e415b2e9384423622ec7294e13cbc9f69a5ad6d92334125498b8799df02e91bff515e48fbcb2a71eec3a24a704bd23fba5325d833bd238078aeb88d51ac9a04c23a5ba21a01ac2b0ea4bd9f4e7f94e4b1b49287a91db6304edefba0c96d39ea25ae822fa82133dd6f71320b314756336409f44984fd67eed821557c4ec500172cf876606b67b45a4c0b06a7bf0f13af06405bbabf57ca1e0b26fe49596db7d5efce57eda0a04c9c0f01f46d624ea1acf81178e2c97a8f7e29b1680ad669c49a3cf086a56371eb84e2be80d50e30051ea0543844abbae915708f0a372bd742e95b7d9bf773e0a1b00d0b6ee543999dc267d4ee98fc09fb417e4a4ca4bdd8a0f84ebb33b64c96bc7982159a30d73247acf92082f34c09cad69520a30fd7705b60623642d5fca7877fb5817e49cb59d7badd88e9c112f9d963b5d19a7d0d665ef4bdae459e5414444d515aabeffb0b2e83d0c2e21db7d008dade4c2cc438de5a54020aaea6b611ebe84b36c7d6849c253a469bdbb9b057054943054650e953c1992125fe5e234fd1ecd01079f6193191d0373a7335789af5685f49ffc4a182d7013e91f01a7db0b5e9ba08c91dae48365b97f36aaeaa40eafe047546baf2fa4cd1516167abf35b2681bd75c22d9cee106afbef4a61b5984371df21cadca32ee349075024491077977a8296504e4a893a9f7ba0b7a5fcf9be2eb6cfeffcd35c573b77559e202768a384de513cc7cfa17ab681ea37e8a6a6dd63f4487fdce407c7edfaf51b302680076049668763ea4929c471828cf98a6693a8061bed7211ae2186a05229e8612809b74b8a8be1087a5b3697f410a82fa1decad017e95f200648c72d547e43de43ab32620f9a1c640e192643e7318b50d1f4d290c78808122fcfa6375488d9e73f28ea05d3555833d2dedb738448ecf32a8a2b88623702edc8352fe355d4dd63e33c3d15777b3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he7247b429657e5db88187307b8d7c1e90b67a5a260af4d99798cbe109a44af205218c0e35fe0c70147b96b74cbb1f7b2e887587bf21118431b5d7492b7636cc33bffe14d7e5ab575084f9bd2222957840fa3295fece6c6b9c0b81954ab73a3215f176b3cfc0903e8dd997daa6632d10df4abed714ccddb370e03ababec0265bdc466f3a678b60c8c50ff19e2043b5f268c49f83729a79a6ed94dcf13c76403c5acd6ac31780a25fa35d3822ab429aa3164d65f3cb691aae025fc0097c0ec459a3a0f3b9f579c636b816e7ef56f2e2c2c88f258d42d610465e5373ed88a587a69040b9a33838e2e0b4030b7e14cc37ac466608a8e2b6a7f4b8dfb55c1b3e9d51c62f1618e96789d54454610cb8b138f28341b6bf9719a2314913f32f93288f48300c7fa470c2b22981193d4c4d02dc1b05f0bf292b3832e648981c0b1ef0cc034a8c2c374b52a43e7ec8ff237a696db167d550e11fbe7066a822e45b918c4304f388eadf4d15ab04f7c4c78d4d34d4584ded8e9b17e5242c87732f211f95bc19fad7749f29a79f09934628aea22febc176472941119fd0556a336f8020d8fb80dd4ebd5f66707f01c23f195a9cea0bd406c08954825c982fa12379cf36a34973ef5b1d7e029886a7b1f12952343a42b65f1e7d427285dfd9d6d499fc02f0b3a66e57f9aea877c875e27f8a1a01e36c3a2c9cea8cecf7ddc7fb3e61c35d37bc5a8f2302a6be6d6005a502e84ed739218e4d7590dd4c1025753d5b81cc3f4f99f7ca09aa12d9ba4d95815612ffcb304d52e887a71c72292bb8c5464747f05dcfda708ab5ac2815d29838f7e19112f5deab49bd1d6568f3e4ce7339dfcf073729c717574221b88850f7f90468a30fa12cd9ad434cdc2c548a43284e0f3fdaa10fa9501e918d1a7d1a447582f19bef25ce7c5ebb8a593562e3cd723d585f33682bef183650f3302c0381fb02159f479888329b20472b20d6264992d76f82ef3543c0aad403b62b27d12c9736c0a497375f419081a675db6a6399edb9422df04e547c2f705b139ba89a62f2d76db9cd60768a3836cd7cca6ef16063db900a6323eef8c65622cede1e78c24a9cacb1bc3f926a5f8e7b81626c73299eface45d9d66e34af7a3798e06a4ba6b69d738efba160938c20143fb6f4913628e335c3a978ed9d8e8182d9a4d929a400629ed4b576b1060712e0dac985a08f11a459aba02f7d51ca80130de08c42acdfcc95888b4f82b0d9d6a5312b51beb998b781be4956c27e11c65d46b81c9b6db0873206ccfdc6c90f0e3e205e0be9719cc0df75caeca5f94819985090ac1d3bf8e2b8d0f92b7c707814e8ce760ae46be78a2ac854a51a3b51a99c84084640815d96818f27f3df8674fbe509df490937d7d786991fee6dde5fec48afe9cc1add6805caaa4a35499dfce1ae8112b0f3707a979d20545311cf02f745a763f9e15548514bedf4df5815f96869adb0ea0c4842997c1e619f7bd074fd3fa04f56cc64f1ae2daf0920e7ff34ed949a00e1263a7a6fb46777e543e0f5f942f91fce3beb492cee5d00ea558cf653d79a2cefbf2954e0159a2f9f80de04971e1cd93b44922d4b17157d3159954fe3dc2a1b06acccc02e6942edc4dd16823d0c53ab151f7cb60564e8137e438f0184b1f01b15686b55d1180d0b3149d843b5546151c6b67018a66234ba81046eab15c15f79d61444a3375cad6c766ef04f145f574456b4fa136de7ad84e70278b00ae455d89b9e9452c9974ee277f4bc4feaea70c5e2fd244454cd61d867990ef127bbef66b9f66d47664871e08471f46e76f0a20e5cfa56066998972bb8033812af2c8ac42d70b18a61a5e9a9d9f98ba585f5be1b0a17970085cd7e2303434df7ce5a8b43349b232ef69cd4733ab8523e83b6251f6bfeeed0b249bacfbc512c2dbecde03d2cb6914a9f654f1b2a3f994fd4d9edf22213b71288ae4b106b345f36437f07dd5e51f77bd648f95f23673abd2c5f2e9bc4a6299685b4eb6469180ee6045a4049ba4b9660af4f7845a78f63f44ed451ea362cb27ebcc50bb126d86ca2a1c3e1cd4c45408c517df8419b928e4cc6ae1b1620c002fb542f2c6a6b0c2630e102c4c039d6bbdc8ce6caa75f1cdebae972e085bd09818cc72bd0be0cd2361280750cd55482ef53b7b9c19fe2846277d8b67810d2ee4c654e2883e5c6b6b81184e92f07a68a217bf3f35418e90eca92d75db10879157422c8d1860709a3bab060096757a4fd810f2d4420e5726c08eb9f502e7b37333389e70a9c385e03e84560ef0d50ad5463609ead5f8692ab6078ce97932eecaccf1d6c63827410f59126188e87a137f6c0104f7af110cc865897e0c9f395e54fcc2d5c88e724bf581128a2199464eef9247e7f945777f8a16b38f0418d3874356f3c25f9ba5b1b9b907d43769170ffa19b9f3e607b672b13cc1ac3f766721529d3e25b94dbe5f8d8e1d52d94e5cd9a7a0277846bd8c2bda2bf11b790719d0924bca95db4032b9f4617726ec601cbbcd4bf716e247b0980fdf2ead913b63d14839e369669fb12e817a120ce755ba9e274b69bc919b1abf2902f488b774f0ec6a596db32f7bc1fabe0013bb5f192f7ed9c3aa33578cd16b9631083dd29252461ad49541eed7c4584c5b9a34bafff239368a9435a5697bf341805b6e35859922782272a5e0a0b1cc17c475087bdd5378dc3fd3a770dd0e80476dd3681666d077f0fc2309387f17f26434c0b006626fcaac1259c6b721298dc1a0f02da54910c3fc631197c473949e0cbecf1d706211f7c0632b3f3491c80bc0108228159328afee1b203aa57a638ce3058e1bac7aecaf3fb2ffaa504a35763c130d33183da0e81f6abf081a4b122328832f3bfa4170e7b9dd998619625f6bcca03d936c020f10853a848b8ea6ce18ab2c6cd7fb2d51708b61a0429db714e7190bb2a7a38f678fc5e9ee15b16e8a45c724ee3d03a3c401b5a30b32cb3835e96fb7d5debf71c1e08071a5f378ce2b2c1dfe23b5112886c4c5d042dd220ef4f56a414852e3fd50d45c904628ec939a538a133dcded68ad5d8748c75a5f6df9f03130870c6d0abb6102d0e1ba67e3f0dae9b4d12bac1e6377d7102116f3fcb5324d519c1f529732ea5a9d3aed9c247b6c56c3f8f4d338fbe79913343143a655e2f6b3cc9dc19ec38616e678e79003db4d71124af8a96822d8d4db7344e99a50b10c9bf722a39b04d60d647b136c3b292e1ad8dde72b54a33f2d21ee2fecfc805f75068e1526284907d582d39b4947f5f059aa7e6ca44a1378f1bbeec336dd54b2b425e1c53b4841d78ad7d6d8a6a7c7ee1f49bd2ba95b927c572b721b0521b223f98eb32106cbb9dfb86c2f879c025c3a7b2610f42d239d78eebd6c1dda1d04e00ac2bc0548b64990eb6057eea01802968a3d950ee865d84a840b798ff465d6eff624d75e4757d64c8e54a44cff91d378f2277c09e4aac2e2bf56a292fa9ab548795549af8e345e3df71eba0426369a98f2d176e40f38510ec3757b37da2594ad4f9b983609a1f60a4c2eee460645879e303b255681ad9b5b11ef2f2dfa7516b7436adcc75363dc8294e33a5637ea7838843045bdb15a2eebae457950479b648c7d4ab9c19e9156a686de103b421c52e0b2a1e9018ada7dd9688af058a739a6fca6b4dc25cf3e8971a399eae4a8829e76b3c562f35a479bbce0b11b1518471b204dd33afb7c5dfb3dd888066c3478c94e82081e55edf68651e52343999ec9dce11293bf2f3f4181b06b0be0606058efb6f2f19a6b6f543a19d815ad7d84d777e66e9f6f9486e8628cff1db4d3aa8ee16de19806bcae1d60418ffdc46ac6a338f858f35689f2646229895c076e0a615709456219449bba19f5d624268fae6c1c6aa039de3d3c76eeed0f1736b08f4341d21521f9614f26a58410e5dfe26fb87daeb79e1cc8bc30ca6020ae7f942791fb2b7674c7a71d9f040ebf517ad71ad76492b34d0ae81155200fe2bc0754729778e73d2762ab1439beb118772e2986bb93231bec9953b6998e7041b86a2f630cf92a6fdcba9a7bbb425384397dd99b124f5dd4226899c09d5e17f1e642653e4db52eeabe1a2ececd0d2be912550d1cc5f071e1b64403278ffb2b807c0b16c5674815d00972a0d0bf89e5ebf4119936dde11333b2b2e6fe2aeffe37608efef0b5bc9d195c1099768851c76bb40cd9d53b9a804466d64ba59f18cbdc0544efa5f23c6c8cc80675abd5086cae22a5bf80d5de4a9b347dcdcaa114d1ccc320a471726e0c26f25c9fac730662f7de98b675b708e7b0755864c8c6f40271ed347c2c1b57f520146ffeb59cb811be3dfb645e1d9b8e32855033153bee60962b8c3bfae8983ea0fec26ca2cf2260609e6f11bdc089a056703db0c532877f4bb6de0999fb46f16b5c9efdd684600743405392c54e8c3170f43ccc7e51bff94403b3db9b6d5ef0f78fce0ba002d930b95b6e1a3d54ab8ddbb3ab8e5c4430c123ad37d86e62e844f2144603a04ddf344aa42f125d9916364ad80e5fb7a1ed080554b1e508054fc533b1603c04287fa6a675c9eb2d2602ce8d9170a9b2cac722ede3859478aa904be2fa32c7d6af69e38689cc3e995f3259f263db56fd7a0be1aae84007c56546866626f751c82e87d288171a79610209d5fb1ce1ee4f2c237fb63757e41191727895c91a5a5306b6bb18406ddc364ec8cf3d4d8a443e1f01a455b41838ede1f461c899b283d53da63af8eba61a5e65cf7e19073d959e7cd1e3f1e49387be1299ebb8a2b6cb4d4763a59a4bf151b42b5ba34ece4097f4ec3becfc369ea580454066901fb1ee0ac04745101686b4e643616cdd7f10cc2ceef6d1efabdb88ee4f679d79f06d372bb9ac261a5c7b41b304c249829cad194a02e1a8eaec4a76d8c3d1ea47bc63e011f20ce961428c3eacc900256836a53abe8ef91454e329c440622149988cdfc7a222ca40b5c0b7abf2aab74762503c874fb2fbab593c877530d9924e43f3f68b289a73290bd319589d5798d4650ff300f1e50ff1872ac61ab17d4607d592af56c68ebea8dbe501b211b5b65e0f8b95d435c59aa7704afb7b582ad960f82fe0808c6aaabdd5e352bcea502eebd2ba9d34dbeb26cc6d7b82026194896ab6756d63ecf5eca0022df68d53d66ab59f6af64f15a5a5812f0774384af2f419f1d0204760e2069695f621df89a1aca0de09894d1b9178de97c24cc09d0a672aba2b60896373b3e706cfcec0b3236f6654e09794cf4952ff8868c92b8959a7fb4f4f08b5562bd34af0dd9dc9793fab48f6375fd91d93f4e69be07659d3194a5d847a357c42e7b7b39eaaabf75fa72a253dfaeeb0ee451e38d934b759dfb6a769a5bf57f92280cdc0812140e3e7387b922ef62f91369663afca152e1cda120ac95eb32e1496d8836779788c72f2ea4336bf15afb9c00df7764656d73846fab0e3d8ce6e6d8b8d76d02579f283b13ff19a5c90b8d44018b1c31d032a6d283e110127530f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h933300fe534ac9e9504a41ee70a4799d242909abed2bc415e09bf33413954dc3c3bc2bb02d6c527aeead1f91c488fcf51ba8bd600e1023f753fb7e2b5eabd6f514c6844f30feced4fde42fcd7c3cceb4d89b3bdfd61c26febb85104b9189b1bf2ee4128fb2e4a7e012c60b5e2d1feef631f8b929ef623cff426ec0590480006b44bf3adf74a1250283b36c7053ceedbeb9c5c34c2411509ca07374e89e1b71c0cdcdb24357d57e2afcaa4497e01c52abff4919080af675861f3c2028ded1c4c624c2f496c9912c93c70daf5f91729f1e1b02dae9224a592bfcbfaa424ec46b89455c6b4dc68fae6259f70f8f1afd02d6a253a4c1a952d97bafd741b84ac42adf95e7f71992630dc8ce9cbf88c9ff4f46f1b0fbb709caa1f9bf2fb0a33e70e8bd7bac9d2f81b6c6de57de42fd0f4ccfa252e9e1156b5e87b205da84783e8e4a715e7a32d2fa3c039ba65cc4c1217ff99aca6e95f7e91c9bd646221263dd832b98a63bd23b50cdee1c5812b7dda667d17fae95a1c611d85f7b498dad6667aaac8374883801323f6f681ea46b415d9a40806e37b866aaa4b3826962cb563026f9620d1d8a3b9ad3ae095ea10be4f50ac2074b902c8a1f290b1cd86e96454a90f50f92aaa68d8f9cd7bd6c8db433dffbffcb748f70f38ec5c875f9d7ffcf15fabb2e28f659393839f839a4af0abf4944a9587ee942c83a44813296366a17fee9561ce5aad0a6cfc17d0e9f0ed7c9d64690fc8df4cc516ff0541cf0f3578a030edaa69b542b390058a3d8d8feed059aa75754385d976e8ae8acfbfed804cf7d91df26a9cc9422d15b54f31abf7c642f9cc8c3f4b97ae321a13044f47a6e6640f2b90454e22138d5626d120961b5ba5906ea901e2c3a00033ecea5bdb577c623fee89b5e08784cc8a780b1b8e1445e9a4f63c9616263a850420f153566628114bca80ff3583af610683d8235523f2dccf3d7e72dcc5268d339152af2b4c5e1004407670bce814e9dd91fa413dd61da4d00ef13f606ea844f9c14569299c94b8e039f50c2b7820ef7ff3c60e72c34c73c44326ecef707642abbb2271133e009e0ec270ca61eb9be6a7921a9fc51184ec114f42ccccafdb1c663608133af0f03a18e9f377bfde71e773f9115cc06c8c5d154bf33ce04425fe18497f48a1d86130ea8008cf2938be66de0d47e0d53a491cda5dfda146f7863822c20a24f8f6ad7629a9a360fe8a37fa90bd9c83e1106aa861efbff58e3884bacf62460158226c661980b059a5e32e946fd28fb1203cde13b53090e5ff20b7d0fea059cb5e1d43535b846e4127de95d3974dfa8dae8dc82442e9426f38a925db108237ee2df62ecb33eb6bd0590e485cfd0c57656c622ca7d3bcc96152a910b959cc70d1f8d6c75d109978c08b5f4fda427af25c0d9054693534208d60b7a66124e0adcd7c8413dec44674fb4c256512f453fbca680eeabf1063e802f6cdf2729bd62021afb3136630388c549cb6f54d983dfde4cc1799375ac5414684c25d7b8522afb32c53fb2ff301577fe48d6afa7bbd87a11cd7fd4f9b722f0913823c40dcfd233cadc79fdca03dfabad629682021fa6722b5ee357994f27b77a4910c2c9e7be0064a25ab760cd2e003feb6876a187867ed21dc94a1b2c45719396fa968cc309aabb8c2bff3147c09c8a7069b90d913738f9f9715df8e7aafba58422d5ac8e3ee2a860cd340b2860eb26fb75dfcfe659d91cfee3318748829d37d299e12a6d2fbf6bf2d4064f1ac0cc2c6754d55ea892f14886ef65e42623db081281ac161ee7e4ef8c3b594a348714a7f09929970f5345be667750303a0ff43b081237afe2048e2294c284a9759066c34251a0f2ecf6b9836a092996ab06425fa6f1f90620d1d9afa617e28e62fb862d9a209621062936f9f4997963e86ec174674d58df305b6e3057b8bb9ddaa059787f4185a34bf1fe937f8463d669a9e17caeadb6ecf3f02f92b4c87d04904e26e1379295cb83915b8314cabbdac0b4668e556d3a9cb6630357b3dda18e3be05a0360297ecbfc04cb63056ebdd3a47e21c84b80f2117642af333207816219c0ef0c25056f5588cd5f1f39a9ae305038c5919fb748e0f50645e70726015c75e022b846828e68f04afa7d4d2cf32032bebb51456b32bea7c9ecec8d19637fc523ed83243afb3a66cdda54c224d89223aa779822633e2bdfeee46af1c5276dba8c14e15b3f50c34d3e8ea667ddd8062381b2269c9c523784202646f4dee614545baf16783a61163028d4364d0fcf70596a1a6f38852513fd4892bf78ba42f6e09768f630d90ab12f4a0aa104dfe1ae64a3d9fd81353ac382aac0af5665fc92bfb0f651babcbc2630b32284598e58496a7844831f19de18806c851d69467b99e168e3785aa27c07da25f214489fc3f46b536cb7fcad4ce5b34272e826fa85404b7335e070fc52345c38976e88641bb582e858ac8ac5fae90d75bce07b2d14ad4ce04b913aebfdaed3dfe9cce526521d0523e89e20dd3b806eb7236feccfc6ce70a040c3eb0d1cf8eeca96d38522d1d2e9a3e4201762cbe5bf7812aa5b2aa30f7af16b77d70d812ced9de2fae645155823f4b840b9c440731927e4c555eb57dfe890de15850e51d75e226864b01c079b0640a8b59aa6862a41da7d7b30a244622f82c5cb24f7c163208c3d4067fefe7b708084e0f8c9d56cfd58d2e20abfa2eb472b19284afbe2e2c828c59685d3d71c94edf2bfc950d78fc4b9b418923ad88720aada30e5c311f5b6d584b7b5a28056426aab9e2c292e49ceaf5e97c8076485cb434b89ab33adce9e80d45525f93ddc72fdc653a6a4493c2f99522d8cfb27d93bd7ed780df03be941918329d0417c5c5bc96ee188c861e5f72e1458e0ee240334ae3208e00740fdecb17ed2d422cf42f9229eff1fd94a335e5423c51090e289889e9916b53db7243990a708cf0cc8342fa78cc99c80329e304a2e5fc2181aee44f208ffa517c9352d6db01bc08a20f4a41a726f72d2007f87ca46da5959e04947d962164219877df849b80662f2d12fe210390994583ac7622355b7c600ff9855fbd9fef7365df60fa7451c0b15b72996076ca5dad29ecaf78a2ee7ae102e20ff3c21a5173fec8575a65bd4abf556036383cb5b78ac5b34bd9d4c4d6c55684ecf2867246fa0ff3fa829a4d37375b772c43dd77c28666cd68ac766a2e13f19808044fc9b1350dead96db61033ba068012e596421b6281179682998202989f13457dedc9a0b95cf8c8528585d99dfb4f761c821429e741dc1c1f1579a85fadd5b39368e269f6b23c80cced388a89867aaed124630cd1eeacac91349f2cb68bf5eebf2d5f30a7f5476908ee3592551d53a06f9efded26b8ab1f3c82d4ad9bfb7e8e4aab2bd2e855e097a4c69c4c0dd09e847c1c80eabef57cec2633a9809b52fa4fe762a5960f44ef8e0242013db06c3317f0518f325ab46904cafc2680ebd02933120cd108c47ee19e37256f7c9bbe593e3fb93c70ecd0721bd8a2456a7454f18aca97af87f076bc65e0ca3b1e40f98ed4b6596e0d7679d235c5e981e7238b33833406968a76f94353859c3b9b789f4b70096305ce06d8e4481fa0fad48848825b80ea316b202f8ab8f155f30cfd1e856c3fade14bbe77cc890a23b084d6ac883f356baceb0e0c56100bb81c9a16a15fbd565e7a826900472bdfef1cc15ff8504258178f70a55fc5aa82ec9b1aff06027b4cb1c9839b6e0c07c731933b777b5bcba17a32fb838d89621eabe19cbfd3f678183b0586b281607995e81b65e0e2efce2255d468edad8f9cc79cb8971cacd109707327ba7252f857cdeee3969952a66af77c5671d2be53b0c4dc610a879479c4f31df15e50f3f15a7dfcd1165ac1fcd3ea9e8ddfa192b215b74bdb3a11e30231b6f78c24b4bce6d0d7daa29963b7296c0093d05d3587a7d99b2e30ca48c12c19995fb369cacbcbdb4b8228c2adb2079f391fb738aacf3bc61cdfc4507b7ad1f29ee94f74f18e85351a9b4c5774aa4cad91378a3abbb76dbf1681a86bb8997b7ef8b1c803d2fbf12979422d3ed4f3aabdc3ec42048e4b7257577f3c53c2a53527394aea02303beadf776f7b6910c9455bab35523a59fa0f69b3c9c9217e8980191bc0565507518324da740ebe1f334fabdce161d1dd4718339152b66a2fb9efab2f341def866904c8dd39d5652c0cd1f520139c724129d91bc95f38ddfb6d6edf26f1d7c5caee1f2cf45f11c00bb225b4db9754d4fa16395556d1d207991cc6651dbf6f216b209a6ef732d8fbfe25c1be4a830006808c74f59e0c7aa0a6fe29098b68765bec9b3f4c1bb39ead1a762598ee0f1f65033125752afb2ec236241ae5cdbe18d493934d85a8b6a2873a7adea230ce6efb6dcbf5a0e964cd664faa863a76b551a6df6aad21c884490750f05d91026b45d96312a4c0e9d7b714a0b42748b4e361443dd05c5a6f36310d134e54a0a6724adf6f9b47e01f96ed72ee24a73e4323a7e08b835ff4d87fb66bf5ae8627ca1ee868cb7c2a4603b19eb0ea2dc91288e61b4bb58c10771be055d4ef1324de366ad96db10ae7fb27a269df1f042f8b1ffad268cf215f0dcea609e30ddec8d0b748df57570124dcf901fb5e36f690bec79d818952fc3ad75ef964b684851005c5fabcce9a17abf25f4fcb71d3300231254b70a068eb6e5346876750d9c6e3cbbf2c94bba8bd34bd3f880c941f822cb945d3667907fc38a71d1cf4a6546ee82830079a36de03b464e5cacbd97917da1ac1835e07305f82da44deda8bcf3893c884af036da20a247d27adf81ca44ac2f65e7b1447c2f3b506c5bb2238e4aaf3faa638fff102ff2c14aebf47e2c0a547dfd745a44a5722286a139f2f5c5da4259c6fa72c905c9961d795af32985e7d2049096bb16b14a7b01ad1dad4ab3426c8ef67a2cbd0883cc64178e2ca33870a4c227c74367b3dd13009f124450ff68eeaf08d93ca904f4d1c1d2c0698190e59fa1751e92d2b2d835a70f7680b9c31b325cce8a09c1b565dadca271274434af5e4871b374daaa347b595005a7daf1f0a3e7617e84458dc099bc486d7ca578caff79081803f74b5831cad7ea8707f68da8aa104f413b2851a70a5cf556f83335fc7ef216f1618f8be0fb305ceb8d8eaaf1288b6a6970321f28812fd3b818e2b99252505905e80bfc110cff0b5552b4c153103a0659ef34dd4d6c953c34ff47218157fa5b3613157d141eaa38962792c6941ef08bc8a5a2f583575e5f857fab3e98cdcbcc2d0aacc3cdb84926eb59e5f6ecc2255280b6daf02c1dc6f2f0774fc978332db3107f86a8f48cac0c4181370694c652f13f47f1612043aae94decc6d44f97b77c282f14237b2954331ba25e1f19e2567cc14e2d9217bc8fcc829964b66e7f300757df99961e70cce938ef549bad5fae9046c08c118000b86bae68db209074366db65dfdf99df93f7e08b69d0827716620b21ccba5926ac22d5f1a73de8f9ad2b41c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h1680beb9f3e9f72e8be9fb8d3ab0bc7b5c2e4a8ba14bc8244bfec4955f8c7ea4ac6a7f4e57ffbcde45d26183d3c984d14e108cccd6de85db85a132762d9908b07909ad4a7357a8b5faf7fe5ea99641906438c5ae05cbcfe6756ae7f404b4c0a06b90b529b4f973d75206d9a0d8d532517a85d2a7cf75d52c8a50490ef5467c51de4b1b44eb1a7799fd2cb8c151a44c3c0caf6d3660b89760a1824cbe986c1b6f72802046bfa49cfe2577ce02e0bba423033bea06e838fe49056e49df672aa70841bcbc836d3ba5383caa8a2a9b83d8af329e458edf8e28935d1b9fbd821f86d345fa82494c54e887cb45baab30ade3f75007ccbd87a74a26071e9d96c934d5e8ed33db8db82c1a41d779fa7e6f766b7c726c73d90c4b781dbf2aabe18900dde05fef148448ea2a0e32e190da8c3f85572fc9f345c5c87bf542a17509597a025f4036cfed2f637165af12a369accfcf55c7b60f05efc8ac9d02a7304c85383568166ccf4e155ee832dc9883dd09ba3a4436f4847a43c555eae3b771f4dfa771a30fd633d701145b31cda1bc8ee740f4f29f87d8d1c87fe9058abb6615ab001cd1772a36e3a6d2a91ad03674a41807517dfbd9be45509b1ed0975e5a0bf9e7e73f327bd0b76c8a9d01445518d0878afc2718d63780bddbf7e52ce4f3e6c56517c6455a8ec2b95a3647e3e2fd3985937e9dec4e1aa1ec86fa8ad3f5af77c90396f4bed5e51901a1366389668ba4a8a4e1e25dbd528b85beb2152b1abbd14f606e6a507fa0099de89215865c49766d0550e2a7d3415ca28fdfacdf40d52508bac75b530f32930a45933e6abcf6f015ee96e75e21620a5a03b4eb8e976472af3a5f28558e49ae7812f59b3c8ff93486983ba5aa9edc82a249363149400d2ba7c96081bdd6d9b6eaeabe6b29aae97bcfe4c9c780c4517fbfee5b1a9cdd13b7f8c765805d36b6334a7d450732503fbcdf23e31ca228577135161da391fcc2e8b363b923a474f4359e168bf4b7ddd29ec125ec541343988251f81cf9672413da2ee25cad6b523438d7e23d12c8df88fca22fdd7f2f381ccc20a998142d91cb70aa5e8bd8ae49a76213fa995de350a8aca14a3adeaed73d830caf4636c1a506340d094acf8a595a07a19870468ad342161f0cf5f69b6f6570658212d9655797ed5dd7fd937c9c9b89b47801638a1ddafa7c56acdc827bf0c3310ae2632e7f3ce1a72ec69455d60d6b5bcf45ac894d90b9f4395dc11d44c0c170c2237fda47e6efef101c8924813317f8c7b8683dfba72a7ddff238a1ca6acb975aba88ec4f16a912c18b3ae46b7186df0e30bc01ceb1c93cc3505abe2f5b643934899f88873b1b2731919be9cacdbe57b1b6fea2fc053604651d89cf29de3feff7723c57d86980ae14dce93ef7c047f5cb63cf61255e8738a0fc49c8e52eb06c3c5e814ee5eddc1803c987d9444358d2ef9869b6ecc254265912aee8ec6bec3eb92e26e91a677debfe1ce639cfbe71fff32ac06841c0167136903ea1c010c51682af5edbed45c960d0babfb42b58357e16fff61904c71c978aed66198c02abb832a5ed5f3daa375ae1c34e6a15c5e7bbe4c5086fbcc4e5e0881b72bd584d1a2c992a2f08bf711cad09f99bf5c2e24eaf3591c5c9bb53604e4a91bb4dc374c7cbb71f1df521720457bf6c0b55e750db5361ee94713bbd47276d9361e0fa3fabaad1af1b757d8a6e82cb0980cf63cfe33a3498fdbf713a713934b99ac22de49a574e98b03e39477871a39202eafdea7ba04f3f9ef5bfa3fea70fc3846489f2b571c2a77e20a74497d2b9e7e6befcae02f6a1f699ba49dea113417cee7075f1d513d68eb118900bbf8e69c06981744eb122958c089f2ee0282a8bec5c219f7ef0857d82b3ac25501daabd199b876f91ea98ecd5edf8997a210ddef1c1d9f4bb90944ef47e40489bb7c595fb401c5714920b6e0ba41fda06703e80afee1fe97a0e1e2d64bcd454a6c3781fb0b811d8a4efcf05fde0b87845f90f75600f526bb7517cce9fa134e4554cfd55f6a89f687c0a84b645611b6c2f7823f67ac6240037b0e94d8887af5d0fcc4190d811d361737368a74c10da54b50678da91748d44a14f084ddc799091db63e98568ea7715e74051ce010b6a26954a438c3a04a0251cae315d5239d74b6af73c4b274826d5b9b28605f6e913f7f2a40c3b5ea7478fa9a9ea0d327dd5a861fd55a02ebd66405074ce1e49d82812bc12fb29fa402df624b08a2045d23858d05dfb32f87e9bc55a432039aeebe6b4a577704d8e76659763aae78e8bc2abdc143cce477f9eee8da105a6148817140e618b73f86220da54da29252f64c97073dc411dbb4c8a93f3c277371711b2fab53e8c41c60c8743342382c0a284f144d5c8b5378ccc1256dd0c3c2a7a136b5f9e1c532aab3f8e1f91a039ec104c14d0ea1066e92004383ee59e5411218348d0c7c87b3a6bec7623ecb28959f37e6b214b3b86aa4bff1751fada6451d80593ade9051c2f27c8672a337fe95650b80c36287a93a65dfc289308fe5127ffcf4d995f163cc947d1c68f71e7818a7da7c7038cd8051db763852bf209e7c7709a971869268caa80d70bf8d1cead87707e9a0128cfc54e50ff14cab3a79da068aecb1df05a3c4e04e5ea4b4c2c2ce5cbc6a8b07c90155e0dee1809dff4b80dcc2047d7a5ff4d45f0ea0af32217eb08bc4088041834e04e6db935d4f2e140e43abe2c4482efa0012b5bf943b3f9d5133868ca2bb37c45462e4344584d239d99eebb964347e0fe27cde533d1a1120d69d9c8d4a05df09f75204000513ea96afc0e54c100a8b8e785e39aee058817dfe13103a1b7912dde94d161674f092a1d85782e6ff743f71ca3a0b92ce224e475a8be5e668dd7fcb0753a2fe554969028fd842759b4e66e25e5b26a5faaaf36ee78c4107a44b116b7229e9453613a1a31e664e9c63c5cc031342597bc2050052dba54269c74c6419a7bcae87cbc9f5aa195cdbdf70185dea7661967561674fe37ae766a949f542a0c7526bb3ca18f59808face57975b0adde02fbb7e2623698870b24207fca3608b74a4c0cefac143330c52b9b3705b3a6a7d3a558b560ff61b4ed9e5bdc7b8db52a8bf9bdd3da01ded14bef3685bd8d2f9ad10faab8d4ffbf59bc5e4aec6435116acae3d93a8006ecb05413c1b6d253bc2e6349dad22e3060350e86d134caa4924b3042cd2cdd97276c145487dc3bce0a9d96df6a273d598a224322a74660723f6f576b363e8e68535756c35695b7609c109a4bdf5513c4693565699b09f3991d5d5711f2d038b071487fb0a609c0fdd1912bc1939f4a018017b98bf23cda8fb451f4c96ef08336d043e483bd9663bf7af45453f16ef616fe36b5a57b8c701307098926b7ed4cfd2467a23e50f1548abe3d51646bc0c2995c744b77af59dbb4c8ecabdc15712bbe1fe10e4f1c98f658d596e46d1d9e02b66362da6023e4d5f1c3c47a3d64ca6533d56122b66e7c79d091456a6d700761d3ff7b728dba8a251e2cccc80fafbc433c8887500952c256c0a1798176eddb4588c924db2105632819c2fc0f4c2faf2e4c191c27de25ae7c71d42e9098b118326c235a965d4d0eded7d31812b1c39c6a9bdb9fadb4783ae1fd77ebdc83cb2a7936769161f5c3da89028cd5d83825d776df9ae559eb2c2478916ba7c38c36e1d52fea3a94d080b722ef3ee4895ea70a5da4a679234d4656fed13cfa61b288e589617752c67753cb6e8ac4d4993a35f6772ccb9cce4ec950170760bf8be312ecab1b30b7d943143f470196edaa548a459951e9a9ada4572a0cbeb741cac2339c492580ecebd0f6614d8fd84d1b47851f3ba08447a64b88f5cdff61a1307b9a46db884d131bfe934d8522640daf9e06375e02c9fb97fdb1dea7e15c313157e00a23173f0d06877dfde7beadbd4dc561fbe4c467f2a6bc5335028fe862ea95982eec3fee7744cba711a55a820e1501053d9802b0cabfe2eee5cfc9fa533819ed838c17e44065e83f2b699d3c0908a4d10da5a8d68ef4873059a7f933447254a28b10752f512ed6447717d2f3151ad5ed9e99abf312785fd4c1df6d8fa9b00a56846a3183605fb8e6d11dc8750497228ef4fb236bba69d07eed4e7c23cebf8c287f1c5b3119303f1e9af029c7097db059d30105be4f7dcc65b19590e9a4471015f7e109beeb3d354c0dda96e1970279c6b8c4829b6b17a9ba0663152b9b473b8655ff39ac38a03aa8582c3146aa4e9858497d91f4e4ae09f1ce4978ec3107aee3ca7c4447d702c37187f4cc0490ac9b0e7cf40f71bd09b30706e0985f564d3b0b759d0a8519b850ec9f608a77ee7f895fc61f9211863ca5b9508844a0a781178444a195102b8edbcefbf0896b683f2ec91e2b278cb97d09b6b083f088b0d761722641fa8e25d4ae551ef9b009aa43a52c3d4097118187b19db3168612e029f1e7d8c3e8cb71294ccc6ca1fab323810a1b2b9af607174b01abb66a6814a4cc9988b4f082b488656f882dca99e2766ffa4ce52fae7f84affef9ee3d767b634e2209a0a33bad8c042634996b6464e320a1f95f94acdc1589de267712b725ec93a71cb7f4e78240c42c095f830e6b0cc1ba7171cb52e49ec5505916ea73a4842a31e602c9f219501e31934ee04566f14fd7da0d4beb94813d77f12ac1557506d67495aaad782c642057c0f7e038bdd7092fef5dd8b391b33234254a5f40edf9b868fdaaa04ed3e471a44ade5a532d6700b307cde6924f51063c4dea5e34ea21065beddb8ffd30478178c5c678d812fb8b2a5299e33cbcc7c73463d5c71e739537b9f3de0795f8ee59ab6a881b394077e7d68309193e6811e5451c28ea577ade1821dd57536b310fc9e2053c3f45167ec21e10c9a2637ac358ed611ca84df12737e52cb7d19c23e927999671a65a9a06a336c954dfb846539afac7ed7af792325440b94d2edfdad28d5c12d963a0f967daa4d1dd2f72eb8b6c901460bd60e5fbdd7f4afd785957092c4c3b2d43658e3449b50a7ba6189634e5208881104cd6e5a3789a2492e2508fb2618e6b5ff261f1c7098511aa570d0923bc2e1d0ece4b5d34d3f411f65963ea2b8045e0640e1df673db40a96b8f9e6be1f7ad7ac34bd8f8a3e18925d7dc1e6d2e7f359a264f6b98ec9ec92eebddbfec0b0a1d48d7f18c190cee55ae77b049f2dcfaf90b8da18c6d9e530a3b1d87188b15bf57ee4cd30e1667cf60c5d0c61ef165435429500e6879512b7a9c1dfa06ca774a141b59580b59d766b19018f77fbcc2982ffc75f9db5c3c833b03be75039329d1d13a0b08382b6bc6f9b57c43e266e408d497bf45a6c4f71787077174a03a5a54dc96ce5be7f9c9e8b6317e0e4aa9074e339842e7dc2cfaa22e14e9f90f7a4ecd4f83bf85ebd386dae90e6de97f52115bf99b0a549c1b940b13f2be37f4531a79b9bab443baabf31f97f79244a5cb08831b6a126d530dcac6191ea6b5babb2b2e0d497f8acb8ba74085f0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h598ed69cdec8e290cabc6889844509795d770f2aa251db2026637c0da0ebe48156c48469545dafc0bb138ad795547b7c8b5798a4c49369770cac8a3fe63d627a34a32630d699847288bbb98547fdf2871f11e1e8152064e60047cda006b972f3ff2b974da906bb49623a13e1f4a37a34fb44b8be2cc8ff96b0cde347d7e6729b441fe9eece76e30d2b46b6f63ad3b77495f3a8d57b92d6712622d741236f0f73af71b1c314d56877ab88305339dec922781a80b0298e7f07849d168da30ad1b8e1571f6c8e5e1f1c8506557bff2f8804a85ea7e0a884308e91df59e2f4ece47b8ffb7591ce54b5a6c86616b1e9954c12d0c074f1f075d05850b3d45408ca6cc87c571a80afcd77eaa8136814cca49690e044304b022e148bf8f58461fd231898ab0194db42c15ea99eeca7fd5eebcf8a2ea6f06fb7b8000be7dbe6f8fad45497d7cde83c32c1d13f36f8355e9f74ff8e507cccc4b36ab8ad387c51c36551ddd8782cfa00a3172afea0acd452667673ce5a17540472943404aa8b66d1e9e20252c26793d88f6f7988133aa1ee6f08ebd1656c64a354ee7301868ebd6aa51af42c08ba2bb5eebc5580aa8c61273121c3a6b9f8565ae718c4960f882fdf3e616b41bb9c929baf5d7f84bd922a4a0cc31b1a3a6371045462425b5ff525dad456fb665cb008eb295348426d115e294ca5bcbd45c9687c96f920eb57dfbfd7c88190e74d2a227017d6ddeb0613dee99b67e7af7cfd13a064a230088263ae5836100790ad3fe824ceb1f8a9f85849489bc0ba5224f51a207231433fa78623843cc1d0e4b99312b5b61297f8194bab39c55b6542b32796affdada6543c3db76ad22a577c677b5150010a50bc815e60b554db99d71885cf2428a55718d96e5f660e61190267adf0d03e136364879f77bb3c5387802ac9fd0dfa0351034f03377266db061adca481b6a2513dafd18391d7f837662852296d476347ac5ad5c86f155649e908597d879a15ad8a909706e48b01e8054a51c0fe8b259cc84dd2b56b49dcb566840b34e6ad7ab9601341c79b77d7fd8142e0f0850e4e6c27e1c0b178f1df252ede9698611abea7edfa39ca8f597a6bc7959b806fead1520a1c163eabaca80b100f2e1942cb8a77f4a22aaa83e5537690ed840517ced56e5639f158809cfb41437535427db0d06e592a1e96e9de626c546ca452cba5bfa13bc2af3fed6783c792223d6a33af6036664421dae40b35a31eb7b424cf5c28632a9f7e313bc271ab1bae674b74ae894ce5823b90e80f2518d22ced97750e6d2cdcfbd28847d355eac8687bfc2d083321eba99b44ecc9b67b845befccd5fe9676377ec504ad91b24801e9eb34f7d825cf29caa3ccc65be1d43974e22bd28b53a4b21cd93feb3f6d43b20641d9fbb22ac67621cc57d219d336e9d64a5d60c92b06416e3b8757f21c1168d573373450c84cb10f9321ac2dc5601806cb8fcb48c3591082a61af206a3afa218319eeae4d4841f79b781ca768810ba4a30731c6ffcac1d1ed35b47a92d4a2e19fb12839568ad8e19fae42ed5c10308532f8a3c846270a6b8399043a6bddebbfce2c6bbdae4467fe79aa5cee230a51ad1e0cc400fd2be29fa591c9fd0b68ae8b6775ada1124a2cfec20767335664375fe376f47577d0d048508e223df1536d1b80e91dd0cc1bf4db4ec5bc434d6e61870abe3a2ea95fc34e897bf7793548742e23f3133b019fc86c1d5658ec019e174005a45aef1e41ae31c39e18148cb106bb3f1dae9252fa7445fa35e45d74036725172d224969e824b8de170d2e666b53f2c0445f30c91fe569a75e0573b574f96d2ddbf50f92505c6322b80af18f601f9038765f0fa3de11e29b8a74035cc828a8355f3f72aa90b9489f9739a9cdf8ae273557df83e57fa466f9b86941f78b8230ad46bc27c51c6a57831ce2de1345b489d3e61ef79f2ec866312a6372ed9a418036a9b5a308efbd90091d15d98ef97870e79e4d7639cc25b9098081f17f76e9fc5f89dfd7f0938a34fdb5f9f7b698b918749ddaa6dcab8e500598189dee30e653cc7b38e3317f3d71c43f4495e2dfa2bae3d2d6905f7ab7b830ee2cf439a99de08912364c68ed2a28f25b661559452121dcbbb422d1909ac8db25624f07dd0fb14a7d5c20cd0f74025ccba61dcbf7a83605a3ad82eb87f296779e8d1e5794c81a4598066b6f673f982d6731370ac4456bd21dce421e9a33f086314211e47e3f8b8a5e3b730f56c6ed9dc509cea470f50ef20ac00cefdcdab4fd4243f3984a69599a9d605f00dfc4c8e095b691fbbb199c0e0658d47059ee11b819c6266154c139bbc4d0464f5fe44d3d5f1e1546c62b9f0f1d40b56dc1213d67cd0ff86b9dcdb3faab228e0b774caec57cf62006ca496a09d25c1e78adba599606dbf3cf333498f85fcfe01c9ef5c6c356f8b74ab87e08228c0e91862d2b06b366715824e0390149fb133bd49810ee40a5c8cc3d3345863ea612c525ba5f0b76a0ff234115d0343f2f7fa6493f664613457a6e684b0b63168c32ef695c93337c8cf8a4364aea309ac5f97c350aab61923c0469d5ead8259d5efcb63b6fbcdcce5fbe5278296999d2d852429db55937b35c51ce0c22296844a62bc63cf49816b9e752735bd2a77d9bfac33386460c171b7258ed01f5b33f0dd6ffac3881910484d8a222e3a42729fe6c7804d741a2f42c6da7a42019808117db9e1f38c68002b6345a45e510a06dd40f8b66d0c8062fa955517d83ebfd58bcda07459838609b9325a83de809190e8eb3558e8d0ef8d829aadcd67d7f238b4055497c1fa5872c38d987c771b6f4deeb07092becad0a61e6215af1396ac62e96eecd4b2068b7fd306e40330880d93bf215bf0182e690a61292626782c570ba994ae0d4a0a969255a2f10dd31a3d0c61b51e35eb0a761a519d7ea43b61051781ca44673a08a248c6c7a1b53833b15bd74643a5a8f789a326eab06a613b145e07ca4c59222c922b8b35bce627dee2fbe10baa352cd1de0f200458056dc79b4e4ec26297be46bde7f1ccfe788ce32fab72a180fcd8d568fcfa22799f17a303fd1c66cc5c5ec12ab072ed1dd62b5f410ef07bb831d13ea34aabb6bc7f6780e6899e662784ef6ad050d2d7817d1cceb0ffa406c77faa81ac124af5d35f86c87d7b72f1330e302a1ef48a64e85fa6222b20187cec0f8dca5caa1c8f5fa4d5f573ea4f278a734f7ebe53b1a071e6f94c576bb3e95377c02bde6bf8120ac13f7075d436bdc1b4a94151b6c9387872d5a7625f1ddafd676e2ec9c1f9c9a5a8d5e0927631d3d0ee62ae67e180a99b1b27f33e26008025c5967ad85d38c26a3deecc688680003165943ba3497002074f0e66fdae11d2051516c7a31c6e868afe35209113d253582b196dd6062b7bfdb2bdb99dc12f6d3e004b9295d8590a94ba9b99bb56dd10c61ec49cbe110fd0a0a4e04a203af52d8fafde6108da70f35f8e7c1665a7a480f938cbb6f95e098f6504f6aac3009f3ddfec6622c96968630b544be31b7dffb523d2dabac0e48ff44612a276af76e0757e3d4bfad5ebdc59d83830b0d2c58f8ddf33d00508ff30aa9ab5476c353f194b197a4ad77b4f84d2fce416c3e59e595753906d2ce34897891b3545e3eedc8ea5bd57bb0604a15169ea8ccba7025af86ed58f98d4df1725cd92847aacc542ccce80514076fd8efd215994589c9ad45bef5cd220000ea8f61245e3834b452576376e4376d3e9cc598644b87f25e5bfc8995f0e265428e402e9317818beba42c66fa93a80304dd3a21008a73d5b156182613466164d54fefbd6742b94150c4f3a40d5e33c9d77d10986dbabb3db2ea464229b7fb829bb6306369071f6ec01612b668bafb5819df68da43ed02a9d968f9389d01e5edb7e5773a7601877ff2fad95f8c46072d353b8daf5441d270dcdf6d7b18f2bf4ac563aa438b5523493e7fd7208ce38808f5a2cb647ed890c15480a2ff455fe594c1c4fe0b31b0292f262f4520d87c23a9f1f0e814d73c8443b14b2787a76f3af604d683aa22623c9d9c79de3b85840fc0cdcec9ae01f56470a70029db1b37574047b652a10cac4657482f744fe08ab2235878e510559153bb2da57d5b557cc2653f5356315daf92ac841587a390a9f20662b2d40bf49209c82157a351a9df1cd8f4fe89da376e3ad6382ffce8cd68d62fcbd55507b95150d36732454ef80be61703330aa0c56b4f6d28ebd7a34e15ea6c36f1d5afd41da75e02e5d506ac46e3d09d9f5bd650e12f72f401cb66e4660f60f0fb80c2739881b49c0dcca497e21eb3d9a9d09de5a5f870d154e4d8c84295aa312b8dc3cd882e92d681bb7b8f64a4ba0b1431e501527cf26c69b7ca411027d9776aa086bbdbdda7bdace3997bab3727b788d2ac6e27d8de914ca33701849370d961e6ebe606700444d5719db703c31fedb59b3f8791a6fe73edd7b126f52318ed5d1026d9fc79aae54cfaa62509e61947b78745c86c80590fc347c33fd1ea2b0d16b82da06124758b5ced450892ede109841c2fc79797e6893911810969c4c538890c169f9f6bce66a17d952451697b2ea00fd081fb1bfccc9b5149d0b9b62771b2d4afc1bed4ca0e9bb5366e50206b0b1990b93d6e21e63df9270425a20c8b051151f23871834273e7b525a71a68c6be38cc9a45bd53b219a3a2d7eb4362adfc08edadf264634c5f3a715ae79dacc9026d9e45b04d394a707aeffe3c0ddb18af1f2c245d0c53de9694f0a70a3fd89ce1a685791c57c29dd409541f984d762acf9a7ba88ededd239d1fac8bd313b55146c542af4d0f729f8e99089244db1509082e235a0ace1bd7dac22e655c52c23e4e337c6bf4d0ffa310c1dc00aa6018a7562a80b7a2b753f596bbf56885b5350390b41d3acdf77078d673c17d29d68ef0b37e6b1df6a7e7c4dfd77e991eca531e720b44b36e428f5ecd105f43b4956b6570ba095eb00a56f5408638756c2942ef9ed570538f86a1969ce566d7ca153f11f153af40d97508116c4622f3a09046b37061a1ef9185bc3b12fceafeb457293e42c6d5f742dd0acd79fb9ae7a3db83d8d988b784c5e6e8fce3cf3c7e5631190c4946543cd731d584d6425f75b03d331030e00b02caa37396ca1093bbcf316c67861ac4442092b743bb05e2c91d693b61e6020505611c19084cce3ab0bed14326edb2736f8be3f655d3474f92e6bfb5c74715fc3e8d8c03ef8583c2482b595f2e2f88e185e3a060ab8b00c7532d51a45638eb0ede963364dd5e572e9f03f9d64c586a9bd73dcf97fe1f05f29aef674b288fea8edf39ce55eedd91a8a9aecb5baaf867ce5b99dd03c5e521b7ca7c6484531825261782bf4197dd051847684280a6f2c3de404cbe24de320a91ff7c1ca772f9e0a9d8dd427c470e3f14e9d406e2d97a1bae02ceec7b3e92bc2ac93be01a1c75494bef7bd6b2228c0bb5b2e893cead09867bfad0b579e1deff4f520e0cdb38afc0faf1448e2af15512d2e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'he8f2ae2976fabb31aaf2df9276be65ea847cf9f13466451e9e9513d8b08af569f25ce4b91595d9d06a430ceb122b3de852cc88fc8ddead6932c138817f085ece020f780c0444fb0a1e79641cc47c12fa5e1a14e1727662e4ba3357ce650fa4c6252e829628acf36bdade3c229bf5f99fc75398c9541a7fa44c4aee42fc8ccf7b52964c25949b56f7c306345c3dd47530749895ca214f9537c97d9847f7c5149fe08e08e09aacac71007537ae980413f78b19590228d0765a0729031de5ba3cf0b6b03b7ecc108eafe0488a0cabf25c92ebc0989a4919e1091074d56ae881ce3ec17a82d1dbecedfd6d6c38fca09a525315cce2b4acae473bbc709f204e7d4dc74c15eb34a8f6d795b4ac99c4c4171864cad7f1c8f2cbaa494a67132c622f7c78be9ac710cfd672686caeb05f1e138579e9e4e6e57e652122d65e54c17fc6b9bf7b7b6facbe1dbe578b381a663c3ea63da4116f32464572c0522838b228b6812feb70367a52a0c1d55663266cc236593c2cd86ef61bc7f3dc0e03beeaa906fe8c6d1fbf755fc3030f7e6de1124dd0237c3adb45b0484530dd43a8be7e72f8190d285d62906a2633936636309a60016f056b101d9a46829f2e073d22db14d461310ac4fe6a034dacc0f5579595a37e42cb3f42aa1771679467e33989c7bc91ee19f2a2e65756e57d8880090a6471813a035b3c2bd1028398e342ac0ca2869749db7735a607efbdb4f6e966976ab3c78ef5599b6285d0741c5e5c7f8fce78d067a4d8f9917e88f193fe4b45ea4efca302f912a3c6630ad8b8eb17445f87a93130b37033a53314515e11546819579a6cd1cf93e5dae237591c74db1b302acc42ee2795e8701fdc69272bde860388da0ef7affdf20dd49d7147adca60fae8481a66e257afd3deb4bfa2a84b066c562edfde724cb5f797b8941e7c10965b06a683db7a69d71c538fd067f527e968eda15a43530d84a5549a82c7d04cee24e05c1146eea351dcad1ff8a6a74e12b3fad6f5ff1adfe02acf79aeb9e4a1aa0be234d9f3f5468fb571ab1c4916732babc3f61b6107cae0bc1c4260c54caedb9b518997721ad83fee757b23d76caba22c6a7e8022ba0864ef8a045da8fab92fefbfd7ee34e78528c89cedccee85cbf2af2b11df035e7a23b6a1f402503a36d82cedc1db8b2d737148014c1f434d97fbe053ec1bc95b25ee3c788678e34a413822f0cb5269f55f19f7f1deb9a92856fec96ec9c969d5c5b834423b44d8c49fb1e68eb55a3a92ca86fb8962001f9cdce446f2fc8a25802894b6f634abee357b25d112c7114b80cea3ca73d678e26072a38b5dbc09ca77103c62b015a19f63538e189dc6b692945f7898eeef8e2f7267107044c21ee428504f59b26495c84839f8e35915f0b6a666ee85feaa5d2752944dc5b6af1739b41a641dbf09469412d9704614c64982a337e4afcae77cde3c0ff191619d6d026c0d50e705e88058b50d0349be078dc5e9f997c8e0d79e7cc970bb2747fe56e4612d643f39b6b2fee1d8c3cdc2e6988fdca4a0a4d33bec4252df3d3f7d31c87eb8bfd7852594a312867903bfd0d6a85ce94bcbd60172e92c588bf3c6c4f8737f9839bd81a8e315d927448754b1b47100dbeb7397ffac45f1eebcb2f88a24dcd0ac2c896432869f335a34fa159ffdbccdadee2cd258f90502254ba0c2056a3893b8dc1782f6e89b43b7951d6e44a418636947010211bcf72220a5e7cbc2c609515b90d7c599259857722c53c3b4b8f6d04d375d9c1831412446d6eba103c122337f08cf837bd566ef31a8b61627982322f4df0786fa8a19041f356098c57bc4b8f4465d1382a073e0c0bede5a9bce24300981d312475e040585c8c5d98d6c2e5d095a10368439541a83fe4aacc31ed68e00400b980a8510b1824ef2619e1dcc3b821edcd1f4edaabc7ac04a43d5b973f47848046700423c22f145581ec834338d462b2f67bcf038097b5bfd14ca9d2feddd459db7ac6c32a61ab032e44c1d00f293b5c31dd24dc6fdd0446d098b5635217425dc00399f560f63d9ce7d422ebef6774a91469047ffd5ac1bcc0b2593129257be17059b3d7522fbeb5a550fed1795670ad3f8b33c8f5feb9923ff804c24be26b607d62caf2d8c78bc4d9f52e39b9eb3271af36f53fa4445ac3f521fc687b41730eecacaafddeefd498994fc010ed7ab7fb896b0a2e4827e4fbe3c8fa358d23d0a96b972cecd19f9368297895e0af09247cd02a205a8c95cef86788a952a9cd1f0c6ba75b0d1c14b874f2ee7a507d023ebbc3d627a21269f201eb1d37ba1fedae313ec343f49e098fa797ca165df95317eb7e3a9efea701c1197d32f71fc89a37d5055ba02c3f95339743d868b88d7ceb0d6e6a45662bc8b553d1c94fdfe501c9911b24ef6da9d2725a25146672d92714896c584eb67eec0695d43235e8f57d87eb9ad25e9a9bf52d67250f8276b6d20799bbc6b2f5d034ef0821b88af69bac12d976a71dfb85c3109c869636d3c1deecddce9a8da1c0d6d0817493029fc6b64031131f055b19b35f2c261aecbf54a7d5ba3af1f5dac65e337e8026760d31c8f4454fff80ff2e5c8f8200432ed87d83614369a295fe231bc751adb401ed17e6f5943e6f91820dcf59b6260e4bc033ee3d4801c13ad701f5bc43e0b1eb77a7aa5786bcedf1a90285795ed617b71b8cabcef7a4b7c043d40ceab9792d4f77cdbb4288ab730afe3e4467e545a4013e5d5914ceeb42aea3318bbf1a837f11ff7d6ffa52e89538de1d4d9e248be983f475efa3c8082a6e433c712d1ea393247cc3a35f1b8d10901a5cbbd46e3825b9e39a96c279b53a8f4893bdb1d3d1713fc3d91a5968137548f159394ae07ab5198300b3fafb5f45039b2b31a276fd83af5851e46c47207ae2dacd60cabc0dab2d7a56b35db935c699960f564abda7bdbdb330ba723d69b7edd5a01c33a451a2ff9f6185fc6567bcadeb188f0f268a0b33af00efd03704a9367ca60b37f416e8ff5be47a517d12f910b6f8f1975d6c6afd814c8015e5f8b13735bed24810664844f744b0b0441c10ef9dbca3a7aba27e45cb3f07b46d8702e35ee4bb8ab7d5980e2f939ebad989bee024c6dbecdadf665f87f06ecef55cc73d8e8a063da8c8d505698da9f7a83daab1c48cc2c78e3132cafd8aa3bee8e6771b0c9e230727ed586b4e55c436ea97370a4b9091db2beb656afff26e9137a062b004c995ab666891c19ecaa6e19ed84e4aeffb9da173097d9b86baa0074c5151f962803ec7bdc6118b1fceff880d68702a46d33ec8455f34424bd569aaf077deb13585fb1c778a3c8e8676c1a85cf9427866ec47b90834a49c503d107e2c97b184aec30a68a1ea32a151e7262c7ebf29e3192a53c2eecdbf81089292fba39e8cb79090d362e1c8926878d268994b6921cd19ba753a22b73a28836c40ee7f3de9a5424b74edc9ff20106e0cd78d9aa6cce21fed458474cba2f111c0d233107b28d5418ec04814c3eecc3dd14afb1f8625dff92483b24a2fb2207672fb72e37042647d1ef8541aa86c4e042b4d60000d8abb539e94862183f7beee7f99d15da1871f98156809e95360f1d820b8c82f56bf2fdaedeaa74fba735a5575194f88a88c442371e5390b8183885ce1a1a2b5df6af9d7acdd15667ecca49c8eab8c6e397f57a80961fa5315d18167819474d3d936d6dae1d8ce3fddf6629e7a185ca74fe8ed3839362df406d27869b39f89540931315b5f1015989d27fda1353ea380caae5a1f51b81a8dbb63e1fae45842a01f8aaf177b933fea16ee32698d9963154d9222ad3b155ffe96a87165d3ac55f2ba320ca9be00df5015c9e085a0c92d536ddcf5f7352d75b9e08acc23ba48e4b3923a820c89eb4ad81c29c934bae9557f3880de4f6040ab4ea8eba7e6847e48011954752875d1067356bf1eb2479481f5ee6993febcb30ff0356bd8e2f7d6d59454517335f7cd315219e30cbcd59b6e5b8a1961d8f1189660f2b358b5a73c89be83a54e62f7845ee875cc452701a3fcbfd4886ed6770e0ec8aabd5c8dac8cfaad6b0993d4028a51edcd517c52486a66ec1bff64898af8c4248bada09bc11e22ea251d749da98c436915a3b8d427f5ac9c5595680201a8a15b39dc44af0077965e3f567dacee0040bfd6fa085f8e83984f5e60f789e91065d5d14639a23d9dc263d4870066e97e7df558993bab2aa4750253f173cf4a29a793967f17f1f78d7dea3a12a10d3dd0ae37542a1bda22adba7076d3620021da59992a05f9052bea18b5b8a5e5ce194f6749c59653fc22241e7a70005cd4c82cbb88bae3f98fdf59cbdeaaf6e251616a53657a64b6c80ac1a1c802437caede9234d11b5ee8625d473e9e406f5ad93b25b4a8fd95c5520a03b337c22fc57de4ed3f34f74ab60816c9d76ec3229c36050adb909b0b6b69e571d33713b7d6b3681fff523e902ae1ec6a4814bbd4ee5e959bb84e0835f632e8b358799bc550b84923194317c42e806af5dd2eccad38b98543ccd4137ffe581dbc40c1afdbd97bbfcbd977430ba35c015e8c3842d1ff92606decb79b3260880c389b683430a8dced23fec30040844833c424b3b163b76208f01aa012e5a0718096a528dc0dad5c218c0e28e10212165fd38238973befafd7ee7d72dd63de336941501d1b448232451d40f7b0577c07bb2ba0af38c5ffcb2f7785989119df996fdaa364c490ef3eef50122b7d24730903f079a48c2014b672208b7047da1a0da1409e35269e7509802c2f619ed30b77e5630955f4a94599a3310623e57ba7b7cb61dc5ed272cc1f59669c71ea0b90bb31abd03b8e98b63a743a5569b8cc89ee3f932678252d5e3236aaaf263eaec0c393ed5d6a6426c026ccd0fdd4d7cd852961910a57af01a8b469a5e433b7733b634c2b87d47d7938e7617a756f6431a8f3ea560f2b8256082d102fd07d676660e6e53122b788dfd9101a9acaf0f268a18ac3b1c36c11d47925c8cd0181590cff3a885cd1fd18b6f5ed8d51b6e8a9f23cc3cb5c11a9244e7ca974bca2b867c0b8256bd58338939a5a7ae6b26c9b903ce1cfe980d2c2845c4b6e2fa2e1d3f33f184de5342adc95854d2ec563953add4cdc0d72334715319ea782b8585624ebacb56b2cffe798be04346c553de2a50d30cceb4cc40f8df2cd3a0aebb9eff0f9c2e34ba52d8e0c148dc5d747b35066cd670238685108c1c7471a7d6c797cb3a8371395eb4a107b8bcd373dc3a730b9244842d772178f874086c11e8238837aa9b7e6c39efccb09f390721c54bc667b63e151f786fff6ccaa031dcc087da899caf9d6f024c7f7d5d98b70cabdcab7bedb1aecc345ac23c60d129bc8e0dd1aedb05b329669d9527c16e96227a5ce67ce39cdeb0bddcba1585227f6d38d8cb013fe7f1638a71ea83a4b060e39051c3b1fb66357aef9e5f684ff2aa071634e75c8d53b2bfd748de57257f82e16367c585799e0fbd818d4826430952cdc57306942fb9a6e69261ec;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h55072c549511e1061b793ed63becd9100be301e49d65e3fd5d28269893f86204afd5ea3a354a6c9e9447b9deffb3c3648b0e43b7998d0b554d5014884bfcddc965b055944bfbe2fa350043efd94a1fe5b9aeb78f1a2861062eae97708bbe7be3fb6d1742deb26fb15b10d15c260dca7b860a6a8a667c744e21502dcc0e67d709fab4a494aa6d2d3aa6b3791adf6dff993c32b36ac364267306b1bfe532a815541a542568458f8d67e1caa07b53826498ee299588428ee5a58426ffb863cda79be8cca5146506c07b1d89273ae6dd883b0518ad3768be02c1dd3e065a7e157888d3f999fe4efe34c4c9ae76892b8ec9ac000e6aea61039e522b1d6e87b447957ddb2ffd4b8564d9c16a800de34ff94b9ee31ac510631bedce7c8be5fe2f19a2d0f337085432bf7da142440c0b54a70a1fbb3008bc7cdb50e2c119181cd85049c922ca5a1c28ffc0eeea98cd17f16e539d1d415bc848ba19ddd7ccb55f01ebb7f04f3cbfa82b3027c39382a7170179c2af3ba28a8f09fdb7c0cb757e09d8fa7814c776783eab5d4b239fe4656a4ab0e81a09cf57496052115bb1f364cb7638906691c217015e180396d2f8b1e6aa4a1abc0bba39b7ba44675c6d535f0ad8f79cc379e3f2c291e709cdcad4fe5d4ab0f7c83879cd3a8cad4badfc862de0fd329cae0ebb4cf6a00dba93496796b3dd60a01d34d7d99dd9a460c97c7f899a8f63952e24508cd8f69d41ff38b103a01a700a80e2874b576ee17c28539346db756eb7bd1f0e824be89c776faecf263c21078946144a6356d58d35f9e2c121df2c71ec7828e4a7edf52c5e78ec908a44433c9dc39d1666582fdff79b64bf4c5087537ed50e6aa05c6a52c724c35561da3df4a25ee9854b9fb71d691576735f4d08e433d154474c8c1245294ad95e32a4ee0da55ac79626b8fc3be4da1f6853e388cd95272dc43d7485311978fd68b5648119fd44cc98c02ddcc126ae1d661f58a432345c786dde49ee82441a6f8c5b5ae56f8319a0fc3e54b3d663140888d6044c3db71f193842251e539bf1cc709df1919adaf6e3104d6698bfb78b45eb1b3c8123b591b242856449eeb60721c86de2a012e2142e7ad2e2074a80b3d67597c86316ff7900177aa05152374c3b2a19a417dedc0103638a8d0bd93c10ffd16073e08cd0864417b474611e498404fc4df7c7eaf62d5ecff3287a9f1a668b04a5aadb5b3d6496d71e19b97fbb5ddce5a23a473cc28ba530ffb9fbaa1864d53d9c18af43782016733f884995f5e286afe81c3b905d0f693a19fafef2ac5ae7aaf9700045df7429002c739524a2b1f3c3299cfc2863325cc813642e1e0df5111536b6f51c722096437fc0d337733947672343056a09e50cbf3c1cb40c5a7b4818dd1a84150e1ec4ca6c7f6f811c4defa53a86cd0dfc58e97397ec0aa4390fcea0cf3e5758b39827b383e192af009ea4447c2f21570e5b3cdc2d4013824c94c3912e003da325460dac3e56d2fccb99e3d7c0d22a06ec8c8838a8d5c8c910e2a359eca30bba4e94040d9e8f6f5e383c261e424bdf85933daffe6ab195d6fbd262615b724f060d972d701f9371197957a5a5b354bd757709ea9a491a28a2a4842d10001e85efc74e91278e0a4b19af512692c07920e46ec92fe9b2cf1b5463f22309a5dcbe5b02eecce80460f00b0c9f05628c7e509c103e4ea738f192bd7d90fecd78c068c38989f6962b429694470cd754a71ecc198e44ef8778f174678dc5914e6694c3246d01a1853becf3270fa90a0d760542622b3aaa3a7923f632bb761336a9e9a37e7c6f1d5c3a21b158a6fee253b2171053b72cb7bbb005d8aa6ace1b597992715a91bbe7137b397dbdb9569f2233f17aab1978b17910d2f58d3a9bc8bdc845244ea6dc66e1a5a398cdde72b41a028452e4d9d7720f4a7af93f00c33d9cf857dd2cae929687f6f5b2e97d5f43797a543a547ace75a6e54374f122fc9bc40d43df300e433bc520581afaaafbdd57ba68e8bb98bab98b61c0ca629284b03bc546cb20fb48272eb5d38684cda3072eb9124b54ef005e933f1b11084b5a959abc034124a7ddb27749942e54bc3fb7c0bbb8e2b0685c397f81368e082462e34255f6e46a6627d7b6c7702f537dcfd4316a88128a8a550951edeac1e3f9fcfa446a3a3cdfb00e3bb80c2673a0cec86539ad1b8b335be45b1ffce49dd4348fb686489e1fff20497cca94b8424044b4e40158b3640c0b824ee1a86e4f19bf3f169a52da407a6fb3d81bfeb3e89e1bf77534c7e5df4e5f5058c528b71d03a9fbb894af105dfd3f185a9254d8e360b46e724520399ee6f0b35fb0dcb46fd8ee266f7188397e693ad0017d36840552bab4d53c8ecf78da4f049d591392447f1e6e04999a8144a1b5b265f45c02d2c49c2417bfd2a1281d3047198b5efc782673d93739ac295c6271f5e7620a0f72ebf6d782ee846c652d4690519bc34109d2a40341e7c6d0d4f51611272032d19afdb7e8679ffbb31b89dcfd65f72565d1eb0f3557992e138a7f85b6e11c639f26277d867ffc53752f5e6150d5599ea79e9156fb6b6a31c5a9efae153907beb2d685d01a87b1f4ff0f90b7c0d638cb65019d2f6543539d236723cda722d451522e628e2538368de5fe8e8e5cd215b8087e80a11a25c8655c1f0058c9eb8f410ac81f4dd95d291c78dfdc033aba3c5400667a376b1e39eea3be1457cac3188df73a522230329e010fd13e4b7e4a90a48742bbc2ea2573dcaf27022f0b1a860d01d75011b49d6d41155be0689e7d5089c81c4f215ac1fc4ece1429e5e4e54939529604fb0647bc48771b8ee7030e7045f68ebf3c04a1f1bddd96df556711ab58da58246520c5cee39832d007bc1760eec92107e1e0bea5d36168fc5e4fcc7273373b0ec58c4d0fbe9f97f5451b2502d8048fdd3734db4156cc77e876472677c68b9cdfdfaecd1a2d54a6dc5a8a0cfa8f6b164afe49bee041f7cf6b8d9ec33e180e71f2cf7e91bf57869140a929a1f2a5ca838e77ac9b0883cd69c22d1c1e7f1a33286aa9f48e6b848a9973f36f6df6d5cfd8e397a894848ec635c16a77b94ac49a9e28a73f8533561faf9ec5c954e9b66ad532a805df9f6f895ce67b5229baacd863c80601c16bffff2eccf58e5c8760b416ce6d74698ed797d7b29885c8d7463c2624898017ebe600bd76f5799e9a0f386ee00d77cd7a3542b10eacfda78d8b15475b8f01909d4d9218c23f8a585fae05ffd6ff6f01a844a033feac8ce51093237f085b3a5113aa05f9daf681b12e8d6cbebd222c48d4602b8a431f056ac5a6c8ca6ebe44396af189c9d3399152c4e9cb09ac101c9c5c984d1de7999e599538fbe3f1c957b0f7172d032bb48217d42fa4ce8308d2e69abf63ad239d49ba93638f36c5a5703e91a9707a7eec080ad3c39ef7b806edf165af7f4ccad624ad998eced5a56d82d42e679a4c9616e351d61f7ec76ef8f86537f7d7268f328cd17dea92172968548bff74a46d0b9298c3a0d6fec0a69d787037293b15102a3932a61256af29961664afa5dacdc572024629c7a42d234d1cb03419a0bf9a041b303e5d3b6b7f1624147001783bd2c1d2a2aaa466b165e79b6eb82be52032430347f85f02135d476aa90fcc94496a673681c3776018fa214036e45e7fa75005c3f69c9c6f9013e6786b600e858f93bb68444065bbc8d57b7c1c49aecf69e6f285edb3c15294c7b5a646ef1ef738cc09b03885291cc4b33b60a503b37388163a7707f477c24dbb3f5db81fcf9ceaace54869cf26f5c3db90427ac35779788b71460bf142952af2efd014ece0e4c3389412e1588114c54a99db8b45e830699ac3dd7f1ef5c8e137a6d14dad1241e4cbf88a221be2b6597c9563380adce1f8a31449f871f755576ff281c06cc3f4627a7050f7428867fdc16af2d7d24d94b426cc096f72fdf128d1c3ec02e312a0945f0704cc183260256f8c2f956fed779a7872550a71509fd2f170f4acf4f0be31ca5e53408739ce18aba93313c18a69ae294581fd62609d01b88374052a8fe0267bfbb12638320fd9e4a192f62cfeca3ea5a19e682779b6d71afa284395e9806bf9f8d1c29015c0f9b76971e6523825c4d31861b1eee5c2810ce610ecffefb708efb996c59a6bd93287ef1ed6c347c9bb6ebdf2393c31d57c40f8cb7aff09855b91b90deb679f7d198ea02b713c858c198b907767cf1594c2f40f7b340864ff1dce1d2e196e7f493c7aba1f9f21784db2fe3a8eebb5c40aa864822a75a387c061da7d0848d32da5f387f91a175e9aa9f408143948b8aac0d30ca26cd978649a74cd6e126c42c3b7929f38ac044ecbca06cddbfb3c7aee389ff2a9efefd3d121c2fc2cff77b1121d3b5f4b8d0cb360b4dd64dcbaf4df30b93c445614534d6fc32584b4fc1fb7f2cab2c01f41d68464c8b2bf3f577a4a0a71739cbb746d650e95082c08ddb91bb76878cc8788e64fb7ddd9e4ff71d454b34346041f0f0b096cbf5664cd47d4cc4ff7d74017f3c44546e1e9f73a5e49c2a808edce8664e5f3df81478d06e8d2b755842b802b4120fd81ce597dd11c70b968c6b1cc230918322de66919308558d8c05a7b01df8cc171d67cca530118fcd4c5d7c0ce84f1f984ae8e83375a93c027a235ec62ee9833d7fc02d8d4d67ee5272f5677c1311e122e6528d33b55be9445ede143e8f23d6125913f9fec1bbc2ca885f133e3e207b0b3174215f3b993e0469fa110aa10d3b2eb1d761fb8941a96d80e1092653001020c83f20bb239d52c1aa32bf2dabd94336448ace6988b80b28ec64f60b6e26f5dd4161ccf4685f7e2ad8c92874da90384fa47533ea3b807f53d3f7af5922339449e9a2b06ec7bda27e7c4c0c8727512178f97fd59d28939ce3e3f6e5a6c4dc8e94781e103f7991b32656729fccaff24d680d4f25c1c440799fb9da85b33b06a214e763f9a55f66b3cff111172a78ecdaaff9ff27884afcb069a5418c3e5448c3e95d1ded903e4aa76ff290474058b9bc388c82243b12ec89e764ee9687bcc430bf98b075792708eb360b9f9b84f8a654dadb9bc88c9d578ece8f1b98123089520a3f0408adbb818ce29a4a462df59223319ac3d2a311511e9f7267d51786b664599c0df58e4b1a1c4f08c21e8ad2b01b51cd3142382df38f290b6026032dba29ae5a072694f37c29da7c20bc26a9894740b724419090e9fa4cb98a2b64fda7ad57dd0e0973674e6fb2827b761bbc10d76c98d12b6f380802f374e7261e113f1fb19a44f3145ff3b782574683ee564eb49b33f5d9e10736a61953140ba6cf525d3eab663cd9cf033b161a5aeb27f052fc86816dc7d3e82ec0ca9cb489c7fa198b4fba913a93c2a5c55e4d04f7380ec0f4389bfe0608ba1a2b0de447cea555afbac099d4efef01e654ae3e7c80b7776088e7969e7d384439f9a86bf0c6bbfc2e7346fe97ef6323190a8d80b50d7dbe6aa0aa8e9e0d6a50af4de78f4637a2f5a2ae9af29db783c773c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h8e9a28494dd201e422225c12a8ff7b73f29abda0d5d578e2e6f20f81a7881f71e2c190ea88a8eef729ecb4e58e5da4caeea395efc56bae0cbec2711dfa89c6989ae1be04623169100590e01c1baaf70c2010757838da7d7a43ebddb5ecfc2d053c9280a48518026835f8b0aaf2534a07dfd5434e932426d3e9f5ab8913366045518fff7346eec81c7ba0f12de14d0f52758c88281711016947dd9a6aa1aefe1fe9e51136643eded120be636378418988df82f1473279f22579f4cc877c2f2a9f45665e1491d3feafadb20c8c78af1b6c877d7f6f32edd97f7d67f7d38223b093fa02d51efdface123bc881bc5c9c7252badcd5ebdd51cc189567b312e123bc3fcec82fc189c4e9f57e887e51b3b08f8ccab7c436a9be87a3053ce7b889867a9abae2a6d73d717702ad78766cd3276d938b6b0009e03f1db4c91197d4f6a285eb3eff00ace161ddbc3ad34e2ff558fea23cb59244af97fdc8ded4d30a38d70760956d4519e0c1174ec5e8ec4b6453a87c6a170165f4ef77c53b57362c19285f499bf7a7b5672ba1c604d99a90bf3cdf2f7c2b03413395d45b2ded64e6e02a837d28ced8beaccbf0157e00952b4aea3d872b5f297808a7c929ca6d7789630cc51ec25ec76e5fbc785d6f5a142d43faa75f3d8ae1b7b5772a8c75f9a1982c1d4560665348b46d4302ee7afdcc79537627546c219dd0bee8a74652a676a0bc78f90c77c0d9c7c33ad4ad2691bac2d5d21b1cf6644686ce66dc4c5c29adb1037b5b5314d5beb46c5d37f53ccc0b4223971c0c75fd54e9a5a72665adfc5efcc39eb69bbfbf70ee17a91afcabc6ca8c15f4b42f4bb9d10ff6425bae094f9dfb0bf3a915a9e51721d7ae21d455ffe6703acc799457cab4607391643004595fdd1a8be077b4f0026d011f3541d1457869b79c346eae5cb78f62cb93c73200325088ff80562a0252628eb7cd80910f5607b94a02f276b805d8d9386aacf2c9807dfdd745c3c08942382be27ccd37d9660db66abee0962b7ad24b46e13c0baf4091af6c7ffb21fcbdc14f4b13a3486613c65eea18118b7238b0cea6ea4da7ab6fdf5e5b967f0ef65613992736ff82bbc0de1ed1c73de01a8273d81b5a848933300f59c12559aec9f5ecf261e43e8e24eebdd07954d97ebb300ab1bb3eb060e30a0c800ddd6ce9a7421f549fb0f0b88ebff7538efee491b16f24008ac35770e77a4ffc2761afb72809d282d129f97423a44492d6267fdaa48bf8a71b6c1d21a14737597dea0714a8f7c7fd08726f863df87eee43198e61eade76f60cb0ca0efe83aeb137f34be4130288267bad4a0050c34d7bde9ab99f0d408eb4a727e4e9169a59335464c8c0a70734f334fdd38ff815754eabee0306f8a92df69da93cc07b545cca45f05c9d0898fb99efb608ea2b54dfa559b4af7ac6dc6553dc0339d1113d7aeffcdbed11a5792a9743900ba2f49fc5e90c5194342f0620429d6a1f9daab5d32178048f22a20b469339a83f580b586b0ac6ed846d9c6c418b692d17d560bc25e5cc765f7ffa15d3b1976e95b6216fa7c8e1c1218a3bfe7fba56adaefa79aca17b7c63602fe007d12cd4924c491942346686f43e5b67b60a89c2dbeadcd137d096d23177e54c444d825f21ad205c07e88e637d1387337b8cbda9b977030f62f72412d82058014cda889c558b249d6a2b2fd3958b8b7d3bbcbe191f01aa8f318a908a0aa9ac62fe88af49c28f0023c19d3162cfaf6a946b1c4600ea0f27af0ffafd51f755b875584396309a2432de3a3c7a101fcf9dad6c804aacdd9837c0fcab280122dbf73fce169cf2426a18c0a0d41bed5852e79e3c297dfdaeee37abe32b9410c053e6eaa3e7c11c4e834a6f4f1832dc85cae126024e5afe4f24e4c17ec5e978b577a306e7b8b2456731fea6dea7a31806671fea2a5dfb93b31f4e4dbc9ae3681158a6ac4451187a1381f9a93d85a6efc1b03f19820a616b284a48f77b2677409b53cd5f317077aa521d384b632e005ecaabe698134f7d18fc94e75f26947aacc371d7287d3101857443d04811ba7e3204df429d4b2cfb67abdca25f1879147f8aff1fac8d0456d53ed2bd4cdde6a5db85e43ed7f1a7b1a27872dad70f13e1493cacd8c1fea64d3de1d9b263e5c3c19852da9b5230f4ce8b9a9185e9f76fc0aac35c45b1443ad3f51ce8b2e5cca77e5a27047aa4e073d55e862207896e91c14c48f4ed64274ff24875519276c9da8b4be74674f7ea9dae52fe8a63550b69cedadeca97397e7085e68c9a3b924bdcbd773b3ea660aaa13d18acfa16ff2899f899ded9c4ea4b25b92113e3d9e6a1711fa50f9004419b881cddfb9e1b0668d4edd43d3802778345a7cf7529584a9f80139ac62e5a6f6014be4831b6eaef899037a222348dffbf3b2c5658e68d1acf20649049670f90148e686f3e3f49d0a24ad64637c9adafb546796340758d66791681e305b3c7a2aa4a28142831fbbf991e3efa472000f067830b5e510b85d9c6cb9b3dd37d4d8e1e7a763514cd99852b7497d9ddef5cf52ae34d3ffa5da9dfead6646bb3f594ca01abfe4dfa0a825d7846e47eed357ddf7b3e684680eaf5fe8bf0674590f50f4e7fd6357bb073a86643c39eb4db96574fea118438f611ac15afe9c2f9a193b29d09a7b03aabcd429dbfba4f575cb35cb1ade872630ebec23c41d36aaa8e0c77b118fded172c0473b6492316fc909117b320fa3b48be3ac62b0517e19b29801d627ecf148764300eb5b1371ad0f52c2f4611a09bee833ee3bb5fdbd2b5ba75efa2a6079f8be11c9bf75423d1b7213f7b23f4c1f2e16ba262a7731d0fe3d9a732794948e017c0cc3a41b89341adbd79e38a2a286e726265d7d1e9346a78108bc383ba31aac93c7f39b080f1e08900cd69df8c2913df75458bc541b756aa9ed1fcc883aad0d046817bac3305dab736c9b2d7bf1d66c02c4e04d96c4755f3c77c84b7ad21a7b8d2892d7058c7eafcc3a76860591c71f2b58135afbaac988304dac1c8c04528edb8f233abf22ca6cca3956e28ab50d76565c5c8d68bf604bab6b57eb21c3a41372ffaebb12e03fd3d27c3d444157569a838e99e14f647a7a0056f791ec6f6b5e7795152dbf9149924b57a828c37dd80d93d81f8eb2c242df95dc04cb6f2bbfa56ba65ecff7714a7982520f6580c448a816f96704a4271b348693ce1e09e299690232f64294f3214795f7d5ab55cf8a35a25df03d77c9782033293111af34d66302eed21f7c3f997c0b34bd17377534ee38369a1b05c4e18e99819ee93922f34a071d31de5069744e782f06f88e7cd327b77b357a889d616c892eef4d6975362525086a6243c880f002ea538eeb12518a92cb843a4b342f9c04f41559f671b9f08e085b979054348d963c0bf71c3094e4ffab95a9f1b1728da10250aa0b88b796b67cc869021b024ce69df183c61747b8da9aa4a23ff272a920f603239d03a938856065f900ca37fce0e4df475ff17d019c28299b74481b7ac88f0881d4ff81497eaaad7fdcb68cee57248a89e788d9bdfc651b53835669cf9f8ac9e913381ba2801ca96db042219fd2dc5448cb5104021abae2d3284ce1742b077e890c2a1a2cc47c66dc0d48042d7280d175d3c48501bffd34cf79875e7f8140e4f21fb220e008179dfa74fa562ada64a3a3454eb4fd03ed3d22ce250533c770f5a5d52369086c77f19c55191d1c576ff347843948f54933c1ea7f4d9f0f7958809a0cf6fad772e17a0c7818aec5dc9e34139893f585ade14c7310e15f5f446f9eb614175286e431c0911b5a0088c49191e9a217380c45115b15219b73aecc3a52320b1013373ff29d60e3f42ddccba71f943c53d3c2032218d7ef97dd31093685c3d492ad6b5eace4354ec5748ad0cc8e248b80976ce7bfdc46fe3b3d3b040135759e97bea8fc3944ec4175f137638fd82e45b4203c18908b2d25bd332da4c8766e2317cc8df813f39c74cce769807fce873cba64c877509803bca453fd0cd24e4778afbea1a1f29e8cffc1d19f12e7dd47cedb4093d47586f134bb15bc2cb865003c5cfd590a53a1690faf81c06bad0511dad42130d80be6afa87fc6d4bf1eb8ecba667a03ed33c1bbf3b864274577dbeabcdeadfada18b399d74e4e469e297346d9ffabfe1e30e860568345891fc94ce8b459b22246f9acac5c873f40360aec1484f853e0cc7624330035df270865815043c37725f0b3be9b77e5a5e0cccb46da155dea16289259eee18f4e6014c8526b87d28e6a54bd23353a6919992497c97a741b5bb81aad27bd243be93fdb75b87df45361ce036424ac1baad4a13ec68d4263e5d2ba13433c5ebf27a038c97d67c2abe11e998d23af1f0be873c8c798f108892e0259ee91b98b5325a01193c9d56768a22a4f4a5c4f09e2fd1f4d0787d8966fbdcd872012155f1307884252e9cb89c028c55df22ed3ee77b5ed59bc7996b3eb49b796663fe11afd3a57485554c625c220c786669be87b124c7c3bfd0fbbdfd1ad45b521c8c5eb0e2319ff3719c0b3de056f3416f5eda53122cca640dc4fe5bde725d0fdaf2cf499d826215208aa23e17cf3fa6e4974cf66a41957fdf8f26ee85c39b16781bca0bba67af380411649f0f46e493950db5a90bbc17a907395cfb34332d2d5bb957da037bfb3bbb75365c399dc90093f28838996e1865c6f299af4c0cfd2f5d6a11f36a3ce0b7d9c57f39f1b651f2f02e9c932ddb96d4f0984178f0d98718e0920053e9a38ec24976390d35793051648db8cb099fb7e2ef68272c78403f72e9d4d7fc358c5794a76035030d3be4e8696b6335c540143a03429897f4a4b28990e406c9b8b350c1d9606bfbfa5c7595f21f63e230c395616135968c272f0f4d0dc69980ed912ac976532b9ebbc8e5a9137b668b6f58141cd87f9545c1fcdca3d8f3011376e7085dacbbe3ab70afb408cf2a450d32ac8b6e77ae5d15c9672866c8276f25b9564a7f8947b9fc9df43f6f4a8810bf7fb56f0dd9a5f2add72a1af01044c251644fe06910f7e3cf635d022461b4b44e1e5773c1cb0baa06429b3195532aedaeea5b72c6adc7a87d654077f8e921eeadc88c2a79e9ca8dde1286eed24d2b9d12fd288b9f758ca355c4966c3aadf193b983f9cfd13b8c031e1fce236eb8f6ad7da646918e4aba2759d092d2c5e7b7be7e285583bfd735b0cf754a35d468e13694c71cf4abf61f458025b2fc328748caa42a7283ad1b9c1ea780bceb6cec6051076ed979e99aae63bb23a86f07c66ad2c19cc18df8ac539ed0609fb91c0b5d3fdb4d61f44fff186e883acdca697bf1f856b5dc3af24b72d880589d662a05291dc76cc23175e8607288677fa723045067749759ef4a0cba56ee50f7f560caa7a8e86e3a90b1deea8c134fa0bcf16e5b9c11ff29b398006433b0157efbe50b6c0b8c89e5a3a84dd726afa3c8fe7e9207b179a7fe44b55d37a5b06fa2ffa818f9949d0df45851e3d55a06203b6518fadbadde67e80f70c6b3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h12a99fe73865d3acef7ad1d1df79bc2c995b1b5a1187a4acea85f2bd9b3d590004f5861a2efae0b9a6ce574555b52ea67e94e17bf86bf4892f0d00dd33ad83ad1ca750a6aa73fd544cac8b14f4ce420220346501090fefdba0a616a4c22393e52dfdf25d357fd01f8e85151ba9a0dedac9c9f97af03f3eb570af365c91aa35635d728fdf3bab05698075bde4c29ac160a6087948d386d061b829ff9531d17daf0b42b9807e6208899d0ec6e1d1ed3fbdce89bced84a7e0e4e93e9f05f573e3cf60bc4efb45057f46f7050f60a3a8d3bc7ba3f612c9569d6de109b07eb8ad5eabcd8ae794e0c5cd437a6f627b213e1e8a7adae60f1f7b3783ccae8dbe2aa6ef6a1da5ea6de402d3635bb1877479f80e6a3be51f0aa06bcfb49b5cef1b54231045cfbbd6a2cd0c6144401768fd9d9ff1a48e813347eb3bef72e82ee0d8cd4e04c3cb491bbbe8eb3ab4d16098fd814b9842c36bd235421cd0f1b2907f29ef9f10e6f7f9b1b69697bd13c8a4ea905fd57656f8506f7236dbe89ca88608b6bb32cd69dc3ce1d4089e5bb82d04c4e764276a3d8fa169110c188d30307488c3ab641015d5f8319cfa46097fd0b7d3482e29319805fa8ae130715ffbd5d10747524abc39de8745e8dbf1cf7899ce6627ab5e76e70e74da832c7d8458d6115c2f7f17e53fd5331b86bc1f7cd6449f1053d9c6fd39bac5a7f4271654bfc2fe53101729b2ea391e503c9b4d50c663f7b47b3e621e4fbb572c853996e8f0733a515cf2dbb73a643aca43e83a3bc8d9e2d2f563162ba68f797f7ddce42ea074054f72e46ba2f43e48894cc4ba168ccdaf111a04884e0513edc2b2a4d361922321aa30ef21c6a831fb76017ce869a3fc9d4df935cddc37782ccc17d312faeb387d5b2da656bb3592db3ae1f6dc29eecc754d65599efd1c24620a0689ab43563a661e5edb553a66b1387477712331b445a69e7c02896c62e4b2ae94370c6ef8704361f88f40dd2e89b546474238b906281ef5f8281f641f3449130f7696b4cfc71875d24fca58edc5130d869bc177e6ab5e2a4cc9a0e5995105621cf63bf75e74c472869f885edc6dcc44c66e4e70ab05a5b49446ec746fcc9fe52b5cd6a885d388b1cd66580573b3b3df70522271222df2b4fd1bb729c42997ecde35cc0fd1e6f64258f2318a2b06b0ce013d220dd12fc343e5a14677bb3879afbfb6ca8c33cde4e204f285b0d42b67e8aa6759e2b49cafdbc4c3bcd353b7a0e4aa5e73230e076f4f29f9a450e4240e9d45c8775e880fda49da3f6167be227f7fc0bb339b103c0e6277c4bf688c52e6be4c91ee3bf5d99025c318422361c18488541e28fa8179b55339c39477e0cf97708b756e793e0382f9a54ee64bce674fabf2bdec335eef8dc4723c3c4cc65b57c38811859c79ff22c8fe47bcccb7d067c492df88675b49e508254340d0fabea334448a9de4fad0fa6f8fe7d5e148911dd14ff7ca9cb2e580321cb3f02d883efcec53377fe0d59ae076a140c1470207c35da57f0879daab43f66bb8733bf27ae343551a95ac14eadf52ead6d993de42896b64a452f4f41f215d1b8ec1583528335d2ec4356f2f66ba33b15704ddefe28262ad0559e4ff5eb455357ba4e2270e20c9bf5aa0e34e11f2fd078d59391bb65cf52a5d34e915df690bc2967c5a916eb442724f7c8f61d437a4a5a3a9ca8e0a8a503876be05a9054f49fd9b911de5313ac636856aa0588b61cabdd8d207d46d82ec6a94eb23c99291e8a0ca730f37f842338f3b834ce3ed3f3f33598b7ba53a8baba1afec440a29d0cd8c8cae1b919e9c849a6836d1adb74218b25df6348b23d54e8ce5b0fd9351493075f2de72c6e126655716d9462120a2145b5c85b891354a85cdb540e1d83749b01d9d09a446b39ff700528e1659a5729ead7593decd3f6a2406cdd36eb723b45ee141a1b34c9d7c208cd5b193feff2c5a9a2ce5552e5d0adfbe844e8b76f792c23a3d4a47fcf8edaa63f60edfd556957669b48d3b0b40371741f5f99e00195db4c3524854e7f71c7f9da365bdf32928e06674c855b3cc916ad2f002bc67a3a990dcb2c7d3d628d626b57ea9cc19853e7ae9a4cf5cd0fd26b50c7ada8545060f7a4afbfb27295b4ad8745831d6c36d70a2f9bd3ac9cd693eed9849fc2978a0f90c28ba564a771389998476e93f733b23c0a6a7faa5b9809eecee245953e235aae49e93f9bb022bd4a4b3640ab8838ef490ff81309c1fc4d9291c6c3e8e5805ab6e63deee811a0edc5f500c706a552dde6042a2ba608fcca32489fbc49311eadf54026871185c88281c1ac2f1c0f5ae9a456cb8dc8e84f18920f65c339f6ca336dd491d4614086b946ad70b1f58ee8664823e69844e319b9c19bb7a78ebfc715e987dd00eaa70285d3f594e173d5ea0c18a84481fe1eb554bcc2e9893dfc0eb172f25fd55984168e4728198ea3f8a5928c815a10addcab22e5f8a8439d3259ac185be674de7842270cbce1b6428f6e2d2ca20b9d3a74da355928200f5456ceec7615f19b52f3b0e0cccf51643190f654b729854c219c2089d1198358788653ec049ecca7a712d7a581e3639f43f3e82b82b058a69b0b167a40dba733b2e86ab12c73025056113a736b59813f14fc73664018cf92574e3990c32a94d859529a61227a10f07819febca344f128a77e751cbd074527f76c3f511a2c9b99f98bcfe5f15f33e950b26f5ab20c28e0edee4083d45065e5492c53729a2929fca819f7a81a5b0882ace85ccfa06fe9384ca69fe954a48aee0d6786624f59bef5ddb369ae1264b81e9610d6a57b5e8416047e94d07ede270fae285af6b5d624361719d09419535a763ee66dbd1c79615152484d62329d20d228d04781722e197e33f62ed0da54d9896d15eecdf3c4c1d701f386b997719c2f049d84326831ba78f3cde1e57b7d4d591730d9c8767d59e3d7cd225a9b76a3a97590d08c38e319434383e9bf31f135fb984323a3cc2f8c216917c7e505b93132b92f4840d00b4b0375b3440e667201f711f1d470c162ddd038b67a863fdaec06fed79f1835b9bccb5469f63bcc9af163295501ed6ceb15a902f68ee8f4fa4226635c1b4b2e3eed1e4eea35cb244a3a9e382c75c757e327a600561689313925d5f0dec8ddf2596875fe493e2bb8d446464902c647c2a785dc9a745c3195335d86f92598e4afa35446a2ee4b0f24cb4c1d33d5a5e799443c6f4c4724a96300f889eb49c7c847dcaad0f14bc3d9833fc09d3657919c8e12af6a34b08db17532392876b7d307fc2a6c9315083ec10ce2728db3b24f85982e1fa534cade494df37122ae956187625d95b8a1a2dad9af9ccc7434e30aba78f5a125188b5506de3fb5f2217f46b221d411dbeea3e63a4d0e548a7da42267740ba29d4567c543e54cf9c3e170a037baad1a271f2ed32e4efb7b2d16e993658f19c8e1763526bfa5b0f75dd73fafb5fe7de170224827f5b1887867f6dd8e93b16804e94cb7fb7b47137f28f230afd363100a3ecf12ac4527edaa26f654c530bab163404e1a70ad94dba9422c7562169473984d11c1006c5d272954d337e41be840b7d1161becbaac4556faf33dc652573b3d0cb7256344f0106e1cadf031ec0a562639b0ad25730d71eb6a431a2b0e77fa06be346d28ac85104de5f66704fda03604c4b3f860ae135649bb771baa4cd2a8c5b0fe49746ec3c4a7140a6ade430ac09fe211c68bbec021dd8ee2f47584b1358ae4843391cf7e5aabb86f7365c52c19c29b0dc8a23623cb05b35020e667a624ceb6b3dbe62d4dc3ab950143f392b075a650b06415814371c11acba07704295b65784c0ce0e47cebc6754f8e46465bc6684a1da3b056b13f36d8d831f9c89b9f6c56937af8417c3e7dd5110475335c862c43e2e0e60bd2b247e7dd8f7661b946413a1bf9e36ad45e05a3c30df03c0184b0f3c3833e5ce8f3bcff5e5a3eb06c5494258f6b5bd8be1093a5d5517db403acb05d264cb357796668682bc3bf665cfcae0dff2384bf8b504ffec94776acc50585ee9312a80e1b70f098009d81eef7b07ce93524ba327c6c6733d5f9580379ed271b4d35e97ed7bcebf11cdc7c461bfc980c36723b8913b4932c90897641af5f7e8b567e432fe39979dcf4e56a73a5a5c91120c5771cd1b55a249abd3da3bca3ebafc061035d8210e0563ac3f0d0382e96b993d15b6bd39784f10ab7e3340f09946b4b51d8969ba658191c8b231b5bc29e92d40b9dd617601f5e47edf4eaf4b0ae4e3bd5a00cd85b597ae00a11e58661b714476b37c867ce0df0eabc95e0697e1384d4e556248bc2bb74daa5b129cf7957159dfd64fb7db7d4a442e79708f246c142e971cf3c3dcbe093727717e77131c9f3533b00581aaf9c46c937184140a0bc5a9984a3f0fb7e655cf828f7aba71bd2a75fdf9e0e04b2551b443dfb0326e3f3e20ce90ffe631e7b931f588eee5df4d094c414d1c106af5c97b900bba929789e6624f1c063f2c0eb854f527876fe5f143f218be72e77c2f1613b500428fc570f4dd619b075c290c4c5f91bee0d00f52d2cce61ac2b3499422bca25e99c63ff4e4a230cd3b7bd8a693558dce63caec25a78cd85eab45866226507f5ef3b0f424dbc3cfdd8cac79c45fac7c942509e6beda5f91fe7220d239f3584cb7da12feba2bb10435ddac0bf902edcbf6977eeb6ab2d8391c19a94c083123ba11e2644328c87c1f70a62b30c3ef991519a071dda9903788a999bdd9be24069514ce9800cc6f6cb1b46e7258aad9bc85d5d9cf213afe2311415d18de49912ec6b1b4199a41d5a383b98d9f2681a5c5cb3b39587f3c7cc5774cb9f5e17e4920b9f440185e3dfdb817b04286e33939662e84df12af781b42e18f6d17fe768174f3d5ebddb37b6db66c776cbee50a2189f08ff2508125b1ac86d055d232786af5f53e4d5b6eeeaaa6c0f24aafc4d3e78dd9f3bbc225d24f9a0502d8daf8e29210c2efb33f1c5760593b2fbc54c14f82bc102024d2c3a6209a505c2f22fbfa30977b6e2b5d7375be07b6f08c84cd2233421494437f6315fa59228208051d9b9cf65082139256647bd777d6ef6bb3d3775a7eb43bc7b6e6afbdacd8bac9d91f569aae69917623505912764e47f1feaff5a876141c6f10bf7f2331a2770cedb26843af37bf78d3b66c3ae2108cc61cbb949fc88f760fc8db46ab7db241e59865c490de4b33f01682069d03914f7bafc88275e011e936003d405111badf53a8cbda24cc05872f5120cef5550594e0d1ca69faedfbe8e5c2916c86586722dd450cc787e99af6cfedd1108d4e2d667e0082ebd80ac948264df0fa4291eb438ab0988d31fe0716a90efc0f256438d4934f44fd1b20ca9018ccb50078a5a2b21ce009fb669012bb1ad62abd292ea5658514c6ed529281b9c3baae1148e7239574f421e3e38520c1b23c442f48f3df6b33fd8e37a3d19e30b8c90149c475e45a719f01398944b295443731d0482b4e8d46efcaa4070762;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hf657d2d94642a653f43cf5e3dee1be49598f468c3cc90b5001222b87da73b7fa2cb1eca8b77e7a83a4995d9d42689272616e0f5579858f0a8cd94e0fa546755e95527f9c2abf353d2a94df8b9be6034e9dd4231cc3c89c5d42b7450ce54dd42787400871cd94deb6b4531b9774f67bdbac24b2c938076bf01d00f6abeecf21cfc4001623087c20fed350fa4c1f38cf4feaced0bfc678a205b717b63e45f81316bb05bf951465fbe932131a98a897f6b09c4b5f84b592137fc6c69b2e6f8c4a2b02c979369d72f67bffe81a8f7282341d30f43518cc3a8cf9104946c0af50149ac625bfa7b98c9748d1d5407a505fcca1d37cebbea08c9454ea5f7155f7cfd3020e66f9748564a047e25849488acc0a0b6f6033b685393766058f1e3ec817ec45a04e8510a608d86193618c51ae5d2d48cd4983aa4b77c7c9bd1e163c8bf192bab97d69f4447a43c7fd96e1d3fafaca28d92ecbc3d38187f1fe5e2a341b9dd7b91604d1b93e7531ab37c3673f88e28d80acd169ed3baadebdd93c79120952d28fbf5fc163dc7c87d76792cfa91fdc60d252cf68beac744f6c1ef93648123a21699bf5072e1fcd0e267cf5747a8faeefa79774bd2ca808444c08cda4a6e0ef07fc9f04da480a36f1fc81e386f53d4e9d2d9e82b2ecb54c3926cd02f215b417fdcb55a6acf345c291ee4b986534e7fc4cc1065e9cfcb0f71c9134de9c940cdbc3becd4dfee94b922d471a5fb7eb8c7e524d866384aafe3d12de24509b7060566731acde26aa8996f155d9440a7846bd0692d86ebddb3632d7a2119fe547416893eb7f525167ea266747e8e9d4161853df5528df6f9f3814c18511da6ba85361fab3bb7020b8fc680c3d6c756f5ae4e3ac48c70f76530c31b2ffa7b7675518421941d295cf9e5c0864ab07029aa589b505262c274c2b68a46b4c98b24a4e69b872667b6e653aab9a8bac21d7d1d40031e8fe87450a8b53b831a67767f0cf57cbbf9e8602ed52a81659b9346da30c85b9d0ac91cd8770f0787dd30c22015083b7edb62d54d0b6b50d31f4a5fa6def752200a3f81e82b7e3723eb2cf38eea665a5bef4a4eb7aa2958e700fc5ea4301a03937534551447bac3d7c8ead3f2f26c1e78367437c77ac30bda99d2c76044ff5264f9675b0f2f5bf3409702ce396398a98e6f193ce355a8586960cf2593eaa194f9cda6accb200f3b702bee93de014234a8c442292f914018dbc763c5dc7c6575ac094dc1f425c0a207fcd39cfb84efed46abf964945c12c5e4f176032a4c9cc1a1f348961390741b3d0bcf60381e6b820b5c8b25ccbaf07fa1fdbcb6c17dea91a13baa4dd2005f1dabd266f5ac89fab6ca1c30b9bfffc51d2ac99b51bde40d85cd0b7d26998f888694ea09c499d196255c7b5e5a87e09f279efc6f4dc026e88591f45272600b221973ee78afdfc6a471de5beeeb0df8ff04850713a3dbdc0a5a1730d797abc42afacc4eba1033b62a376672737f4056fa78c4b0f5071c0553d31ad244bfe50c9060d0f02bf673348165c50b14f18c8ca684a8253776d82b7776f30b1786f08deb4824ecd7dc9b5dc5ec96440fed1d72a5a0bf97c3bd7ce8fa7724e44afa18226e7c664f94229dacfa9d49524124b904c8ec65e84a28ed302adcefed1dd5f6bdd5f626c24add714f5b0b358b41878bf5fc4b35302e5829a6106cbfefe7fa5582c41f8d9af21eb947587b36b356b2e2d18b707acabf79961ea5b6c758a1172f4435303b8b4b623fad5350f77ca5fddd1cc21291b02c5e56f90614b58af28a161536a678aa61c33ab769aec4abc686536b330ddb0d8c408716931115d798f60b391eba3dd7e9a85ba924bf32874ba48eac2aa4e71164a384f3b2dda4467fd8973aa483622a761c36d3789ab080c797ab62d74b83fc591c6d2bbecd220fd4e5af0b01070ea4ec94bc8985dcb273c9eefc04c2a7aef5650de4540bc64b29a1afcf74b277722736d099590d1bff70f569c3e675ca39dd7491bda51495c9f5d56c59c5c12c41c8b260157492b4fdf77aaa089c6ec3ffe3a38bfec845f2286ee90ba38ea9ca6e882ab0452de925f4c4fec98b21be75199935b1d29b5b27c674aff499b7e9bb3a26be037436ef11095b9c2557226aa0ef638e488647ab69849246fa06a9942da3e632bdb33110b926b45e27b444d6d58f8e5c864b6671474b2ee04c36b214bc0433e1a23bb26f5cab2d60ae2cde29f66d889dc4dd405a0cf27722645945b9eef6e19ad19ab8f32bbe243456bbd14ab96282089dd6bdf5f2bc48336dcb6033a02f646c64d5065e12dc97916ee1f3c61194814645f7131b52357b506229e1bd1d1a227f452dfe47d43b6ca20d40ea372d3db6f0dfb15ef5d1380c8461e0acc6a0a5dfc9f6405fc6152652ada8037bdc6d578a335a82f482898b9d793cd530d852545e936e5efb5d93903cf73a4fa96c279349711d13bb70e1b10edea9a6f4b56545bd91536fbd2bc254eda04263c2f384119f4467f694adc72061bff570b101135519a5a711f93e93211ad4886b9cf7977ce8705cc1f5e893810e7b4ea3bb9d3c48d9584bfa94266bc2dbff05d93cce6186e86370170b30d405c0bb8560e52e6332d22de7a5d767d5a41adfeeaf7a70e4296db1dd3279d145c5d3e8071665f9387c8437a6523cc54ce0d3b82c7a8c8a1aff8d35cfaf52527213c2803511effee684c1442a647c3d3afa6b69cd7e92f0a6e293f066344bd869618d207782b9cb4ae5c2df642f55e172407f5a3106a24b4b3196f9b6fd5af615ea229735b4967ae5669bafaf570e4361424232d8f9ccab39683f44c12e70772c4851dfc3318bd7e2d7f4816bf8ec373b20f3e4fa13c60c1d20a771cda1945f0020ade8cc3fff3a356d9384122d647e0e7042e8576a9f756047979d1cc969d371fcaaa37c673bb44d613f9e6fb9a09aaa9de8c9f743280d1438ffb3e43f0ae5f13956f7b3e3c120702d3f94168d950890a523180dac7fe3a10ac2d31be0ccaad2fc2a8e9a21f95831fb93aab6382afa07eec981e8308d542ed71b784e178c2fc31b7f15d1f0590bf4678506d24e496211a171fe473949aca0edc0f7baf73a6ad5b18a1cc67995914d5c42a677014ed230eaee26b128b35109041b0259544fd6e55af9b471a24652b8b5301a99f6fee1c7735c8f3787b50804e06c310105db94020baee240636acb1a72e13b3e442064f20dd8fd960bc495256ae1deb9734b99f889ea3a55e435050a76f76ba4bea01c72d9228dcd16dd20866302dff925f1e1155ae1b26d6ef7ab93539dc551e596b8e279e2340b63379130af0586d460fff17b771314f10ce9d86ba89eab2c15c1f18ec0fb99184a8a047a683f138eefd070fb9eb0c4f2f351dcc8bae9fdb7defc6ce2e5c68a784d0d9dcbbf85cc31d279a61f4385ace056caaa25ed04ba6e435af5520ccc21100971886a054ce9b325f25494ffc3c524b2b0bec9772f70aa83250ff8af8fc98cb4e982a24be8f3e67eff5173a078ca77cf7a5117a512f8e059d66703283e3f1889e4968f551d748726a32a3c115ae33a2f34ff4cabc67462ed95e3ee8a85991eb91b592dac7f2c8a4b06b03e44947ac2f617b41a408536903cdd3006510c9255abd243c2c8f30dca0d343028f7fb022bd173745f2069df0ef31e0ce24e86d171d6416cf08b2412802aaf4792d9f2ac1ca82c52e89b833c617d0e3d793eefacc3628651dc4dcc0eab5aeeb5017ad681972da5d5f2215f5706072c890e319534b01a94c70e0348325b18964ddfdbf0c16443f2d2891d68bd4706b47b4f10d72a63d44cafe3b492c74158aa27c4fbaae34f9297e30bd7e7732cca1c8a28d49cf3bda4ebd2233ba103b6e58bcd530c52cc4d52af55133693013967ec488eab7a4c7d479ce5d26218cd53e233f4107383fdf7b808d7b9e1701828e1ba0bb9441faafca06ad040e9bb3e57ddcffcb05670260f6fd21c334b27d75eb8fee2448ba67cbd4d6eb03ef446c110c08541b60ea480725a20fbad32bf011c04b0ddb0b5ec9d1c734f8436915bbe3579ec3ace7cf961e7787e68ba1770d6a02e872ac823e21082f211a288c32959626a237365be20ec099d1640bcc25948dd1e24286283e0e821033bef41ae3dc2c65f28e091d7469c89a64cef6f14fc18f685bd3cb3edd5cf5edadc6ad0f82ee819d221c245222828d2546cc4eaf2003485f28e41b8bb44229128211ea619973668706795b182151d32d0900c1113def044e0bacc92203282c724e939fe25467560451368f9d3359c916f6a9c71a4e640f1933595e33157bfaaa3251da1030127754e110b55ff3e6cc2165bc02f902638eaa7a3f1f0a6f0e324aff456bfd87ba7dab79afd0ac1e131855af738959a51d1731d0aafe456bcfacd2fd192dbb4fd81b602fe552699aebf2d186f47d82ad6571c381afc0da6127cedab8c6b64b93c4954a128bd98925ef1790a1089abb32cacb525dfbecd1116740dae936a7b38aea9ffe4c89ee7b8371a3125bdbb7a2c2dc784d199b869805119bd9bee621ad975b39a91e831ba7701954858aa6c8689c8f87cef11a34d15508c30f160ab8e22a2eddbc31cb9c1744426bb7808fc7b3541864c173a9f342c76ae8e605f62fd3836ce7d23b0427e688da1085528b10f90652fdc32589a868620dfcadd3329e73616b3d557df3e6e8f6997ac43e26cb69084bcb0436fa77f8dafbba196b86410ef8a332d4d61888c3d0f0a655bded2b84c98cba9d15217613afea33f5cddc65d721794fcf62e810b760cb128782f78a968cea31a23926640b25e5a4ba8f28cbcf7ba25fe18446bff7d9f1a8267f9e0c55b75836f5f35a0fdb90b1cc994ef166e7327d7637c8b62e618e9850bc4fb56b6694dd46cf37d0fbcea486ff3d68123f7c909773e3da1231d26d32180cef17d299b1d307b4c09b17078055a7974003145da4aad65258e67701098c8eed4a0ad0344c7d3c2656a26819f02f8c536d45feab72b99d592900703a1f5dd11d8f06e38497a2ae19d81b7f9ef1add6f1e194eaae1774677d703cb713097641490a836893fd24f83dddc4bfa80aaaf730d1be0f9cb42b62603506f3cbc6cfb135369469fb12a503c2daf200049f927dcba31b09171178670349ee20557aa7b467245d25041ea9e50d5a2e7f3a8b29b99ed3991a1d1ddc41ce6d590d769997807fbf4e94a386ff5814c05a58b88b7bf16fad2fdfcb8e91b58760fe1bcfb80decacfe19c1778c836706f5393bf0e18f33ed56d56d2e82bacabae5703e20fe39dba1f16b9d9ef9d62c6ebefd849e7eabddf22f42f21a4656004e3f44a3f7812b2e372aec6a786df360885037f853babd48be14f08c4c32e8338abcfa6c537c56f384332fa40edadf62f8e61f1cb3de83d9dec83b4b2048646361f6fb19a300c0e05f954cff2fe8772b2fd5ef7a340aa7383a768293501ea789fd99814c10a8475b961de230dfad2155ce7bd6f07f506015d3516b8dde5f27970e87e363974cd8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h99f31f538d9c5edd35c74e2487cd6262d27836749513c03dda4cf598a5fbc748c093a8bac86fe789418e313a9dbec40f54f97ed676d2d7521d38729eb0beb845f30433457b7d290f618fe1dc8d36ac702909fabcdcb303cadc4dc9650a47eb374dd93499518a036ad9d2445f00c0eca3ba24a5ea6580097737eadb245b0075a774ef83f77cb207e80689cc6dda4884c95e77eca4d40751cd21e4aeda11cd9c7ec4d471023fa1fc4026277c1206f92697bba7e58518366adcf679637724a391ac1603fd1b0d81854fc01f9877090c848defc23fff8b25037eb275da19f423c7fba21f10d799b279551b31ab82266a00de21eca6efd2995b6b9da4c555853a85adcba27f1db2858a9c40a267f36cf1dc241fee3f71583501ed81730802be99a22697316ae35095fb490c7e76d55542f1031d9cc9e1aa85b75795d99f2cd1c97fbd18b88101d5180315ec7b86c10155e9577a9d0d7109295eace1e86c76338f15b8e609506dd1f0de5a07976a3ee26455cb95098c57b776ed9412314a91d8cbeb789fe4c43ea8ef4c41a56f24dbea85f6c2d3ae1344d2e7507269c5cfeabafc410602566ffdb529d815697c0c37634ccabb0d7dd89ae761077e9949c03f3c3a4c0c7754adfb6a73bb59346dad89921904402e419bb2dcb4607840a1339ce612e296704e6e3f558573eba0de691d48fb75327a73e8182064360bb5f5f91cfd0c25332645ddd34433cfab17abf39cef2006040af601ac2672a292f7c3271d68e8f21f7e096e5eb671410ecf4a32a2b70ba8dd0d2d1f446316e403422f39f61f9b9342386dc2547fe54f0241748ce1393eda6969d0a1417f3a371390f2510e82d50b8645fe3a675a25ff3edfeac70ed9cfce8dee434642a2eb78f6d1f1be8ad85345eb98da7f28c8d2024f44c220a7ab89e81c4a0e9c4a69afb58bcf44f53dd534d62fb12be21fc9dc6c16a729666033aac4fbb03d1681ac588776960cbf64fd0520d46c55ab9e4eb4f3b369d043af7994c09e1a4e25bfde3ed9494a3ef1d9662cca0ca90ca4141c4eb002b3562970e678a5097d143504f499ef9454ae03fdba62c02f1144a477969b7afe052c1f87a969509071d28c850d03574bec2a973000b9fc8210fa285d2d5a1b0f7cb993e831d07e7b18d3258c2d4b5685f87e040d6cdce6cac284af7463bfb5db016db8e24b2fbf7bc2389b805e11aa7f44add2733093a45330a3dafe2b6fc9bcfd987be502694e214630f1de44e161e09fe3d0bf3a0f778e83f10883f7e4159a4f9f025ffb0f19e9518ae115a6ff5f675025eb8e803bab3796e6c5d0ea9ec4f53bcbb4fc9442175417bf5900b80e82cea73c135ba011d8f355db20f4c13188a765db2d1fbec20b8de0209002fdb6d0dd89beae07c89c974bdf667991f98eb44ae759310a1aec1d6f231fff6894c6d5a80bc8f77cff09a96ae47e55077c5a1525d60127660f8ebd8e6068fa745f486be098198d94f5d3d2d62dd2470ffa0edbebbaea3f46adbfd5ae023e83a70d4739649295bc5f1c0fa5735a819fa9516e07c830cd6d099529263212e3a4fd9c2ad1ae598500b0cd6f252323ed67113279b12eb1b6fed17c8ca0df0a0c4ce55df34a3b30a18475267a05d139e9c33fd9b36bac83664568a17a4c86d3fddb21391e5430e3ae2070d41552bbabc1c83f6129411b2645dcba1758e283921170cff8197de457ba4d25cafda87c23516c6610b9a8a123bb90cb5ffc06d3b730701439f321651ea14093b2fc53028897ee6f0aea1b33ca5429ebe1453915f0dbf551e02632c0b9d97370e60b160b14f7d3ff8f8e956f34ac67f2ed3b3da5661e208aa949e4cbc03053efa8f30c47712cca2eee86856155390601389fd65e99950ee0bcbc3fc7d49ecceec0ff1d082ef0dce543817733cf8a178b4c6b75c04e7955e78e921e715770de8543b19aeed0689ed9d99405f7c6826457919453ba812977630b4be76e390c60084ab23016eb74d386ff751c50a09962a56bb22a5204dae5ab4870f003f1b13faf82896bbd8685a9338364f1f2523d67a281262cf9171474112a43d5d50d86f871940e0b9f30b92950030be6e600ca58927507fa33fbef7d298ffe2b09e40fbc1fd0e4475ab63e23c8de839b221a6b0b9dee920866e6bf83b06bd796cdee8bd67c423c4bd3beb117aef392f8aaf155083882042b137b5d845bcfa6abc727136710d35623e94e9ed8f0e8c48eed66a9c97a3457a90600d468288e43ca97f61b37ff9d0a405b288ddd8d6eeda7ae842e425b42a87f80415d63b7f435cdbdfab5fe285ff20ad434a0eaa6a33165f762bb258fbd1e980e290f03a475f252e838cad8a8a45fc55e251da2b063161c11689a259277c9842d8b694931c1916cbc9364de8dc4b207a88685a16efd48b43aa2f823708c4b0b8ca3439963a6556dca1b988155cef41155cc4fd1f964ae35bb399c4314e8305a8dc09e7a454c26208a1800312b43a3050277a94eb033acf3f44a6c2aa72c6512b7b9f35f1d068039513f7632277e3d47c1b1a7c334c6315de60208a7a2ec23ff1e731d504546de69a9a34fe7ed149d68c630b61683f1f59522a190424e1975eef38cfa8c4dbc6bbdb78a6632a5a6dadec4acbb0f23b08b97a83c2014e629e900edf01e0d278329724d1f80f36e948e56480075b1468303a604bbe83834afd3d8a9c32e05e6e6d1da6f264d416be49c761ee432663936078718afb8e7170c4d8f7b6b3c5bf4dca1ea6cfa34655951f7f0897630646d9c28a9b0c4e1ae443e2d39b49b67d71546764341bbb82de153350570255e8ddb454b816a4a24b0a9397c7afae5b531fb14c03bd8edc8c6e48872708996664befad9d618b0f613fcd2df2e315508d34e4a7258cc023eaa076b7f7325fbc0989541c55b8f67e3c811135d2dca04a22ee0afc4a50831c2739d297b601973f825cb451d8a9997d97ee549196883463f87e4f21bb55425d1c276871e0a2847c701de9e4d060b0741063414613782d014bd46c5361a14fec605da31931c7ee1634e36b5017468bf51738a60baa5181801d9f7c8d4c3ed9298dca63d58a47cb5d4220f5c29197f2efdd25265e5641d743d1de4be408bb6884c19f5228a9bbaaf5e1b265d54ee442c5409b52e605fd5ec9e2845027b59559a88ab1566eaea20c4ffcacb6a5dc347949235069e3c1a7a50811074d770080bd4bc6b91cf9d52aaae8be63df06cb3d8b06363ae40a8c229d858d08f8acd2f21aae5da46d597b9cdd81e440ca6269fb066eb45dcd11448876f8843cee3e92208d45c40378e510fabbd1e5a3358bedf27814088f9559eb20cd56340b24fc7e19830bd922e786447227190590952e6890f097c93bf29bf23e478e403271e7508729bac12bc79b2f9ca9edf022cb0aa7326a0631ef6887efb1669e3710df68f194029d841e6ccf0d0fb8270b85f68359fcdd324382dc245378ae69d5c1acfb686e660ba5720aec88ab7ac873653bed233bddecb2b99eb90b9cecf25ed5f121de5d2a90e9cb859f7c9a549a061d893e3f0e07ba5027ab0a4542372aee109b95ebe55aae9fd8c4458d9ed77b8a960b17f2edc7815563bdb4e8e39679278081fc991e50449eb132b3d72115eee1de8de2b89fb043d0c7df9ddb7dc07dd440a8937c1761ffb4e40a5e90d4d2eb89d82df73b8a2be8cc910992d054a35a16651a21e9d8a0010581d17f227f0bcedb6c63aa8853ca339915e662822a17d108562c941ae911dddf55148c16cf7b06b903bd3b2d5805193f2ae963dbb15cea4729a0c474d16879e3570491f7b0bb1f594290e19936ddd3dd8fc9316fb8a635ef2bd220bfcdd56b23e245de98f36c5aa2ef97f5ce37f3ce4ba8a00a347fa9b46a839871479b2809ebd25f19fb9e37edd5a8a09100d71826ded6a28af2ac55b2a40e6533ed067782d1d9f1a4bd03dbd40c83df77b6593cf989df52fd1656cfab6efbc198045aabbd1c0180fb5f91d16359a752f053db195f01f2b2f4780e49d771bc0572c086ba1226a1420dc19a3581f6a7ffe5a78a5e82fd7385061d943ed79813f0089fe205ce694fbc6a309b464b345f23f6c12282344fd292b34d9ce997f9eaa2c28f5e878dbc28022c67f43b0063612dc173de4fc104460340230f6dbd9d8799decf8ecf847d675ba18c16982a9a1ecd0529f84526daa61ae7b02d2de87830a08c3821c36fa567a2629503d1360d2e57994dfd7f836cf155db89a41f645e1d96c7693602aff8f999fec70ec895ec6b0fe6c99bf2e93faec310f09ea1a6759537a94d7f5eece705a8e5c1c8bb588c6eaf1f60692087a056f6a2033d3456e47dda4ac155831b40fdcb7668f261f87fd25e2e4f690720cbf3d4d3dc95485595a1c363047833bd48533a2f86e0d4a1cf44b191f57677707b75ccb62389871d9a9dfaa1296ea817fd7b496b57545f67fd3f119e754defbe0f5dd706c6204866738060d720e1293b18db2309da94fa006814e2522d7050a22fc4dac2f898115b942bf83b13d2b2e7a281e34c7f8ddc659dc41af182e6241aef23d51beb19e1f73067dd3bf7bba66149679f1d4a6fef9cb5a8c165983c8559e80b609338c34cf35f6c4e563233095e945531d6115ce4285250728e2ab7a21a559da92035b566e31951cf8b055d76f602d257b05d3f7f741db4d33ff2e45cac1e1b6ca9f91b4c90b1e3d7c8f69d39f9ffd563c70d9fea4692ee9a9cd90bc39cc109067e038248f7c5c1321203dc1d8b31c9dbbbc5c88018bc0330cb16b82125de2ef5c377586478fe43a7c769ae80a9973f3f914d158188068a427e070dde3416aebff23d9f228813ebfb314f1af00b123070b9431fcdb0182fc502a2726f9a837943ebc017d942dca224036118e47f7833ff8e67af216a26210c2cde2c6af3b0cd1833cd5bb06febaebed4c1ebfa138bc1a69adfcd1ceb6544d1ee040d9c68e9f7f0d982b6de8391d7bc89df2ccbf4e2581bd9f0e58f2677f41f72f042ebc32aa1ab8d34b4f851812fd503ad012991ad7cc43c79d8859371ce06dd28918b76c24f3fb9207971e58b7d10e6498984a75679f4963415479691f13cb00c41268d5e5719eef46d0e4dcbf057b6b82cd4e4a084f2104e6b87bc88855e34c2d35a222f357828410a0a9d0540e22682dcdc8e5d573527e221da25e66aeede080343a2381f884d8724296caaaaedca3e6b7448285707b4b42a11708683e1cc98c33b0b64b5bfe3a6bd9468a76895871ae8d9b95a0649250e88f41514c527ac65a16ef0dec019e85978e25711fd3aa1e83210991feb69d7ffaa3cdb9989834e938d5f1bc1c4f9348db0bfca4743dbcae196990d903955deb4d5bee0bb185b0a1c83f245496940b654569cd9b756f7ff68cb2d36588f77765c8262a423b34a46741678e7e636625c3517c8c8c22fe04994fbf818deca1b157e9dc67e4e4026c79230dfef7a71a3100a03cf884b284b380380417716f700b5a2228145feac6d70795cac8a9410fcefbf2abb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h4900afa5078531982600ef0651745b746144694d75271ac757618e6cc363a02829e3e071de21d886556819991649d79edbc6ae964f2d84a0a5141dfcde0ae8ca289c0719bd2fb319ccf677e9b131ff5db1653978cab5e72d5168b9874fe329a44c23be48ed3b3e571d1c347bca39972d0fe6270169592059194928ca6322fb5e80d600c95b538e855da515f0836526ac050d6a28329fe4fad7cdd5a07fb04683d567c555d04a49795670b549f8451a3153b74dd9c6d03644abf924160505501c2ff6ee03a0f123ae17c13d6643d89f71a4481418426c153ac283a81c10a63135531042c903f0579fecff0cee8918fb1234ee56c34b3f9463d8c147973efceda33757a1558c38da93d8081d43b1fd2e8867ae1406260ae4ce73f3a67ae28b4f361df2848ddf02f14b26517fea0b0c9043109d0fa2bc15b72fdb23ceba6b4d848f3fe12b79676a6404aa7c9c8204f0bebfe5ada62e1343ec46159c9bf1c36aa55394bc9cd37a9f2c1c8593250d923c67993e769a15da43f032ad8e8fa8702be91bd84bf26af6f194664610c796d5d3f5d2c50e72fb17f31273188827bdfbf7f9597e2e97d25236e56be51f3770ebac4c8aafdea61a3a418fff6d102f144983abb53fcc5ede3006d3817e3fbcd4383bd12c3481570f733e0287336a0790f320104a845a657e96e4f4f777cd38598af3f2d146d0ff187994da744c66775052e4e9325dca83598be91aa870a5fb91eeb8455e6cfeafe83d5097bf3b43016b7f000d8ce03bd10202468d542e2f337af141fb546fb2a8de1e39363b6b5b9fce32e2d4abc2b4e19a974f8b47d8c914d037828ea561e1dd66c88a159fbefea637bb34d9303b2c91e64fa0da7c63e7f72c4a20c7b2659087b87ef07727de99b279e86091531483d5e7a6540c7fc791fd138888bddc2cde3e607a70be0f86d65419aded1abd7a21bdf3749826ee706e22b3506e2c4ffa883e2a21d0e37088ad8ad30682f41b468ce1315f7240c37c649482eb34176061ece152494f77901000e781f7a61b676856b636ae839cfb2b9b7632a35a858c84f71c8a76647db665eda6b7664b6ff3287e2abefbe69514e5661c3dcc4aee140f1a84bba3d6379b81b74ae443929f2d651fa9625ebc4227a0e1a2d008c5c22e764eaa4f21f153fad8845ac9af91973729705ea4ef0bb35aba23e7bd535e8da369ffd1cae9b4da1260c1b3288ed0b8e0f35961cd2fba1986e5e15185661f996917fa6e20c95d486073985ddab5c1f9a6ac7297fa814b421cf824244e86b964d259458d96b115daa64fd70ef8b3befa18356013d3da738efabea9c246904c93510cc4ba83e898bdaa4b071bc23f6a119c892380ca2c97b0fa36d6ea3b2e4bbda82dfb25d7d3e3dc9a1c52694c6257a941fd196566ebb22fc656db63273d0373fea0c9ace37b4f6fbd179e799dba16bfde0fd375254cfe6d1714490780e511f58dd52ac3e4c04d1fca585962551e2a03a11abc5932e189de8556577fcd1858d0cf42dc17a83356d371d026153bb0937f25783a20033f81e76beb5c207c7229effbdbc4d097016decf55b78f1b0d17215c9d80f4cf171335289273eb8fb5f2eb614e7c7123895f43631be9c617db6e53ad388883085cfe86dc8358dd0b388722b7f3b5ec24485e1bd142ae70a4eb754efd7a87f6a9cd7b218b562ee7a5c0a24d67061f0192e06218396ad4e9529159642e9b9f43263e3ff39697425ae8451d71f1f7bcea43010eb4bfc34fa239f69b6210b7a3ada5e2661c3d6bb5fa48fe791af0186cefc89ee83ad3c30a9af640069462e0c62b33d9ace4de8ce2835ab8317a18444d713584576b45b2196354ddcc4da4b34f4ccc644fe33a36eaf8e4ece6ead1c652834b738e47c752e064f415292905b9031610367c4e31b325092a70e78740178291ce36b27ec30add79185ce8b2ba36b641772915d1b06f3c21c9799e645fb719142fa32e6111652afcabcafd98554285f94f7ae2379c0d16c8ef80794886c6463f1c9145a7dc54950655a3e10516cfcb4e4cac01bd53d9c629aa8c063c5c1206311818bb6ad309d7fde82f6e9aac912d88a2cf35fe882322d41ba2f9117363841c9c29af739b9c1daeb2922dc622677006f679b45c514bd7be725321f000409374588f0568b6871ed9efd74ef86035a58aa5b0907dd96aac36b3dd173958175f9c866bb1ad0d82c5aceb2b90cda09c8f81bdc565ed8d4306604acd742aa72aaaabdbcfed15ae9b96d30fb9c836bcb7ca92d5609bdc29dc3d6d536ad83c7a46b2c9f84442486b03d1a584a122a4787d62a239d15fd57dee85a752f5b3aa6d2a34d02d8de21859c0d7acbdd30c21c13d7b7809e344b00cfc1f83a3bfadb3299dc119c28df4a9251833a352e15bf80d41a9ca81b1303734f964968bde84bd73b4e5d01805e0aeaa034268f40e21d1887bcc2a0e981f51903b30f2b0aba77c4bd686689b0ccaa99cab65b2412c65d2f6f4fc03be88305233b4d6818bfc91b94047f45a91c7bdeb1f4aad9e9a7d1e5f972ebd9c27fee175127a67b0b4adef9c446f10842dce151a01a6e5fd7f80056cc8e2d92e506c71cd3bd3ca0e753f16eeddbf6ecdc84c8274a09342cf2335c8397e83578fe0bef47a1cb434dfd89ab56532a1d24fc3831d7444f86aeb67ed7cde9bde86dbd4def9fe4d73f78a6065dffd237bb34bd3304e8628199a7494fe642cc4574c795b6060778e6276746b843c95707b54a197d81084d43c9e21364fd07829dbb1c681ad209a55e19f5fd9256522685cd84ba438d95cd7418b838dedadc00beecfeeb4d9d7af2634758426e4f3a9eaebca3b093144cb33d57c2be1cff9167b523c2513e52f4eb47b88fffa900dacf0b3c0fa32dba139ee7b086c4d94b2d4ebc88647bcf3f93d72b8d5b0c7784f9dd3c59cd150c4a3dc1543ec91511bf135a65f5039cdfe926bac223442a9cf4a89be076b56c3d70a24208ce546d0f7f32272c7aae015a5d8fd7a42adc9f9a8d2a401717b47fe6af2798754b4cde807908c0f9745ee3cdcb14958f31a2b2da2e0b1a5b1f14af59eac82bdfd910adcb0641050394b5be95ec511e43ba668e0891a1aa4de05f73e27401108cc854895d8d353d5c0e718c7a94b15944dea5915e89b88e6d4b35ceebd4e17ce56b85a5cc3ac1775369dee06a6e4507cf9709a6fb496ba3457899f37f310321bfdeafd9cf04384d91fa4bc7f9714b47171beb85a159d7b5a0e5f24f812ef197babdb0a08024d6c51c4ec0ea421dbf0281583fa1dfbdc6796910886de90b24436af3abadffab79e5417d7e0085435c6bbc2d2716a1da3bd62080ec777f78cfad1a22d0f5d3d2e17555b7880f2e3dc6f0f35243d64bf5680cacfccc269a156f3bb458e61b7e84267bdf76620c9d0eb52d5d6f4476acc0e36275e0c0e48dd7e8aed463be5cc8a81ba6fca6e179621b0d01a5fe5afe087b2f88e9760f27d4a5ace2487ae72e30bc0f938f1c6fec70227f4db07afc97ae777e7c8281064a35833b472f05963305206883baf2ffd1c379eadf31ac06af490cf8447a73b9cc7679568b70e50bb8e8a9d45b62d292215d1c2fda14e353054b0dcdaeb092e4266b3711718922cabbbf3c9f792fbc073176feeab7c58d7f90cd0681394aa75d961662e079459ce8f7a0390f57bff9a9f57bc44384260883e813f25774d3205e4babde994554c7a7f3e1227b61751248a26c1fb41d6d010ad62e3d3a914f8194ec778acc9fdba59b9f1b3f8a1348155c813e320f607272d004900488a448439f790ec1171f8332e06954a5936c691fb84f1539019e303dacb738d50974ee42203d2ebd4e1933659e5a24e70b046610b334eadbbe66d592a4e22748f77a8b51b5b77ba1f66657c1da87eed81a7dd373a67c74c83bf5543434090d846fd5c5bce65c35f2594828741cc4609303e14255caa0d350859c60abee898ec72943cba27073e7a96e5a8090934d95f7c609a65781025bc526faec79a07d3fd076bc487e23661732f27d8de1ae56c9850585607fe0a2e966562e6c601780b5a17337a59ef4c932a2c52710e727ef28f0976c44edbf5f8032acfa839006360ed614c912d1bc8b947f2e9acd58c710a0b16db875bdb70c5b455c122019b442ae739a1cc2fe02b4d2560451e61d27c996064efe7643d743a671c176a646be080b5d5ab90a0b66461fb023bc2d8510598e7e42ba4427afc6ca77b6ece799e2408cf05cb60b3c56cb761bc988e325afcca9455deb006e20da1c31c2bab5aa39a0e0e6d435d80dd48dec9036121e804ae4f9f493361cd34344e9f2ac19e0e2c41c82d902bfc26d8ead2e4e8478ba9fc92f37f18fc628ff7eafd2dd0aae0f5b59dff18c8177bfceb9e008242d7782dce8ca36c0cedefd440cbfb258d96c7528921d5cc7aadaa3f0a0a5161d60bb48e9752d503acef60659de6601681d7547d41db8a0eb792165a376a8adbeaf35f445f4901a657e396c7bf8fe51ae498e6b3322b120aa8051e78fafe99a074edbc73eb457dc64bf101176ede99aedd621b09c1b9057dfbd63a74b4d46e9968b67639c1ac7683d128c3aa9994047a52174c85e5fe63609f9aac45858873c5f1a81f770f5a7e74587a16ecac911a2716c1d0751e3673559ffb2e08b40f0e69e6e1f974be575352207d90ba1bfdf4207fc24ea59d4c0d9f358a8fce84a2a3ec2436aaf02436c25d7c0f3d25f0a90a0c455c42d95ec970987cd42e80f7b7091aeeb98ff3fb11f0f222927b926ec02e2f2c22ade9412d9fa833c5ff72247b7edfb60f3e496e4a82fc91cb6fabf92c644fdd0d1f4121f85a129d99f5ca839791f4f967d994ca385a2c120464d22a2639bb955ed0cef29b2acb2b024d92378b86cb05d9325cd63cde19d800b890b6829864967fd31759356a9e1cfbebd7f68f1b278007742035238ccd972031e6faea5509e3c275a9d4498e09e81a63aa10ad1834a1de22faeb9adda2814484d10aa13a52e74c7bb56a4fc917058f8f27325ad539f0bf77dd43c691559b447f4f919c3dffffa9dfe4d6d6a09032270e45806db2c65137a5aec5a03e5161ae94f3470d3fd52722f04d64a9d2910eaa847723b164e6118b9ef87f239d12de648f49f8789b6d4d8e498ba257c5588ae77d6f66e322ef7db80dc2c92b0333df090a4fd752f55b2babbb89676c21d38a94e4e54957ed0a48f515ae39f33f87ce079b951d6e466bd99767aed73cc9ae81198f243622315f63af975c6a2d678b21a118177cd90da5623c778f4186967a953f936d6574fad76b40668f49a859dd30c7443947f51295018f0fed3ef273c3074f55c54782f56f929ab78734c938a8e553c07bf4cc48f5bde28ad496aef480fcc438af57e881e455ed3d709f9fff6b2e00f4869ad5d1f4e959354a1f8c1ab272fd8e444e5d09bde7f7f31cb30ff40aa66b1aa28cb75c6f53cf1c499860d05f493b0dbe979d4e8b789df09bd2820ed414d362e02f558f665938027e1c78a2cb4aa5857;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h72196ce7ee2b984b65ce528fd7343c9cd1cc8cc54ee01277fe79503cbc9aa91ee72dcab48355c3b753dfb90ca8da05229e0d0db6bf185f505ed0e1ebeecd3894766f43462db47b417dc396b71185306c81ce6b86187bf31440f35c57b139d2744d242c703ceaea93e729fe7b3bb6ca78d83bc46eca72c47b371b5dcbf9aacaaa358b363a8c71e0083a226d96a271184632202d90a2aa6a8e4d6cff78c45049eac32f5428accfe23ba101a1fd0d29ba3e3d99977dce0845a0e3c0c219bcc3e49c81cf01d082176b28497fbbc7eb2687e00f267080297becd7c4de04d4ec649c3005a95370343d464eacddbe6039da0149a08d4b6ea0285f57e3cb5ecf62c0aef9cb69939686ba00ec837a317750815d469c8548678e2bd47250a3344ae1a4b5abe29aa4ed188ad93a0fd1e7c21359e9a225931c78ae44dff0e4465aeff3879956b9844764ae0887d56c5dbcca74b1c740375fb1185bfe6f1e94550e2e410ef3f88de2ce69cf6bec7ba3d9c5a782bc5e6f26a6a6da155c3091a2f47a4d133dddaf5ffb7992bcc66de75b8cd5aa9c9877a996f80fadf84425868b7d880483fc4528c4cfe105979e5fe94c22d32d87b72491c78320d9ec760a32eb02214664fe68952caa69e3a5ce9c382d90fa7334d8707493601e5ff6e8c84f0f94ca1918dfa0df4725ef4e0f8baf8a91a33a0aeb6bdfce087bbf93038e4a570a179be5d6a7609e27a50468fdfc68a70ebff2f5273cb5ed283d7b425f1cf58c94da6eb1bea761a954a9a96542db509a7e45d98e6b41e1962fb5c21206c6c2ae993c6fb08de0f6dd208754d7397c91a8aa480d96983b8cf097f68511c1bd414b7ebb27f1b421f8ac692657d8c09a859626ed7dce78827f466a78851dac71e509c00e5ce75ab3091ae64456993860ac10acc99f4d2dd62b54caeb45afe9c5932734610a436abbbe2b4762bad966066499709313502f9cdaa9dc1717f2ac9d169e25a249cb6fc78d6c08cd7f2013a276c5ed73fb00a93658e2b5190328a66a0fee87c361f4e7a37f3b4c41ba1e24787ee775435fbb6ee1e9d463361c5df00176bf65f0aecc8fa26dfa7a1a85ef0131875c3bcb645c0b89e45779b2c1cbb1e9284f7889578de0c82fa86ce6693ccd2291588302ebeb74139732d1d21c6688df18ef6fdc068fffd37a4e04c198d76780916b29764d2a4818a2fa04303dbd2441523f211b64c00f78e2d30874823a29b0d34df6f823115e79fda32a8720485107bf18b5c3f9e9449f89cfed11ac9c29c15e8494108e07af812168428fc3f4a958de76b8e48618974b6f8ab38f507e83f02b18e8d10311371ec6f434a52c5349221dfe0dbc958568f0e578c11277feff15c6c465df0251d20a13519b44f8312c42669655499c6565e281872b6b8063f06611c1c05a9dd2316d1d414a90b0b5bd838f516eeccade1146d06cafc980668eaa039fb50351fbcd34351dd7bef991b38c3286a677bb3fbf6661d63e963b416f6eddac8ea3fd197c7b64129602af66394f23e88749c5ea875dc76e37ce92a04d9cb4c35c577587fade2a0d4fe8d5fb91ce3a07e823306a81d476a36befc9e65c0cb345b32e2c1dfc4d67a9d232a1b6f1784e918a3d132ca63e859dc71b9dd14698ff5879b664a7222f99928e8702f4b71cee64092cdc37867eb59d8534cd33418068e183da6952df29e423b3d3529b013e9f6f86f7ba7f552af4519e190bb50e5700fe04e4323e954326a09c978f96361bf15f1095d4b750c8b9e076da6bf075390853c7550ba5f17073ab90656d6c05ffa6b3cd26ac73c6f2095579c5f09a6fa1f2920091fadfbabd81ee2fdd1c124ec8b12eb9899c6318d1d420ed764a26f86380a8187d605b2b408fe9a8ce7c602c87d0f7e58749016e54dbffc2476d393d9853c5d056168e7fcac1bb15828d194c497827aba76cdd1ee5fa2ce5353d616569eee3e9e488912a7d38061f67d2c3408983373ff91fd4274d5f1c334689ea650d5240a4d5ce131becd4ac68ae1bd45c54fc4fe0aa2bdb03e4a17dc723d1e1b594d0aa7adab804d570614374f3d44f4cb58591e743cd865d20ea9b308cbf1f5b67838fe7027b2dbe51f9f53a1b8a8a58c521d48ba97f9b72ba692a5c6f2d3dd95176545e1d44f09d868af40620dab2ee8a3b1220ab8297886b605d523bf188420e8a1d13b936fbff88c992fc630c62013b8e872c487852c5ee3fea800781b124890a33ff8d73fa308d41c0667a8c624a3a6984826388de90ff41cca5294a952a17a4a37de5a8e307be798deadce371898c824f38b63f2abe1bf58ad76374db0bbfcb477629be90259ae4e95ac5a96504b256e0c3191acce227943a1651cce192caa12699735c44a30ee4c3f0d1eaf8e3d30486af92ac159ae99edf790f9b1c310e9abfc81b982f5ac58f0964593d647b45b02b871604e831ecae2c3ece5f41a53e1bce9c3efe563dbc8c7395fb1b6be399e965ec1533654f6374dd73282c324b81361a17c35cae55beb643a78d98f5202693c37b45b27c93ef97db65d54550a1db799e952edc8769f031cc801ea35b30b7c1094e3d5741ecf30a3e79adf18f28682036de197ab61332273c1cf0b83f7d71d091ce24dccaf32f64ad49a3d4c431f3a8ba1070311eef211be83a0f66e214bb82805c961c74a359f8c7645b884db2967ce552c92c15a61d4474d2cd92bc38b5baf37b26a98671a47bbd983bd7a1c90b6e6756c3d11e067cceafa7bf26acd280d12ef0f1d048fdab11bdc495d1e1e24e339057e8fdf71dcf8edf74cf652d1ef883d96cc0590959fa7ee0ac02926dcfe7eb8a90fc952e2c7841a64b59a15667d7be70ef75596cb470bdfd6a19c98aa4b8d5bc4b27476c788e394d8a432f2ded9ce0bddd96bb91b78643f9eb5d8801261c814a290bbb31dc899ee24661c0f3cf755a5a2d709a0734c6d33b16f2103638ab939fbfb3fe3423cec9539362c29ad1506e9546bccfbd46ef53d3134bed4d8a5ace0cf709bbdca1517cd9cc6ce1a994956887ac7c02c114dd12a1c878f92cb8da0c4e9114049ef6ae426dd54d48d2a1bde7e9ffcab269a8efc212e96466f39f789c58208dc82ab59725f43cd7af702b6dfcb0069b8db6014c13e995ce7647b39e4f9c20d9b0ad6ce67af46a4a3d84c8f31e2ba3a59aea9858e28bcb33ab0dc179b1ba2aa2e027b079fd908fff9db71e214d788215ad7d7497f6803bb44e49b7c8bc12355244f95fc8936e715ce9b957aef6d6a7a32bb298181f2a5b72a0fbd0e5f6e81c0420fb569817171422d49686f56e5c2b11ef9dda9e42cb337113fec26623656e10d94e26f5ff35051ec1c771551a5d66092ba1bc5df078659565342ed561b5b3cedec0895a86008944ef860ea8a397069c884f76a89a08abb39527328502399f2c61cafae450018005fa10dd524a5fcbeef6e03825b336cf49f260647dbedc42e37fde6ecd7bb9dea9134e2475f67d77682ac412e1f32b46a8ca14b6dd72b8719e81ca53ad253839344205de564f5f3fd13def852bde8b0e2a7027e1559f6c5d6646aa59211915e8b8920bd383dd7ffd3fd8f41d0a3fda6d5ae4f478a0f02093a3ad95382f55e94e9b36ed6b673d76ea03e8107043879ea96edcd0eab733aeb0b36c585d47bbc4fbc6f2976d98eb81382f30e4bc64d05f06ac365af77072dc70b0c7cc57e5e3501f072d34c8e989d8ff3ab7aae0a129aa95c451a56a5178f08e211ff9f1cd12cf4c0c3e83c2d3570f554d92cdcd62678699332802175c2c492ac8f82a84ee7efe33ca4c03ae605802ea575268a78ada51d800e64be24bbf4af056fa1116a93606d9fbae45ab924bbdbf7f1b21313fda1c3ec548477c942b879eb6c295c9fd7740f029c01fe4756b9b356b97ddae7c9ab4d6a8a684f7c393658da674cfa8d79cbde48befbc9e739649e1abd2271d703a183451bc7badbccf437ccd234c33c567ff7a4e9fa55535a6f5b764d32bf07e98742a9d807c063bd414a316c7b8b2f29786fb79618359ee4837109e9fa21af0c2e2e209c52a44c09d8bd40b0c773db3bad904487dda4ad5efa12af6568b0e51284ffcf026db8468b331a05d678ac0162099c6080c5a39e6cd2eb79039c2892360459858a72d51d85011f4afac002d7d7af9f2d4e63a65f036b79980318358428c8253493f24dd06421686dc25dabf5db3f31a07bc338cb9fd36d1621c587dab9dd738fa8eda4f83fa8f3ab8bd40dfe8c06d461b8519af500f019e15d2a784222f3679c572ad1021539a0c9b0f014e3ffb1dbe7c49da56425213489971c3ac74c82f0928a8667c329d4a1cf76a8fda1276dc1d9127313988fda2c7dd57e63c3f0921141049f2d8ca76f0369fe938d6c1f7e11ca693acb22a0734d9bf68c94b21d2c048b926a8853a8945b4ada11c313377453191aad03d6b992f35e275bf8122092a30e23fcf2c31af73ff4b1b03678d09f81471954228ca4827ea5173ac81b90faa606e4a4167688b2668c2e0a19973cfc6a28995fc34dfd1bc4db6d2637f85879151032896cede835761fb54bcad33a18828a43746dae58d608b4ac3d2fac5d5a096f71ce7b3c3c62c6644a84ecc26a3dd85bfecfbfcb318f69f3f26c8444735d0332b146140df069c61469a5806376f9b1e836f74e9995741e7517133c1fbde85da163b52d59dccd6a6b1ec1ba0fdfdb5e2eba5fdb9db6b16df0d6d05e08315c5163a91a1e22c86f111c08e5bc111543f20708cb25928feb2efc5985772cdb2b6542f15f7639e903e267c14bf6e1d6115db7ac3b4e0a5c3cb8012c24cbceb3f6b8e0047c38f5f2f8ae82ee406b8ee5803d2fac3364d62fd51ba4b2b519ae271e32f00629c51de723552b74f5e9368cee2a7fac2d9c5e27da17643cb9d1cbb3188b2c20d633826dc0a56e9adad59ae7a08afcb8bc93dca2d8f479c6a449dc7a3e549d5565a41775b7a752380e258bddc24b87e1723c49b6ba6139836c01c4e6e5bd81c1a6ab287af4a70abe8e351d7f827f970810db7045c11fccc12a55bdb2466685cecd65e43132fd62195f19d3af82cfc9dc48bc851e2915cad73e988f7e2eb12de0c7eb4d7349a71bc7bf805932f3674e7ff48c8a44c5b7764e83f5e250c6f2486424523ced5795bfdf4e2721bc8c25b606cf9649a62e9ed09831294151e3994f12805b6ada122b24b0d0522692d24b5152896ec92f5b61fd056408a69c035b8a433bcf7739984195705b09b69be4618a7b3440462b7a80f552fcc01fe4b82b51cb4671746d91af8f723724c61cc524e6c17cc06b10ef96b21895b4a1fe2940ac44b893c0075ffbf8ea0a979390477eff2cca26094e9dcbd785d0c3968db3c4dd559189d5bcde43c5bfba797e8f6c5cad61a770231d878ffeee1e57295ec5bf0b6ce72c06914af0f073427b694a12a20aa1f851d8d64eaa3eb7fa24d7b2912ea2194df74a745ec4e89e6520d061c786cad3e9be58b46ca42b0234eb8ab9f4a444fa5ae6ef38a8406f9402b246e80e5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3161c8a969d36d7682d795ea9e391fb82fc235f17035c27d82b7f6ffcbfbcbe8a531428d93880dd0bdec43ab89230cca4b9d5dcc046be0145e75a0242baad1567aaccb8dec9e9b0d09a1706328730f2623037c1e320ab2e08ae2539294038afaeb63e2e77240808ba9c631afc2b23bf7facbcdcab5143f9691bc396a87ceaea568530395466f6898e9fd2faca2b6321722359f3d9a15152da99e85bdfb5be9a8be175f704bf586ce8db42611f2c89ab63e1675340f82d826e7feec465e2e295831a63b11916ea4bad31ef8802d4a22fd49511947d8ab84db7fd9264b238b9e14a34170ea7bd3c65a15a16dbaa300b47995d39d00c90ee62ee8adae75181c7db753453d9ef0398242ae5813731b783e519ac70f95c1a3f134e19bef68b5812f6e6866674dba44b62f5d76793c9547510a806206a3f0cfa7961edb7031ef1ee068a708c15e8eb2d4c6825b85f4e44d3ca3488ae650dfcc594f3e469a7a2c019063f988097d025482944553932a1d05922f4322d2eb85ef21e86aeb6c5834423f4329b411e70a5ea4296671e6bfa1a78e87ecc2a0faa01c7b5cc500e57796606883934d3b82022f7916f82f5b3763f49f19ec85283080050ab4766ffdcd5aba513d9e76fb947f6fe43ac83cbe1132377aeaf25d125d50843ac22aa1646ac69dba37764e0a4db9b8dfc459cb1b7782bac699f8c8d7eec8d09145d158a76221aaaa1bf54e45c63ec1ef4d5619e42cdc70877e7952dcfabc29b8f36eae380c46a3bd727d433348e50fd878d3e7424bbc7b7359bbcbc7e0d3e1e0b384e5140eea0a584f422074a20a1267fca7e5db1daa2963bfaa01df2937a39b3bc3d99d4187ccc91d8051e2f7dd9f81ae625c3c27fa54b9711ff9b4a87bb64189bc27ed06cd35fd5697b6e527f9f992b5464d65ec78d3b9f7b9ba4504894e2d73ae28b3fb29def3b403ef5beb2b224629db59ebd501d9ffe5247aa78651ee9e9225cbc638a4cbd7ad171d0cbb654224e291a2e8912b78eea162d6a3f5380f56e35ba7d70b248ead6ee08644a60c72a1ce3b80975c4edc62feb5c8f8f97b214d2badc2f77c3148fb841c1e6880bdaf2015137646930c8b759eb65bd8b6fd242f9b4653f75dbb9805abafebcace2f16cda848e8371838986340baf06aed25c1784bf2f50ff88035f27b81213f3e9ef3bb99c6e0b89951bf8e7b67d1fbf26c70bd5bf2a39884b6e43c5927ba524f5bc012be32f415741c3d6b1d8b7e80d0bf4de2dd08c8dc5a49c5995d2fd8beb289929f02208ac71fdc52902c4e1b8e6b330012486b2881d7b3a8f06db3eb300273cb08c918f7c89db17aa7e16aa6743e44cb37d0f5a43a8eb63f037199ea9e6758ddccaebf55cf40b35acdc2a591194d481bab885bdab24dd0f6a6c4043fb951a2946ed0a5c2862ecfc75f33871927d0d32ada96f04e482563daa16e54189478477c918e06edad109ef7bf0f2e02f76f4ac6f6073427a4b68dc0d1d213a7b7002a8807b0953b69311e6af1f2b3b9d238e5a5a1e216d2b7780cdc37d274a56bd3fef3c6e2de6e4f800458f5c8f42849af07fa57bba50f9bd4c02924de903697699817e45d0b026d621e3eb57608a140ef849d80421224d923f472eb16402fc32b5eece8a6b5d321335ecbbb356f9f71f193b11d6ae290dd17e40bac609630f206f7c4b2cd57cb4f861b4e7fd10a960726822b770bc2d224c9eca760ce08fe98ececf11cc8ae786c860cb292c5696e7f50da43317e27510c82ec4c152d36ec4ae90512b9d4d185c795a08e8040bd8b59d21899bdb11ae5269dcb393b4d2585d36847978d73f721984a09ea19d353ddbe6b8220a0f2132e3587ed9898cb11b5f1add563093fb92915cae5fdc6f0f1384363277ce7366b50c339a18b17f38510f28bdcf60c8360ee69ab270b050e1651409102eba8a3a9efd1993487b435b7d9f0071ca678066da36e25c3615fb4c7fcff57ba8a97546e8445640c335ec84f146c8cc2fc5a602715fc8c88e0216903031af7846cfd4c9294e3f1e44c49021f58e68e8a7456158a604485b4b6c906f5082a0a14aa72dadcc3e34b4cb6bd1cef42ef85bf7c0464f223276b2e52b8097689830c2bad66730266cfeb7d877f02d0650bcf12445b4fb01d5234981ccbe3dd72eb8e560442c3c1dd43bd694c2a6f7478d3d80c7e59072ef9e74c34eb02c4b559984c0f0478caebe30b7a364698affb795b1e38f181dbce314cecdf5a943b530fba2ac65c0ad41d7b244b84b152bfb9701675650b65f9a52c6a8268666a1adb0377e4a2283c22d503a18cc9a8c73748b3e8aa8cec06f3a5a5e361819c4521fce3c03f0ef338a71a8e1277f2bfcb58bb1965d548b846ba5688667f60e34ca5f4ba2eaa72cc246e39c653d6f95d1d0dbb180734ddd8c33ff58578c142e57b55c4d50cafa799f55bd7bdc599d81ddf52cd2b0da351b322516aa0bf2ad702d6ca1a02588dc180e3b62f80ff6ad5ff574c16cf80876587190858d601ca7df7e6a399e398c8b9ac12e7aaebff972028dbc5eb207f98ee7c2530477aa5de726d08b8ba668d9ee016b514fa38634ece3d5be465f78c496502d9f4658b7c56ed0d16526e8e3d9f300e4770dfc7cc70b8da298a2e5e00b3c7ae4fa3945ebea1890e66b73e3264035f6590c224df81e7fbe23afeecbec39ba850c3fc7cc0aa23b4106d708ac7f99eea631f18b638cbc584466e59d182ab8eedf9329093f5a39beac662e1460f22a87a4c39a5a635f677b200b8e221cdcb8be6dd230074072db175fefab0738fbf811e6b25252f8617a0ed9e1473b898fd804b4801842062c946876293384c2c9deebc7079ab2f7acae6088f713a5677b4dae5f002e09e47edc2fce159d5e99f35d3a3418943214298a9e0f486bd1fde72410bdfd023b452534b534f9b02915c6c3c5c7e801531e15d301aeab560d41ec23b55845795bb782ff446f8916b5225ae7af82baaa891a9ede20c4724d4def7773fe761e198e5538e90c2c284f43e1d5531805ea2aa8bfc0631ea93e7978ffae964573c4e14e98b8e0b8267a750e34a4695dcbe9cc4e0e908dff73ef2734d0b761daeaf42a7ba348b98394a89b8ec825c60e5667f0b3726f514e68254888d83d5a3492fb8a6c5e87f828c2b05e7a2d65843f92e0088bc3e74a8a5eefe7dbe4306c63d3a29eee996c4e9b902460f8dd9b5792e61685be3f4f7b8838bcd59ed499caf9e865d98303ee852631082ea879c87aaa0927f146da9ade2a61e7f0d081dd0ffdbfa9d6080b31c21857d134c2e3d30db41e3fd07f421adfe08a455240160360b522509dd67102125167a4a10f92846b9f5148dc0da5c180931db039eca1edb169c16fc0f9714aa6f9e1c697714232cfa405c46f6f117c74aa7be86c7a82b871e6625fe263992255c1858115ae0f9541738aa08997ac3a00eccecafbd6e21cac672a71e1d532f3e989b0c82084fb9cef0bfd97498199aa6ceeb3b886c808ff728563b1cc3436ce1044712b94bf96f51b0f48b429e580443755b2dfbcb6298c56b6b4d1e7da2cdc5e5f1a77be4c9e13fe92c9205e5f16ee1378a1efb68fc7ff2c772abd9dd1249d4caf3e4ae5365375b782964f0985a52c9470e6d3aece62af91e87b5b7e7e6b37b2fabea26a7c985658b07e1d7550a25c053f5464e399fc8f9fba0ef413f1750128f5772601c54d51bee93954eccabba14142a2cd8fe37c3ee28b5704d047e93f82f716ba7ecf3429e41600195900ab6d6bce7232d7358dfc16fe6b571c2127ce58eeb3795767f377d34ba1b77da60c85da286bf0462fc1ef49c189b30a38b604f3a0d367fc316aa1780fddaca2ee6739bb5f2eac92f928e9ae3ab0ce9be079a1041c56897a6f36d985222d77e2067388520d545f6400ae0931f9350c512672ef8a0e4186018759781da9eaca54e538ade16ed1661e9979ac50ec56dc109a3afa935e2f29a85f0c72f4fbfd67c92b9ec47062bd4099e91ce8223f25df18fc3cdb0add991cafc9f89fdac9df5e519720dbd3f8255666d684bc270ad38311db44c6e15d7270289b57c6178da7ef1641fb41a5cad99ebb237f7542b9fed635a9fe2c9af75f1ed2063a94e5d2fe78b59448f84878cb85b818bddfc849b7760776b274c495068cd1ab205a475aa8816e023f984ebcd7bd3d40a099fcbd958fd58bbc257685cffe2025289e00753353d854c62d4b1b82c6dee4f590c40dc824e54835fa333f8382dac3f918f15bc10d4401091f147037c37d6260c558585e56011a2eef4568d641eb5ff56f316102e01551fe2b2e4f18e7c977c0e6377a06f0b8c6dca5019827c0dd9d3ef4dd4802a9593867cf942cbd4cd09a5450cfd247e2ef49eae8b36faf0bcba8f2df040769710f65c6b63a0f0db822bc9747d6b3b65782ee79e98296125749de08fb9e69496e599c9937d246758d4ad85d043573d866108dc02b910858d8d4a0de95528dff48ad1e3fe75aaa830c164d577f9cc1d88e8f1cc5308189dba756b25eacf6813d67104b3a9044602180978005308aa11d565d74ca3a25d3c93698c464b37dfacadc9fe67b20466fcf44dbf740194b9e0a23df4200cdab8292555a276c7bf42865ecb35a4bcc9ab69d47641ca60f1edf631b8b9a0d386110bf0b79a940877c3c6a1f73abd65f8111801cbb0eb65beb6605df0a8ede87249c6ff6bb79c3509baea732b7f021e1feeb3c8cf198a58ed5433e5a9043c0448bca23afaf7317bdaabe21ad29e95aeb255d882eacd529ef8c97ea3f73136e4a7d4827b600da29562196aebd8340c1655dc776edf06972cf88825c3c63b32b9015e5fcc1dec6ce3b4c18ad8bc65b8120df089874ba0e428de855b922d516354c228eff121b9b70cb44f79eac624f75c7cd5b161bc8ad30a277c01ad26e5e47a2a96ceab93e7cd448ba48a3508b99df1e1bb50d6adf3eefd5b0bf91df17a5073080e8eb0eb105c3246e9cae1729abad3ca5bc644cadeb88932d6d468583373ccdae2b65f969e54db72b9b56e2058d73ac07876e497f5312b202bd833481e2b75778fe24d5996d1f60b27784bc7266430aa69c195a2d07b14ca3286a3b7628585cb3fb6b1f9c7b5caa265c371a94b27fcd463ee37991e8549528a97430833f288782308aa5a36a401d3a63d4b083c4456f3ac90b38f5ca40735ed2a309684c158e3dbb300344b65053eb4019f8de9af5828d4d8ed2096f1681c4518974989694692d78d6746c6cec9fda7a6bf085458e80e6f156928673e19d490d8d99cfddb7bff9014602e7b8680a8daf1a5eb6059ea9246496eeb7ec5908cd966e832845a2ac69586575b8dd7ca2371cec889e222caa08d2b18d2008efe650061586ce553e9a293a7eb16132cbedf5d21831e22bca24791e546559966ee91184688d824121807c5e0e4a07c36b5b9d35aca42ba5ff70c462605fe002b4c03a2416b846e06638f0b6edbf0ca31a79033e61d61315e4d07932b48deed0bc0b1275b29c8a22bd1593cfc972de0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h868c4977e2c5c8a2e7bdfd33d7fe068bb2a1c96efe8cd87673a925184c3da9d7f2cdbde6f679c58aaba683dbf19c70c189dc73e861c3291b737cc81505d485b93d385b608f410abe6abf992b32cbc685e094c3a5de2c775f405d6557efecce85e5a8b90066e2ee06e91e4092045dab4cdb61faf270b28ddbbc143b187c678c1b5540b3bc36e18b2b3ef9bf6d5414f9aed8eda1442ece72f16b28354e4739d8b4b5711e06b7b3b36cf12d1396c0a70caed1aac7be3fe3754eb41a60bdf5f79204c7644c08d40277d76372c14eaa5275147fdda019b975101ac6405477babae53eb231a71f5e5fdc1cb140f42a37c5d09221afeb9c5512b1c40f54a0cf26f0184655270eb2309b72fe33139ad52e06b535989a36decf4395e4f50185606c4a333793040243e7e99a2eddf19cfdcca7032e6e8e5b122a28d52e05bad8cd880c4d2a9b7fed1d8572e946496ffd5fb9d66f5d06f8e76ba9eedd08b03eec05c5e883278bae9d77dfc4c794ddfd656a1d447c5908e5ee8eb393a87ba29aafd07555d9532a2b6837b5c85dbdded597d3b18480d86429195d62562d90a341d25125c1e2080ce4ec23b07fa852df426821e435542789cdbcfd88ea7d49f35ad199e70136aa1731d72faf081f9d110de8122a29d679c6b1da4800a616f559e6fcc9dbcf80a888d42b203c50302ba199bea8655fd5ce3c1289a343674a9618027c74d941a7d9fc0b97a52ddb1e6180c1413c639d85d43ef0f5a877ee6d6beaaa3f3b1b9425ee2f636790764581e1a5363ae50ad4997a54af10ec02afc295ede258207966c706846243e3090b3a6d81c47e5e0bddfc94455228dc4bf2e59e4e1df3ac7ccef512ed68b91ca4de85d04518879f87e006a0a6db727ca7e797e0e072997eeba5bdfc198896a03c79b961b562a00d31a3b8bc898b30fc51cbe5a85d12eafe42d74b36a11ad80e5c2cb6353d0a3a53c538d500653c6b1f2b0c96b8d7790efd98fa6ef603066b5da4cedd281a53730574a87d9cbb1c3627990e3419139bab00908d436b35a05c09f102e3a1548ec4427e34e2699a698db721ec41f39baca516ce6aad0ab8d24315871c2c7c0651af1257fe48feeb90fd8a8dcbf04d07d753fe740a1c597693026b727371c12156c5a87067b4f7f4fcad4d0a5b6721dd824ab65629fead734b5644520d7d3f3dbc77cc01a008417cd30fe72c5995250f0f09d5407da8d41d99dd34be9be4af69118b5228397f950a210f94683a9974de177e50441e2ba6c19937d38e02a8f1bb35499665205b177e781ca80cbb3ab8de4ae61fdb01d6479326f7c93078328f6991a913dec80ad8e9ca4c9e8aeb1a6338dbe5b6a5cfb2f9a88e816f2601b29e934714c932ff5c6ab274f255d9c963cab31395bff0e876fadea1bcd86a97c0c01ac5dd097363664643db2127ef1c3c652436b1928910e3593d66393d9b37cb0f75db7ff8adff00cfe3aa862441195a2548bf0c69cf363f02ea289ae75bbc3061715c060d441231ba23c4edea8c84a5028330e0365600a2728906141481168a8964382cd89c8c5fb6d511d30a8a58e56512221217185fab5cb9d80fe6b2bd3f5765f46b66ac88eefd1fd8840533ccf4d10bebb83fc07ecc12437b8a908159dab787baf2d59420719ad70bbc33f9d80d0012bdf2d991e24435dd07e0ba50299834b5feb7e692c5f731316b59c5679aa4c66a47c361a68da595a0a808c1b2a7a160cd7dba0f5f8f2c044721f8362837bafaa6e5bf9699adcade95715a3322452d452ac54a7bfde66c3c229c545b5ca7905f4e95777688d81ba9d43dc3288f38ccda20cc8e5ac9cab9ae50a338986f7ffe21a9b0aa2a507d3cee0358e8996ba5197cfd88bcce34c2fecc687c7269b99150779d20d07d362f564ce6aa14c8e27dd3999f228c5cf4dfa42893f73706034659f1e09b41fbdb9fdc203f48a453bc3ffedab0e06b2bddfb4cca973b1158709ae45492b6f33b52e3684390364e81aef20bde74012607f1e3f4445e1179a13c944b020c66be8a3d8e33a06bb1038ad1a9e2a969905dd2ffb23f98a1ca5fb1acf03452fcb8b7be1d009859076b87f0afa6f9712e549888b214440e1df9d093c9e29e8074ef69cb9ffc6ce4dcaeef6fff3eeaf271e85b9bd37b9703dc8f3f8a0b94c7081db6ef7e544a693b3463067c2908e7c1b3f2184f34056d15de1711134a8c0542558cc7672d6506465d801fc2d440000414a903517bea7c46b1b5e2bd69fd8354198f92d9682d2b014e57ec6693592278e0e282ed5c07ea679972343d23f8cebc25ebe1b0a9545606d409b0c15fa7746090c0eaa2d4aa0abd8dc0ed3a447d0d8b5274d3d83f3cba380cde2404cd6b7a862c364ac679ef57cbff74f321d760d200cd1e5182912c755530ca7fe43038de44e9e358931fa9e860bd6c4228fb460526f03a28a1d20a9bec5fedcf626bfe8e6a54d76b197bcd57a45aba161a6132418a929c45cf8edd430d4f99b0ddefff528f6ae6d85dcadd7da85201ddf929c514b9c73081ca188471c077515b8665be296c538be8629f11b4649abf03b6d95c2ab042bc452c27ea2b62917a1eb5a6a4c7d4295dfa20aef7a2edeb341eee30874f69872f1308f659cb23f3fe7a53efcca7c41f5e64d509f2057d8bd74d10ef00de8d5288668f0760642a1d30afc9a17bf5410a2b776b79b865f67d178f5d81303b347f2eea27b4a45b43ed390a92321bf2d4a3bd7105411e12c64ecfcb93639eba3893b39cb4673b577f67240c40b2ae586264751bd0e32c8d71d9f39177224708db71fb564961f037aca7d67959375c3418d3a164543e40b28203b140bafc30a7d7c72bbc777aaa7ab045f00f24b8b402ee4ed08f44891d5153394a1737252e254feaaf24e56c06de6a5eed310283fcb63e6075543937a98b788b8496db57d86496244f85e313473124b261b8ba4b4de84f5029773034828f088cc62db072ab41d3aa16c7a599e1033bd5e3442260ba152e6784e064f6aa3a321ca1c9fa8d6b1281181a54539544de944271bd6c22aad86661d244395e29532c3eb604caac7a38f1d13342bb54977fe777f46d2674a922f07fcd6315cd4041f156f67b678916443f28dff40daa6d93214d80d36c44d65b272de38640913135dccdad8b36c1668c303862ef1145c85dda533ab046bf4cb860d2fd2aa8da0274017fb6720069ad3c546575cb718668f61d66dbfab5c91d1a160f41629fba00f43ce2a0fbfaad92110610b7eee11c36bd0ecb84c259a885d6c6f2456e22a5a8ec895236703d02e5d1b7e958d41bc2b6a121f69ec08b8153ad2e6593a8f75ff6d9baccc25232791c96a46ce17f021e6b328c59aa09da7297b726e3afff67a26ce23d30ccc5ff80afe990d26ccee8cbc74040f3353b487d267f2f0c35f7925f2d62a9f0b9987e93ae13ff90959a51b4424a7b349cdae1ca3d161ca5285c6b556e155f2badc6b56f635dfa3fa84b63fb063b3ae4434d878d3a54701be3ed3e375f5acb8d92913bfb8bdcc893e05a27cc410e156e9b5c6d67d0caf21785b9923933a65ce91761fc4d839db5e0d6006b8ab1e153d07fd1eff61575d2bee943779db72247e2becc73c98e3dcbd4138cacb3f33d19245d445bf012cb6fb99c80ff1cd92537c8bc66749bd6baac2683f5be7a40786b08e9656559b21f0331c6e9f9e26491763e5f53305aa9be9545457a4970675e20d58dffcaabb16f0d20ab847150b793ccfae444f46066008c719b9a2613c6c3391a40ea273f9ac5885ec7164b8e42895dcd1cc900a70877beb351320bb59467eda3381befa490f467177e0ce1d79431af192b09f735a719c50fc4187510cdb3b80ab5894e8b9359c637dd03a817f8c08b784fca9c8494e9d3c845f612eb612e19bd2e0b0af5219486bf747cd82810da6e1981cdeddb9d27494d45cea89be5cefd7c585b9347521d96ca6392763cd1953a405c469a78d7bf7369ec4c1b5b01570bedc698385f36db2b44465f0c97ea513af2d4571fccdd220ae20eadbec079b02dd61975b4f39416b111cf03d69533a71c9bc718925466a7ddc1bc5f30a0d4786594fb05520bbb724c91656535a12db8955147e444abb9c8c6fd555dee891af90b540a156727c4a8b400e5af073fea2ffa2e871d90cdd6f6e732cadc5d8d272fa294dacaff57238e2a96b82660fd8e9e2525c2c9d936e5f9e14384d9e315aec129f3ed61ba472e74b333fbd2724038df24b4f76ca8f015f93a95fffa63b0d99592fa1199723400ecd73e218ddb2b3bd4e1f26b7e656445ed3460078be9a42daae1a70aae36583dae9011a19a4469a69647a5ccb15b70f9bf3f8bc19767eeec5fdac6932c208f58f66b5b1073700809973705de7dba70c7070e50398f0f5ed84f01f2c93e2e2b089c2b5dd021f16f23549cd356c4bd3e9794f5ec9dfeea87ce714c5a015e52ad2acd31a59d57d479ef436a2fab811a57fb2e23fc431f724d46a5aa9fef7134ab854814cc5e227e908b9b85a1ca67e3940f348b02dd7d0c6cfeaf597e53a96049e5265e078b699b2d66f13f0597375751540419ea12d02305954d1b60fd73fb8684a8d96e872cf012f0e389ff29baafe4a86f7b3d636aee8d79186f31f42e61843ce9326113c45ee38a07117918550602e8a22bfab2494d2872480498c76fff2d0bedd7f91f87c55733106630b03fe28ffc51ebd890f421bfdc69753242d60155fcb6344ec800b13aa007fb790f0f404865d5c629c855adf2e6bcb171c30b8342f3d581759b8fdd3411e26cbf28ee8981700171e85874c64562cb61005334459149083913c790dbf0fdb67072b9804723a8878b324fbee1e455be27cd3dd7b9cd640bb5180630d27e1ca526a98e270832c8d0dc805f59868ae6d0304ed0a2d007bc19d78d35fd2f59f0399ad4bc15c7ac13e05e2a72d5de95a84f28c33b3ea6f04c1e01b08d4046ea93edc138c77b5f816587d047c9539d40a37bf1fa96b7e0cbfc004e2222a44b593a6e221460504d7adcc0a95267690fad9e5348090f0049b9260a69ccd98cb62f10b6c0ef2f9d54b2396f6583dec77825f8bf62cf617cecf6b9ee35828081e35e6743b002cf9864cd101f7d1be05e0fb43d6b14be6223a25e89538f1538c07f2b137ce7c43ef42a314a54db115cae1635fcec461560c36f619ce443507aa5c932fd7436bc1731ad545d85d0cb44c7be452b8aff17e658946bbf75ae2c75b54e039f5acdc0f9d2ca42082a7190439f6547b2ac0a91655afd396417dd6f087aa672f3e058255ab0588618cf402524f32b00ab5d2ab5f72008f209585a9f6bbdad5c2c41774db8b6a686437d91015510b4fe4ad70c7e83d63cbab01e99140c0c4e6a973ab10b88bb87787ab9a5fdd53de7b88ae50eb82d919b4b8f4f7a83c0749b9442b6ac4bc9bc45890d02dd2bb051cd7e01c0d49bea233fed22680d4c8636c62e77fbe4193eb29b8de76bf34146ec527acb265aa1bc0e614c1018e6269553d41f786866;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hfecabe636a88fa27b186e22bf179dac12ab07348dd5756196ede92f26227e2f3bd99eacce36353e18d6641aeaa9620d0c0ba497a57ef8d5b3c3884c72205e35520cb364dd2b089457d0b4460055bb70900e623185c9fe82b13c13a71d268806583136cec8df1b6886e40499e7ec6f8f7c3af6c18cb935d7404ac4f82e25e5f990c90d09745dc9f79da65a4b875399e60feba399195dcab5e3d310e6ce3555962327812d72f8340455045ebf2b833f7be374fd1ded19d38769aadb85924d27faf08ed9ac7ef2b0ec2dba0e3d1a32c2b7154f1bcb49e9859801f1558144f6e778ead5242218e0cb6576716f4f7ab0c559a89b9bdfc26e98d6960bcf297208439855301d78fe047631e489f5263b219a553cc01b6582df5b8cc1b8e5ec5bb6721a5c2699ea3e5ea513f73757aa00e26330db84e7ad4bb3a8895fbf48c7fe20282cd46a78d62affef1250f73a0079ec5bfc54f08fc9c3893637dbfa962d379c4b9a8d09db78899956b2c665288518ab671aeeb68942b3847ff62d61530f4aa850c43bb8899c0967ead03876f5d2bfaa10e245638443893987bb2a0bb4b4692ff18c2435964870f80da4bd45ce61f9a1cc11d5332d864be663aedb5ff3b346a878114f96fde291f7ba7960dc33c8428bba573403f7f205e6e63294e292b6c91d188ebfe5cceec12b60d1926b8dc1d9bedb1db9f76ab2e26b2bf26075f8bed8f88095cd72b5db3bb41ed2ed412bbbe145a982b6962bbf464e93f27b1112ef25b5913e24e6c10537bf3a583f7004396068a75cdd459de84be204d16bd27e1cb77852d378134d1ca794c5cbd0f45512378cd00d524f2ddff3cf477c6c7fc76a46ab6c0a0dde726cdec4ae5817e27d42fdf56d7ac991c4124f89994a62dbc5e01b0b659dcce2d800e0714bc71b7030bdfecd123d69fbba88360516b9e404d6fe2abff161ad62332cf18da0858cadacb3e5b2d8ad0befadfa1b156af862ca0d4e4f3e08cda8684b04da9fc87b29b0a7317120311db49f3db937071dc7c74075779c0d9e548fbefde381b66d715f36f865d70eb38c033b20ea5b45aa18b6ee61a6a685a8cb2ed3ffe6f88e104245d61585fd1f8b9fb74203a8b8c3624ebc1e758a4803b762a6cef2c83b47ed94258528b07d8a1cf96e7bbd8c65f554e871a47f6cd4aa25556f87758dffb1945973951e3607b9b9dd1ea6579f28b81de0c94b294e2b67ac242035995262fc236efb6dfb45a9c4eda5b316fafb9b6e452439fd4ef9fedca18d6d578017ef2628c755a8b16721a910dde147329d543bd515714f57f22df27d80dac2e8e4d2dec4a17f93d1ae8918584b4a3783702d66a6e6c7df03516396180d5aec61c9a3549a80d48c61d92d920ac227f103bc400ec57e6b5a14373498a9005cd751d21afbaa2e1302eb26d6923a7d1da0e7dc48008438fa3b97d6b42d6445214d6d49868014d6d385c9c0d3aa5e775d57389c51c2979dab8bd63c18c5d2b8e1c6bbb99db2f6830ccf6d17e95f89f06d902d376435a77c723925828486581b6b62e8000aa60a425c234ba6766f6b091fcbbffb19b497e13106b7eaa4a0a785aac144bb342cd3a4818c379f80261abb734daa48558664e5c1211c46456abdcdc6b941f339ab94d3fcb78fa0e705a8d03be31c47ba31613ec2132d02152c5926936340346494cc622d10df034ff4f50eca0b5193d8364d0df24445f2f21723e90c4b402277ae8523de39d4bf5f0c3367614a4dc4c0e35a1fee55157b58c6fdff1282cbbc51c95ad12d8364f74e191d22f26ae6a433d2c3ff3f755f283658b1bdaf6f68dd8cadce5ab623a8d6bba4e960a55a0925761da3886b36d9bf79f670484db4a11b8bed372b26b1bde0c8d9c50628f523211ee688f00031b4a1c358c576564a31ca5920f3101fcc725543b3049091e8c3cabfca9d29b772ccacd407c7c87045bc2d72feb3820cf2d91069ebf2df5cdf7f7a8b32db92da5455be6626cb52f971638ebd7a1b62abcc0ee78ab5da4af8eca2ca0c96a25783c19e369a0e74ea275b542bff798621a6e47c7b354616f67005adf857a9451fd60bb3d44363f34eba6135a297d8f232e659eff9d7eb3a59bb319c0933c94e5298e9b0f2e86b64c8e4d088e4b850e50b22c7a217301fe7162e7a21e022c867364057a08c9d1554d2b533636ef27b8476376faab363f0ff8cfbcbd6f9b462150720f700eda6b18f9d32fe0a3862ef7b0e12427880c468f5e63c01db1846792d4da19ad81a61bb98b454c3ca1ddbead373682d36ad89c34db8fbaa3c23fcfeed9eab8d6eae59b97585fdc3e9292bba639460fc660675b00e9b5d3954e197b91304b1cbe612401b91899de490d9e16e6c6106d547c6f856445aae31388eca4584feac1e8d5e7d90bd7bc6a408fb9b881e44216a1da389cc1b8d9efab36feca1f78efe770b20531f552e223c401bea70338db38b73a6a8dfbb0fc0d1a9aa1b6836c7a00929a9c53d63d7b7a06cc9c8256e7b7ab213acd792dd026d4f69827bd93e18070cc20cec1fa348496cc8cfae4b0784aacebe85e9e747265702c5c2db0737d7d84138b66091db753d48068c22843c155eaf5aa61944242dbb97902c48f6bd3c405d18c8d3b0cef15c52874a30124274de0487f4e152af37bf34253de887dae58f2a43c4e8556f1b60a6b013182b0390230153b1d3f560f4475afaf9048f2101d7989bde8435a60a4c07883b966e6725cf75481c395ba2466ad895e22ec788043679d67ab671f22d48074660177b6f2f59516d82e308866a0ad53dcd4a7b9d90f312c4c3e358317f719893839b5d1f5b0b1669389fd0a68473b675d6c42560143ada390b5ab977f57e71082a74a75d80b162c4335d6b4ab9a16a0c72cf09f39a51ae1ad08287ea4c45f95c5285e56b0d1aa677de66128b990d0cf12bec239c5df05df38f9d02392ab95500fda34d499daae2aedd33fac3be91c286a106e17ab70c676a9f17a6ff07318607325dfa047e41853a1629bd3f8e71abe6833ac938acaf2beb298182ec7793aaf9c7f75bd8bfb5388b0714464044d49724a91e08a8346565e76e177f58cf40eb2d074f9c2ff0e7427e06ad2e930a434fd6ca888c4ebf4e6c43698b20603fa0091fd3254729ee63ee0b99de14a6d73290da229deaf326afadaa66cb6273f1e42fa32854ab9799355b7fcd79a408bc0535dd31b3b94d78924649d867ba57e0021a8ad9bf1eb42665aa83c5d6f47dbe283c6d7dd243d72f1ed544ac6c7daa018add3e568a62c5a569a6257e5d6522a9df7442fe0fb4ea9b1310ea4914260fff3f862c0563c4a569790e4bba8f21fae058b3572e2664b7df6d158ae5c25ac8c1d706f202569761ca047d4e5a69e4a21b45d9a36b97fdee4cde21f4293ccb8e09255800d1af5274974ca0a49fe81a740036cc15e6543b0d414076265fe4322cd255fc233fd2ccb68d332fe6701749926e47c7ffa4e62f1184b48b28901361a3bf0655c35d9de1b22e4e35334819cc698a86ed0ea2290e87c9c7c0e155146792f49d24887190a21efed3b4db7d3f6dc5265e2b9babae0f9016c284a8d3a956577b4b335c714ec1fab97c362eb67cae8e79a76b949397cc4d09c97867d9d90c49e89c79d6b3573547eaa5f52844fbdeb2f771b72b72f023a868144f77e9d6e26aaf8357983b96f8518f48eea66ae2db20bc56f94bd0d225afb1e2ed6928eb433d140371b187a2e9ac057f1ba027cadc894bfe7e7953f55419274bce0bbc387f5d89f43423d647edabfc0391d66bb93f57aaaa7ee935db704c65f37290428af5698f43cd7f71bee6cbb78f4f0c5281450b0a79febe9c9a83d89c994c60b0bfe9e828186add9762d17922acb93749644973f7f5f9cf7fe11d7af27476ef0205ca8e99e6836e06f82195cce554a0e22598891e3a3f9280ae013f3aa335b11c0fda8dc75736e7f71ba4e9af71fbe701afd61135da189d3c0f8dd43bc6bb153d3d0a673a1fdcd609fe4d09264e36aa7e3d39ea38f335ec56be113fc58b5e13038287839d6f375238cf0b6e4450613e8afd8c8c4b31d97f45a40a83e62e72abfd782a167cd0c7a3fd95c7eaf9e7fddb0b7a6b7c4680ccac94e83ea36a7c29c91da3a9e508e0e0c9a4cbbe910cd393b144f1a90e2eb80167876c73c7f5de66689ab2aee154798ef503ab0e22a20673751e90004346f688d874447c83f0bbe090235948011f0d1a02c38c4ea60905450aea81bd687fa0139f706cba0d99923544e2a36594094065f704f6c5ad3b462e4a89c576a4b2691069cdf9befb5fd5998d5d826a8c94516cd47f92ef10032b7a20e6311df531aeaa4abcf9818eb0a9d2fa3923ea94bd9beb62ac89b2ace25f982303d3e5effc58c2879fdfe9ef8f3b1e9ac3b31dee425e18a50831df1033b57272c15edadfdc3950d9607a76d1e0e60056772e22bdb8bc8d0aba6e807f759b406e648ecc9f8d1487355755dadb731e385a3212a8a98ac1ae013718b419aaf5242f1bdb54505ab0a8382b143282cfaf4bee021b8edfdf42207b326fbbd81e6e965924f789ac21ef5668f222984e24eebf0dcbe936fca259e9741444f25929bd57ac13d9048ab6e656406e973a8810df5c427dfd24524376fe107905c2b5cefa45ce1279bdf538c51237ad6ff7341a24382d01a22ed8919e6170296daf6005825500e9a157b49b1aaee130037dc6f6a79c6c003dd8afef10e8217df72cfafeeea7b61127ec6ab7b6a1d55f753f011a50d5fa5646e74b526a21eea9ec20017927b22cf3046b4248e5b70eb28dcd52d2de36339d958936e063323a65e4787e09017695f6b28b6038434c70c1744b44a8a773b986cfe45b30a61bb52105892e5c48a9050fc8983d474d30e937cd85525da1d74a6ecf2c7a4046bc75f536ad09e6fc7726e544b3b980803bfb910f5c6e31b8fd5b28ac359679e4f4a94bb00a8d8b7fec29017e808fde991efaeae9b3d599d4f42d0a09eaec4f249ecff216bea8b74ea75853c29838f744921c8c3f6658af4ea1640f320e44628ad178232288c8de631e212f0ce408ec12ba8f27ea17c53dd144bc57ec7d02dfb1907b4d0bcc9214aab6a7e38f081bf7a18816364811f620b112a3e8643528f44c2251b776996a4f1b86957b6b7e728bb40fb8daf7dfa70b7811195d791b607e71ca485112f66715a43e55a4ed830fca4711e1c09c8ca29367cb9fc3f0f9c3ff4f190c62087f5296b88227cbdc95a16b55383a517f0492165aa4db36677803d400752dee26a0147f96b8880926c96b88ad896746b536915b1640250f219abd5df55a10a9c17e518c38cf4eb541947821243ead5a89c917067b2f3880a36d59ec2ee1e3e03cfe8ab3b6b61c5b86f6d0bd2369154e9b4afe5947c474de1271945c293c5a6a80ee70aafcf33bf72745f2a21c9465d8138414d4cb14bf3ab502b1cb0190c8bccc7dc5d772ba7f65df565888835f5be6fad5600f35a627146937ad1bb9cba3fd183b3218a783aa01dea374869;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'hf900c3dec6aebbcff073b2ae192dcdf1a437fa667231b0b53e97c75fb8a961d309d7f6bebd9382fde187efaba77a30a2ada2fcd16e0fff94aaf06be179c539fbfbc6d5949a9b36aac1cb3dd51365fd25dcce963cfbf01ae6e19ea7b6f53c2fbf47f4afeea13bf56e38fd5d5f601c5b756a4df87602facbde13a667c184a3c8cf54aee0fa51cec636394aa1d80079267de2462f4ff4ee4b0444ca6fdc7bc44e3008e706557273a71f024a2b4a141e88a26349ec4325891985137c4a219ab9dac325239e91df6633b480d9a965606338386f3bd22dd9bcae2c1ff40a230a983889eeafb3d5b827d4e5e8ef17e06ec19b3cd126cb531357e8f8505a5a0e38329d813f5564abbbddedcdba7abd58cb5351d3e13c3beb0baf6347df1343a2388a94bd0998cd940d4f0e0e1aa858034563a7122976c416177f0215a5453953bfa59bfb040d67d1d1fded670f9f298d38c829ec59eb8a9fb08f6a317f55484f576cf6a82e0e7ae3e3bfc5d58481eefb7b3d89094b16e1cf1e231ecf3b1f7c3c75f8f28fb53e241a4f9ef9a39c1952d81e6dac7c5ad7a6e7a8a96b79c9d526579deff5a56e051b83db54b051016f7b6e2d526baec6eccf4393d4e6cc25559a6df019c1d07e0e09f197b4edb841c9127d865304b758b04b8059081b128e4e7832ddbd41c19ef96ad0eed855aa2c2dbcfe59e88f845b0c4fd6cd4403f43f5eaace21a4b844dd137905673642626a71cde6055d682d0a0696917c1c03a415cb755a42bc926600bd2f952496b9d88a854feb5ea7e06df9bfe97ccc424763aae6b1c858b2cc528782abfcf885823ac2490453cad157ac06bf73beee2ed4e356825e5296cf24d85b1cad3943fd9ee2607016ec65dc3cdb445e682f1a1f64c63692c4ab0b86d87ea7b299cc30b7d1ee150588ecd2b6e8a67ef0047b24e2944c1fb14d3b320e695757321e5acdb62234a92cd48cf409d374ec7b59a22620452745b402fd81df8819b914cfe0b87e38e624ba47f40eabe9d84022e5d0b5d4976262e7199c7c6c5fc1d95821da45b424afd7a575a235a00fdd48eb5353d75c9869dafde66539fee1566f43b58b926eb5edfdcf83046009d65be6b75bf0046f4ef34822d03973e0747471144cd63b133607199df186fd9a10d68f6ebed757e55cfeb695dff0eadf52648be0ab73bf9bf699a82778a22c71ad6013e5cc3c98f04a71d2bb4fa58241448573a5423b5e1263cfcf9091c7ff6bab0d0ffcdabca40544814853cd1e3e8e158ef01a6cc72fb8eccd0725333d055fcb4eac82a09eee6500d776356abc28b77ab376088a0890c2539b4c3d3908bf8c144a4b84f58725b52a13ce8d1da2b6911d0c3bd7a5d2725ed1366593d02bb32446dfd53803d83d68024ffe605b0c1d62f70a83b676f6df732b740b0f28d3bc6279a01b32951eae8bb60f7a21103e13ee67428f858fa79d6b1523da65a72f54e58fe37573c23d282aec17e2de5906788d01f4b297fdc57567ebacdffee0f377a69f38fab7b49a8b14276f05ca1c58f1654ab142beedd21a652c71e342fc21af5e755604f82c9b0c2da64ab363b071ef5d14d8ac144b332ad1920364005788f09a1f2c5b9d7457ba4f59196167b4148daf5246a24155a136345526abf3c21dd7a10382cef58a9bd091835d450f14b5d9b175ba44b38cef85ad0e196799deb9e15bef8b275137437f2f74539355a078d6f609dbe256c9985b71465d343c5bc288718d9e03e5148d040b8a482ede760720e1c406c8e8db5c107cb743ca294d525ef6577dcf692c1b6620e580913577d9e4335f3aff98d9ba5654b880ba16a5c0267a673a5ad7fb429d970777d4764ed2632e7bd9cb0ec5509bd516e356396657f3066742f5a49ec9d31f68e2db0d44c3375ee9014ef5548bb9a68a62a08ac42b0fa1853833579edddae1fa2916f6096e5241791017f898835a1a5f0b7714166016bcc963cf06eaa3611a0712aa8d12fcf5692aafcc58418c0728aaf226b0dd6aa09198204a67fa066f1dc76938a54ee7d6f1cf798639a2a2b108f8be09c683552b80c5c1664ba62e70b49939f10eb4c7fb8f6a629518f6629bd798db26b2b0c81a4c8c6e1f58e4e72b9af8602d7cf810ba0aa49f5e31b0c0e8b3272fc9dfa5cf9a9be6ecfc2cabe6b2b5a3c964515749845517d422e83f34ac7d6bc96c6b63849f1f7078b1c7aef7566914851f001812d1895feccdfb39dc77cc06faf87eec8710f6c6cf93f7d898cc1400f4f7b38aa23731c64db13daa2305f5fd8e5b4dbbef88d2f012338adec74c35998a1f57a11dce652dd3c8298278a564ccd5e86013baff09c3bb87a0ea41aad8591953dd81ae849309e9e0fd91b41ca826cb992b4f95e6908ba617ff6c60b68ffb6b01e0faf7b0c7a79207bcd52998fd26f91f039a884325e0dc56315a48d9d4605bab04a103f1b6ed6d0e17a9e0ddab10fd4ea16f79e232bc7b10d1fa922fd10af8818d8611cda7cf126bb22b748eae9d05a451db137d1572854136f1cda30aaef9e1c50257e28efcb681635230451f7c23e2356b4d882d24b5f82992c4714e02dc5cdf9f6f6cb5f2f329fb3aceadb4d3d0184956208c285c3205cb103e6388c29b964f0d8f5a9ebf286c3ebdca3931bf7c365716f97556139e55272be42dbd75740907be4d2422669db2f5477fb25bb7537c78a4b2413c436e6e0773afb3c2e67608ad8b041f6026685b4d87b8d5aeed146daa4a2303cfc7f8e3fa822c932d80eeba410840ee29f70b3d5be24d3139dc54499f60a87112a4aa96ca3f82fcdb186016303c04cd0bc0f6d882264a54a9db917ee5abab1713e4f64c9b91db339b49fbad92909e934b90af4105e15d9b9eeb85441152dbf841d07c1f3594ad214a60438f14bcfa5dff8745280521df40579b65df2de6f7c2f8986cec99795b4d8380ae666f2d617d2a002d7459ca48edb98d4fa2e0c8b4ec9d3a0313e22715ba2b9e2167b359e8267ded51159d95f5d0c32b8b3691293bdeb7740e23d7be3773b8a11a2c1ad7c0f91c99a0c07fefa2e88209738ca135a8ad63d7713deb8dcbc114c6c2f81edb981ad0d9cf3d9c87e782c197fb4961fe2984c2f02d4172f61abc7e486c5af711db78cf942d2496105681c432a372d18d81ab6874e22e1f84cdae0fdf3f28ab413d3f2b1811942ed410e73dde6259ceb6baa1bdaa134ec61dd6e69e0cf96cd70520ccd917c18e855d6d8974dafe314a9864c4b9ff3f92095f22c5127bbc305bf9e60632d515f5db197307f3f842ce3c557877f6cd8bd85ebee956c38484143c81e47d24177db767c5837dbe00bd3559fb066fe861246cdcf7b1a49314e3f872c024fcc2406107b104128f2bdcf81c42806ce6d0dac84e8f43629959e6e27727fcfb599a6a5779747e2d04f0892ed2e7095ed0df6eb50cb6e9449e61d7d014fc16bd81d74ec513dc2cdd044d6a57f5d84d30dee2e1667380d421ee7cb897fa5cd335c95f7841a0210145a0b9ddd1db64648c558bb8f1881bb95618e5ceaeb82e4eb1c6ff3e233916d770c045a368e92c2b4e115651ac1c8043c7a7b8e55fa6521868eaa1c66c6e07966cd2e60ec28ce1d7d1fdc3605287e48f995be294131aaef932f8f0acc9fd3ce87bb9a3fe1f69e42bbadf232f61863c448d1007fb7221f1faaf767484d892b328da8475f5877f2e4443fa0b643abec8c37f604a6bb065db5bc7e49b0f236a6e20d3ad02ab6e03185d62d0fdce3ecceec59623c58346c8fd74247d0b2b384fa8c003198a28073c6725864885ef5206a2230e92e39d8786dac80fbdb7e55c5fa7ef6a92690dad92b954bcece51e609de1261317d3c626c46198451dec4201d3395c767b7718ed35b815ecdd72fb2176612721f35a22b01209f94943ecba525edb981cd79b240ab81c92e577ff8c89cdd320aaaf8beed9c38528f32548920c2b12a750964d9de299ce203c85fd6ca47212d198fb0ddfd6372af0673a4eaf20aa79d8c731be0d3c3f85b22e619ae2d0d1ab1a823682653f28a67b6c9190e724f613837277474ae5dfb08e5b691308bd9f2a216ea46a1fd5dbf84f96889bffd728f355c8fdf33ff72dcce03040449582982b8b0b8cd338ce5a1fd7080721d458d5633c03a4d47715b2b0f358dcdd4a78f099bd384340cd379b1f3deb37baedb91ead0902d10b33ffe06a9bfa86ce69ebc5dadbbebc4340da89b853f97c89bee75ed703499b38351ee98c3bb397293b19c7516d383278b15da165e91d2fb136e7e1240d3ae27f9c241580e60832ade393ce81073f28b3938416286b507ad5c402c43eee8df8aad7044a26ac88cf84c5d6d303a96e227ffa3277c9a2d59feb242b77a0893dbb3161c3bb3ab2f2c8f0a9b6c93e8286cf118cb487b75fca723e5be72af2cfdd403ce0b5a05ded6787dec78447d392793cb4268c289cac365d16a0685c2468834578d9a8b5a1f35ba5b963ef8292be1b86b45811247e4c158dd9d13f33bbee174567b9b419788caf7a69f5e0a6e9ffbdcc250e4e16325da9569912b3db4604fb3e703d35401550e37ebd5a8b186af3d084afc1f80a93cb47e1f4fd055dd300a2a5caaeba3954aa9ed690466da671f364704545e607adfe07446ef028bc28d4cb13c9899f9313fcfa41385aa1114e7b9d2fca9e8e2204401a8e11e0880bf26ff2009a6b2aa8bc7359591fe5cdb270eb4b012b69ce7fea35fefd5b3ebd5c6c01a99099c37b7641749fe709892c7a10f42e97ef8fb157d0484206b5161ba9742959f9ab0d4997a9090847b27940ba639a5b0f106e8a9caadd71ace47c462209954ba26c8b6d53c05172875e85174c959dcad2acc02185c0c8a933840c178213ed59c3a2c98648a16751ae5bbcd6133a57ab3d4ae3a261ec8f72fe7b9cc775dff3ee2e8e5618e60d8fb7bf117dd1b33bd173ed3477fca73a44b38e0e13f7377905c19d1e1778dbfef9c21bc700352a8ad12e4270979c0a5ff4e554280a11f34a651629c111c44e940223e4f4fe7c8ca037a5b161640eec0cf9b26d7442c0ccafab20d2258ebcbb36e26cd43da61a7928f5cab1079a63f4b82148d377a450cd0df269681892cdc07301ea503bff3fc0c84109678392e41ebc0e8e80e1668ceafd1d83a29b1f87255ea32ed7eb5aee3a278532222f9ce2e5128bf47b02b594c758d67a91f91a33058c94c282bcce3e22326bc2e4cf0d1c1c2af9ad433c2912ac04293fc1a74c92154973615a857b136a4be6079e3f03a3d9a51d88015aac989ebb2828e7f5560e5351d14f67b60e593f3ed5a08d2edd8d8d784fb09bccc7ecc6923bfffe1295a8067b902041ca481561a71aeba843b8ae95d091688eb7ef3ce7691fee214081ae33cf7e64e66ffcdb0d55f305e56f11727daa3bb641d40b30754a58f99ca9c861e01a892e6952ea308aae2145c80e53cb9c1d572ad7cbf5e7c8bd0ef7fd4c3dee5cca042ae8404ffdf63580b68786da12b2256de53729a0014b7dbc968a271aa1de551efe93e2448f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h7764e24e30fcf0c1eedcff6bf0314c3f3db742835af3fbba4dc5596dc6b8548ba9bec8ed81a3a9df667036bd451fa28f5fa3021cc1b569579fdd7287d53ccbf7a0dbc5b5a584a3306ed8a5d8fae8ca8ba0f86ea34bfe001fa9238c8f7f43ea0783190c860ba446ab8eeefc8ae8369f15a0c5faceea8caabb8954be009beb8e92e3de4158877e4e124fbda93a320dc345714b156b7f9b96b8f0d33280ae3fb1085606d4461881463f5f2a7e2142c58e7fb2865873dbb317f1d305a37f30c208ce25a6f7208c466996c168d763e40f27a02ee20c44c07c8ba6fa7da99ba7c22532d3571c49306ab8fc4a2ff00123b163e6ede0e6582237f215e26205396bc659885a35bea0d826aae945084740686dca7bfe8f7c662eb54292edfc499e52eca0e77da6d17bea63ebe32c4a0a8c79d90621ba50f46b7590e882c7fe910800524296de188d8f2cc04035507a98a8ea9a5d851b35942ebb8e5aad5c22fa0c4f26cb14e42d7d455bf59fc8c4a8bc2effdb37d89eab7cbe0fe28a97f1236563805df1d8663df4e897671a9c1798cbfd826646d3dd16875704c06beb8917381e3203881d7bf4249565667528ed7d6c76fc68254080afb6f65442dccb0d43939a2ca3c793101a2d391e76f706e5ed2b5a85e6c4b74788bd6b56ceb8a0a885e102e8aaf3e62d652e44d47d32fd1941f9fdda4c7bf5c123a55cc1a23e2fe0aa43c0f68ff7f5ac0a92c81549945e1966c579fc020fbe6aa7b5272a2fc9d38a5ff64c46672262119fb45b95fd4799b79eefb0467787a3b6b7fb08404fedd0135e2429c093785ceb4d6878d2c9b96943244111a61bea7da6f605046372c41831cf6d0864d8f70bcd20794a89945bc83adca6a9bbf01c55b36152454b44b55facb62b73cc92492dd15a24e48b9f2928be7feb71bf28ecfc1a0d7ebc28a72830210c3884b4c1d33f3a38e3b845f6351aad08443360c3939c5a9535be9f952439f3116a61cf5f3d29465b250fc83783cff9b4d01a1fcf54798412d0942d868df1c0043fc18a80b9d05090b75c9b9a0fb571a02a1b86a2c67f4956746e1395eac7f5995808218d29b04c9caa80d9c0105120838432242adc23bd15ee6c8951d3ac37cabcb4405334cc6720326d7405efc976a53a41d8e75f3f21646b8f6ad3716020cf08785db579f0b4f2b1142c728f6bd201281c5e25e9083c2d942349e0292f3e428d71b05aef28dc2a85317297d7536a87ad0b81fb66045ec37f89c7392f7605bea154f26fc1bca115d0dd0a6d7509ddf50e74efdbab9e3755d16058701335c8d0864ea2b281b7460a6b34c0e985919878693e6ae7fd00a630dc8d6bf3914d5429ae551649ab0c08a046d80426d98172b5e010536be5fe6a46c267eb62782eca2a156738edcb1b40cf192b0f8cff881fdad0e50a916b60f34c7acaae5b7933ffaa85817d15273fb131f196e70e473113166551e21138d74df916e1e9de2bff5d5431d7684d4c714a0dfcdc4b4da4a4f1497e852ee76d179ba5a446dfa4567fbe1f20ae8a47cb83eda2c708917636d7e4d47f4a34fae4de32c83c7220f086b443139215ef50f73727d7b4bf7c98543f912d77ea3fb105dd224d9088cf1a951b6944f9693543bffffa5481b7eea462c16c1679fc19e899a298bb718a0fad4d73c2c6068f9abfad87bfeb08cf7a5b483926b54f200535b5af6915a1b85b51ff41b7ec9f41d1fc36d6622846e7111d6364793e7e96b6b7de49a39ba58fa04cde93a648bc557ccefcec2b76fb63466df09ce5846cc2aead8b37f740128c8c49e6bb8f0b7779f18cc2339846ed1d3f51c6340cd8b18b6d6eb62f702c3ee0056dfd3b53f4f4f6581db41a34e07b40f1118547ec5854d57de0017609b1e3360405afb60a106a5f50f610906357f797ba01e53e0b4a6ad88b2d2ae383f3703c7a7ea63839163a7827ec98c81b35c458944aa7d131fd108900d2c320e68b7f95a78bc36b9950feb2fda4e9b8395c2f0f0e3835cff576c2973bac830181835023ada24cc642db25371f7694c41a0b55395190853d86867572e1106b846d4b393958e08ab27caf8b64967d01c44e22d9fc1744eb92ca6169de2154028e46e88af78cbea107ea0eda6d4b3658d021bf412d08688d6d4265458ab24438eb34848f05a1e205532720c846623be5061b39a24fb25f1d1f7c59d6d4186fccbc8aa38a7eddeb424e4b4ab3e4e8c08a8c5c632be35b519d203a7345fc49301c16966a4216c78d0c821b6cdacc55b9e58e5dbf006d5731d0a7412a7f976328d7965c0f820d1235e55df3d8a4c8bf12d1ee1372ca69bf06f834d77f98182c4c2f031a80dd62eef7a989904531e99632a2ef8b85835876c42952e4772c9828f941cffa3ab334e9388b884aedc3600af177eb20c25c3d072d3c4d1e608eb97e279cec33cc32819c8cccfeb532451007157b5b212df69f374a0fbcd353748d6f4c3ffae1001419c7fcab79f211b5061571960ed34acee1c674cb6c943f40981301ce24d97b46eef2471bb77174728f4c60a2fb8eac8f06986aa1d3f7535199945504f20127f1fc163c52d7c4a7c5691e39b5bb8814caabc3b88fcfa87ddc7bc8e55ab15c1a7c8b670a740b1f55351799996fc9fd652cb562988bd9b46730e04053d90dc8333172906291c3d02a412be978f1903a5b3905f8dbdd18736e8b0fe70d63268383af32fe95977d4320a73a096ce1426d48cd0d9297c00e36e248ce882e3cc1c617c9cc7da64445803ead8a8e2abaedef9e9f73f16a88aa68e0b548aabebd30b76374b0e9eb4cd34a9afb8c62d4ee52bf7ecdff5d8a331b049d09f8c64a7daad7be3030ce75cf96071eca5071bd24a56973f74411e6dc02306925846b2fef27cdcee94b8f199fd24815bb35ec1b18857db89b58a21252bad6c63061a768dc20db0febac8ea1a67d1489a24d2ad9dada1bb27cf74c66479fff429c62cbae94e39525828ec19a4bc0af0e0a1b91ac9265d96c6972e2ddafdecf9f88c55bf6d5e6190228ef9df330d3cf746c9260842b73a50a2b7060549158c028bb5b15f221594ee183fe027122fa8b2ef14bb6725d82f0a6ff54bcb3c23fbf7b06717f1ceb0932c64c72b4ce7c415aaf22d6fdae335c235f0591343e69cacc1417ca77cb1224b51d4bb2d159c487a59f1293015ad2fbd5c1c1752d8c0acd8cd0b5a5e2fbf65616dd5e43b6a6cc748c7576a578b1ccf522a61dae45ef5d71885f56d22f30d36bc2cae64554864644c0f35409ffccd4be8b49d6cc8a342be50378ba296157b70b5622e85a009bd44dc00d3a556682e747a4cf04d50920a2b6812f4c2c4e4755f2a49c7acdd38141c4db3c0ace6a9fe925c8458384a918cb2094e0c20e7d553d8fbde2d79ba4d5346e1cd234e42035000d7172cde725c346d6100391fe1341481adfb8644555c4679534a95998f8c987452dca456dc8dd9062f2069c44e43954848d5d278c93fb9c54e85e89aba00619430732ebf69dafdd8337c4735940f9db1eca509a27b24a19754746ce773b63c935cfbcb8f8cbd9c01c3afc2cbf11bfbc8560f787dca1ffe4907b20cb43e49febc33b504539d2c48e82090963fe2e0c744440d7823358eff5cbae35cd1552416dcda4b1ccf05fba154c932e38e1bff71106e989960036e573f220f5ee2753f37c66900efb340a6f8932feaef24d3d01dbcb7f2c464fdfa0b23458001eebd2a23fd1b77cabfa0b9ceecf7b74efc74361167d877f0d4fe668680f0cede39bb07b8bcc68be4cddcb27b82042c0336d2630911f93eb67002f5452ae8c0bc4923e2009daacee1cb54790f307773f57aaec4c553e47270c3c7ca45d813dbf31bad56059020f5140bc44ac4a85b70e6c35970b92cfd02b66ecbdc3cc70c53791df100e1a6880dc952d4ff3db5a57cae05dec1aa04e2196def001d3617ad14380732ce16dcb452925d4026e381fbf97133f6c4bf9bea2cf74a5e6240532372692fe7a3587c51fefe3a2d90ef02f4b6274037ecac54bc312a8b6de48ac945af815d0d4372e289e74e15c165ebd4cd5c3fe49f33b3646606d1c4f8f3b4958bfcff885d6934591383bfcc07114833261a1d5ea7ac8b1ac55c60f377e2101b99a2ec92481a96934bb359f1a87782bf15410f1069b541126c935056c7873bb664e776bffd82b8437d502cde5fb05e94ccad4814039a2cf1c55672b4692de57770ca593dc149740b6c17ce2f5e7675003f8daf6257cced9381006c13ffabe8e787e2d8fa033df27a46a9c70abaea3e835158fd78f57f31c4075cb5f35f1d835f32a0d8fc0ae8477cb7747f6596cd39c9dbfc7b9819a1c5ae980db1f4b260ace6a2e4d74fc0162c039fa44813ce5756ebd552da1f339f463b47bddb7fbd080832bd5e20a37c6c0f540646a841bfae98551c0b416704892e69c64d3f7b8eff08a50fb3912d9eb1c7c7f66c5c602b8b0f48bc8039513cd09a1c53a29b25da409ece54e68f157468adc69a001a7c5681aaea7e994ae13a397f49277f98d5131a88264500875c5ddf0e2e5e248b90ad3736b001398409d9b1a8333158f57bb2832687525ff3402df4632129095d086d0bedcb2f9617106bab5b49c9daaa3ddb1668643ba921408d45ee0a84afc3d9a44b5d9171398ff025a5467fbd0246d71828bf9a39bcf048053c8e6e0cb991192317046257fb447d8db192f45a1e9027ac89a97eddda8aa63cf3aa1df9fdb5daa851654e305ce6c75f111352217e28423ca1cd2a74d33779f081fcb2b64eb2d37c3dd99efa8d5b0767b197772c48bc489dc29e9fd9d900ca3950f6c3c7743b29e5a361bae70279f4a12fc59bf036fd854fb1ef3f06d545eab2b6777b6af46d60fdc181bd438ff5f488b9e92a87f069568eab5297f19ef83b51e6f75c862695d764dece3366547905b30601268d9863dab4f92baf0e4f10fc755afa88287f2ff8e72c3cbb48575afb0fed216a7cc7dc06a89893cf1a696dbbddd3fa1eec01e6562abfb841c2ebea19158efd74ab41e3c2ccdc80604b39eafd03ce15f2ab9a76bd6886e30668148dcc8e17dfbdcaa00fc7e465a1736b7aec462651a42e5d704ca6b60d47f4faaddfe4a2ef411a9f826692955e40a2ddddb040d7c054fdf1e9ae77696ddcb5c03b9c7eccc66bf3a4c0d5ec607bf31e33356fab97a245339abd1a17be2b0bde78e970259846a859996d84f31d57c482fabc4e1448f4798abc226d9cbb4a4fc7f648a6ac4fda4578f7b13cbbc02841807aa795288c00c1b7dd3d54c7f7fac8307579a04a35622b16cfdfb649b7795cd63ba45169ec8838297cdf810fcdab9fbb650dd891c379592f3149ad80f99ea9eb82975dea3b19291e0f30aee16d583b9fe1a5fbd85f5cbdb587517dd090c78a31062b2a41b52784dc2fb0f73aee4f2768af473effba1643c36782d7a7c8dd8009c84413d686666f04cee003286faec1d87d0437ca29c49ba20f5c5c631af00682fbda67596f818386215e3fe0344709dbb63509404ba526d73;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h40de208d3a1c9ba7c86891b7f7b13d9303f094b41a9ccf16236d8d2cfa1a745de5bd1bc7f5328de3c031e8a26f54aebebc43775a8ded827234e3436e5d74dda157b5d0aca5b15942bf976eeb0d3d14bd3c1b405a1a9118034fe1aaf0e50c61a2b05fbc4272eaf626d572a7237f43cf3b9ab8e5ea2eb2e15ff51656468daaf87a31fbf1a46aaa9329593458dea1d04467bf49e92d90200a3d728931b6a6444411403a5e17f1c984a0e836c946084155b45775e2727a9653572a5a9e2975346197c08ab25276c42a632d0b68a1e8e87e6d47fc2914b41780ab071edf1de9d40afa975b7f5c27905dc59769296ae5bffdfb9dd5e27b5218e4f6de0822f42fa20bda1f303ddc431a63f69f444c27d4ab8828add6feeb83dffdc497705c97e43e8519d6c1a1699415048c4c0284425fb97c2db1d0d36a5daeb056fcfa30fc379ce799f074efcc7bcac6468e39b020900723e7454117db495e4a32b5d4e091b43fce8cdbd75909c41ed22997be503222639c0659269192ff381bcfc59005828f9b50c1077fe59cdedcaa30c760223bdf671bf16f2d8068b6df309aef68df1ae16740dbd1de17f1b15bfca25a5a7a065d01d36b57949d7253011ba8821d77278c2d520961369d59d0cf38c9c2a99dd951496c487c39895d0e777cdccd014e339d6f87f30126802bfb22005c9384b9bd95d8904ca08671fb80b933774d4cbb52c8bb45840b9c0d1d96911870876a5719d1f021213de1ee4efbc93f66f94a186c9ba9854ff0a92249df7d4dff820094ee859ca750c475439fbfc1df724b1e6502354bc6186529f3984174cb3aac735ded6aeea4f322fa3ba2638933ca24ad8a7d60447e2de44142cd9ea7fd36ea67f49a362addc5fca405e4c715b3f21244affcd015e33f5e6ff6ba4ebcfb4b8ad54405f9b8d3c42be0326edc932e893659bbbbb809e2a533dc321e2ad7ad67a1f29366e62ada7deea3c4ac5cdd7b3ceed79d786d854300b22e34c2a5edcdcf35bf2067aecee07418eec9010f40807b138e88df1153ccbae0e38925d9d0dc4178813f3df801037f03dbda9bd138d59869505c72e12b3d3a5a0b86c09d45fb086a5002921683ee40d600558d6dfd89b2e415c11435ce8040c5b9231e3bdf7aa3beec334218eb8ca1225a2de4f2a3816a2534d9ead92b16c0be2688bd9a096f2d7daec3b3d7baab46a3f57b6025359e36f7586edf92e3458cf31ea371f3361ce64ad42c930739ae4fd50bb5ad0ade1a4ebbb838caea7dc64f8578e0c08003a2c4d9b8b0805fdd6ed47e762c256ddab1db893428da68df7e5d69da9b13b1badfdcc9be80d02ef5fa7cb9ca923a88115349b007c10cd4f3eb23a0d4b07113fc53e874abb558d33278d9d06d8271112306b17b301a8da77c57c42b5aa9ebff8cc6c4e887ae8636a40b508d7fe29eeb21efd4023870ad8bc3e776e89115ce99972aac001a72e4b8dbb1bb891579fe3c65f4fa52ce8e49400a8b1133e0f25a71a363dea8fcda0ce6fb70a00c43ddd7342a400a9aedcc58369f111069707ae1ff3348a306302874f73280a4b552a540fdcfa2d7f2739a0f6223689a8c2e509e244585114004e95cd48eccec47867f8b9a0dba73d1090f2717797dd683cf97aae380426b971d7f3ce259466706a3a9db5d94243aae416e363db764a411a3f0ab84697ae89e9ec47ae76ca7bf8c976076e93a5fef52d1760aaed2f192d9b8210314f226762942420ecc456c49025820879b8e5090c3b79724d97137021cd5d80d958d872dc32f5244d8bee1fc080a97d4569328c8c00a40f86ff0d34ee929dc8c709fef613b49fd0725fcd6d4caa69b187e9f94ac631a8234fcf233c914a7ee4c841faa92e388c2ea874b6141ab856abc63443c83f3a0ecf43bfef2dfc2bb433542016e502e1abab747f671cc64d4de8d1d8d75ef67693a499c103a9c0cd880a244fd04e749850e160a8af844e1bbffa294c092ed11b92af3ee8b802f21b0f0cf589f310e938edb9c7ac3a77529a833a403833689017f1cef83f72e05325d54fe145a6557bd4410371083d9fbe57e5d60822ad7005d80c21df49e1186b66e65ced6d485f8883f92db74800d65dc59e157f2735f9e0e5b3cbaa7ed3ba17b8e77d09652c03f216fc67be16761470f5ba82b4ea380bf3adb0722b00ef28ef56259a20721451b440e864ab7721d7e7ceccf371efa7cd03903e99d85512c919f4a39b6a3329c41aec0a5f50e921e9fc25c1f53e707295904f0891c7a4378c3630b0e257e729614d9d810261308a2cc0d0f8b950aad6a0196a648257333b695d0fa7ed47cef3e374e45c74b7cf223450c3169bf9c228a596797ddd9f03dd45d83f277245131e41b97e70313d5688c338a185c0bde880e26d1c6bf1c08ac7f3e645560923892e55dabb7da09cf680e2703338850e5d69456d771ed3c200ff35ef004d92e4a626e52d9f45f624146e3805dabaec02b65995491fe627b4b81d0677328231b3a4b94a68764bb6c235ef6c99777c4cb941a4e7c1441daa20de8fce3fe8b3c67e47601708f5f9d96cfec4ea52bc252c312d0097792dbe9825d247e1d40e0722de61f06f3ff8536537867a7144187dae7e6ae9a47a50781741ed47c6771344bc6b9748302b54e502421dab011195274fda9b663eb646c261cfab46d14ba1d98a4c8228a9f4fc1ee8f8b553349c84185a0bc7e63e585cfb6d8699143f40d527773cba739df3f33a582a3de71f5740d17cb9eeae60528b930618c021ec66306966a10583755326cad514a05e7d466ef203880d305797f91e655710ab6197e889e15e0764b6c68536fff673e89d64f902930811b35dfc2edd8881d1d8930c563cd69f10fb00e738649e2f5ea0333ec5d9a7eff9bb521b503f13b32d7c2ba3dae0662a52bd1217319ac20cbe5a481effb4ce182bc90724853faedfcbf808a596f711f999d246d78b8a74ea0b8b5d9a4a04c1d8047329ac11689daea1ed2a4b9c2605612971fd3d2b829de7a1e22042f631333ba6d307211a45ede5e87b66d9f781c1bb8a54a877807fe42585546b233c24a84d0be3e0d5ce4b39e26120d5dac9c0f5c2b65d76834bdd731ae9d435524bcf96cf6776e26076f5c69663d9a6c53513396e95a3733d67f59ac2e5d6234f68288a0708f6a19e0b7b18abab7bf29a1c68b9767bbc3f030a65a893c7251aac57c381d0be40833c527f19955e00db4dae34cb9b98cefb3bce2666e4d099846cb7548af59d6fdb09e477f3b91639a24c73475a72eeaa42c078c9fef3ad55d6cbd85ffbe2d23512ff3c4d828f05cb98ab7f9597228e91fa78f58b2750aabb3fcb18186b9bba5e7200839ea33e14ef0bb4f933c15780b09542dcf959ab5227912c2e208ec6b0b1a8d83b0b3d423e8e68368d5cafc8eef67a923bf12f56f041a7fde9b89753a0eca2e9370521c2a1784c6f6d11840919101c44eb8b0fb664a1920049c8cb4d6402c114f00fc42f2dbcd4bc7bb5363f832d65941ee2d58b89bfdbad3ef12dff6a93542d99b8487936dcdfae2bded9fe7934876b406d0d1e29a99f18c6b01a1f2bd72b77d798f9664ba356e1c811efdbde31f3fa8439b4eb3b5f1c60739d9c6175995c63d6723d7a85f68bf6f1ab45df84da9eef8882a44e0dbfaab3f0a8d6404e349751701df4c5608f3c91e31eb259c972971332ce6c940b0df29ed384bee117801ca5653b470f1f22b53d2c4cb5353870e80d0d5b0660969329176a4cc1577b1793aa8e7225fa754a4db11573aed41d3a763febf86a0ef5e9675ecd1c9b943f307dd51e9ff2dfb1858777cacc1b4f888623e7c471a99c285bb4084a926ddb4b8521bb6f36c18685b9d1d3b82b176846e220973899281066f79976e815fe1574fd0bbc2a2ccbbd9a1bd38dd46214533cbf7b3a9a57ba0f62592a6ee6ffb6885793ebec27da71a40d63c4ffa2a21bf5974f3887c1cf47c943c577f9e4d17331e8fb5219b8d42a3d71c46476522aa90aed7b90fcccfd8ec381333bd6868ae32a4885c766c6d118272daa47ac44024e0013dc33ec500fa1a0f74740f2c46ae0d27fc452da2f7dbd8308df0e031d2561808a3db79ae76ff3a1ba97ac754c9b1a2b5bd41d64966fedf483d263629c661b1996e75df0d73fba06962c0b7be35c6f90aef4348a00a78f6a5c221a8ee75ef988dd3e78a726bc11ace2a0c0f9e0cecbb3a56f4429ed8669a4f9f057d0aa8cb09a6387d8c3611194bd05e40aa063d2cfa2cbf3d7fbf4c0ceb34a2b9c4dc8f4685e9cc11270892787fbd473acd0313a92db1fa5b8057ba0c7b28ee5658089ca5984af316e6ad36c7d995f7592823fd2ad0799d197729c6674d15b1e342105c3c5b8d967b02466b73d304fb62a1f47741b962f1cf558f7b6be6a7594cc236da8d7273dcb6df279a82c21996ed77e957becfe0b15dd1404300e5ec1ef893108c9df3d044d5ad6f439f2d8d849a46a4dd0cb66b21dc9bcdc054b41f49f1e45d151569ed89ee6660469c3e5653f43a279014bd62ae87a09be9080a111cd85b5ea2adedbd72069933dce872930c0d84fb520ec453f77e9da4cf42c915801c3ae191bb684c4f430a6e78490b90d598d91608008da137b52e2a41b4b77068e5cdc9cba75b2a35a81b0176c8470fb7424f163f999a8e026dd1a0a3e314b8bd1b2609f1336de51b8073ecaa645ddc964368b62596c134e2df70a289c91acea398f0d7a5546248025d2bdc624dd2e74062f766f281fbdd4c7fbbb0afdaa8ca4b3a508b4f1928a363b9f27db52f99af07c4bf73e61200d7c3c3f04a33e5bded0d82c3cbe69785d85d89ccc7fbcad032a851f3bc79066ee6075254e27b583d92163c5579bd3f958555b3614be451900927177d3e9be3b83a43bf276cb056efcf19b3127826ef75754b2ebaf18ec8c67fb2e45983f0f05b1b13ad685e7b71d7ffaf7ba94d4c9d7d762f743174d56d10bb5dcf75aceeb1df629e7f8d85d8366749e617a939f0837eedaae742e3a3b1ed457147b52f59ca55ad7622bd5620393af9585a3962eb4642eef28853237b42800b1d10ec90c38edf8b25836c9513ccef68bd5b676d3bd82b59b28f2f9fd335511608ea44d50f847ac721dde64eeec81811d047ccfe7fefdf03e71e5f8ec9bbc98bf4e0a5dcdf65446becf5750528198570039c51d755dd6f0521f704ccba742da199b6d97b3c2d78a3176c8ebdd3a32665b198965d934a788fd193d96f5e2fa0c06316f82e025f0fd8076e035334abf38c85fd6fc835075c3ad8905931486c0d96941c8d60fa315217f7603306515aae0e9b0798400281e6a279b3d7b0d4ba5cad48e15f0c8ca28c9c65b68f49c69f2927da468de196bf6f37132718ac4cd5325f44117531659d4a05e05ec41b6805569650810bd4793aa62c5921f34db9b10610a9fe196541a6382e341d89da81e321309d9cef5adc6b9372b47348845301d6529ab9dcae50338e5bce72e790fe4722e6b2b80d788d0864d86608efaeb727b49d906404;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'h3ea880171ad808f56ce5e7ccff450318361bfea4a06238144bfec9f01fa58b189789453f23c9c2dac255d0e620b12b9f0de54c1c7b33e4f06efa611efae07a3d16b4039f3033ddd567c28e7e2a0d2d9fe0b525f891afdd32a3cd757c722e1bca92c66bc20e385e899f97228d2faea107cdbf753d02d77cfaf9e81c9e99302d08de30dd90cfdbda80033cfb1eb5d49b3791f7b532e2b21de561e751ea67e14c68d5304647476edb6f7bde49b14ca62996079cdbbff31d174068a5b474274427e596bc235cb9c17856184d882ca61543aa256de87886a5e3a20990658ecc70513adb4903266d2f33f8e7a4359d82eca7595ce0c010b9c75581c30fe34f1789b23bb923aa518948d3be704e8f7de088566d1906598220bc79b3b0825f1e72d12dbd5864b72e1b1269d48aaee38f593806bf2dfac5aeaef3390f4b4ddbe221026629d053b06a4da2536cec61bc794b49a58f52f758aeae3f42382dacce462641a5debdd0ddd23520b50c32343ce3e7e449838ce9cf025f629eb541193147673f93140ed8f41c994ede5489391d1a9e2cbae17016968c3bd412f0ded03633a9b81f7fc2e868988102e56d2989f1bde2cf3b62a958521f07ab2f880b40c6d40e2a8327413562e0a74003451f9e79e512f3cc0ccc1ecae5a52b62ea108e3afaaecc935f1242b600900950040f408be735faab84c0e743ac20b72459ea1f8dd234069a59d154319bc9608e0c34a8546a04ecd5e147ea27c8e28f651c1b2a55132d23529d5ad41bdc7e9d8075666c81155420bf62ca06930f986e5287fe832055fcb1c16ae0db38ce4c9d0765315a665372be793a4eaeeccd599000046de3c4073c8c1b4af916f9f75de7db6f5d7382ec09822b8223c754e4ebe4c5de77bc15556a2dd7740991564836f13c678a61403fca602a42b9b6aa4246406da157764790c555f5f88cf11ae2d2b6f154a5a73ac7a60796ab3bb85fe0109981fae7bf8c123cb7edb3af4d3ac35782b8202117b45923d89d0bdb7c7878f60f8c23a75eac6d2105ca4a75ea11b431017e30bc67992cb3db60c92fa7ffb45b348b140b462d73098c4f962a526b0c85105492e0ee7871c23c38075c0cd0fb31ef49eb9a8c34bfd590dbf10258aabf116daa834d4b10fb3104c80094992b693888c5d684bd9198a1060871c093e04f9703866ea219504786c1d1e954584978a2865fe3116ca9d7053f36ced7053dc6a8098db749c9cbef44a98248db3bb55f64b6a477ec20f3add90383a49f0657b9102952ec665fdc56130be2debbbdd9c281f6ea7e1e6cd726dd703522f776cf3a0de563421beff04405d08d1c8f8b1c1f4c71977eb36db9ef1128a2f6aec11c442e75361a70bdba5dcb842683b8679b71ebe044a3e1ac2b47c006b619e246c97a37ff068a55ccc1a1d27d84260acad7bbeddc9fae8f9f5c2bbf67bb9a50a4d5ef1041b2fff31d618a4fc6ca337c15a47844ea6c5c47b3b2fc634b509057f7c5db5820fa9ba8db043de1fd669936920a4b8cf9f79146b612e98c89bb1366dffe3a0dc4b15d497f8270fc6de28d454756d622c330c6cfc9bd41e464773ab47503d83f6a7a1416415ccf801ef0cca76023c74063e039fdf7856385f9921eeeb506825c169206356ea813ebcf66790b9d66e8212f36fb2acb4eef69eef9b2979ffb5f71e56f061088b98241dfbb332cfa1535364f5610878d8808ff23f796901674cc226179b5cef3c1311460cdd865d21418fab62ef21332c60de177b297b72168e3b5aed5ee5825625a7e75643bbfe7066f2a5fe3a3d76c14aba959d42557b8259045859d39a0fe6404273148c40306ddf16ffbfae76b9411a04fa5af32cafb97ec138cfe7c273a02e8ac3a6efb781a9909baae9adc7e8ee6e83959f3d7566b78b0f3ee54a091208d21e3672f1396faa572c6cf9b7ee90d007a7a10e96441d86ba862aa192e1c9003b93e9241c6ced8e69acdafe35471dcb50e96cd11541ac0cf3d3e53c33941cb58fb3a4942badd19d08856568b82f45e02fee6e79d40a517077d68d7eacbfbdab67fa078784e4ed0fd702858246c9bccdd66b96a56670eafefad903c90f2b0cdcb30a88f4b78ddfe252ea9d822a5ecbae607fac3fb081b2c4f39b73abfeabdf074eaad380cf6e8f2f0e2193449c81644d38a9368ea8d73fd73bf3fb8efcbda904ed01bd69de3a69910511986080fb98c2c21aef60946157d3793b5706ee911bcd8fd0579494477040e710082fe7284262aca6ee4eb579a64ae8a0630391fd2475c94641fb6323a8d70ee1f282d6478da17d497094fc447efdfd9dfbce9a390c85727d247f97a2ff94fc14d7cf0f55220a2b8da2808b5c2fddc8fd2b99d3b2eda110d9317369bb92a7998f2e3f82c2661c6733a6903008f71da836165194bab6c6b4af3d2c5b0eb217b9ecc85b5b3873f7fa9d6c19aaf46024a4f79111f32ee28adc4e2b4d23ee4e895bbf49c5a8965493d94d73593b5e8a7a777644095f93b9a04fbac1e5f501a34a1e812ff83022bdec41bb5fb25fcf90cf19bb04a4e7f4637ac4b5dd2d25e4b09761b5c8176f81cc862f23934f8b0387c3ba2d80470a74acf76392b87e1f7a80746d785dc014f66067854dee6ae1ae2870281a44a267e7a730be37b51afa62ffb9bbe3c5632a2f24204d2ac877107b02d9ee8522c8a029c79bc44d4092f35b6f0e0838441c4f2447f371c0938954fa27046d49e970e8405f5f511b6b40e95b2ac26f70ea1c4f97b6dd2f7494ea6927a04ad4c63bd85bbec1e6a51b9da7f1c7b342283c0dd7c9f618993df6cce5eafa2fea1f8e4b17cecce4cf06c6d084494a8feea5242ba974acbe14383c80ab73c35069879a2e5321f8b7fc2b00228d015eea6a55a708b366bae5cb82e2454ca3352ee0e45fd435a5fbdaa537419bb4311e116be0c6c77ae948db025c836127b8bcffe43458d6763c8d909634b1e5c4be862b6dc4f780ea408d33775b053ce715d7f8c1eb511365cfbd6c3fb5c8d3cd5c89fa3af8f3826b6b3dc2f56a7edd0057d092b5de5b0ebe173890f8dfe28c445d4441b9bdae6d86a80e13e5bfde262171f9518eeccc3ceb0fda063aa08fcf8af5ef2db6737abe60117594125dcb6ae4ee2eb31ddf8efaf1cce7df848889f3271c002b600ebcfebaeeda145062b72382af5b3b327522c889e1379f597cbf1fe6fdd172ac5fc63f42cbaf8ea116c828016a8a26410c3ef18e5b40aa06f0a6480d751e2190985ae700693446836ae384229ed9e8a114322e743efb0170e73da4cc951692353c2b468bf9838ebf1c1cec308db3868e6889b45463a2b6359140c763d5b4541098087507da8e7ec646e6ab64f1ba12f4c2aac7dcbdec1e79a5a57cc31f7f7a1fb1b278dda32dbf834649aea9615a3c9ed8e39935d1dfb0d865c7495a09e4e65ca1be921a5e97fea8b8a4f3a61ad3dd0781a66e317d00d9d2c04a9f7b63ac78f41cdca62a0579eacc740db47ba73d54a4a0f45dda6f304241824c6373f0384c5dcb18c48b29e546ddee57e118ed558b58e70a200b76c4537b924c51ce86d8b978c3331174a2db71df04829e081016a86c318524b2ea3185f68989a80cf01ef4a0bd04dd83eb93a49b8fd28c71d031efb9ccf9642c42984d11a4754bb6bb42b80a98471c9281456b0c299f5ea6b7c24fb1322c73743af59779c9c3f8659d0331f7e54893ee24a29922ff77c35c123b0420387027b3e71783f05b81ff53ce734710cc2de5c1e0521cae4c5e2720a4620c42a15e3243508898e2a1473b671be8e28d20cb706e4a2a02aac2f28d43eec679c1ba583e585eab5817c582777575ca06c5894df13501e6b29f6aad20545ffd345ba9a1c8c4d1b035e83ae19ede579876ef7650e0fc60f70a94b9a3c0bad24b93d66086e4ef93c32b44a89fcbb4dbb63636690e54ef8d1c38c63a2dde4d09fbcd935134711070b2d456365cfa8b4775984e814c8655a2128a7d3606c2c38f67ce8edeab9b53a11e3392864657eae7f78b3bc86e62cea5a0ce249112cbc7abd497a80688e89cb97d85e9e03babec1b84ca0919c61d19b47e68754e0a15284827776e4b3395d7bcd38bb8970c5100fe0b05aeeab8872af3fc0e2ff56682272275995d3b3c7b1652e465a1d30e14bfb43a38ce6733a50ee39da74a5940fa549b5af3ec5ef2869e8054141fcc3e5ed44edf998249a3ef0a80696aacf5b84872a449f7a2c181465de9b2bca16f40702fda5fb578c2770b4135cf0a8b19bbc785ed25cfc3a0b028c3e1e24200ffcfe9551b2163582110919e7081c189e2c8f37432d76b8ed03c20dadeaa2b193c07dbcfc1a59cdbd47dcf40a3e68cf8aaa151ae5816ae7e60df86629b5ee75f2e5bab48190fec97185d97877e82172eca205c4a8f72f62cec9d10f312907c2e490f74d5bd6e8469a4d99408f7dfd915ff30422c6ee8edc1befa466b98bb7d48044ce12cd3f8de2c7821a00dd70fdebd79643c7506a11ed6168a1730b25ff5c5c974c6ed3499dc7147d69f209b3706f122d48f6ac64e574f45420def4c1c938f2e29ff92caf34511303ae610de65de56fc4288b29e9665abe08580bc5ae9f5958c8e3faada88889cbe37f69a035dbf6d2e02e4f4d0cf2a31b32e241ebad2e8a05f6ecd9cdf2ee606a154f7b5cd177cd43fb913f08071514334a6ea0c94cb202d8dd84c133908c6cdb7ecfe911f9a3773ea09595cb07a1abfe277577ab117e2cce273e0e8abcb9c881d8a4f88af48e22c0b0cba5f95a816af1faa6cfd6612eb43a30b2a4ca1de8065d84feb9a2bf1f3a350b12285fbccf498f3e31a2bec8dc3c8ba4c442e2310c9825495d1ba070c20a0d6a2c72497f474c61882e56c609cdb2b2848cf13501ec3c6698351361f4cc55179348679d15001c7b1b0457771ed1f84cbfa6fbbd22f6931cd4637241042aa8722ea5b326558ee286be148d3450ddb8c388874fce51179981c4ba6f89d31e6d0f570da85f04556d5f3dc9751e6593eb86350d19c7ac7617abd35a8f49b985ba0346d1a01de3d0a5cc93d7bed32857c407d553dd000227565a058bfd4c65f533234267a6d14cb0d40936a9e72dfc65f129a63747b1a3a7565a5a0cddba9c51e863f15666d0bf41757fa6d601a23e5fc6e39466e532cb0502ecedf34a70e3fcfddb425edbd484d9a9196c0bf2627edcf0a9e1641e3d077b0feb45abf788763eaba2aba3554e5b15a81043d69611f3e96d5729c63f84d684e1a600548b2e9812c6bb54936f22c6c60cea0427382ea099b31c35e0e4bf72063e6eeeaaaabd3b19a1dc14df238bc696861813b21e83cca93169775469eb2bbae0d1c4882b1af6ed8220a67f48267cf065ca2abe33d23526806c293d4ee9b2611cbd9ca5b572be85e03db019bdbad33e2ec0ab2ac0f4c130e7b3b524751b74097457dc05c1c016d4490d6f1602f0112b35b317f6a32df466d1939f7a26d093f99508ca4a66721c76d408a3710b5c1c198464ee821582b210c6051c5562c268;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 31104'heab6350e71ba340f16b697ffd9f87c03950a143d459d01610c715f535e4e8678906abf29786a6ff59698c13642a76f3b3324bd789c06a73236a35176ecadb7a06bd30af3c27f9b4bdb30cd67b24e1ed0c8d18e4c772dd49494de02415927d33260501594b96fba124157af9345708df6286be60fce15f79cdad1887563f12a222e1555d7234a1b7554de99b3c20d11dd5c2c68d00df6394986a8d23a00de4ca87684ba93977fbb286baf33f1d3cfec5c351d059085f0518bebf1110b92a593f0dbeda7c76351d34a300721b54fd0890485ddf6cac510d06f5dd11de79bac47bc1ad96ae0036b947e0089f3b59470f54e45f9201d3209bb76f85472f9051afacfb63b69b11d85b58edf5418ce09f6d7d79564412518a1fd8fd175365f68706bd0073e1fca6770f40e20fa7b8e518faf44df16fa0181e0ec62668ae31148f86c181cda7c1e56d6ffba7cd7e3d14b83ece152848eac69cac6c467d8992267288cc63f2dacc7e592c7cb0b0066801e0994c7b53a1eec6ab43e22cc23145e3634bac5a9346d322cef6c17e398e574e23489063c54b935868a505cc4d850f4e8231cb3ffc76bad93ed5970f4c2ad5e4b0c787eb946d06c112ea7ead19dc50e3c6a02f10753075b5522a853748e37d834876856db62ece26c1d1034be03e529e1a922ea872508d7c7f849cebac04af0184bbb1c0db83d270639b6e4958de1283bf20afefca820e15f73c48931e4cc956050ef2dd44b8b7b767f096f6b66c58339ef7b10dbaedf28ce6bbb35f3519b382e5b50d39a769a13a3a8682d3a63bff88b3e9818ce258d8a06ce738a3852afb8ecca6ebff1926b124ebe01f96f60fe50bab4bad1be3793fa5a03db4530febd381dd8425fde4dc371c7eedaa6b7288557504a640d1b55f0ec9e1b940404549c34aaa3bc098d5948885754e89dfe479253886d9d1a8bf832c63662329f65752ba43e606aeafcc40d3e6ab27a20cc853c8a7083d94286a2dbe8d635be3b07d691409188bef2a6f5b1ea274e0d201aa463d6135203345b4ea9de9654cc31ed71bdacbe0c6ce86b507ddace28ede8ce0f2d7f4f52bfc463465a7953a810d908a04052857d8866b1aaba68c358ae9538f58c70739b5f321e4631706b00363ebc6a11d2c6fc175afabd86bad6d74058e0d1017c0ce319a15b1a68e536baa7c1f91b077a90d1ce42afcddc46b2631a53a74b3c03f99d9e25a649edaff1d2da0af040cea78d77b3f8709ca9cc71f357ced2a4c84f33c29730d3341b6f52b49d49f5fd95d39845c42e7eb952dc369909df23094a884833fb55b25f842b90696219e9e135faf2048e69c3db44ea24ae6cce4bb6de7d2777635cd644e280c72d5bea16db8c00b2b2bad10f1fca623857a9e1b39f9495d3f82bf6d48a82abd0d12781117b858d6109dd3e7a627a4e5af6cce6c8fed65b6a0c3834113a57c4016288c7826f04c204b46198d32402d4d27818d40beb87c686d0c8c687eff200065d6fbd00e64551b32e9d1d46fb519f53c8cfceb0b8dbf83a0d3f3f04ab552e6e24734554ced9e3aeaa972a0397fd39aeb02d83b42ea2d70fe067e440d990d2f62862cc964daa1017fe6d781a2057e6846c0814d03ebb0d3f659cb97dc4e6e6cdb033634c6381ff0a322259ba35ac0103a5f96c0e0d95fae16abc821f4f76c1f19db38aa724f678bed7b8da68a9a0205c23e5ced6c72f7b0b57a9b6c2167ef0c95a5c59bd05292ba3fb327642bb1987db37dad9054f979b0ffc964f3824d9df463f357aba009bfe753a7e501049d781ee79891719f821693d6418267f08342238fb845de7e1c7e0a856e0ee22b5903001bc64f0d060178f6786e6bb160e199aa363e320feca3207e8eb32167f47ac48ca95bdf219cd90a505153a846e9110646de788a29dc69541b11f4934a2709c1b4b3e9c1a04cf10a4b43705e49fd3507016b37d3d92dd3ed1af9fba03cd9dc6b33be397d1a5959550846fbb07672a92f9416d9aa38f25e06f8cdc79dfca5737fda545b5ce941c387d9f58b234cfe13e854782ac445e6006a112ae3705b1b1aec1804ef41e70deb54cf14d8c86c889cc2205cc1312c501d6061dc97ca71aa740eaccf81c09e2e651979fc2a29d165d8955b25576b93f2c9de1c267a05a300d4e467f4dd1bbf169787bc996d0d50ca33c718cf0e0bb9977414d78e1899f61da5a5f0fc63cd437ba4c3adc227a94d2102194672a30514973649370c539c0e75b3d7a8e630ec72d4f8635cc5803a1c27fca9e0f1b945945efe7a56533aa3d14a8271468e798bbc8f0e9eeb5bb64d9541ea0db447796b91377c4b47db4e71748b857d9aad426964bf162734022fb0d32d2e70c7ec4f98029c9edc48db7de28712fc45f1542ef02ab2e573872e37826b0260cf583be7377d0061008eedd85d97a1bd106b67cf579dda6a080522d6d9307c21ca92a3865655caf5da979ee481aafd4a5be37ffc71eb521364ad3e94b15d71097a0c3c0843130a46eff160c6d88c277ff2ccd7f8dbff8732e11f6d6c4383dd230f1320ed00f404c94237330d67c269906f08e35950f431bdadef247eedf22ed05a65013bff906c7992d65aa1ff14b610333c81ba6219329745f95b5dcd725a951b6965ab570923620e946d5ee93632c47a210ad73ec1a6ccde48d2c51c436b522bba62dd01d2b31a136382b92961c1db2d68783d709056e27966dbdb92527a18088fd80a1d35fcd33eb45f3d54b793a226ccfefd39b7d165c00d02fdbde24f918878b946c81c9c37c29dff079aa459dc0ba0140297550d75d74bef27f6fe5c70d89a168b5a64db572a7cde8069c3d114bda69c2e8d61fd1db5c6c603a52ac183b33238eec39731ab58b6ed71ab0876e4cf33deb5b9cf552c1fd7f7a2454eb97cc072bb7733bf210cb174f71041b23a9aea07e89f4cb6c3d8e2fe332539b6408da17ee54c74f9e9621555295d00a61ae9192aa7a6646dbf852615b8db62d4211ab421f8e3703432348af91e3ea752faeb40b0e9fafd61eee0c7c5d45f235775a9bb0f3351264e4ba3fc0b40f6b26e08fdff8e1350c0ebe96be7507d56208ca7aa96247313b111a0db77f0d1e08276eaf47878648a83ac088f0e4b040cf60f25fc260a3683c660f063b4ca6e5f93b42553fce6d32a007d4e9f45fba2aa563e4efaa641de5eef7fc5ebc5921f38a95316253cdf0326f348ce4982025c0aebdb9bae20c244577e53af814534ffef1a127051eecfb65805866ac4ae7227197326f3b6b988ac55ce202cbc6202695edc413f210a0f86953c2fb63fbda3595d41a8c6a27f1b8175ed0d99e87e4f737645fc10b9a3e2786ab7e810a9bca209b508a7ede6f140ede6e98ecf29e501bf3db16d491416a42a7ba6cd8fd37bedaece0d1d32153c9adfd327792937fbe2dd5f8c425401828abdd5669a4e80be162a8646a51dd2d7c88f2bb021f114dc6f350917acd4216594e98c691b0c339f2196fa7fe388a29a455292dd6c276d726d5e0f28e7c63d2055deef9f9857b4541223828247e5725211432e149b187ec1c24219b44ba5c86f0849b3e2c9e70915de58552c47d1304b18a5ab26f28a60d3e1d10e2b627c285b4f44148fdb283fcc932c97ac7f0d76a4514e305146484dfd115d450073728226616b82fa9d4a01478e71833ac10f5fe03961d94aeca2209956c6e474c8a7e7daa874c17eedc5d7a8be103459d87b6d0994294f8ab361c44500131049fb03ad78359a1971c8d45202d79b7b037d00f5b2eccbdf5630d56a4a7e929c08f0800386747742c2ab37ad24d23b6eb1456ba3babbfd063c24ba410300b2c271ba12ca0d56c26e1227cb71285172d3e7ad27a16197a6050bb1288ea02323ca81b7dab033ec8b9ab7a162bdec4b0780fca9ec2a47643b927532574ddfb8c2d42432f1d2f2cccfc20737c41ba6b752a068d644d0db0d3e144148e8a6aeaaa74c4d3ea23d5d7a70edb297886a638bd952fb78c0ea45c3fd0de14b524b5db9e9f624f2b7b1f8c2ecc8163936216bd323d9e2ac4293061737bf84c3f8535451ef37415c255a658a745c2bba84d8b214c76eb878251eef6bee5d422f2e50000b8bac6da8aae9a6541497e26a14b175d9cab8c58dce4da8f0d91e784fbde4e3219ef75833e68dd4bb9313aba78445935a003746a8af8a986fc1b5ddbb8a4276868eecf0ff66af7f4c94d6e2381fac3b204ace94df79fc6aef5ef2e2816c5dfd4fcacc5923769cffa2456a7f2a64c6549057e2819548100db7d945483a97b3dd8b8d872a1ebf00067b6b61251639fe1506c9d467c7a116b9351de923421c2b51fba5b8e3368a524a790afe32907eaab59ea3800318a4f53f5cc2856ae0dfe59390fc85f566cd3b69dc3f88c24a0367620b473a767be49b092e96b4c16f86e340b1db07949a1cf807b7aded2834607d78c88467b2dedca90373f154bcd4b002eb880902ea022a58019d5e487d8eb2363d54165515936dc51e1adddd5280f3fc3e78fc3fd934a572e0e972d25a31e43bb7a881562744c47c8010cb09442994585c6d0dd77f7bd5fe6099dbedaca0d93857606851f5cfe88d7968d7e066bbe7dcb44112f975da2ce9907d42b8d9089241705625b0ecd976e5d07bdf9572e2efd682bff482178ff17793aede0aa406a75efb565f903e188aefdc49ba0a3260c7e0a9513ed0f60c91a532e8fe3ce2cfd4604e66cda093336e865f20982df48d9d1a49c791754f1fa2d3c54e2376aad73846a5b485a1be847036a4d32b8470004e2cb7b8335b9124af449d3622a325e37afa11847d8aac12c5db4f2623d6dc0f70ece0c21b50e94a85f3b4de130bbb089ffe3e64ffa8f2244ff35fc77350b0625b734976dcba2bf5311b4240239a9f04f91cc3d652799b5d97a14cefe193264eafa82ba1a595ac270608ccf69d31a2e09b599893eb2c8861d0a4818149ad152ed88ae13e0104e2f246014effb5e9879e9181c1838ac7b4240ae2342d92e642abbd3fa077bbc06edf1a4340eabb3e4ddd48dd0f4ab005b8912906bd86953685c7901fc6e2040db75278c75f92ecef5e7dc62e5f450f435f98e0c29276399759841caf8a327f922d236bd58090822d6043d8627d0f86a3fcbf7a233b58d7a1706fa033c5d06d4347de8d88fffa690779e94bbfc5aec0fb7223787806b30ea7526db0c4fbb9216cf20348d8b104eb78679d3f518ad29aa3b0383d55fcece969f64bd6f383a9eefb1203093fd373efc716aae89cdaa2ab7725dfa27f6d620cbc70424a4e0b7ddf24574524fd164ba55bf57e124276780721368c4c8fefc7b50c63c602737953007065ca751e9acfb7f8cd9c4c21c2528bba8bc5363734698d11a47b3d7e29cbe16b1defa3c014cbfaaea3d5297c80bedbada4be77cb00b74cb8ace143e3d0f394d6d21680b49801edfc2144cde0abb5859adc53b41dccd7572b4de45edc7af1c9908a1483dc7f38eb21eeb22190f9d5c41e6a42b146d3c708736ef7bcc50b05401d866;
        #1
        $finish();
    end
endmodule
