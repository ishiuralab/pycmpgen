module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [22:0] src24;
    reg [21:0] src25;
    reg [20:0] src26;
    reg [19:0] src27;
    reg [18:0] src28;
    reg [17:0] src29;
    reg [16:0] src30;
    reg [15:0] src31;
    reg [14:0] src32;
    reg [13:0] src33;
    reg [12:0] src34;
    reg [11:0] src35;
    reg [10:0] src36;
    reg [9:0] src37;
    reg [8:0] src38;
    reg [7:0] src39;
    reg [6:0] src40;
    reg [5:0] src41;
    reg [4:0] src42;
    reg [3:0] src43;
    reg [2:0] src44;
    reg [1:0] src45;
    reg [0:0] src46;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [47:0] srcsum;
    wire [47:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3])<<43) + ((src44[0] + src44[1] + src44[2])<<44) + ((src45[0] + src45[1])<<45) + ((src46[0])<<46);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef6eef072fb95bfa1e4a7ce2e0c6ad4de5baaca80e394dbc911e97f2a8059b940777a670eeaa43b5fe8d0107df49ac9c96055edeca68dbb9b68651eb74ff59c6c1419ae82316fcbf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h120a4a0069e21725677ae26c614bb1d1d68a34ee40c14c2d7cb4ad756c7d4882e3b60d93ee109e46dad30feaa5d1f49b0a937adcf88abfd8751eb39309f2fd64196e3abb632f9324;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4c592383618b931600fedfbffcd9629c022ed7c23e85f15cfc03ef9393a81112bb02a2d9577a39e8a769b8c6ee49f600d8403dafd5c94d2e6083561007df6e699e2c6e195613342;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6d06ec74d756a2e3c03f3b30deac07923770c613205b6a7bb4777dae3bf9323fc49ad3a11a036f0d321f9a59630d9446e8aac0d827e6faee56e7c20a172654e51c03f83d9d4aacd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71da9b9d9172d3d5f109c9d51ecc5745d7ef92e885ba024ee671d012e73eee7fb1ca881dd7c1f1a9c32267b7b20b33ef166e0738b6f22f265304a5fe8c6a08fdedcbfd6292e0bc3e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf96a3dd9ddf54fa8ea957d269a34f76b96215f12685c9dbc179511826fa67278010d6854af58b35ccc4edeb9798846d2d52b2c6112620a8325cb76f5582ff868b252d42fb0ef696e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h763b19179ca661a2cfd13ae16c699fdebae01f44428fc609d12358369d84b28beeb85d1294d8e4bc16c0071af7707dc53db3136d57c318b447f481d2f97692cd21c18b6a2ed82f46;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9d0d829d7507015c49b92d36d33d031d4d611a7e25f2255ad3b0e7a8498f0e8b669fa315626c6ce42180bc5559c0c3d4bfca822392b6dadc4932e96922624bf72837fca78a4598b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h228ee9dc508eae9c374522d2bd0c268aed0392fb399f49df9f741b1e7e17cd186269047cfb9130eeb7f0d2bc22c7c82f6f759187e7eb500e258bd1b523bf0089e7d0ef4f175c9975;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h812111f5e59d459854da08c5ee0f8c1f0023b37a6b97c610255e6f40469fa924bba8c4fe5cafdd3e7e36bd536cfa12f83a2566afc069d00b4e647ffa1eada520172896d9e368793d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha51fa5950bb328948c1238795446a317af72f006995029f4835eddb616f5b99f55afc97574d9f84e9e73c0ebae393fbdfe2ed2beabe7b4873678ce2c12855aa020e8f640af597404;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ab17629a715ffdc37ea3fe902fc25b1fe28f654cbb013d15e3e0b611f84f8548755eca00b706b2d15c611b3ed20daebfc9798fb57ac86fc0ac8fd26bdbbfa8b6f2d46c48aef16cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed4785e03132243d690a0edcdbfd9c37f26bbed8d812b2e649745dec978e5245cd74d4299235ed7ffc043486492ad9b60349e7046f228647434eaaefb46f3b1b3ddf689304264a12;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3a526aa90fed06b4c6f33c02fe08fb8aa8aae2d1c2dac725b851e2a763303028b46ee0221e029161462ba521118a58f261eb453164ceb1196bf7605aa032905682412817256a5a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f7faf57712a7216ca9ec8c482219d903e14c5137e4a23b49f8c2134aeb490f6952b4aa57429b17f674d01aaaa21b0cb3126c074309780a835c8c6aca266d91786a68ab3b16a199e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he36e42019bf32db3bdac7130e9ad32cbaf84e36fdca64444233901f51cad801ca89f26b8ecd831f77b34d6cc1338f434447d24e38e7b0746b92b1608c2d5dd7f607173b61f3995c4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7305333fa822bf929eaed431a463de4d2d4a9df265b42275f732c689348291405778520e74dbcd6766a5a6be4245a47cca767e96b2205492e2849f27f992fe7aead219dfd1b5e260;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8704ee81e97820a7b7574efc505257ecc9caf35fa0c5c642fc43570fb916173828c424110aac5fa9e66d294b6802347392f80d8fc661aaf0aba2ab28b1f6e139d62a4589412f5213;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff1c61273736ad0ac8cc7ef6f3a51b1b017ea50221c1ed940dfdba239580b84976fe0294ca19dc24974df85eb50f5811840e95baeff07126dd708967a7d3c4a720aa317c6a5a9c93;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65d24430ef621ff885445e5528508176651bd0597aecf91b9f6ea2ab9e4e19f6f47e94917b856e99ec1abe5495f53cc108aa1a8bed83827478eb4a62042cd53390ea8a84209d0d1a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78cb5fa0337f9b7a63594a7c68758c3f38183f26e7da9a50214ddf9d615a09230ea89dead77ff8239198bd238453ec8c88a44886462b1ef7a58dd5c9cdae0a0b3bb6b8d79274f39;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3b22362981e8da634577c5ffda20f01c626f352ccd942632b22c7443166cda3d9c6ea3fc8594c005bdb8238b56d8bbd6c8c568fd990c724d69da033ec2b497d47bd449b0dc531f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h238c4bd67e8b7965b9410cdfaf4ef3eb7dff505d72af4dbec6bce3a70496cdcd0048781abf9aa157d602466b23da3652ac1c2efd9610e85cb6ee2cb6676fabce7db1ced541a19a0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habdc44991ae12319340ed78b40e9162739bc5557f0f5bfce955fcdf37558e9f2b50983fb659b441218727baf1698c469948d5d798c0b47e309c08dc1ab6a5096262f3a0500a51192;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47f089a27d5b99343c6fddff32c8a29ee9efffa1b418c8bdcfb9c102a3cdd552e528773dda8cc7eb6dd63890ac3ce67d9e2affa26c4dd5f2b7269036065344ba6bd0aa801e9c1ab1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd00d284066071725266687265d7520fb93679763bbb3229b71f31a99973958a816fe015b5807d776f61db59f30bf746369cefeeaed67366c4e829266e09a86456b9413e301d2cfa6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48b2f13270c374659d9fca1c88bae3a16e1ee149134242e42fdac6e23a355dd6083a7597dd16432462a0bec57cb51fc23a3ccf6e2ebfc8530d2106dec9a9420d96ade38a95e5b388;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a6ca4b014f34925b06579198027cf3ddbb287b8789e24e3f71aadf4d9276ad8e2cde0f0b416b274a0a7f257c687583b38955c460f9f27811ca0807ff9fe387a30061a3a8d7e788f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0ba9acb43cb6e7a62ecdb2e9436add219871f0781e0ec57496e2c533da39cd9e6162e6aafb3e762d4b1120f8f4dcb42a3a5ac14c3c72dc79bb0ac5f0e28e602e6ad2d98673e497c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h340c54b1672474ef414ebdadb21803b6bcb99c276b108d842404f961dc9ec3a0c66e23e8888e874d57dc4fc5b8ebec8e2e12b7bf2e7e4c04cf0cfb87107079ff1b52887b18bb4195;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8e8e694fc4ecb66b44f542cd014644e0ab0f658867c26d29c63d415de0a50ece0b800aea0043c217c0991cf4b6ab9f85527ea40f74a3e7de3d7d26fe017c424aeda4a202833eb3d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd96b011b780e8a880dd3414c3f945c8f1d0682893c106d9594b65cfbd02ff9d3b397eba4fce9fe0234123515e8dfe94d8390161552120cd18425223a27c635f731f9d44dfe7f608;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7108d7f6c406578d2e9ee609f3b76253384149cdfb4c5aea9b18a46c6227c5b3e7636e36cb9812e757cea7db21af05bd1e69c133ddaf16489217635298b117d5919cf4f543b27067;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha236122e3f43d96193da6b1f1820356f16149b216a56b32afa9a0f18305b8cbdc4625d11e4a4955a2ce3fdb8ad5f449c65ad2f94dd40bb71ec740cc91242bd47929be9e399a8d66e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d3e98525bb847b0ba4a98c17592d12bb8fc7ff55fee32ed325f1c8bc0f7d3337e096d782c45ff3279eacaf0a3e5a16d19079fdc32474643057888f06f8993dd31beda10a2a2889e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a1534909d4fdc52fb7334d5bbe31c4ada0e98e5c3061826bbade50fd2343ce58128e85a59396e520e9fb9d2ff5fc1c787879beee792828625a54e8b84f8bc4e4e145c367749b002;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc14c7af6f946aa6b9f27ffc313ec93a5e46c520f475dda6c2e308870b9c6e70b741164f197a948aa359fc8a408293c6e5c0ae093a1fffd714fd3d617565ed1fc5c88328e138a0569;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha745621391521f54901a66cc4f1d44bd81ba2e8c009ceda710dff32e76bcc8c21b2d7b023fbf795597278ab8023074e26ea81e4972e0b7f5db88c325a459c9a8f79fb49d1edbf70a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f1f084bd0d5570d308ac2c0c66d10cca1b86f5584ea946db8291e656a52d3a92e084b02c65182e651dd89f9d2fb9ca77d58066839692e820dffaf568a8c2610ba948498bdd38a46;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha856d5c83d75086cf010fadc3ce3d4ea1a830c34a276b398ff7063777609732ebb607f4a7b477575054246b28062f8a2b5f6244433e79faa4bc8315e4f1073608f1cb95ed6eef8fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd223f62b67a92e358c1c89e74b786814ead80ec480fc1e65dedbeeeabb11f8a15d9425bd8d31f278c411209f99715f360d1cd42166d434b2c8eeef86a25fb0339911c77689cf0e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81f750ef0b2072dce843510f7bdb922c55ab08af8862ad1ff3072688b8a2b843c9a29700e207ae4b3255bdded3571523c82bbb491787955947a65a6554627ca4ccb3987d326613c8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9bce8b8743693bd3519c2b9637a0980263996388000c9699616da4dbfe2edc44d3d6f2f3e06f4faca96ceac538dbb17903db764d621648479de2beabea4fbef1c68a0ec822fb425;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h101bbef9700db1c5bdc36954c0e606102b13a567cfdcf493752644d13a61860a197d7fdea27294e2ea81303997881cdf923e7095a14d2a1c5e93ee4bccb54f41da2befb07ad44511;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ed96f018ade4bedaf74aeaa498de10977495e401de8d97ec6aecc5f09e0dfcea6c33a5d56581e89b4c3fead5c68ca962a88770668cbbce4bdef12c9fded09843a074232660a0e40;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h545c62995825603b243a1c8a5e00e82f856d0ff5148df04feed9d7b06e00aa7ef39c7ddb4e0393a75abab47a9db52dcd05163d0560297941348564119ab6db6ba934c5485b83cb57;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cb812ad8b3519fd1263b5f53a7e7d50c3d11ac1ecf4a8ccd0750acedd9f5b45297c295d5c503f4b52154014f30a7b11a45a6f31cb133264660264d6fdb9c03f0f68d2dea199607b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68c864dbab07b6f0109bfc172f68036b57d9b661e9d1f43e274e4e1f6a135ec4281dd98c86f587f60f0f8912e024e474da26a3c73509b85084a0bece352053c897a4089ba404b845;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd68b8182e10377f618afcad26b0dc06caf14e90c0a83fef5af88ecdf71d525ee601d2f8a230dee802cc6651e1af703ec13e2d2916c7c880039fe04ca5b0bc76cecfe2692a1d786c1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cfc31e24dcb13039c3f399693e82cc53c135c544a76ca6d4c9a2f3a13fa96a6b156dd72279f3a3e73cb44ea6ee7c14b44536c8273442afef09264d13fdb1ba8a881fdfcfa13fb15;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53299463c591d5412192b2c01a71f7354b89996b94b228f860c62076457389c8f9548993be1eeed6f9486582f87f8b3e9814f2a21e53bc22169a0f706f86e6afbf9da45426961c6d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0dbc9b602885da8ea15ec886386b2c10154d6b4bfd036924df3504748d8e02d5ae9adb30aac3108d9b7554873cb39193b86566f2cc3415fbebaac91485c8acd58fe09a507436ac1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7eb84ca812af03cd52ae97e294be7c151e867c80f43e8ce3a6db0dc704bee07bd68f0e025ea020bb72017715388574e4b197bfad63acc87b2f179d475b97980fd189d013b18f3cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3de6c2067088d082130e0f96f30607ba8ab1d2ad40b23d3d03107eb4b2a0a7b5af23b2193d02c1464ccfd3e5dfe1c781f32b75d26e7dc46d5435dd6315969a440ef96f85c8f192f8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3a5a8443287fce64b8bfe1cb0b44a674deb8b449afab2899babcd8baeb9f821aa3c129c261633e4ed0863242ce822b118186ef6365b81c154b62f8cb66f1255f80473de8f25261f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a91fbf4302c658584fdb38e5d3f201efe5691fd1ef78f5cd4c5a3e3207256a3c9ba5abba8363ab9c8997f969fdaa01054cf76284a2c672a378e2071936419b58eeedd57bc6f62e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9fbe67ade81e2565d973ae645004abc20e677107ff3143840c6f2a645b46827ae9e03266095e95bb035ff1b755b7a4c8f9beaeddb4719c1008a537aa1a074eba11b929e23031087c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h213391847834f14b973d86529c2908475e482255d8485c5c1fdf449789ccaa5bf3a0ff68a8a246f9b84edf33fdc4f33bf200e9c26ecc394cc0b3ae3fbc12a596c16e272d16f6613b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h265d24e3a658e87347222f10c34c24c5d182f25d558636165d6a291c22a4f7e11c0bb3421ba5662c6fd5be5a10339e570acd982ae3f62b1255648e49699293cb873242a926bc3b60;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hadbc8a9a9e9a9f8dc35e6dec4061936685dd3e1a15f8a1d46ab8651f1617ef17a689f0d9eaa88288ca2006d81109c0b5e5bcd51b6a85665612083ce742b2539a39cf0be4a7aec0c8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff10512e0ecb59a868bd6365fc61c0cdbc827ad9a0229a5b275eda20e35c3103b13b587ea2ee06a02c765f832ae804b3ef40c3fe4f794db947862a736de39000e8e90adf63dc98c5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7726769aad8959ff33a6c6647a6627f922dbc2c77bc54a847349d4db30af49bf921d6b02f1acdcdf26b6afe1a0416ebf9304c91dbca90caf1a3f291be7edeb5bcf85102180b63b9a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef861cf5559eea445ffbfa989c559da7ea602b22140db8ccc9064a8a296119169dcf7024009db391eae5732b6a732f5e01f9d45dcb2d72f006836536cb65d0fe98f0b6f67ed8ef37;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb32ec47d2a215360ce5c903f52c7493a5749ae4df746ea234527c5ef87f9a0d88364b7269419927e291a9b32191606cd619fddfb95e1e70423de21c869e272d8165ac16014e889b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h726fa1730a6a054e8ef513cc74e78f2a0e6317b81bd00b2776a606a38c804d133166dad19656a8bdf681b0d8e8106bea3b3d51afd661238ee0822cff0b88367994c87e7a99b4478b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7268ed7d450b124d7182957cb3d677917dcce22e8b2edd57651e5c7cd795475b5656ec99a346203bf6d48af3adc2025df5e32bb40e79c0740dfbea1f7254746e3c4bd6f445252a70;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5086c39e82eeb8f360814e7266169e360e931f6b2251adbb3b9a891d67dedcb872f749b5c8c8185a5aa08a69af14a82836952db5137f3f044387a746b321f994fbf58cc621b2a2bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a27558579aba2e2636202d67892acbaf5312b825b787011896ece5237b6f148e260687a7d07a7a2d5c600f96e920802c64e2cdf43b668da301716b7ad1200f4a5c674a5e1317eaf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a8e5511027b75efae29d5e2f8b81ff6187bdd896b8a3cf805e8de2c1d51fdf85644f0fe4e13cb10572168449a4105fda6944f313057aa24a24c8465bb745e5976533fcecf88507b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62d753f985cad30eea03dc36848462e1010adab729b44acce3b9f920fb717f78afa79d3c011515c453063a2ea18b35fbb7e0c1db8da1fdb836ba8ac3fe3db041504f7e1ddfed1eb1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d51a4378f39d9ea859eab1bb47fad46fa5dabc5c08a832f2a3e85f97b433a96b27a532959999da20f4ffd48c9bba5e63d426b9cc00e950531db1a77e12f1556c5c06c4e89a4bdbf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7ba9229f79f183d0bac52557b09ccc4d8fe1e25432fac29bb0a62a60a3637239f090d6a0577480ed5bf3829d810312a334c0220f4b706e6c8e500e551cd5f8ca04eb6a1d106ef6e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5324f72200718b9a4649e64fa4dc833fd8b8cd7a196dbb63d07622502ff5b48914d7dbad39d3028f64cea69c778edd4b5a4c9eee026a2c19541eebd31aeed7a8798d9db00a1c0d28;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h209b2fa3aa6ee5bbb27b4793d1e48291786dbe9ff10f6f30863683747259c1e2ae65c6ce7049551157e7385b18eba361c89bc9df1a793b33e19a90510df8c1ed0d507ba8a6d31828;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb880adbfb0861bbc38295838c690f45bb1bdfbaf45f6e59a50bf7543d1ed45a01a3609e9127b3b431788e0bdf45f326192432b7236a1d399aa505c81365819fbbe06ca2477ebb00d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8e85677040a658c460857dccdd8db31559a6112afcf15be6427934b823fc1bbca937dde7a4bc87c4bad2b6dc5c1ca59f7edb28f9826fd4d834158bd315bb81aaacd20f7dfaabc1f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea9d67f59c6042361a7151542a87ff9c1d99ed048dd9141a98a52b5f099c07f35aaa7711a7cd75aeb565fb6e8fd6a49490e4cd74aa7fed295763fdb766ab4cb1391cb7cf11d6a351;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56634b108221aac1dd45ea63068723a5bfc73800e25dfbf1b21bfaf85186c4b904bc8f22474b9a7dc4e51c52572592cf906192d81ab844d2eda6b87955632eb624a0856381eebfd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5dd8942a1fd6a6c4c524a7f98eb888619adeb5c2a190e8f54bf8492aae5c6e6b47a1046edbe463f34f9dd5d606eee98a5575c44095cf4b830f22c8f97d918310b4ccfb8ff34380e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71b1c9d3ab92198628e35bc06a1502489186c79b6b7807eb8c192d356a87633f0f917fabcf8cb3228af94c1fe1db374c74bdbcc729d1ce8f49963a522ce7251e891e61cd60b97f85;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb9ca655be4efc626288c63dc492328fa019fb24054cb71565cd91b65a6214f7aea964d0f0f3e6d045c45211a863ef48aaaa9206a08acc5b62ba54713ae0fe61b2e5edaa17457574;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h881646c2ed31af0aa85838b8271635407bbf64aa16922a778a4fde6b559a17532ac0ad95595c996f61cdc1a85bcc081b399a4e0ce086414c8ce9336a096916d271c029e2958c30d2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6498293da8380bafde800c10ff6527e6aaa762e93ae13464fe652af09ef9d07ce1a47e25d559d32cdb6a570f4544c15e3703658f730970db429877c01041092d93ae4e83f98e49e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d75fac2413c569e784d9e948d2206275f9376a43483b0473e43391c44519f62d9203474b397fc2fd93bb358abc312f176e258168870cb580b96f99ba5eae4dd05ecd94e5619c947;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2a3cb8a9c45820637fb9519572fc11c740974d03d098bff55e6115b48e63f713628b91622c5ad5880c293ceff7ac169c64c36d7d49d6e34df29cfca79ddd09f6191b7e2102fd65b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b0ed269607f7add6622c04425f156203d6db0e934204232c210d68b1b3460b8087d70bafc1709695972e73b15116fd95da2265956936eb8be83c3690db548dd13f4dede83eebb83;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f6a5f7060bb91d4cd6df2365a02a48a4496c07868299d307553af8e76f17414c9ca6a933591cd34b6570c132b56603f89836a7423b46cc403ac42ea4a389cfe9c4436924b9c635f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a498ee3c99cc389a3cb27eaad03bafb16355b0723d694b0e6f4bfe390aacd17fead4b8301f212d5539e21cce4266db5c19efb4b57c92a036c77d990d9c3b39ab1df916e64a166c5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefb989ef0a88e68e52ecc8d4e59728d734a73c23f55b041c1047452ab3296ca7fb0534e0103cd0df67f3c5e07eb7fcc2a03ee605270cfb31eaad40a5c740cbab9cc7863b59716ab5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h283078a4d9db85bcf54ac0bb16254100df76751c92acfed420dc27d21b4ab4ac9fa2863f51831e598d81ddc37f2c5b8ab6edc433bcc21b6ee8044c72168376a057e8d6e9b900feec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44b69f0ea6e926d6abdbfb6970c6b12e15b4e792c708132a71b6bbd0a0625be7b3fba8357b08a1cdb0ff84e36b9ebcd5f5fb12a528081c6bc6f604b686f8455f31502c8311e91d57;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ce8aef5467371a736428d739d6670804a437ebf7420fddb5db142032171e74606953082cfede54f9fdc807b13bafd14fe3ed87878a9ec73de54841c8db08a7a6b2992caad3864cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4655dc62f6957f5b73c0cd1f42de0fa23aafa4a3af333e9af20d574973f6edcd62271e360ac58d13b0daf09069b46cd6bb7f53e124dd9ee5f73b6cd4acb4143bc51e383986927fe5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cb37787225b3c60855bb58d6e9a39fc58890bd948b4429572f13c835370aa7560c8700292afa03da45ee8cabe40960e20714b7de08cece1dc257320351d97bb9841f71113ae4b3f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3befe14eb95c3f1a9ce0afbf599e2540561f04a74c5283d9eb1f94edd399e92d311509cc534dd5b47feaaf82947d25f601836df08dd534ca88b1f1c3cf5eedf1891e8028e70d39e9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42a5b7e9bb5d021c2c8498fd4c6d6352b0d13aa8a4685f14e5bda5e25fd1519abebd55528469a690bd9c700581cb55611a94ac3ddeb65f300c60be83e1abb9ae81bfa31fc8ebc8b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h818238ad9102c8c47e706f1a8b9c8ec704bcd9e96fd8e750ba7a736fbe428b5da03781436a5f1c75ee4bdb3cdfd52e15f05a9e09284d92b305c8bbfe7e62434e5f74803661f84a2b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7f9a2681c03842e434867b965ae829a697ca66afdf0714f71a08a6dd6361bf55e46a9edb70b69cea72d0ae226d0b374147443574d15f33b008fbda8a5e1f23c05a32c5684c9f582;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf76322779eddc2192dc7ae9f123a00597dce84b5f05ad7c8a6faf26382239b3338976510b4f10e8f0fdeeab5bb4445be356ee6d93dbd94141df3aca35b43873428ad64e1701aacb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h146cf7c6e221b8b815a827d8d57b000d723df7666820cfcc2348c981f5da6dfab371459ae0b2cc263a5dc898a9afbbb08f6092c000377998b89ef15a3c9473f59ea7448d27ba410e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47f070825e363bba2231de41c38bedbd6d52a69ec694f4ee3af5b8bcdff697e67f50e628184044464da2933572c574ce1f70866146f451409e371180681b058287e5697b2ea7b7e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb6fc72aec6b8df0a2b4df00d42baf313175ae580a433fa9b779a719f73aa30c743b3f05f5023fb8b1deebcfc4be077e9eb953293bc5a11b3bb04d056997eda3ea999d6453db362d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42d6de2f95c0af534cac32da40e35c84b8175f417d3a5b4716fa27d22a59661591e1a625a826440f14aab7dec27d723c4f87a1d4d50a520f271998d8a6a39e2157a246e579e8485b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h535ed93ab6a0df387c1caa15c917200435aaa4825eef7ef3d8861baa7ee4b606b40b9e987e140e3d67552487a309eaed212910100fc67d7bf4955d969cf113ef49223587a532cfc7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f36a3c78b5c332c867e8406952bb6b6682038c671d9ff6c9785ced440c5be27c1b8d4911b01d5654b6326c374409019e68cc9840a6ce03bb7d3a5d03e58e73b2f03907c9b64d7b0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb581a1d8ca728257c967dd3b524fbf938160b806012c7710ee07bef245737440d002574b6899a4e5d16758c6630983cfc73d61e8e0c0fa37a8de0f4488362bad870a234be7b60c28;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac74a6f578a193a4a126f573e4abcc1fdd14bc2fbd217e29b07b1b5b06f726e5a95757704fcd0de9e6412d950e3362158f38556215ad1589362cc2fa6ccc31f32d761078d365ea10;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2226a26aaaf63c5952ae72f09b12de2b19be2e15efb47396621e8da64de69a0ece82f61e55c815351af968172476d11f808aa53f32c2564a781d1ae6b78f4254bde6f33e81b25bcf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f836ac5eb67bfd4482c4ca56127d0aed97a3f644fe07f81f135c8e5475a98f1b6af634f465a033420c8d527afcf6dcd5d3fdcbee24549073c0b50aaff522fac1d7933f1c6b50cd2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbfb05f77d56f546a8913c6448067f9dfedf7ec41a67b0f0ef4056f83a06cf6cf6e5b2631541e9a47964fe34d6e06702293c918276913e053694cd1f069ffdf1ac651a71615e39c7e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66fa10e9308ccaf0cef4fd6197a7398143905f9b7de3d0be3e7775da516ecbe4dfedcf7aee3faa3ed42b71647ba801aeb7ee64bb80d40e7ccc28d8ae90a07256e1f19c2967188b35;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83ecaa1e798e258d253a6133a9a6a8789b30b43d1f1f17dc1e094a9da1b81fbd427230ceead21bab6eda2927401e09c4a3f35409537b46c6c78c9162b8bb9518ce77f3cce27096dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h337358a2f0f05b45a6122c6376c20fe7181f32b75b7c960540f8924b43ee600896eb8f427b774efe752c3a4cb2f3906cf7d0c2928173f57a7286ab82ff41fd690a7d109f1bbdcea5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7fe72fb8edbf4b3c01667a5c44438d8477111a144a8e2e7f17ad6a7ade74638a4888e721442526e0f1a1556ae297615e25c19e0a268eeceab4576af3fa20c3912b1efc36e081163d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f23da37d04d15a10d3d1bbbc26dcc1fb64304f6c897690dfeea99236a0454ae0c4a6d94568f7d335df3ce05f062636fd8e279b5a64340c4dea2447d4b52d78d15373f28b513a5ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e93458c155a83d6bf3fd66b2e553a6f563d3d2fdbac281015e49b858c312e1b5826dd5b31f080f9f5d399f8cf4930b383f7ce876659eaf4bac34ecf86ffda855e626f74d971d092;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee59f2fbd5f167bd19902886ad494e336f9936f1bcf0ddb8d98a162a9c2f886f652b01352c1a34f5cd12051b789f13d7afdeb1971f88d74e9ad9613d0277c0dab3e8439d443f5122;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb1f78f876731a9de6ec3930fd6c22341f9a08409178c078a09e1d165c18b2023d0b10621d915a702019ddb5d3c5ea27b14903822ef20c492cda09d5ebbe5fe7d7848f9aff7ea556;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b2c05bd2ee81c6ebb9765b3cb1313e1a992df77f2d026525dfb44106ac7935f33a69d29475bef146ea485bd7ed8f352389255d9efefe408166a7b1fe96922f284467ccb388823cc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce93f192665db0678de283704b733d6f5811598785d0359bf6bc1346bb82219c734efcd545105d0a8330929a6648197c76e7ce3dd241c6879d08edd041cc95ad88780b47f204944d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec0970348b25ea1af3c050d3f5e16ea80f0ce32abd04087588b7245ea58fb9949802ac80c692c1f02695b5d296541b8accb20e0774b22f8b89fd0b7c64778f691907bc041f2c4221;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65013c7ecb724b9f22dbff78e753bcff61310dbdfbe91236a7ef1d15de44741149c1143def07f8a4de78e0259ebe0bedbde46d60b25fdafda47e4d286580cbb3ed6718d2d5abc6ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2aa25d2a032492997f05ed2bf84e0863bc1566cb620f3dffea4f4f14ebbcd63d9f7b15bad470fd4c9b79cc0bcfc7f7a7004ed95e11f55faf451e699e870d59d3c54b4e8b603c399;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8a3f1fefbadd0e4e00abf22df2bd953ebb45c0d0a2edd7838ec581768f358532dbf69ed0e2f509d3998aef57295165a82b95ba223bd78f43f6f3efc169265f23064718473e2ede7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11e1ba942e671f816d326fc83817ab77f55eb6bcf897891bc40a999caed74093338a4044aa89e28f3df28f172e4f68a104082bba871eeddd8ead956d660367bbbd576b4ef01f11d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h472b48858e329c24c37a27fec0b931d8db27285ac4594c0423ba0c01487f2d58c48894387f4b6ab6e86d47957891992f61969c854f3bf9a6e8032fdaa810491f09245705e2d0afe2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h450a57689b0efee1d38010859aaa63bcd7f642bbc3590f2c4d68740a87c39f9bc0dfcac21852b392e9cbdcbf39c61f90ed3f2ce7a8546f9a502112a3b09d9d624187e238afa4b965;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b4c258666d3bf59db66a6fa5e6a618a04ce0771df513b872343df92adc7a53996b5e72089bf251b45a0105168f2edad765ff588363980e51cf953415aa88e1f2b963bbf028ca9bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6598f7315e71b9ddd399dc398a816bf4f89e537358142c4f2f5001d646496728728aed3ea9ba0195602eed1135a502d6f215bf1e0ae149660fcd0f76dafee723f4b6a18ba4574191;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ac2846d07c4c3a564ba35d45aa9392571f7a5dba40ae02ba7d8f73a23887426f09d0c70d648849728f295d16ade422fc270cbcd07d68105e5b519e84310dcabeb4363298409da42;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha80891b85faf8aa5438b35816cf92a590ece3bf2c22cf1f957fc95263b68c9845fb194992681cd114c0b167f76e4c40d93b69493c73a57528466101acd5a2d2bc98772ea3801aa1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb40e1609b83c163a74f28067a6a4e6512eccb6f02c7589795e55af4d356e9f493c1a69dcf32f9c3d02f360c94b4ff6ede6c94cc6220e79161be2ecc4345db39754f42ca27c2e91e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6cea242432acdda530790fc37404a924fe626b29fcb33f4724db6bbfc3ebc2230e70e024ef82fbfa3203a79888c27a551b4e1ecb0cc7c995f2ca102cf9dccbc709046dc6a449cb0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3e7761c57f61ecd73505c8f4db39ca9b8bb14cd3809da06d8fd5ee1d2522e046243af3bde813769ab48a5cf7e155ec817b71a80499fb893a5d96476d37257c1ec15b3baa00fed77;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5e0626369e9f0936d0e1e81b60efdf66e2eb0c5b79c2945a3e3fbae0675f83bf9efbbef91ebf9cb2dc63d228e60786640f2fc9c139c297482a2999b5a0354f50a96f5b657751cfb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9274519e0f91a1b18e305cf3fd8c2bd62fe6fa0371585cf534722d80f2f98945d0b8351b431a4fc79b10e77293ce82d01757d0db0dda0c0e5e58737646893eae43482b50327a1f9e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb25bacd9d276cfbd7df1902c98b6fd8e090844cd1d0d378b79475ff5979f0916f254c8b346b7267df977a0658d4a70b75d5362c20832ff07d2f5678d51f522074df1b4bc7750d42f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h888afafc1933360080cc9eddcc8e09c42b9319246f9fd7a6f90319b57fb3e5fa87a60cc431e3fa9565c02708954bdd3507fc03ecf307fd7605ef907bb0130e65957c38e7dffd47aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha687f48570943e58d905fb54d1dd7bebadb464287f87a7158d238cfcb333330e733f46bf196b535d025d0831bfb846793b0cc6556f98235dba59160a17499c68d03e4dd138842e7f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h977170b6ed412ef83f5af2b209e7a86f968487f48159cb7fb1ffd9325397fc8bc1d9c22f6c18e31ddded1de1cccca94c3b98ae055433cf0dc4356c28749b3b1378bdc8a469f54a29;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd74683bea60715e635a19d299904f0d96a1a9c58895b056b25fd424c6dee1da23a94656787eec6bea7ea81a4e0a8616bb06eceb0a79d10e2495a49a7c0ea192cc1593695764d6f95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde6e216eee343d0f1ac61e7bb3509c8e0b5a57a70e01a308091a3b017b3ddd02106e29b936eed0c631d5c8d8f3913b1a492b9c80ba53bf1f01309ce684a02c38b26d32da66b75833;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2787b23f7db6b4c9717924a3c2b762f871cbef8721780bad42b756239cb553edd8ddd04c6efa6bd717b45e4adaa6ad27d22b55f4962876b70f59e9a544a3ea6d05d3e180f5f2ec7f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8e242b926a2559dbf9007ec8f06da4053d0f37494180112423d4a1799bd29a87859bac00adcd59339d7e32f0bbb07bc1a6be8f0e45f0dff44c5da882640ee9c61df952f5cc432f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f88d240a87fef1ecfc8ac80abd651f658bcfa24f71b5f9a5d6c4a06b3e7371c49133730eec61b7a2ffea8a4bf800020435be5e191dfe90985e3d68922f2950e2c388415a8cbfaae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd098b8c8f179a27da8afaa05cd5c9b7f7ef169bec6543a8eae180fd9899ee46575a7914a388d78e9c57657fb142942c829545b15676fac52a6110f1b97470f1bb3dbd1b959232adb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f55b72816fbdecc79bddf9d94c6e3efbb6182f416de456b37d31251179625604225c947dc6faf94c18bd667e128c6fe7634b71618bdbaf64c3a16fc66a29b87c5917fc95cedf65a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97b228f375df0bb7259ccdba0e639d2b5c685b94170c546e471e7dba9cf49ba839e30165de08645faaf7bd9d7347c52f336c0d901a7ec76eaebce1a241ec6f01ca49b999a2af17c1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc856c0b9f3f43bb62ab685e0969075a4b8e5bd641f83a9e9f6612503fa98b32dcd0d2a5a6e6e3851c9c74ee5140a7426b24823a3a484f97b8ebd94022b35080fcb2984b04c822861;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d8a0ce984b16c4958a534c44430ef9c4e43dfbcb3e5f2aa1a98b5fa84c78cdbf4debf32beb940e744ed9c7849d63534c2c2979a48983c8ee1137d2d4e88530ee0614c084901a362;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8e780726ea7f411c37bca75bf5ca3fb767f3ba595e060bff63f47bf8ddceb16f79b38802132acd2af9f557efd26c3f8173c42c44eace0ccdcc098c2fdc100f423f288cfe86de6c8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9653db643489732450f369e27777ef2892eac4ab62612df0b09479a80aa3de6a3ca5ef0e6b64d5411797638d345cd451513e258f5d2a5a6cc350fdbf48d7e14ddf5027b37cfd53a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h434c0ef869e6dea78e658dc89d12cb4f3de7aaebfda56063f7865f5e033bbd65b809f244cca3b3cfdf0fe98e1c6077daa951fde2b4219cf80086b8d5d1d39e647cb9a6f765068d96;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61d796ed196d7ca64f0a05a3430c872ebf8e570fe41cdcb3e4326d3d121658cb22b678d04a18204a9fe9ebd357830fe4c75e893f80541aaa43b95bb0b1ae2d3640ea64e3f7c19b27;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b79ee2fe1fb9d69e6fdb3b6da02cbb0e46b4be0481c7d71284b359fc73865120ded06a4b06910a6dbf8c57a8db886d0a28caaa050cace9d30fe06d49da4d7f7070e56ca7f92d562;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc40c331af784d70bf77adc5a72d2d603357ffbafd2d0a1fcbf46c7cbce232830bba7a318e4bb2fa52f1dd133a0a48f14f559f8b82c629fc27843d0dcfa2869b1c0481c25ac226e0d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd4d4f3a748f2aa1d263756e8e841f9d7bba1e742010f636c1938110341b72557c280cebe7940aeaab141a2d7e8ba27e98c739359ead54859e222c135aebd9119b7f2d2868b970e0e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ff68758667a577a1eb64f6766c5803b4ebab4d1455b545c4e477e7cd4a3578e5121950b1dbb530b329dad545854b694219650f2f535ad18a87e078b56c24063982a436f7c37c606;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca3e783009762403e182ede0be619df263bf77934bfd2228f4de5de556978eda305b6421ec7e3ad9e3439c949fc938766b8816efb48b29ab16ea7a610fc0f8fa408574d36c74856;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29e5ecb6e3c838a0c0b3877bd4234e284c3203c16a4ef33e2f5072bf9533de561d2c826f34da0f068896b35189f3ecb7c9ccd61827da3509fd5d40ba848f19c8cf908736eab47b53;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdbb9b70bac9bf39b28bc3cc2ba071b436b7c812a4581f1d5ba4ee247e0f5f120d9513d4a7a8ccdd39492b48c82726905814170c9592abfbaac5dd83440a03f71a942fbc10e49d20;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h386a2a670dc744351aeba895697af338456dda2cae776cdb85b359d4e99a8852f1db30fe6e108f5f30fd073edfa8d1597fa0a2468533ae376936cf3905001c021857e4b4c50245d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3dec7acea91cb1ee5b55eaec237f5f79be8ddd0a359239284a38e3b707c9f64eb0cee3de79d227f4e8e41d6423cb055b41329623d4de23a9ac950f04dfce88ff9664837b2f4a40d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58953fa27b2abcd3691bd29be6042328b73ab306d78e771739393da7e0e729632fbf7c281daaac3b8c6866856582f944ea83770a6b8276abe61b06b6581eeec8d9bfd20635f134aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23ba94bf3bbf66dfdca5cdc5086ac5384980ba2062a749aa38afb64a8d57514a1864be07049f72082e94013eafd933675d84f53dd10ff34feb70efa931159e698458daf1ff95ee10;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h404f1b37dd9d6359f92e1081acfaa5a30e55683dffe9ca82bd9ccd765f7149b2f750791d02cf76dde66ddeefc6ace00542b8c294fc868f103fe3cc4e7ca2cad2347d5a9637746330;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2b23b90cb328c498f770e781614eab79cf5eb0311a4785e2a35c6b94efb5dbbe25d03e5491528e8e5e153c36b64d02f89f86c3cebac77c79c4b8e379b9ccafa19b49a860310c5b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2da1fa9f242e69c5d354f9e80d2e1279dc905c0f5434618b09557d6ecb029ce2bd94b0e2da57334a99e205ddaf231fd08276a96337e0c1769169adced35691bd5ac980837b5328a8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1ec4f03a5b94290a3760479a0e30f8d2d08ef1832919b5e41f319edb906f1fd8bab106f257da69e35a36b60ce185a6e3a74882dcf31e115f367ccbab9169fec6aaf74df117bf1b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5933a702bba43aef6aabf00551933e12be9dba8bda42bedfdfb10a4e19f3816f943b1a9b2c7728a758c38525ff17befc03a448ffe5d45c763b9ead8dae552c45d9517335f7583715;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hadc3c3d25e2e554d77ca2ffadbb0aba4725239aed431e3034aa2e224f54ef6effd6f137529ce644632d9cf65da68920a5a593fe3f9ea48cd93d732aaedb8190c745f7b7d0143cf60;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce54d6f426b7f925d5dfa7ee517c582b6d4f9f7474db6a84d8dcef02d3b9d7c7e8cda73ab7679b676ef6643cb1b25dcbc20f485070d2398cb79c89c3be039915110b58323826caba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h825e09de0ca8aa62de179ebeaa48f710cf4daa28129a59d0b3d68e0fcbe7328eb76ac34bc540290100fcee6ffc29bf6421e789f401b02a17f46f4217e4c695af76f2b3c098d116bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f7af5c0bf1c35e602dafcf5644d9a7fb18118fd8a422fdc7946155c719c91c82163b4d40cfa88bee4efbec6ffb566590a7351ee96485952f368ca6bceb83909d9a8932a5e8e36a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc109dcfba048901078c3a5d559dfdc980c407064111db5143b6825292da493b536ebf8f5e004294005dd6d975add420d662d1b70cdc77e6c2a1e73bc7bce13049f40628d184b2cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8bf8d13d8b80ce95efa12b5ac93af52da6d1e3b08563ab2f96f30ce961912c0d2e1f6874335e85796990d83189e98f3154aa7a554db26e13b524a99fdd8f49dc665bef87d029dc04;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c64b8b68d8869dbf3a53786c959022fee3bd915fe4cf71fb56ea9d39e4e86e8ceaa5d1a31e1f0c293c32e34efb8344188709561069df2bbb49ad1640da87f6abbaefc8fa910f21;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f6f6662e434ab7ed31a7b3ce9b96878fc2f600f55b59ccfdfab4af460a3a66f4c0748685417bdff0b7bf7f4fa26493dbe86381e282b7d06fe5c2b983ca764f1ddf326d372e6f259;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27017ce8efc04de9d7dffb7487fcfd422696d324310e8860bba92e173c4c9af54edc545e3fb62eddb2d4ed2f3cce1afdddc03c2621a545e1e0098836e4f6a508b938e54e5114f259;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a2b8e704b5d803eaf080abc480deef0e3c11fe76618dd46ac9a32fc02e6e65063b22f69189e667040c7ca26513f010405769bfbdaae95613a3eef9ffa8d7d534e88c35c157cfd07;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46913ec6225ec2d0d42111255447f4d9f0e0bb92f73a541f596b6068e21e8e6d0a1a2036aa17adccdca404c69a5c0562ea53e7385d558e35c93f4dcb83d75848783da125ff310d4a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdfb1e5b5ec542c8f1284892a9fc825c9afcd27f8f9219a199d2963bef715cf90a18d545bba9f1cc1d3d962d824372b820e952d0fac08001219baf1eb808c2d103989675d316e5fe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc921bc9caed6b8eddf72dec837ee2895cd8cc308c8ff5b66aa44f7480b3c77c75b86834f3df9bbb5d17b3673563714a5e6d668066300622c6a2eaeeacf971e57d0e0a5ee4278b7b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf19a857df8a5a3f4c4813cca5feb1e278017c4d81b09a8d7ed1726d6df7631d3630fdef0e390642fd99267e3f464c52f551e30f17c326f76372c12d447a9bb58d605c8224cd816b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7fb7bb990e129d7f40229aaef0408a96bad996db6344b48d4f0808902579fed44de31e0e752f3915272457cd9ea6aeb59057f0670240db69f028265dad5c47f53523791934d26715;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h147107a85a30e5a0bb9fc96d354ce020b74355c63436bafcb7f3246ceb7e665b70479582e17637c68081028988f7a7137f39919c32481e76303c0ded5d8993199d96ff8e6c429c8a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b9477eb5e3ae1933a23421ca37663964696b04fac633861291036ca28ef54350343812da93b3d2070807be4e21b9e7aac17cf15aad1dc0f6171b4f6058496d3b0df19b49382ccd1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha81114e157e9d8bb680f5d652845c677a0041a8b95373d89c153929ac15804f2b2733862895a83841612448424fc949160ffe8d4347adfbe8c8e095aa847efc817e3c448d6ed82f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b840ea094c7e89e225528055033e3a1a1f4ba109b4d499393448675587840fdcaa9a11974b93a1478e7cf66d7fa607b0485392fa03f008b9a027a07135aac349914d10ed8b5372b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h768fb51689e1f2768a72e24489b8d88dc8e8ee54964a80fc80658664760738accd20fd6e2cacff35bc9ff75088ee5fe084d6030f65819b9f3012804d33a6d25b555ee2079817f167;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3676e9f5c2efef61b980189cffba6d1c3d3eac70b66ba5dbc7c486cbb658d369f0e0d5a5458cd1b9222eda49a758ff67631c759b5346e239f59fcc325e5e6e7108715ee160fa194f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h818e1bc9c274935d06ba69b7dac552100dfa59a36bcce234022a9618db023e520b5d3b1b7432e6a01749a85950d43d9b5eb0e93bf227b25fcb6db67c348f88b9b26ab3563a454965;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3925d91ea134fd44b5c7ef30b499f366dfa077a6bbeaefbdbc11e3d552dd9de455448834f535a7790c1fc4292ed6633e3362353da97f40172e901ee96f16ab570fdbcc111b30f7c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1dccb483928c066255eb2183dcd04266e44276b63fd8ac55654562c67da17b3f543323faaf3921326cf8627a1b0878ffb757687db222ede24a0bcd460a7b1c381e1a3befa6f05ad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffb4d018584cdf91f82f34082b7ab65673b3ed04d1dbc90aa177813b7a4693ee8f42ac9b3e7b3f477ff4043ef32fcc6fdadcb3a2ce37c14ab3049d465ed5222d2930455882652038;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e69c5afdf12ab33994f83d0b66d61990aa1d87e8c322522ead2060db1b438b98046626c179df4da8f4540807c66321aa2ea54f0cba5ee85965ae196bb36cf872c46fd3db0d72943;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70bbd8ca61f6b39c271f0709d482d6ac012748c31865248c29fdec211d6f30856d70cef6105c586b9f7a85d47f667ba7427e2e3f243802ff897d9480250361e6e16313215af9def3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1d9d979d902ee9342a6ea77cace7767619819bd8bf87379b23f9b02f74f8097760899a67570f4aa061cfcbefbc9b5bcfad50aa8904bb372305ad00325bf29525f4d5542694150e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb21f91e04bed03fe9e5dbf11911ec043e872ed281eb85d4a86129a4a51b0c69bc1095ac08faa9ae4b9ad6b61cca91ba6644c913984f3b38a75c5ef8e9f6d838812cf698a5565418d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb45aee4f041204d0e343cd65f62c6793ca6f1369a6c34e6a4a39c5db7a4f47a90815d6e4838d9480368c8def875b88fb8ad7770e4171523a1ce85c8f377a869fea9f20b65a14db7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7591b02b78584ed9bf56914dc357451b64c1035cd81f9ce4c0e7b1c28eb1426f06b39816ee11f22b4205bb8e66a865e8e30aeff2a584145038cad153a6258095dea0760587cd714e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h455fc49f6ca2118a13950ec80d0dbcefab3f4133a8b9bd27359c703f9a17643eb3013287d57a82d4f2b145a5ea4b5ea380fcd195e0faeb8f43be7c51c001c43c75f4414ec3978d78;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a6f7a908eebb2aeb46679f700a6a84259eb1b8443be8ef52210a9b50d9176a8866e52cec84597ec5242296438b3d2f4acd0108983b8490b2b6fc9003551cb746c2a1479f6f26b08;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7912e2f28a286b5c4248ebd74b611e3aa690aa780d4eb955f6fa87aa2d42ac569a2189510e4e4cb22e200524bb0a1e0a66f44d518ebb613b5e7a0c7e52b9e1ea5c8edf617dea95c5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h144c1f2d4459042d60db0d0de907d0ce6f343ce28cb72b2b22e3d5e4e8c2c81046ab5c24ad67be5952c3adf7819dadfc1151ca7ff69e0ac9f40e8ed34b595a56f5fbd9ee986b7b4d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69269cd9ab5fa9a9985290b99c1f90e700cbe9bc35b13c21c2682711b06044a521390c815b9f957bf3a8e09ddd971057212c030cad805c70cb2b3cbe785f9c5ca9da0cab485860f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha974a84d0b3070d57d5ac2080ad904c83ff29fe08c7de858caef440ea5b740a6bd830beb055f46aa6ec91f84da26a58cb9021f329e26a0ec63f9d5ba097a421141ab33787df72df0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf18ea64e1a06f4e50aedfb392f862072e88f718ddd79822506011f2b05673234027a112b690f6459aca29ad54ede5e40b3b0d5b7721214a9f51a9d18dd1156ee91bbc5bcd00cc0ec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he72f0807b6d3029d5951afc73d4b6bc8aac8eaf43317c8048f72ba6874f73e460dcc515cef2451731f9934ae41b105475086feebc7d251aecec2451d2e6cc4f918254a719911117e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8061b103787dd2e8dbda5cd7aaf8d31df0312e62ed3cae9745df321aa479079fc6d5594d84e053ee348b42517e96a180c042f8f9c404d91e80b0ebcca26f0ca9bfbd512327f7c402;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3010fdc3a04ba9cf62e62fb4acdfd21267ba0ef87dcd5ca9b6d44098efbe5a6e876cbd01787e4c636b5c7d7ed9396905fed4d2e37ccda52a21f0ed31d64844180f5f731091016847;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6501fc59297e93309ec7073897aa310675f13ff800dbcf1e5e7a112e9ced4e23723532303f3ae6c19ace9124bf75d2d8761fac31e7ac14a97d55a48b35284010597cd529f8f3f09a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h173dd412e25dbfa39c344d860334480df3b954b31025f02f9052d655270a3bc1f582993c839b00692ddc3d3fd8309df20922343616e5ae52f97884269d31dfd1ae5f354b45e845cd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca21222406f1dc28b2e2c3bde28587a9098c652cdc923b048bf04f4fcf08b6b65680a669ba580039f0a8531f7c3ba5cca9d5771307df4b134952c994e66f11d54893a26891946908;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c6d84dfbed1821aa5bde5b7996f6f63bae1c00d2c91747efeec15a1d3915ebd37ef46717ea9c9017663a491865b89c41a7cdb8f416d0f973cb7516359a84992115ec0104f68a7ec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5094cbd0700f0eba0a50b3cbb97eb17a749706b78be788ec3f3fe51ec0ba293503a0df4e4445ea77fc03ef0352e6cabaa413ec4d902a3e65e864e22ad7a710ac6688244367b43d6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h746604c96ede59548e3f1935034176015cd1ba33c2455ed2e084e68ac720af0e63f08ee015de70358409d3b109be70c6b3603becbcc0244ecec53ccec2632731f12b6f8292c6d345;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd438b08b1912e7241f301f3b99680a5aa6fa514cbb0277b0c34372ee4352098253b7a644ed426651a5d359f2436ad7c19e28211d60aee5171382301a36888453d4bf42dfac1b3b3a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4300ff073c1ea956b3c49e5166c25349420659266991128c6928834d392b059eb0cde974cbe829ba476f7cde702d015bc3e55fecc5f0b3a525606ebe73a815e06dfd5e1b48d09444;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h162318f70c01dcc72e4aa299e889448aba439796516fcb5951544da8926492c625eaa93ce3aff69429bb655a4e12019160287440ed44794a4a5e7f159393176b31e0e3674685d550;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h253746f58be806345ffe08aa5043960f2e28f98543c94f32d397131325611cba81dfc9e0805ca37a5539dba596f5fbf0629376ee845821d23bc1ba7a08ff98d54cdf1cf3aeb70b0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77cf86e1e3a888e00737eef5fc95bee6973ae0d2d6abc7507f0b684e4629fe398b0749ef0d937199e54b40c238f7a4ed98f4fe6fb974c0c10851081a951e908c38761633c805488d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6aa664da02f52efe4271f73f83541ab3354167ca7c62680a9c1f8e7d10a02f957e76a76ad2394e207ca382567b065db3df8cd01501c09fb407cbf98bb9a8fda1f7a07a342f3d943;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e98f44f5dcbadd4ac2d0a6b10c729f499ca1379affad595d10a5ae92bf24164ece80b83bbabf90a5b1c1122635ed8d9668db53dc260b3927cd66a2c84616bb977c28360b487987b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3926bf118330005343fec6e3d03120ef2370c946bbf33ccdfe9d252a3964cf9093a8814ae1087e4129d5a640765923f1cc57a20fc3ed4bf65c65dc9f74cfe33234b2f7d4a3d4b459;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h179d56c977f171e715f382fda1813c05eb8f6f106c5765a6a7c23c29cced030dbc2482ad7bd68801a5df5bd623f3e3798a1c3d2c51fcee23856f9f9f2af2c507f9acfaccef01c328;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7631a98d11676f086d21442f46bb0547c7fa4f4cbba8cf51e105ecb84abdb0754f9f238daa28ec55901224dcccf109d1a0f960394b77c43fbe4a7d76aea3ed10499bcb3c48b5a37f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99d3263041ec147fa169d06c73a9249f829359df03c4513b1b510d13ca099dc1b6736ea32e85fca4d8d2dc205bb61274d350fdebe34b4feb4c416fcdd5f42e438c65f8b72615adae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14be2389f118f37c3ddb299adc229a2a4b896cdaeed8104e6617fecb7096ff21e9e89a4577b9bcb9fa1c3f61033b03c2762fe95391a9d3eb4988b06cd099a4e6f72c06de69bed9d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h363e4ae59ae54e64b19b0235c92d7c69b65556c4ac32b591548f51b6f215d66971fee3229337c622101d5e50fec331c42c99adbf3c9253d39c304d58517ac63344dd118d8d46c839;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7836156a733aeb438ce26f87ebe04fc0f76075d8b188739fc2f440b5a998432e6416416fdb1453d793b234b8913b00efc127837cb2bf4b63f76a609efa7f0fa73498bdf82a627fb4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77c887691cedf32bfd14041702c6337cb8b8e52d3b0d5708fb70b3774bbb0450c758c8b4df036d98a1a6ca11181c4bf654fd88bcd9674937a557153c3e3a3d6e1b270f0edad4ea98;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36b39d31420daf196d7d598b26c7952a525638631583837dbfcfd0170e92138e29cc1e4c91722f6d0f6d73f3b6178044810307451da55e9b85c52feb4bf869d3005f6463e7e45e6f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2423ef54525b52d9cbdfc8073d85087d1a2703ce86daf6d830b273aa27115a31063ad465607a9ede5f059cec4b008d3ca126cfc874756e1cd56c0140694a6671283e48493a037ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6105c668c755976506e7eff6b50637e82ea1b2e013f296b6a54179364a06bc19a731e91cd46857d8e1af4c686cd9650d96b384063151fb3b452f323030256ff9bb897b89efb4ba88;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45be2954047565dc5257e5db116ed699eceb86676591095f3f7a704faae9f97b14df72d839bb5e3240a28379c95206ec04409b8e06a17dce69476975c133a31b49ab33eb303b0979;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ba8e8cc4059d6140d14a7794b2717d6b964770314429fe80f665dd7ed59f793ebc133b78bf4911c547f1da534309cd860904bef47f0c1dfe7f9711fcbd0239fcbac61268d1c1294;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa0fdd63d4f3e6e1f4c51ca2c9c0752ccb6872fdfc093a6a4b42fd5cbfb519afb4deab6e6cee39c07e6ecb7516a2575604c3c3fd18d0da45c5f6f8a876fda8ffa29b263cc3f1dede;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc88cc12635abb8de3af8d8f8ea8baacdc98520d73111bc32e4d39c530adbc282898bf048228e2c5208dd496f939a2837d4c7c7deb609c348fbdc3ebab7f3373f89bbbc8ddab2e4e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32ee7e5246012d24c36cfa1974ce3815997623a31753244a36a81ba8c820809f3fefcbdb7a9be67910251670b48e4886fbd24a1891776383a96b9f83fb0643c93a412278afc2ca4b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9810a598e4a4893afabe9bd4e72fdd6cc9c7993eac3fa9ee53e05755bd4d9a00041232131f806b2259a8406449f49cf960faca537731c63a7c0dbe1dbb9347e105d68c69f5ef60c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6603e6a5e5d77388412fa22f17ef8b67939f94f670f62c25de6a99393e0381f0548318c35509ed530330ec4fb8e6db20c1748d8eff340275cabcc7b3fd8bd4e46093fe95a3e6882;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7169f113d4463dba45f67e54e79f5c19040be769a926d2f36f797b21242932b0b80a3a0657d6cbcb7734738d471ed25c2254363bd8304989ccb319e7a211edaa647b7f16adf4f4d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69034b698daddcf815fe2a735328edb634f6e956d9f64c7f07b99fd898c0cfa8dea3b2984d9554778f2c40c807a3221d7b6cc945ef5bd2eedb8f22f5c5c7c5c3032098b4dfc555cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hafbdbbcfd75273370e023ad9a6c24b92d83e6112abedfaea29b3356d7a9d048a7d4c830e6837b98081ec325e143c0e16a73bb5dce5918849c66917e5da64c0a0ea8123a18540fe06;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c001f537b6aa80b5d5b3f3c4c26f5789c111e10488356befe4515feceecbb5382d91b8c86dc3cb5a2a99a46970b9d987b169a7c5dcdd083a096de312958228401c9d17fb34958cd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h838b00403dc21f639e8e2347e14b211033aa31c7743e272a04752702b9a6f6d88950b2b03ad0bd303354b3093a6f87443d6aa2b6e5f87cfeb8ab3647f2b51ee74a8a784d02deb0a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59b4fd2ffbcadc591b800c97f21ec58383596f361e599c446fc1257721cabc48653a88218ef55bd1a4f3a5efecd914c70d489b9b49d2101df2c2d27de36f470d3b5b7658ebb4f8e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedd859c5f0fcf15226af2cd23818c398ca68612d53254fdb73a70a4d6b05266c1165e6272f111d4a699d67a6d6f71cfcf970e488945c03885f68501ef8b9ec4c238fd9027b44f040;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h297b752b494a0170c57819f02878bb14e58024d4c94f6ebec88f12d820d70af7284120f64862859bd99f0f3d72add47bf6c530edf3ef46290904af69eec60357b83eae2de676fcce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1c8d4d576ca137db646070cd5272a90fdb777e8ab54debee4ff9bbab7d64cbc54187458aaf892cb5d15763ac0379de6beee260e3f93cecd6cc46de3e5f52a951372881a5cdbb582;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3fb077e76bc42b1af67b4f74ab02454d1b38a90b9d85aaed766f66d9b2d31165bd3dcf040da75cedae28af1797b6cd4f017054c5356002328aa59866a5a4fcc960a0c9f57ef900f3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h745995118bd4b30f276d0361d0597e4ca1b1c7742639bd4fef030b0b9844e40ec8a4f46ccf5a99922a56f4089bdd6e80e4faf1124a942f4fe042173ac28cb009cde43c87a42aacc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9bdec95352b95b35a13a3ffa27fff66a73a5db52b2d2ae6828a298202835fc069aeb58c0b7de6fa959a0ac28d50c792b5a7a53dcbef527f426f02e0048f172204dc496e358400a42;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1066f715c743778e306b49c26b9eb9abd7e3d53262287ce09e8c64c877c85ea6ea2ec3f2685c7d4ddc821f15ef4f9daf3dbbbf57e1ba7d9a1548f901360895e01182be2f3973b87;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22d04495f8d7e62b43d4c277ad7dcff38d2e2293260191d1c9fdea1cbb35ea4a8690a38313d5c1ad19f9d49e7eef81e8be4e1d8d42b1b3c833476a1409128508537ecab7984afff8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52a3db467efe4006a108b7608abacde889e8d21aeedb6b194d03ec8dbbc172121cee63efc0a2c6bbc80946790a07940b85fc94b8d68350c230aa7bf0efdc5ecbdbc17330432bcf58;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d78894d702dfee7a85bfd7954757279b4463de596f8e6a510e078eeecd7ef0a8ef858e6b23811059819cb3e2eb39882166fc0d68347a8810e5668d272712ef27287ece667a72119;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a0a061b5016f97feaefc66169c105225c3b14f940807ab4023a44da4fd88b0a3fc452a2666c972d0d5925cf4eea989cf971c1ff1f7c70e0d817200af25d300a140729d89c16cdaa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h643482af6516afeb83091caa6c3557f73c0da96fddbcb70d77fa2286ff0f653d811ee153d97836301952616c873e66a2b84c41d2c81bc0350c328b77c3e64299454e5b69795ad770;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65a68fe697f8eda825ffb8b72dfda505bbfc7b70f079fe4ad057e2f46fac05676e768ba951b4260625caf5a40d8303d4df0fa930851f24217034e652e5c64aa172ff8fcff90109d4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8048b2c8eb96e97f86d44e67e643ec869041848c746111d60af44146ecfd1e376292213383835ca70eaef2ce04af46736e2db343d6741d08123542aa34e0e2c7ecf2afc236b19393;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha173cbbbf8b539f8a2c45592f2fbf1a528098bfc6f8c4c673e55be550ac4f77f152fc5dad81e2b2ec3a26979e1d9fff3e2a33134a4385d5398aa38a711a37dcd9f79ff81217b9711;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3c6ed1455a1534c8c46f35ed24c181375234221663249e9602f7dffe01fe7995e7cdb7feb481eb28298ea28d10f59366dddb70e93d3fdce50b67721f9d5316df7a19c2cf5fa25d1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69bc16e13f568f5c8c9c921dfae0f0fbbced971b7f1e4b40fd452d47e715887e00e11ad58977736b499d48b1f6f631d7cb2adfcc31fb0ea71175093796939fced7dbae1a8d3c52b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h246c8e9bbce38419ee00d879be9587eea18a0d54fe295b80a96ec5421a7ca538575b703cf0e053db488baf432feb8368349f1fd8355d3917b51509d84f9e0392c4194f56c6a79590;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c940d15115947ea12e2bdf163bf8a8e78e34339da31592bb32a331fdc0292e6ae3ff35e988397f1a1229c3c04412af9b29188f6618aceb2d27b215e91db99cdecc57b14c0d50473;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5e8d9566581b2aa117cac3fe931d3d184c76187fafd6e126e89c483bd1688985f476dbc7f1a49584e5fa2d77b7f55c4fbefe9a5f77a1b436cdc3e6898a033960ec9762a2c409a29;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hadd9f89c2dc2cfd6d965343095322d4cbf31e3922dc7c437c43519fa6d45fd0fac3172bbb8f496811cd5ffb5bcc2d2591de06341393675b3b5af87a22347c389bdf2471d95c70013;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd779c2eb737a2e2f58397108689c017f423a8f2f0c005272e09e744e7bd8502af6a81c40af0091391b427b1cdcf6ed692a4f08d3cd197435b612056ad0a42432c4bc783c8ed1466;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf299d828c71e3b1e651a934ca10a65bb8384e3b11c1eb3f41101acf428210bd4e36beca44fe466fae632a6de906c5a355d89e620288df3fd3722198c5e29bc2282c958a253863a4b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1d71c596141ae12ec85da9eb0aa59801d88886c56cfb38406ca9866fcb4956689d87454c704c9e3cf6783a9de6f3d22fde29c6522f29fd2deea8ffa0269f915b789768e3a6bb87f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7375eac4950f579332a2bad76ee263c9779515810c877f8638fe910fe25f6f9aa9f674105acebacd9fc265206c9804b7c0686ff1c2055f8f96a80e0545f4ee0c2db6d022d799dc5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a156e6c0a0369baef2ecb5686c97c8f70b01e1d31a1ca815d129868211bfe3afbe64ab44ff17d8149107d78ef4e39472526e078a4046cad632661434319de6a1a404bea846d5c19;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75c35d583ba185b91abc9ad07ae5e35309f06e328e5abcead835c2b8a5522c5a5ae3f7060d902682dd6158d89b9a0e9952ab869fed2520391aaa5288891c597409a8a8c86daa99f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h146b8fcd7baa74e0b2ed883a4e80e0d56293b396b6a8c9fb42a7815aaf990c9db0ad2e88a1f4a300c5d41ca33359214c93c6e90704b921b64764170cb38a627fe0dc57c6c70d2661;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ef17a160b3591bc1e39ef88496af9fbbc223ba6950955a7539e72fd2bdcfe94e8226c4d0f5dc534624b181ff73ebfcf39e818cd57d21986ac58afb30fb9187df388b2c8abcfaf5d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62ae7a6d14c350417460d59d7a7462a47e403409459de32cb9d4ed5342f9ba6a11504c4ce5ec366cfc1d4a7b8c28471e9ea7b00aaabe0e3ed788a73dd54dfb9da72d5dd20bc3f68a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heae8612db5af556d99726fafc5f9eaf3d2b4dcd1b4699a55f6ca42b6caba20c2509010070cf36b181e7008bb460b9491265201ecb623c485b96250a895cf2caad1caf290966b9a38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc74f05970607e696b8ee25dd1b3b5b50309354347458a9238434abe4e47e9341c13cdd72482cd2e2e91314e95164bc28e6ba466d483efa3eaacc0fc03f78f5b75743635d05e1701d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8afb7762ee592a22b928b5e835372c7aee98963c1e1b17ce50cd3e28874e57467e3f07b70c5c2faf53b3ea071a44e7a99e4853bfc9986f664aaadba34937b460f9c79e3aef215152;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h361c41e4610e3c244282f6712431f00e1673be46ca20159f86c3a10a14ad38ab61004c30135b402409206c3c54ddc43d7a2692a3f6e7f50d4cd960b72d9ea53ca29bb4b2ee82ec45;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3e2280b6e246018c84c5a890483c5acb5b227d653d04b32a814243e7c0d3aa85cde74d360de0e73d259eb97c0d01121235be22a7f39c5950804ab44da8ce8d2130868d3362e6c15;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc91d91e480fcf67336644ce09d965a63b15829512cdea0906d2ee1adf7a3f64eb9c720de9d253cd9416216c138d4801554b8f6343dafbeff0bce43cb0045b37d7a966e8bae0feafc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82d053b6bc3375e026d6f5020cd1005b7e07c5b4ba3b3ee2d403d5fc3f805dd8ebd0849c25d223f530cdbe4eefea890afd74c13b1d415c4685d6da781efbe70e9f50c8dae9a39648;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7496fdcca4e186f0bb697ee2150f17e14df49cfe8c0f688d07d20d389b4a8485ea361841e6b658c8c9cd5e9741a7c04272b81567b6385dae64090519c521dff62cc7bae332c215aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45a133b165914516845ead399980222bbb3dde97679d5c3435058c7d9d4899f6a152f795e51d80f929bc575a1b56e3429993de0b0bd7902b328247b341a3414bb33bd6b0ca118d53;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9f9044df6b85ddece6b4c45216bd162942c2a841d6e0d5838524168cef036479947e7e1006ac42faa2752adb6d7e44269510e093bbf700d4c66ed5b45b8cb8e66b5243573b62480;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a0d91345d372ffaca7c72f098fcc17ce6b84cd427e865787a111a00f411e08e9fa4fc38c9f3b4fc5f0037c3121cd5e844c7743486447d9147599fce4eadc808114de4fa30a3a812;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbda4af18f86a2af9f5e014e5321d2f81ea7dc69a4705ff283196b718babdf76fbc4767c6614b391146de4e64a7f48808ee9359afd9123742641ea6651aa3099804d290cdd87f5a02;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5058f0fe499d2b863935e6063ddb8bad61d2d1c598e89df1441fd85036678e7c6db30fa5df95f5ed2da52eefade4f8fa3ba054f46e7ebdc70717519d6d4d1d6cef5627fa0ffb367;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10098fee0cc33bc38b7a865c40cc5a9881134540dbc53633dc9d1b8560bbc4d9d13f9a1406ffcce2b2f897ce259614e2f791db3ba73bd1953364f745520ab1aaabafaf6bc584c84c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2044500073501ae76209e575d98206608a3416442e49a1e3f2f7813ff37f189de7813ee5b308a9c054ed59634839fafa6ba6a15e5d775f5e1a26723f89ddea039f0e8b4db3b431f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha923dbcefbfeec96c5dfa784c35f37ddbd04be4bac6237639d8d57d31b475ad99c5db0a70bb20ac74c68881de01fe47948f7913784d5e491666cce07e0275b632c42c2c31f14aca2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc89e3b2b6f5054ee24300647ca87d7899b34e30fa4b1dc25e505a25d638dddf52a8c903a3e35d55d07f815c2d430c73777624180d6e6ac36413a77a6b666f506c40d32e0391b4d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7d5e9bfbe060a90c1f51c0a991fe013f9120830139224ac18b08597ca4cc1aaebf0a531fe7669792b4c233dd5bbdbef48145c2340a27eac64141068a9100ebf4bab1cf13d91c089;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93b60f9d3f78981c2b8f7eb4264255db336e917bae5ed1e1be688f1e58a8a73ad9dfc8792528577ac8862be32d39a519cf19f1a7645debe185a76156a7ee591337f4367f2bb55dd3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18dd67db11d99a44a7b20fbd9805c0d41462e8a649c4b73af23fa7f13aefaff16f4d70c136418b5f7180ef45504ca5423571a1049bb819a39e56c6ca2efd545ffb7011f8a497deef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h28b3b0a2a1879867edfc50e7296cb3422099b69a99dcc056be5bd702c3b4a130d616319ff7019f8e5b4cb22e60b680b5144a421234f3be64e9ff3f6984f8357796ba5a11df967a34;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81259197b535375ff72353353c4b6488fd5ea77f2696df5fa84076d02726efc0d05bb305e4e395bbcb1773fc31ab05483a537b8de247858ed6d7fc3b072ca54345dffa6c71d0a5ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a6424051647f04ca973477b85a83f61e0b96da36151a8059596e92cccf091da5bdba9fafcf7b8e7915e0c2785c7bbb0c2aee4eff57c2a79a84c3e3561b1ca687b5d92cc8c0c42ef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2f82156b6dca152f7bd4b4952c052a8b29e4c431d2e3869fc266e9da0e19b5b1b8bf86b28980320e6270179a370fe66261bfd60d577530274fb8b29bd2f896a5a4da14e45e1c390;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda3ad210716d85041fb1089c26771f4b392626de777b7d87128d94fadbb0e77c3d09b3dc6281e2e03c2d152c8f6214e6ed960dc408856f37deea3aabbc0f6c2900f0b3d2dc613097;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7bc14bd190617efea212f521cdcd6e61fafc69c57869d07ee914801ba52b147b0c66f9ee78007a1c2830374a1f77c44151543204a513693128bbc7e426c3ce1ad7d8dd1380407004;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85d188b6c57e92559c86c9663d9d452f6287bc9cbc3bdd19af24e28c61daa0443ed94e1887cb7b622a69a270cfc6b9691911c3bf721fc790a5d34c529d6f1d0e9769dd1bb61e4a65;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb773743764375e90ae008a92702ff3beead1174e0cac13aee37a162ccd0c0aa1fac45fb68de07c5aa09815d898baf5c7fc34a90ba0ccc4d7c265def5bb3495f6801aaba95743e1a8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc46716df35ab915565e08f7937ae8ea8d889704028a0a372b1d0c4b76615dfcb8ff522c5743f2a7696b217323e1b9f0f9810d6bf8b6e3f0d76d4123763b639da1a02878f0781be0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0369fb372cffbcf3d37095f4ae8a0bec8906b3d5d398483ec27efbbd4c7f55e8f52d86e301a0423f887c8ababe4f53b2b07f5a9f8c3733e40c6e524ae7354b39de9cb755c5b296e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64e9a5354ba5c0b8c2f8049e2cab53e9fc8490e71df0441577197f5e5345cdf8543aa04d5c8c1a2b69d3c49f3709a93a2efcccb2440f234d0c391be924a6c6e7ba42e1faed733581;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2db1c7957cab208be4c58643a689797d6689fbabca18706b81e3c9f6799a42a63a03afadd933b1bd4bd71be7f302319a603fd537dd16f72e0df5499c055a74e4092b5a1058b7a61;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95e48ddb9ec2d15c1e2d36927a300435571a51d525e8d6b93468b74d871cbe3001f2492abf58c5c026160701960a58acaaae1aea838b206cf8dcd4230cc225abbbdba4fe965648f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a731c3807abe28a6d10794272b6b19b94984882288f0d9f360981273e1630eadfd689fd72905d2ebadf793aa36395ee503d80313b8bd96bf85d5d3e3e0b48ed15a9c4e57e93f127;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haae8ff1c9298f95283104df1892d6fde4ebaee1d8024ec264ef4ff3062a1ea8e01b357dc43fd8ae22f7831912a53f5a5d1286c275779e6f35442e34aeaff51396d480bfbf26c9921;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc73ffc25bac96b723b139eaa41ee0eb52621ad8ce7ae4faeacb7ecc1e606b69c5f163cb2d1f4da6e22b109a77404de44dace94c6501d13ad553bbd77a9fc5ad4b68c54a4ef00ac4f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb38d1702757159f34b090237608b7e818519c407a4a8daf7552d3d1a2498b13372a198f2670cb650f673c85aaf77a3a500e1ac36695f6c764136f0b7582ed755570d5fd65461047;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50f3cfdc20f53e064b267f08355b81440a9f42e23a510f42f85ca76871c70703525bf900edb8898de92b1d134161c77561aa606ae19ba05b6adfe9bf1f8b5a4eaebffa23e3564e12;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5371832c6e80ab9e124519d22b87a04131b1951451b1032f6d6a16fcf48f9e436b73ce35fb4a6cb221f91f905afe29c1f22d1f3b409a3375e5aae6db703ca20602e53cf4e6c16f65;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h420cf9e7dc6b4786ad919161e1b0ba8cce92802312a4b8bb99d8849777b18f33d545cea693607eb105029ba52285400e0892e65b80c025fcbfc8bfeae425f5fcc341dc939b4cbaf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c504ae5aa8d8976c1e41e9eb6654fcb99cf4461be8d25060780d56daba3e338ce9d46dbd275b9fa39b48546899bf9f8fb594ccb06fb7aa0c87da8239a5d676cd25f7066b644f726;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h888139b6ae69ba3c3a43f68591ec0295ba3a0124de61c0404b812df339764051faac04fcdb078b31b93d2133576f639315b4462038d978a55b5f7f771bf0422b154679ba765c3f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11b7759165440a8886d66f627c47aa86cd1fb9178ac7b38d19f4e1a68f5130bb950bc82301436f9c72a1d3668561c4c585fb218c33a0af35afe9a7f456c40bbe3a3d648563db6c5f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8925f6b446717a0d7a127aa2ecc3ea1dae604544b7c5bb7036f4999a8b7957c25556c3c63d29808b9bbb3c69175e67e665ed7bc61904d19895c3da6c7736dbf54c12dfca3ad338dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85b4619bfdc09fa880639d9b959152322236c6812193ea6459f71d1e18c62f7ed7c0d2c8fb10bcfcbd0640c33c4b7638e065d0e13a395473b8f4d456a6a1da0f1664e7cd8ef59d1d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9ec700edea23516367708d35d56acc5ac76d6276c5f9f1ee0f17f090317f9d7b2ae1dcea83cce1bc6019681442866ca6f6405a38f7e07deca6a931bb03d6b02fe57dc04215f5190;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a3ebfc205ad929375c9c33356c143d35f7aafc97a8fdf8777d13b0e52226562c2b12f4194b8005d274f3e45899343e9bc58b5f5ad9ace1421858c8094f2bf469f58b693bd8ace69;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h890ef740fa20f290476539ecba54b97fee01d770e716b8fa44825e5962938de9a6d4e859c6b828c38fa46d2c57f90c6a36ba2742f9de56f0da14441fc35c8a85b785f0c3a9fc66e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83296da39848b48b09a99b3a5ba5bf155501f2a8d7db22b8e13597e32573f18bf92852a7340aec8cf4e4458147a6713bc32dac55e0c63b7f480334c3175448c9c244dfd349dbd66d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8c36787cef3b64e1479cb761184b7daea4d7912c732de0d3adb4a328fb577daeb0e5baa88a78dc7d66bf6dc2492285897ccd4f39335f952817c46e260b91ccf2fa951764349361a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3da258cb5fd3479939922b324cb0cc1d31659b487108368e2c00f96ba1e69dcaf034cb01a25a164235f95aab685482781b42ba7fa8c06a8774ab02a62010df5233750335e69f9a54;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf98d5e21ddc23b28e9efbec42201260d2ede1a759f13734ec686852b0bd28b932470afdcaecb2140dca4c966f8d9ff40f06914de4dd398025c370cc3a03c1a95dc46b783460a5997;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd576a47c4f24184a934b53e5452f8e9a8b9057eb259210ca4e8eca90e3952362c2d1351c6e60378330d3aac601ee8de45ef75502846e3616002cd705b5c820f905c66f39615a2027;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha83b9c3a0116f075d82ce59985eec07395f812f73245399907b3c715b6a669a9ba42054565e1aabe364fa3a2e450636288fa2a97df2e2dd5ea510cd635b7ee05ad8e0a05a4a5f877;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59ccfe947fe87d77e7748db864a343d4ca05d437955a9e8577fc07d8c2d9f67d9c35ff7f090d8a844069c9210ef07f2bfa6a39cedc406a216860fc9bd8ef4b7d22b5255e8fbadbdd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2be29d86a885bb7954ad327df0a3e9de645e39d7ecf4be748136b824a4e74c630c2dae9486693831a46e10abd5db2b14256fc79fc4f91f03676f53b1b875f79ac07a2da44edd748;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b8336f3608ee09b6caccd5d0670cba9490ba9df5d79da8180d32050ed6d65e5d20221ac3060888813bd913fabfff1a64d11ae329ca05d0ae7ac69ab438a937077d54564dc06c51b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h650d6bd89d7add0e46597a8e56dfacce0070dd06f656a817b0c6dc4fbbd7ad18f1e7e662b0f45a353acff83f3af7439917a639209e9f024b58a2ab3b54cf17b1334a6ef3e65881b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6f9b9ea9f1741225a157dd74f23c46d1094c96f4653cac9ba46f17bcde50e447f30ad8a7b8a9814eafdb530a5ea2791e8e2f60a67f232b57b7161b33f034af7073e60308e379ed9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h483a0f414505e4a02a3b9901afcc95ce6be4e541d2e36fafadd35a589002b16eecf74c1b0fee50f2be158c5785d9918d6590429769985c9e8800302ec17793751057e814240e8169;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f49e0abb7c0eb454eeefb3b4853c9cf3ff68d615ff848710c224d07e23e4a1474c777a6ba358bfa86b3cc30994c1e5c323cf7be5e6b7cacfd517e645f00ede57bc383d57fce0d0f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd875767163931469bdf3a18dcdaa610c330015dbe5f8c0be5faa599e35d4e126870ac49a4f4576d166fb3eab3174298920a77c29f8f86305059133921f2e8f4c51e11838b8b01a1e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a7f1f51a32a571bbd51797ff8aa9f85dd2f513a91c14e2f7364e54881bce364c9d97be3980e040eea3b177a9aa8be89179c51351ae94f85abe1ec7faefeaa2fdf21193c155e52f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h969d7b13daa937c580618f19027b6839c1b9231e4275c34b41e19575ac4d5e6089e1225b55c53b03626e884ff3d82709625b308c35ea928aceb42853c06b7b8e5be735d350d45bf7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c7f54c0d5644d4fb7cd9c919d235bc5610592873e6eaf7e4d020ce46c8147cbc661d3ecd8cd77161e2f2df2beeb2fc445ea0014981f053c0b608e970478ee341f35eb893efcb88d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b184d05de8b0bfd734bc63f97c7aa20dea0198b5942dbad90affc1a94a3ac13aed8624611428a9e4737ac8e864aaba8c1196560efe4ce20ec5733c5e3eff580f7ce279f4c54ca57;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99905db6cd1b95342f374c569a90f773bdb954594c70bd220509f2c95e4d4d1412a55b2b520aa825741a08f9a698aaef4a2885ca9788a036c191f925050f31774610b0c424e0fac3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb918e863847359a73a9143fb3a68411aba2906ee08ef7d98785879961a300a499645f0dc0406694287c31486325e8b5a873f837e1a3cf260f461198f819c0b2b73ef77a0a7c8378f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9adbf1f146787353131db2f6a420b92f70b37cf5d20c2383055a11ac168cbdd8166bc7564221160e59bbade6ea11dff44696e39979d4b685c994b266ab47879e35fda1d68013911e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he70ea94b9379a7a27d9af1a296f05a96391de977a5d96c6bc8e2dcca238c43ffb6a08e1083815acb0644a3242e87cec8e1b82f0342f7c986a63b5efdd19cc75b0f98a51b51b3eece;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9273fa2b63d95e759f54a35b408a02a2818566b946fc5503e3ca840b6b6d76157a3fd35b68399102b33916e453ede55c4713fc3e074777e7451df408ba9060c38706da1513b9f9bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4defd603285de815e5e8ff8586616b2acce8c85f04035dad05d648ab30e839d8e50ad411bab4ea450fce431bb656777bc1a299db274f2b1fb37ef0819b6f988a0b8cd61561940ff2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h84c67e84bfed0b64388802d118f96d525ad38f470165d2ddb79ae37708a043a04685007fe558bf3bf785a9a0c01e221d37c1cc6b098ecaeb595a7b51ac953e6a5ab6be951ee653a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac8a181e6818d911b020947194645f40d67af40669bf1a06df434e39c3a5bf7ee1435907f631de8ed3fd9db9a2ffe3591269e70844fd57aa2fc6e0c81b5f82497ae5bb563be21bd8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47eb626b16820dca63457222f3f29f4e4e8d37d3cf277bae19bc55c2f22826ca3d57b0d067cf2ccb4112bde6bfde140b7a72b043d8003d1fb6637425bd9ed371845729af32a81941;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d3a77b45115a3cb3daae8dbb2f511130102b34a9d50c6e9f9c8d96ee54e7281d36f4441f681ed5eb3aedf10c7146ca68b75d669f1974775bb5cdd4e42745f3b6708b1c4ebe32db6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1aaa981be2406a1a34025b3310192982dd210687da788189834326c8534fb03320cc75137d58e4950210865b31d99ae14e45e53f6f3ee5c6b4b85effd0967bb1fb060daad706ae2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h707bc8414e4fa7e2e440c53b20dcca2297b90d2af8f2cd53f31892fe99e750cd5d29853e86abca1e3b4049264a22035376ef738690092158da52bac2dd57ae83b8b63d4b62cdff64;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h700cb999a8205bc503aefe83515b132bc6f700a2e565aeb28f906bf67b5ceb7e300bf0ff23840e607d7a810a6573afe15da220ea016b296ec304035d1b83a7aad9633908137f645b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac9a80557fc2b1f54765a4b6bd0dc2ce8998231effe8558dce89c7fd3a2ee4caa7a799af317556b46ac039ea7d5a1e4df02a7a5d28844a1dc59cd9933e0dad274d8274edc7946fef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9fc1d51eb0d5c7fe0adbd7cb6d41c55ccbbf62a6fd85efcf4967df99784f0f3f49cbd27ce446b2385e117686764a811ab0de83be7bb4faa024faa7c44135438d190f5a9889f83432;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf3609ffbbfd26a1841155da261bdfdf6bfff2309f4fe161476ddfc24725eed67192a301800e02377f37c2c0146f3be24754c0ec9881007ff51dd05211de8f6d0b027934d9cb1af8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h492c470b61a0fe7bc45990b58b554ca655632d814e6f642394c39167b04bc1e194c494fce8c7ddc17f26c9030907cb0a735f97fb327f772ed30398e6dfb33f3275706767425db72d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h749eabfa4bec41947da2bc43e65ff3bedf9d821e6a7e6e1e6abb61f621a699394787d17631eebe2a27d506faa4152a76352193a9591b36f260f3e40518ad696f62bd863fcc19cfbb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2669de9806b6be35cd998fae8e45dfe41d7ccb02363b75737de8581581c2650c94023886ec2b286aafeb6f0d56da69ff8b1893f021500ca570d57dcffc9ac0221b74b6cd62d390d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94c2ba96fd24a737389c7b962a3a1aa7bfac38e01923f7315ebbc33e39393933d5a8eaacb02191bb8be92650ae63131e759323339c67638ef8da820bc90d4ebb727fd105bbfbb18e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf72f288327ff94bc5deb816f270bf32fbc9d8e7ada6c46d3ff420f7c49cf012be93da197b4988cdad4d8818e2b7e5fecdab319ae17fd8d768e35176761005ba5ef59558ca39f78a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd37666ae140017f9821161f9a2b2694a87bb40eccb9f5f807ade5da8196016a531a66e638d0556a6a542fe7e6818775c0e88b099f0d12257448f81f018fd31f3cfccb821007bf40;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6edb4809ab4b9f65782a0f20356fd861cf878ba6c045590e98aab56e2b37c19a14a8cb8fc85cb83cb619581865ca2fa646e204bf074a08628e7a996625c4828aa5ad729af576efc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42b0aa2827a16c9d99fae45324ddae72118f11a5690e49c22eabfcb7fbf001ee79412a621a1fc667fcd30330f48ba47702acd7e299fb2045b8de50f8780ebe1792c204e3c7f57940;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd52439c61916ddb30e64b2ac4c2984869629a149b2f699de0b990f14e4ee4fb383baedf6e9256ded40c34cc617df7e65f3689969f8538a07e30762a414ae4463117f39a75e8d8d38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50874121c45fe39414eb5402ba5290e530bb119eb8083ec3db4363bb1223afad82c4e0a0e263ae511b5bc164db7f660d9f534b5cd9bd8c4bf30a0547daee7eca18fbaa7429f9dfaa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81337c266f3fc516e4046fdc8c8a75591bfb7eb32679d6def436affaa5bce0f2d69f632eb3f84699617033e73294597e1440721c6b9061190b4ba6c70cb9589fe3afa7c036c82610;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hacd0423b70d926f5022af6cad1f6fd96f36e769dc8fc3b07cc688786db9b5eee800ae0ab06a691387b2f6b99639de5835e10a3f2ac4407cf8d1574ed4c648c828c590ecc7398e83f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2996679ccd0b60a748437de1155f2d819ff3bdb35c8d7d300c4d95e9d195874617b11c6e15688211e23b0837b58ad505bd7a1565f68d617672475532dc713d355b15257f93e55df;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8150c4b37cf2c728759d545b89a15e58f6ab7b16df32c3f354cbbe49025ed3c261621ea663b2c8934aa1d690264721cc0be121d4ce60161ecb82ad3c8f9c5d75ec6fa789cf1d6e98;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3dc6e7d5f9005c28dd43f7fb6bc115f6cf8f408fd8829d8fd8c62d11dca1d645f95f86a916d161df8cbaa15565dc2be22fd802b3f16aed477d08419b31afa15974573c007622395;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc80c960fe09ec259bf29293321294a24caf70921110de0e433660d6afabed4dcd75c65c2b9dbb761107a81b72aae71fe8cdf3cc53ce846c8079c13af2ab2a6a40da14b22c77611e0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha55ef963b4ca7c537782ad128e3ed4d8ef7f041becc6385f8a7ea54b43d7e43fa6ec74e05d5fc358be180c6a20401b93414e436da44b7ecae69725a96ff024eb51120c45a5722db4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85b9e9188b90a0a3e0552481b21361bcc67036dbeeee8335bf62360dfa7fe8d7aa996e5314247a2b1c85406b2bdcdaa4926199b824eb65c00757c3b1a0c11d01fb4b3fe3fcae9570;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdddfa0a0e95d640131bd2e92267d6339f99786c6524879415e7e2122ccd6f24786dbd838736bfa0b5c0a9b93a7548276df4661dcd494efee074ef310a6ed6d1110ca1ee9d916196d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7762c4744db511061a768006e5e806943c51874c20ac0825da9ee6ab5f36c6bc2e037c5a188e7fa6baa06a1f6d3b412bd35e45c5670b6e7c7b903648253537a1273cdb5ba3eed4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14a4585b9dd1a7d2fb1665662bfd0caacd71d5fa88f4d6d9b14d846be3fc83d282ad254455282b99051eea1a4a807e599b4518de2501b307eb69d583d90dd5d3dd9875c273d8f836;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce822d8a49d5eacf4abfd291a06b14a63b4e776368b65a0a91eacdd2a4e181bca1299d9db99e5cdb4e191f4afbe1746d733f6f27d042ff7dde387e2bb42c7109b1752b5631bbba4b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h112c5ad11fc7bdee55baf6349c86e5583c664b66a8f2bf7a0bd03b9e7a55fe09bbe99280a71a2c7ab777ddc39b6d6db3cc0fa1794c60380b25afc880a5ed5a4de996f41403c7b4e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25a5131713a26e8b5a7bea1f1acb112519212bbbbae57a555086f905e1f78ed6033384a1f15d9c61ef47de889eec0cb26fc8b19d5680be290733204856ec4fee55f4282299eefa7e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h383d0c481443d1fd2ad7e227f9801eb24d845f0fec06f6b759c96819fb02f312d7d57391bec99028be1a578a187678f59f4834e2a949cb6b2ca9894cbcc4cb951e697ca9679ebac4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8dc3bb89e04cb1eb955050cc7d1bf6b57895d33c76429a25f6c3cac3b60a1e47cfd0bf9bbc8021df11a6573edc55a1f4164b58576ca0887a161d6bbe0bbeccea8a10d74ccd39a09;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b48df8c6faea1b12acaf703cdd7c7d84477265bd3dcc0ee441cd65d1713584c9d5d8bd57b83fa176a0e20b2c75db9ac5db408506d87fe7c472925f278850ab723c636816de1ab88;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1808615bb562d8fb3a62b0b9c4cd06060016a0f3219851c88d236624547efb358eae8102ad8e0350eed8673f94a8f37916c04fc132fa7b2bebccc02ba54cf05bddddde6613bfd5d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48da58ffc6ddc0d86c16d076127356602bcfd670ccc2b66cb9b246941fe1ffa15cedbd1b8c8f2f365b7b1bd7c5604d77d1004a66a3c58de5e0b438e6f0241ab0df81324de8ba1db;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc924b28c716f0384241b21ccc7bf6018a149438486f1be5e12369a20b1461114087ebd5ec5ccb3f959ce53699df93b0c38a761b55d987b511ee28860873bf501639b60f1a7c565c3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha70d0bf0428a1413f6e861e5ec92ff1c202ffbedaf560726a7596af242c9f874a0b24f90aeeec93c20dea2357cef7eef32b54416757d6a244435ebb48967a3323c4c14a55bb76fad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f9f0c945627903472a6f10acd2d3f21ebb102037cfd767c42ece3a61a53a8a54a723eccac5b92edbfaefed5dd5a66470fdf0f54cc4d482a831990be0889a4eaa7e71ee3fd22044d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f63bd9abbee68ab65914f59c0e21deaf813a79d1e73aaff6ae54b07c775bec82d55d4c830ab8591d789bd3e9c44f6ebc65dcafc838b139a08de73d3c367b96522ed1c521d1ecbf5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd926825707a91d04f7bd0c82dee3e64ef9cc5009252981205ba1e1b362ca6a9b4add415b0464716712b132dd92539c8faa41a330cb74f2ee4452b3a5df7f6d86f237d3667542c5f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf26ad7b73d07ef6582c998a5708018c08ff4aba2f93d053bdfe02aa1bb0e1c3c2f0d5c7c70ae43becf1b541b3f09645263a7d37b6bd58491735afd3fd05b9706a35d0373670811a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecf6e004c2c518d440f4516c23b65d0e9264b229ea2e9b627bf9d3934abd68b13225b67ee80cc578f413f28599a7251b9dece86f5f7772784ea4d70de6fad7030825344c8746aa9d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb19840afdbf3402f6bac5b287a28483288f8f032c9a3e9f79c47f15630fcfa35d83820f96c1de925d1ee39bf63755c9ee615925f14bb85c97fdec9ade28baa7daf763a5665e75a38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76a5f98e12689850f539e16c58ac82fd01a34dbe8418a641845666bcf4e488664d5a7bbfecf45f27a43d2940ae32d6c43f5d6c8e2be10d2ecba7d606923492adf3696977dad59995;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3891e120e5a812f620623c4debcb16bdf7749b446b23477314bd3f9c261254ef6c695bc761c372fac5646226facf3de51502e44f1f492f0dff3b323d14e3770057103ca2f8c925f8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21c4d8927795a18698a4f7b6c6d21d7fcb1c894b2034e6137d9d3935b4e3dd1a37143262e387cb406257a2099a4f025af4d4f2bb6477e53ca21a5a510a4681d2a03fbe8c27839ebe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h134f9712cc5075f7ebc21ddcdea396c99fb7278ca47eff132e204db19f8d23ac8730fb74d2b048aa0b1efe67b541f1296dc61fe1bc9b327934e7fa5d358f61ca934352cf0ae6e954;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3998a548c26daf8a1d53efccb779b4fea0fb6f0c6773c5939026488f634d054a1a2ceb2c9dc9088ca339002388196f9ea71fd710e7d8ec474031f1cfe5a3065b76332ad80d579621;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb36b189011b2513ab60b960995ea8cd08c9a7508b9b356de039b68574cee75b5cdc843199ef584016a479b016239b66f07d727fc222c707f320f62ab1341572eb0af7aed325bf643;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haeabcde611d113367e85ec1b28376777f4e994262b6ea390534b2046491a181cc90efc73fe8bf2c8967184964cc693ea9c880c665dfbc8ab17cb703ac2e0e12a6862caf1c5978688;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a08b4942e3cfdb23bbafa687b47fec62ea5657fa35a56f833821883da00769a7b550f02ed8663c0a63a828672d9c8ceeb9100666dbe90e3f6a2d0f09e44e925d743e202e58384ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61dbe365b0852f9fd63b1e5b1d6b2c69ed19f8e1cf9ec6a1f8063e810020ae9489a2c938658348dfcb82d79e9feb8bdc3644248a51c9fb64bb3c7afb9d16dc8f76bbe0c96682f52b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcef3b6b1276308027e9020af166e4ad443d7a8ce3813265f7459bc673ded69708144917648a4a02c75c928575c84e66c51c7e2383c862274b30bed082bda692d7476994cb5ca74d5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf67bcd4fcdb3c1404bb63797271a2b8aaee0450c4a668568b61eb495205dcfd60b6c70e93f883425d4f8f2010f0e146ddd1a0a077fabcb1c135f8cf785923d4280ed87c4dabbd0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16c8ad5df0efcfa91b4c17a663f8ca2eeaa8b168444e7759d3823e9f55e7d965a897465264114162abc30703f76f516dc282381b9babbc3e66a75fbdb6ec079d7933fd6fef65d75b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h346a9375f316da9d866193bd0463677efaa576611f4f6f3badc57a7d25f26744b8851da2dcdc1f1c1601848579019a248e02a642e21cea30cad296f8c23905798229678001dc9495;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h534efb297921701d5d900fe50729e6bde4ad6c3f1f6b69ab21d564e0d85ddcd10947d34803c18a99f833b4abb910018fc28b2b5e5e3dc56f49bf0431db221e6b762e7fd2cd872ca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0f76ab0b3a5adb1b46c41a457e1a1186879e2965bc29af13d4cd3048db1bee613b277401d75150e78f22edf3ee83481ec236f4023694f169480ee90e5bdc5fee4bdb81f812c6d56;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c5048adfb03d2c800d36bb44e4794184e7216764700b6c464ca7edf70b646a5845b7e761a4bc21b73a9ec5b1ac9b7120fa508a5eeb1b5229376ae891811b626a05b8450b2983b32;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1321c61e3fc1da9b627da47b6a1f0bb0b1c3e4573133ed048a44b7e722c9572d012c10afddfe3780a2d56cdac83ab717846ef74b1d7abde182948e363a8baf321d49477722fcdbf8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h900fe93f3db961c0d5ffcabd5af45516f8bff3db4b8cef7ae3fb0589003b6b861a9bc2770d409b23a79f46c737e6a6ffbdff3e935ad84986a862fcb7c6c46241b2b07ae6d1661ef0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcaf849e2fdaf2763817e0edf5ae3379258fea4c9095259f347fcd58a8821ebb93470f8ec59ae29e39c5df4d857c99fff6c5e8298c77fad53be5bdc805c75970d6ce546b21050697e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha414c670d90c03e06f9439978792b77b168bc746671bc786d9e07c29265e8810b4dd3026d5c0b2fc0581a20cb4fb5f945e2f4e7e2e92443cd4b2f401c7c3ad3af7faa4aaeebdc327;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbe738696a55b8b03c7a1111890eeae240a9c09b9371c65c1e928b32b6289c15a20c5ff461c5f42591ee48f389021ed4d708183e7744d8e9ecf57aff6200b25426d840194b5bb94;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h169c1351edccbadcce3ab32e29e140eaa4afba902b9713a484814f9875927264dce016a065c8aaa210065b4f29aa001e79c16cbde3a23c1b9a6db842d97456907b3ba2049efb6d00;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcbe39899024bd463894f83cc009f49454eb9c29f58b9324147991c2a956e71adf88be0112b1bce6d44f4f4779a6c1b7ecd6a6a10d14ebcdcc61d9388c4a52abe3bb4d201bd65cd8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3979f3311d0bd78dbde1b95f91263998cf4a4b7af377b7e5ef18763a992cc972a103b70656f77010038a15946e04b6669f54a7079f3c3c4307c7b0513fc41516aaf1b6c0e1130ad6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd385f6f97aedafef34be3d6047f50e076806b6cfc6b67b443fa7b4c7b82cb858f36b101ee0e69ed9e05b0a61e5d0f5b46ebf03a1dd98c8fc766fcdc0124e1f732901a8c16ee8de88;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d23c7df96e3b7253fa110a8bf4e40efe503fdb84e50498e2d617c36528789248daf0af51fecde15326b5a8675a8ea3aa57a1b15a49dbb2724e052f5cad70bc1cbb9971ef051298a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef0cf8dc946b76e98b5960ce8f5db30b7b22a490796985c2e5dcd2b1745493047afd152f98eeb0c25cde49b9cbc64fc2ece46ce2f72d24ae61ac98d6f1db5a44fbf043651f7e9b18;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb640496f72a77c24b46a5c449c8737cf570f42fa28f956cbe4bb99e85508219b7c28ee023e285302524e394bd179eee9557570a3d48ea797825f5594e33c8d858b839a0a2c3b09e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba476a2ed9394680bd32d310e75e7c5be59db1f10243b095d5a68ecc5f8daf2f7f837abcc9be90af41955d26ce403b8a305e2728b9e256f35920d1ff9a77132ed2a1e015e628fe4f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27caa41734a0ad38050b9df160e0d39ce9f8fef5b3773505208cc7cf7d760e6c71eb72c1f603de525b5ca1e0eb1b39d133858bb8b731564e75f301a3693c019c7c92044bb9de943a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd711e42fd330469bfde7f23cbc935f243df4bec1b43ebc4161a7bffa926cd04ae85d2fe3a0e4718ac1097aba500d07068220ea20f4b3a4d91756b04e7a87ce6dbeb8994d21f1165b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc074edb7dd4817485bd537f782f8da82847afc75b899093749dafc144e24a527fa5285e4e09dc55b39f0a07ab59a90e60b42f418fd28086b432ac396fe6bf1b53aebb55c2db28e9f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b65a0d06ce541008db8022f021b1de80ec220d66f6411360530ad1087d28a7644f23c94966fd82e520d62f3ff42e151c47f5d7f1ff42530f1643b977edb0e58950c36481d79c59d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a909e685caae2c6e2c4c93a68c75db13f9519a4028e5d7ca7c6afa195ab511613f9aebef5062d588dbc2005d5a671f1a3f81cca82b9ef183b4e3e006598562227ba689eb22dd1e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he11ba85fb532f452b16f18d1538ffdc46144e11a97bdc1477809bbdd572d1137286712bf8972ea0271c3a1e5cb83abc7980475c6110517182e66cac03fd83d1e3ee12704d6500a70;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4111f99e3160ba2fa8b08ed81be1feea0d5d8f317948a9f4e17392d5fdeb71a7777a648aaf2bba53df43620778967aea375aadc00b3d42218c1b9a7c2b77224c754db09cb0ccae9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h235c890c029b97ab63880f5916b02694521e1e84160fe34a23444a8f8e7199e820727366539665ea472257d700897f0ce3544a1b8e8c710c552994184dc8b76a7f20040f2d2ddaee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51dde88c03baaec6e5d3f6497e382a2bdc3f5ede42056a967592e24935d4c0da61e1c4100f264a4f46d907e629796b099e7b7abe290fcde7e0aa9493a819f7ac9dec98d5e1212f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8653866f9923180a375953dd86ffa5cb0f5c29b4fd63d247929bdaef1b7b505ca8e6352d5c37b5267b1e697bc667093f2ec090817d0dd84fcac31d4148412f560a467655339b09d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30d394c17fdf064dab30f2c1d29c0cc62d8f848b075716105a89601d561bb8f02dc96db6db4f1ca6d42d23ba70f6d29ceca0ce256437a82a347790c6d5d2f76d5f4a54809d135c4f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h747202e8a9c46188446cbc031ff41b9e58ddc0c344ebdc1ba1d137aea8671f5e8588729e5ca382f5ca9fb86440fb75d3a596e2c375ddd71606007ce65f9066054b331916ca8de9ba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf3753e463e34741e24fcca9deab59f157c3095c1527e5455df8f93f4c39cc4f92b72b648b1113ef4004ef219494c27bb0a3444056268670b5324552a68ec752f8b525206987fbdd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc6e66d895149e276f64b24b5ee185dccbea3bee69918f67c5681b435e66a907c2b1df794f9be5a8fb9e6eb35e35746cd23462ffd4ae426195dfdc10d349e299e2729a240cf71cea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heaec0e343a3369aad6c138665ab664946cec0181c96d8d0e9ccc3f53e63fe13ae25f7b62508a8aba878b829d3da4e5dbf90fa8dacc03599bd4af71ebb9fcf3cc5845c227635d4f49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77b9a22fab5812075d36bf0d31272ea855e4ce49f9f793cd1199e78852978899c462b3408840cfbcc9c63affab53b80bf23c699a55eefc8d7bf0de03c962d443dbecf42fae7a8db5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3e73cde6249f410cc1c9392cf978be75148c22677fe986465e83098f422e9e7f1803e94f25a58390a58ef9d4bc102e1872156369a2c84931d74f2d96aa9c8e80639f58492abf01d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h450a488efe99f2d08f264b1828dfb0682d9218b50ca981d6e937e0bcd835f04cf15cbedc0b127c9d61e6935243b0fef726f0d7cc46c48a37e106c47b69c75615d6f926fabbc1f86b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76f4a1f50c566fda5adbfad7c8f281ea65512828e258bcc2b633989121e9d6998290ae99faffb9b3a6a0f9e944898bd5b4323e2e94953b91c5530f02ea4f932f141ad33f7f175947;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h515465dfbe41096aa549e96c5cc804c0343c82018d16e29c42e8fd7d0e4971e29178c49162b0db179fbc447581a1090014b3d9b7acd368bcca170a1cfd418d3c8decceaa2ac24e8d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd92fdf6c13f6f6a6405e6fd512ec767ee76c9bbdb9ec96c37c2d868036af0abdcace8dcff466702f17ad8428e642bf0aa1451cf33f3b20facec6ae3d312254e1eca8c75baa86002d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7ce69bdee98ac6b2bca0f2de4f08846068d79c2945bcedfc2786736918769ef9f1d0dc8039b1ba135e49697016b38952296e677509b471317d3dfca23e28e90464a1b5408c57fd2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5098eba0a8f25aab1ebf4d581072efd41e3d22961bc3f2b28496965b85463bd30b0891265415a6d3b0c75c317f751a5d2d76641d307f428a78a0820a047559bb720a3a6596c8531a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34e187dcc900606bdd1e229479b0f9b5ed526e1f576ca1efc5a241c7e0ff53b37d1992a835363b64c16b58fb43c500b7c275b702ac23f8563f5f2c1e0e997fb2ee63455b21188b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8912baaaac8ae14729361f17fbbb24d8c9824afc8ffb590143c38ad9406aafb9403f8a71b6cd67a57560399af9eb08441dc090324f66d90e18413f23b9ebf4a95c6e191ea5d8ba1a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfaac255260c95175a7b506f347fc551551160b362416d59136d3c6b5646e823aca013e0c6b83a6b4c27c00123e43c7aeaab9d88c8c76b82e3a8da2ea5d8010e09baffd1228768654;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c3bf7047f120c31aaf2e5f5b0bea68271bd7ab3db6fdbfe3f1bc397ab6f79a67360eb8aac30a0891e14ee2c5a58b0780050638c6b3ce1c1970fa1a222e8c270e02dde4d034817ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef5a6383ba343aaa2d848ba02b7d52ba29b01fb4cb44cc1d7432a05efe337ad0bce22bfc3643b6d31effcc7340a829e1b86cf7f2c98ec820c327f4d77e45743893734c8369d7167a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c33ed1e3d1a0d522a829947dacb70216b53c13b63ef7b335d000f3f045eae50b72afd619f7e06e1e099a4fa106ada759df30bd39bed7288b2e07c551a5d7ef22758afce113e19a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19bf174795dba6a733b307b8f6ad4d29d6231225da20fce7028826ba7db1aad4bbf78953d9921a72501998fa918877c45fb5f097a0cf94abe6cacf46b304df36a9db98a147c56c98;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb56c46b546010e19c374b1fe9757a8d7617f2a312aa16a44aa3bf03003ab3e5be87c0430ebf6af704414df7b92158a27a275df48bad4eb0825e0a287686cdd502215bfe88167761e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6daaae7a29e82977ef4fc84ecf0d9928950ad57d5ff95436afa306455d6a6ede1cc6e34071ec5c571c5194193610788fed71c96abf403e84b9f6d895f11f4f0126efe616129fa263;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc8d304dc2fda22a4fc547e2e958052219f2f73c55d3da7d36abb75e065d26fef10cf1ea75a5343d987ac715ea7c18a956782f832d1a153cac223d387e219a4b68e479c2b9166b21;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea75c91fe60f069b5e1277c79443e3b6c5415492e7fd368149d36edecfb15fca2f77caf14455b0756457e182b7df217c447d9c131072219684b03a5183796967edc0133075246485;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0b52693c342a45f0ea63a04d3f84f567eb86002e9c46b0035f51380c4bab517589fa0e40b61765aa2ade8058f6fa5e6f360a9c3aa6fd5229d607f2df5a3be8071462cd51ac9a56c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf90382f662a2f8f9190d985194695f25ce7e368f7a2ce851bd30f646498a234b86334932f695583721d436c013f8fcc1e446f9cf07299be2eb8afb899eb722ae2ef527e67a5c6c6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7db0bf4c444eaeb03da43f30ce0e878b603d1bd3ca84cb3629490e411431e35abc4200e92ee44c4c56c15b454a2cd53ab6aabd0e0d469fdb286c0bad9f57c3ef573019cb8086bef1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc484a28eeb615cb2174974532f567a7491ec5bd016e69321283d0dd3a66d6df9df47cf08c90e7aa8ea1102b054822d7e030fe1340ac1e278315d9e8c8049fcfe4a9bd800b3c5d0f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30e992aeb9a2a3098c472d2ddf72a780e651d21b10b1d77fbe34142d0f58012fc406dfc3bffb36cc39f378961eb865c7bf982ad5a32367cd01a0d74c7986a632b4d4f134376a3477;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f323dc0225b630d71e32dc0c4254b27f10276c31214a9b7698c8b473026e32f2a3334ab220e6595fe6126d19785d3fb79133984494188c693da186db38d7905343646a691883732;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53b5eb6a851edaee98f08249c2c9d76e67647b7f3ba058188858eab7b2fabcbf7a7053b8d63a8b1cf576723480e3a35359807aa60635656dabee44a1e2cbfd03215c47eff0bbfbdd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce5a562729f320deb9f714bd678bbf6b86f786e84b156ab1eb7ba4e4832f5a1084b1ef0ec3b3c81c5c86036c00ee6464a98ea0bff9c899f991604e23f4cc0d2491e78c820d5ddde5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ef1c9bd9a1b31125f29a1b9b804ca362df6df0b374d826eaf6071ebac2b89c3e40e10af05a995a7fe65fffee7a96b81afc8e74b629661ceb815cf74d9bae9fc9641651c78d64418;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e7410bc9c1e066d4e757b116abd4ee264a3780e99c3869bb0e61df9e898aae9a6f4c18847e841eaed4ab7638b2fa9dea26c5d7843c0a936aef567c2c2c5fe50e2ef3927149586ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h970e17b5b74b67a22cb4bdb2f664dd0a6309f5f6c8cbbe09e3b5f5d0509cfa50002c7b417f7feadb4dcaec92b56d283d6d80826ed67ae2cdc8dc1350668073542d05e0d948e585d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9eeb4dbdf56dfa52f0ce28d7adaa88b59404fb38767d9995584a92eeb8150c5ded306be2acf63bc35f92265d48b016893da7f70d9a69ffb2af20d84cc45cb2929d680bf8a2a91dcb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb0f539d035dff22a4ab609063d7bacd9dcf7b0cc4852c345f7394af5b1e6d5c582bbf56c83047e15e93d1f639778f19c87863152ddc766ca94824f8ab0164885eaa9b4d44f180dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8fed8615ba2a97ab22896b07f45ea18bae6d6b5d6fb010cc588876b06337611f74b512edb101d2748f700bc8cb094647f02ca9cc06bb5010f7b5b1a69ff2876dbf8195eb63bf28ea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb41ea4516530502670cf06fd6a6b0368184c7549ee54a3066fefd25b930ea374bd0656c2a2f1a55e872e0ae21438d08ad23b34295c3c2326c640f9498f74a7051afcd0d242044e9e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f15a8295f4a9ae12bf5862c2912d0a0cd05aecb2cf8855cc13a55f0d186a39050d4cefe74ea14e50422e607ca06d413c2d49e159eaf3c247191428d4e7d2cfc2bde3916b18c4e0d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74e71632294a35b6d165e9672f8065fd3ffab7ff2d12dcd778b80f9de720bf0e2ed8f1fb106d1bdd145ef738f50fa1850f2929edaff65d7e00d90f7b0bbfe798b29e3d624cdd332f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ce178b0386d604374efd2f5a093e7e6f1ab507bf0167d20a1b5ae3642c68bab08e825b87b862aa9ffc291eece6d4337b16566099997055e8b3d2b08583d843509d006cd66a96294;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h516d02456d9f9165505925d41cd4ef7461658a3658429b4c37045c32fc4782519ba07c7af6b94fd595ead9dcd32972a2fee54f868992e9f941997146afd4883398d1c0ff6237560d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h511caaab26308fb80e33c4ffd2ba7e1cd37bb928dc73615bc289e18e25f7beedffce2f86fafeb3d5e188f824c30df71b71e3045eedb17bd6dd182b43d567d30fb81ffad4e03c2a8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e04438572b79888a0e1d3358ce386d4a9ad1112ffd96d4c45d3d9c9c3937944c9d68b8fd49246474aac24da5887baa972e2e12323ed0409432094587145947ebe14e64b3f6bf178;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h152e1cafcf8ea8e0dbab7e5a70063cae5971d37a0e070d382e8931cec77f7c715f9947d65048477bb0830a1ed17843db4aa795beed78e83f1d91aba56fb1ae613efb7bc457d1a33;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcedbd6125a3eea0ecd73089225c19cfe3298c3737dd40d98fd1d53ab31392fccf142d05fc707790fed322ca35f33d62af458a596a6878a0d190f612b5f24c2e8fa6f019a9db8e3b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h149d01495c0e4278a0e2b362aba5672c68a641cde4e440eb5e82f618bdf6ffb1a5bb9adf040f1b54b840df54026f73c514f27f926051a3d4d56e30fd3e6f69d68ff06730a4e9d5f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51cddea6d0903074c2fa640b1b414fd05fc55ff224b816ff3197663e391837728fe64dd1ad5030c90f6d4a7d3a9dd1e0a2abea04af7fa4889a8c4a66e3da5a86130161841366f3eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ca5a7e4945215fe48807ea6f28a320082e866064b439de53d00fedfd7baba98e3331da85d988f9319af9bbaeabcc95bc7e89d122711b075f4016e6d80c1e2f36ce7e3a2f9357048;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1649a4869d8e28969d195017ec603adb8a0fcfe1d409b654c86d4d450a378074ccbd81be50b42f4f0e5df798a19eca47ceb0f0c253038166dfb7d6527212d41a89a7e3458d21993;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54cae63905b2b907f72c2474f5705907480af4b01e0168b4d999b72659ad49d4f5a97c45cbf619959ab8fd79ed3d0262840fa5bdedda668b78eeb4f138d3b0907b3063a2d7df612d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2166278e7e707a5c8575397c08711f95f5e4cac6c162dcbcdc524308f76146e2585af29cdc2c49794346aeb2912f70a5385e52d76fffd0dca931b5fc165dfa71358bde41d52c572;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcebb782263a1976c4cb3f4a390804af1255a4c86244a588f4fa439470321e0ab672abfbaefd370d161d9501c0c22ac42f2e87d1084a914509effca52b3ab44442ca4effa28dc53b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29e06bc7b18501a230171483007f356c04a96c96b3bc20a673299213592336912954a1254f0f5c85c74549efc805385ffb712bea1202546b3f6076862823ec3c48150d0801b1b140;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h226b2329a43adb1323f25e0a7b05a03cae92ff5f3e0678410c2b58b3481a096a728b07332dada14a7d2800ba3b7553f44acc0d9d20a52eddf241d1f86557ddc3980548d210139d1a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27ccd98ae565e8aae584ea98e3d2c6e99168a285871fe4f12daf8a33275d3d20d96aa020e981a50004ffd5c239de16f2f44b6b1c7e712e244a024ab01b585a46d36c4c1614659b0c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4dc7654c6363e0cbe396012787df5c9dd605b5ea734164f73c71f59b1e4ed1ba93684c13093ecf9dd57b52e1eb46046d008ec542326e040fb588847317c43894cc5c79dfbfb21872;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1894e384cf116cb4df62284c99dbbf5b1460ee03a19e69ab4c552f620355cfe129fee494e8b020d387172a56002d6310d0dd6aec31cef87f6a148a8b54baa4e5dea901248131baa4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he87adb7e5b82b869010385c69d9a459779fac4e889207334c3e1850e74f8a397d7d53a790601597a604a967bc0b70aa733a6908f625edb66fca0dabb2da44223b7e8500a4812ea00;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6d34fd432bdef40bc1c7c350e22109d01db58633e9717d2d5c25dd99bc4e2b8b929fe86c8b14a5df55868c1c6b07247890aafca31700a66c9815af1d9bcdb273faa5382911b333b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d2641324a979de908274039a2f3282bc60105bd731d60a275be700bf69b01358da7b441ff381d5fe396bd80d59a0be5f66b883f2fc91b2f48e4ea2b665d10981be1c76c8a7f6807;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ba8ca5f4eddbba56d577dfb940a4969ad6c8678b94bc0b2046b7994a657c3a0997a870dc8365c9ff45c1ec5a67e00cb212d4c5a4a81be7e99f12d34823ccaa6f65e9d3201bc21a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he209dceaf67e405a60f433f8fdeb56df89dc416c64965ea93d35da6c1220de0d4f3f4858d722cc8f731dac653026690f22e76eab42e49a144ccb247be6b5596667c664651aefd57d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5642eea10a49d2e4d3ab395f14f141c56b76f43bb95336a6ad5ee8672633d286d9800eedcb8b82a824dcf2f717a3ddd85f15077de18189329623de862b919f1b4478b76b6238982;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd4be3cd4e510fe369d1b2a844d376eebecc2cbc04636cbbac6e7bea5e053f3573f946721d79767c0709ec7644e52eb90200229d03ef62b4c1f50355378c50affb40a3d651f93a02;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd59c828eb7c35b4e3153bcc63bea702845c7ecd07cb51fa0ab445309776a0f57112442d63e524fd0bb961f69471d3b373b5d1cb869a48e16da3f9741d4bc93c1badea1a17bcc970e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f917832955d7341437df3f7fd96993583a680777400ca3c835b363ee43df92bb32a1c6474c055121f8ba90dbdd1fd9da8cf9d6d3bd54da8e009b58a1fbfbc919ed3af2cf6e3dcf3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h587e3124f95c1421a640462d9d4d72b47964277547f393d48e3fb486662a7e6deb59682a0a36af856d077e08465a2287a40b0bc55766f34994cab5daab652b70c6b89b4f71939321;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h513d346bbc4f0bc9cd3292c0d7941febac7c64ef0a191a0acb70ccfb1848552b205119e5c5a95f37adabdd6713a10d5bb508ef5295977d06415411bda42a215d3f725a2c16aafd0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ec5db41a25cfed5969a7fc087118c690e8d10787aeb018cc050a94c738a31cfb90d3dcc0d5045de809413995805872f5d42d9f1eca17c375a9220f326a60b213ccd9b99d165a947;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd11e0f74c29dab9e6aff89a71d4168062932f78def1a12b469476b2515a3864dca22527a6bd284aa2c320dd88d0f09014dd84400e45d3946e8d7042f36d807df02631b89f812040;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf87736e9c06e0e74db8016f1826422d4cf3d0c473d0678e950f1b3a179724fe76e136e02312e284e61ef674453da50de9000ad0880c10177c2d1e80ae69cccbc107960a58c7fa602;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha476c671294de55e8724b4cfd4b4890da3e421df5442bf20ae6a244ea365deb316a526602a123a5fb19d5058a6731e5d948ae73b27f4f3f5590aa7829d73555b060d231310c42bb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7427cf58ba76133016975210097e22635ec48b7161a79e06c491599b479277933efc0b9f77d3a9f5fa220018be1e2bf2fcf48261bc675db1b0277b1422cc853faca72bfab01a0ad1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2eff05362eedc8e2e3c83f9f8fb42836fd8ee894e3a8f55704de6fb14301c3df8dededc09fdc43b8460cd8a559ddb76e67ef23c77c664df44797e3bbfefd83924b85984c8b569fd4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7017ffd50be63dcb40159d28cb77e4d725ea03e77782a60c15b97f419d4b07898a7f53b12891a850bd0355de8556408d730781c06a1c545e1ee7fae492b26bce14b921620bae4c95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13db3e4659d70afb333f26a71a9a08094e7c1cfb9489de1389b9bcf4cc88ff2ecc2541c1dd3b3a26e0a05ef63b90b5eb57043ba64bb7a31f03e8d9158b3d2828523c01a9e40d79aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee4341bb11bc5995d95c8d8122f45c6041d6ee8dd93d03132bb00ee585b7ff44109d7682b1a02f042f459d6c3d0358a7491ebe93e209d36511fa12bc9351806cc68dcbd0739ef90;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb55076baecc3e70518aaeb4eefb57a8dc5b642337037ce85ceb623fe28a302b4358c4d73717a796fd09b903e7baf252f5f47bac85b6ceb19590752737a5ec90fb644822133271e9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1bf6b1cbd42d3e5b9faebf0641dcdbd45b76fe65c58900b551cf8facad2ec74450fe875105bd821c5ffd305af7d84a3318a3801ec7f5f55e6a79e2c0dc389dac26e69329ec1d029;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hebd1c14b4046bc9838443965e7cded310ef5903653a7ee5d10f18d2c953d3b67adb17c84d9dbe283e1d28ae21381311e1b2bca17900fcdf47cd8024c6f5d6cc1d74d51bb8d96db02;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8b60ee933625b528565c3f15d4180e7ee5cf4c04d0af2f7bc4a8ca844f1d6306c58df719952014a475307664d61f5eb2ca22417030e4c1509350662ec3d64a59c75e939db30c534;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd45c4e92edb0d3e9bbc346d06a16aad7a40b95a42d8adfdb5a19fb6682ecd0d0dc748909fa8b2149cba198667e26583c71d5ea59a8a931f553bf8afbc1a83f7c6c4f4cc7acdd68a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcea8d227236c3d72a3fad89f92815d7266b84081d5065f064390c3fd1a9a4a80e7cf354068f6cb10fc70560ae4807cc2e0541c2969b76249405f77f494503a73e49e7bc8b330cc87;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd41efdbd19b5c8e4133d02dd12dd25b664f520c85e8eabb820fe50435acb1a3212c47977fdffa35a15a87b34d6476b35b021e99b391cdb4b6b3bd8819e98c61532c8d5df79171a23;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h492cc0475a94adb0b40544124738cab4837796fc2bac6dc6943097eba4e07cf88f52bb8cba7037b64ea115584499c058096d40b65902919c6da7653e21565375f491bc03c3af17fc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72af0b023dfa63a0e50ee400e072c2cdd65d76abc60eadec790934f5cc34ddbe1f497563dcb8e5a6c50c8bcae8600cb272174ff312edb488f4a3eb781c7d71ab27ab611df5f0ff1e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4306bd9dbed1d62c3e18fc7f8fc535f1ced5d9b0411b8839d043c751de3fb6cb40dc265d1372b173912dad03520f0360c3f8d4e5e1fdcf6c1a84b6bae1eef2d18bb618b24bfa327b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2e517ba19496149205449cd16a732fd966b99160b9c174db571406b3cddc91deb13be90440e0efcdad2ba6b9b8f57e52535d160465d218a9e6d7d6fb38d104dde4a616841085913;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8fc12c781d320fabd1e791717fa3bab424da0e23ed8d7f2d7999776bfe4c80f5a180cceb50983e4722b8b70ac652db239774266a24185faaab364fbcd4eecda0ef629769f6e2d06;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h28ca71ca0accafe60a20531e4186ffcd3cd51e1c819986eca887bab95b92a2954d8ac6df2f12316f3bc2dae9804de4fde7e64b0cef4872a8baba6baf95399068cccc8ce6499968b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he34c95d009367f394543376593ff1a8702e5ae78b90a309dfffe3e7b406d1e2c6454c0e651757dfbb4ce7ff6af06b96a8295d7570fbc5b5899efc477727d6937605a1163e3d587fa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he067aa4ecc9ba6a16688a6ebe2ce7425a81b5871ed52a11452143467129f030a54e59ddeaa6819cc5447053c992dbf16aac559a52d2fa18c858c2c03933f9ad88f749a6d1b893b70;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8112e7f564bf98d77e0910bbf9e7bbf29f3463797274093fa192dca207535838ea50facbb350bb6f51a2b26c57d390ff275e19ec1df5fec27c3bdd27293dda253d45156ede91c73;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfe59ce59813705c55ffc7302b750f34e8a78ab1e5490227e354ce6eb3408231a51dec1ba3dba2e7cf0f0addda6548a247d9482da1ac28914264a309dd6996980612484dbd179ed3f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e2971b3d65f6a3f715e63543ccb19884b9adcfb7156d019fcc25a67d361367228ab4a99a940856a22383c4bbf75ff36fcee1b1a96ca3d49d9772ffdd19d03ddba867e944ad8b698;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h288d19cedc39d4c12c1a1f158665d6eec6659564844362f0f78e8ba5b7357e9394bd3f971505d56d709ecfd4f625ab672b7e995f1821126f2a1ab708ab8e00c2035a321c560b9f65;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85352bf85fa0c5e7b0ead50ccbf1431f50994c26a5af1cd17be630f9f3b3f1e17b6383249c3936edcf19e71d8d1f44cc0879037d2528a204397812d75053456d981c4157c179cfc2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54bdf4cee9ff505078db08d91d4c4781df6d970a7d94313294a3561438f21467b467e57c1cc083f1030822350e626516e2499b2f9385f4886fa108a6cfd09d7403ddddfac5acc97d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde51eb176399c03032712e621fca93983fa5f2949e8f602d1f145d1ff004339e77658eb1f024c0a04a82554b2f13ed43cbe2413fd4a64b97a9ebc8147d75962d5b1dc2a649d1a8bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd36a86c92de547c42b905b280b41a3c69089fc3b2e76216dec727b2ee91dcae08e09f1bafded0319e4db06dba653115189b59c9031139200cc63ffed8f44ed9f1300322056a5ddcd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf632df6236af1967642460ba0f6fd6076d8b33b86caff72b8154f91fcaf66d58edabf127d9fc7c66b333874732045a14f7606f828b4dfdacfc54a449396dd4e3f8d7d86c0778491b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3d4b70e869af633dfc75bfcfcf15e5adc18f77d0718ac7d703a3d8ccf996eeedcc3b17336d0418a8b27e9ea751350dac3e065c40bc87a9b31a1fce5d9da2d7538747d6d7114d6a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf75766b0e99e6e238d5e1be1adb180ff2ec2d52f0838f7a4bca0db28796916dcfe198beb7423b161f05871d1cebf0183278d0bd07b407ba1db48d7100f9650fb3c591b7e42127b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1915cdcc579e21a4757905538adf528d3661d0355dc1bc6cafa7b73828f8f5568e62bdb44ce7fe794d10e55aee915c9fb1747f20c6792c79346e8f273fb0c603939d0cbbbe46b894;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6cfc8f9cf1459c384260f1704ff68a5df0d6641ecf013072e3023d62496abcd8bfc21a97277af2e4401323cddaf812cda7a840455ebc6cde50fb023c3e8295b6203487f0c26c549e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d26c9a63a08939163e0de2f32f76e54ade303acda18ae9d1dd8f968b1d6bb3da4f1c037a32f6f31c291f4d6eb5842c1516d2af94f3bf4661676bfc5b0988a57e9c0f98f2e56353f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63a4b83f176e9f273c2687ff0470e72e8af8f59c76dc9fc86b317b9c4b9750e2cad7888e0bef9109b6e4359ee2348a68bd12318bcf76ec8e3256daebbbfc5cdb25f58398e00c8098;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5970328e78e2f015d08246efdec01a2b7570acb5f2f1dcdc44b193236bace6410d9cfecf212187a58bd626c14c257aa272535dfc1efe7b62e5c8807fe8fa790a479a3c66498cc80b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h180422d466f99f01cb04831eae44c89f98744cb1ece2de005066698ce6274c6d1487d5515df9cdf62140ffb01717e8deee267e0a2500220b7d50a3f15c59cd3d3be63ea820ffa19;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb97b7e21c428baf104d5664036accc76dbd6afd2e08a0a1c894602ef8e33be10c53ea719a63c62542272b04fe24b139116e10285f77584c89cf86b157f6f5a4ea974c53546ced10f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea08e97c88f909c578a14d8525cb8e7222386dc56252cbbc9c7f0b497c15cc25f335c3fd12c96cf5679f1f653dfdf6207ac1e7703e46ff5c2406d326b75a823af8628dcd9ef7b9aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12fcc7ea57f5653855f4015fbcb0e61ff261c201fe59e1f66df949c24e114a4e25fc2c4a2fdfc2098c19c359fa17591e11ffe46ac34d231b103c41d7319ef812b63433590771744c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b3e12a0f5b513042ce5d120a422b310f9a3a64191ce35d59e80c8f78d2e4d2a5a43d3ddaa38034619757a84fdb55541a52cbffbd27bafeaacb2b40a6f1ba0a80d547168167e9957;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd107167a3d975c4570ecbbe252304c3d70189b73a46c6118acd7600b986a8f7b51b2a084ad9b424a96f7b70e4b03daeba1465262b16f4f6372f2fdbcccdbb6b93fea113ca0c8e3f8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11cfc91700649e4e84874947d9f9e109ce3878287e0ff001f952482a44d223056fba4938aebe5d5f9e50629312139b8e24713b76a042d1aefed407f2de83c700f485da7054971316;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cee9e60b640fd99c5d037171bd038161b3662fb01174a9c62bfdf0ec967a0e3df23abdbbab101ea307b443921531390b8ebe34be972ce03538334b224680b151eb2796f069588a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hece7165e94cf31a1d47e2bc63df3853d528aee6b65f5d728e624660e192d6a5f267712f11e2704885eb3863bd840c101afcd37b0d27d4beeee880dd9b08c7b265a18ae1dd1d78ccb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he17146311d0312487485472359a6884683e12e7b0bd8a4cd9245af93959478293ab06e738508d6ef76662e9aeeead2542935345ff77e268f49f857a4e301e25264b5dbb90709bb8d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2cb76b0434d05dc286360f7dacd5074ea414fb0b97b1f5ff26a695c60b4f6c15c1eee005a6a9c3cb13ad681d2158d3c4c88ea659cec0f83ab434b3948c5aa58109ec44d98b4ded3a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5163cbda4a715fab2eac27120a26f429efb1fbb7dce1535fcc1922a3f037c25622f13298ef63d88936d651d149f536a4ff2f6fe9423ae9fbd2e583cb1b7c58acbef1b6402b4f41f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8921a23e841f646e6797442820977d5b509d769fa8eebcad3fb744a0a2f9042d538b856ed0423c67aa3f70fea74d51c4658309805a722c62aeaafb886a5e77d142a0b10515e0fcde;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc029a2a40b11378297be6448e36bdb4e1eb02992a3d55712339bf6092ffd1e8c4b6ab61036c67489dabc0c35026d0145c42c495c7ee98c167c3961b8a9b54efce79af756fda6d4d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97ab3937790616ecd860836d3e862ddd632e9049ee1a4024a66b046193731a891c263718814407e10ddc7d04bd116a4f4b11edddfc3c250dbc475cb4dd20c7c6caf4c51291d72de3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f47fcd346a634a88828d57fdca8028d3a6ee576817c6137a59e3ee0c95036beef82eff81a669b4c9a8cb671451118a87be4b0c65881ee865b77ea4d134d465b034d0b09db6cff43;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45617d80b90b0e810addda739212408af6a86ce82768911ab53aeecaf24a8d50dcaa04d496ff5138bf722caeb00a9f56adb6e373f008c8a072da898fb60c1c99c15c8c6478daee2a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0dba937e6ebc98cbb9b2e8fdaf254f3132a714fb47ff35fddd46e4c6d89fc0504e18cd110e7fac50b19602cf0515e097726509c30765af8de6c489eadfcaab237c8325a156e2e86;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h102d502d9f78b5661f615cfb3a3ea6af6d6737a90e27454ddc830bad754a1838dde586b3ebb81d0309100227ebf4302f3ef2e50249c53082c1bc7e9e9ed918d662164def1cea009;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5714b6816527d596b9c74e2e4a3ed383eb56465651cae53a3401aebc8cd7d54f2444afaf598db5791b62f55a69064f4f59773d2699c900ca2abd2364685844f87a0b98b405647977;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd34c98b28044bfca13639727e191baa5fe35a1779833180e225a8d67d1b2b6a0e83507f3b753bb401c647fb1018522ca181424dfa844a430e001deeb143093db6dcff0b5fe83b1d6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf638aa30e04b99dbb83b541824c74d5b718873fadf6edc74e0e9e3ec3b61b30be11cf923214ccb9647510bc5f8903af5137e4eed7de60e54b70e9ee1a8af5d6b4a0e3cdf6fb60bc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b4004c17f3ae8b9e9bff2ee3a518b9ea0c23fbb9eee004d03d16753ce43822e6b10c0c577384c8c39632b835bc967f1b991f889e83fa1f265b0a942e311223ee4357b921a66618c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he77bb6cecc152674ab38553a6e77f0415892f27c0ed8e27f52d9eb8c7fcc1df58180e92a508b40654fb766beb0df846c7f7a1e8b6810456341e79ff31d1e4a77831e39a7ae14d5a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h160305d5955d77e625d8ad42bd472e863ef337c3e4c15636fc019c6e54938089049b25ab45c72efc4ef79959392bfc783fe0036e984f28d209875c10906c3d9a38c6236ef1308d0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3f3047cf27d2b3fb4c01d6cd556bdb13ea6d254f5f8e7595a78b024dd4df8112ff6a0c9912c3ee3510c1949b7ec7a49f7f696421f4a98b6db172363cf18168f5013c135e3b9c350;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbabf7db2373e2265c000dce2335e2ddd6050776f9835c7a8987640ded2b2f77771b910874b67589030c09de72411ffa0f0a0eef236bfc81a40ccb1b7c8f3e92809582175fa8b16de;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70111c1773b9a7accad12b4c5610944180b726e5192f25ecd5dba7c8401f736aa1ad21b91a2d1163c2149cbf763792a376d2a17a2287bd76120f255bc1965a5281c627e506ae580d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd00659c9ef5a51776b01804808cd84940fac4be704bad548c10264c697f6529784ded35cf13510b555d3291580ac611d7d30da6150bf24ffd1ea98948b978e0a46ba2cb9d8bea26;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e12045779495fd67c5eb0b0a610ac29ca99ae212608ad4cc2d8785706c19d5370b17e882359314dec329c2e3fbe0477600bbc264ead2287c6260cd60b47ad65013bc0536cafe75e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6daa0c344f922d8175c07f7d22c35e25cb938330667ae3d4f837109160dd61142de708dba9b968d784aeb4fe624aa62cbcac13622e6f8f267fe877af59a6ca867559f0f753a40c73;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h864fd43b8ad4dc6d6756bec43677df70a0c80b7bf891d3c3bb9aa6dc5ec7ea68bb67011d884f6d7de651499c03e1562b3a71f7c8ab83cf1cf8d04ae618d5bf556e8f720bbfaff7f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf21383aab41916ac2b246ea262dc162ebc11e88ea0ba4bf1f882629c9dba6e05b8f257f33e857ee54c2a1a32a131dbd3694b7c85f6aedcf127b5247179e2246a32fcffe6bc066f3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ab036e961baa261670690c10dcd9940e51c5d278c6565a5f08576e388d5ce9c569f7957184a1b3b6bd65013316498733ffeb58ebe4dd989ffbce69db97ce8d8d2ff195dabc298cd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cf57b82f55b9418165904bc64ca5b430f6aa2c1546baf1968fe6d2c15fb4995e12b68e4846fe2ee332fcea1195c21a86ad1a34237428385ff08830c07e6967bd3b1ccad65d05634;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34b4fb74157a2c626e9b777e544288afc416c750ca8ca3a5c8b0a55b108f2a5845f913df7f6ae3585ec2c09c7c9cd5c88a300286d9cf1d0d1414dd04c8c5ce2a18b289294e44194b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h730a91309249144d3a41aa1ac3a14d0a10a73da78ff21764106e5d9d56c7db944fc474716ebafad14352bf5e00d7223ef8e4850f1401759d723ea4191f6ce52bb308f87f86c3b6c0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a0d20cbc83ac2147513acc34f5f15b868e323b6fe8e21c9b6191798103a21e2ee0a1bc9d8e886ebb1a06f1f26242e0d15af409e7380a45640c8ae1a75022aacce8f0c5f028d1446;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7c3203584fa6b95e182aa300b1c7ef28349df95db8941a612b5814c8935489fbcce8445228432d36443fc564ab6246ea81fa02dbb3151794e623691f36dec5f66a30d298e80db54;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e94c6e26e9d6ad1bc9ecbd3fa64e7e619e6b912746ec1c7886f6bc4b79a60471c68fb0573a1653a9f442b59a62e845a9e61c04a7f72ebd2908178ee80a04cd5ca1756aa5a11e36c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7353ed5d4c6173956ca0ba2624ed5c1ddba043ddbb20ca8d2ade5e5ffe4ffd2393a49e6b8aa2cf31f3ce389b714c8795b295ca257655d2badf26d264186e007e300f43ec712e91f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe85b01af3ed94f4c0750a8f7f0a62f32052ef8d66ef7528feeaa2dcbbdc927e5fbaa9e05c0a60e7bc0cf88da49b29caa71a5db3ee8d283860025bc6dd073f10dcaafee08f1b5240;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ece70e344a87e056cf2eb9a45a1edc4c4f3b6b98c9e74697954d869f4029db0f74b59c7beab22df8077a04f3596d46dc5a3aaa8cc0f084468b203ef6e31f2bd3dfc8ef129a3b974;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf69138d8e7fbae555c345906894dc20354b168819e6bbd74c6edf6bff2f439f906edc3c940145c622c319c1cbf2e81740712b40eb91bc76998dfd8ab534fd479c7e652e6f52e7028;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1241c9cfc0aa507aa461893220a69d101c325cc37c01e6ffaf81688c4f374b541597cf70e0840e4a070e4e2c3d981659a12f5ab10de9b36af4ff46c0c55a140bf5647e63f8ef2e7e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha472a1a3db08427d7f1b9343bb70b629d7933322022315c59531470da96f5ed25e41281b26d8c851bd565cf2a8a80818710cec240e3723b76d30e2df5bcd111ae98a25bf92494e1e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62e845d86c5dfcac4d57208e1202539fda2b83a2299839df22219a8431a5b222574807ee21f71fb7ea2d673f749ef7c7dd5befb54520edab3e35a9ac1a17a1495190b8326e01b29c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b2ec87f7f7538d71a3531e420a92c03769de8d21f3ae3f6ab304aa98012878c02e9107fede80d757a768a77b90f608faf0969e49eddfa9a93744e94e23e3f7b8635086e4d84b172;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7aafd090fa9e51457bfc9f7baf6b7dae57ae7e63c5e080df822829aef3b47de9cb513c817aa28b01d00c7126a4bfb4620b42a9a88c59798e45d51a693224dd99ba555948d63ae162;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h625db3d89089e5218ff47a34d8d7fe7dc22317b53d30bac5447121e8b6b068fbbd420023434f294287d80cd2b82b4adc31416746b3a0ad7dc891b9d78b8518bf288ef4801a709fc4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89cede089514ef25e82cb865ce36049075d02874a636520912f05fe5e08e5c3ea4cf4cb2e6d122c67fbb3a0f8ab9016f5cbbaf29a7557dcf4fb0c3054b61db394557834f77092b1d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48f3c7dcd919fc98726c9e9ef9838e580915a35b6057dca1a9838d4658a7dc432405f156f123934a48fd7e070f7eba53f3e5d05d6f4e940eba5a4fa4d9bfb3d2b1ee05055880c08b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c5c3e3c43492fa1aa7e9d9808f7b5af2a77d843522ebc7407f00e33791a605144313d70901effc88ab411df2542975754b33b851c0f88c7dec8fabbb8111ef1e10c0ace97e832d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8da600a243680db73f730672736611634b16c8eca06f0d508a134aafc25731e0c15cc8548ca0df168657f5f8bf66a3d2a1e4d5063d3d62b38eff289c006c4f42d55ae5e704dbdf27;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11b76cdf44b13e8d5ac5e5d3ba50ac5d14f77cfd0fec019999194378d328202fc3880ab3a8a468c657f89e7aa6eaaeb4d93f7e0075ed75e762df1c505709db50206afa833769bc87;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e350e76bb263bdb7d1e7746028f7482f47e26ce68726057066b8dd4ae4ff32549724edb145bf861890cae62fe65f28126eade24a5eb407c5435bc05398c507bbeafd7f88b1d4cc1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h430a3f3edadf7a037f3a79be89237ac363fa6711f3a07572bd5c6a47959528bc3f065fe8e1c0c1067e7397dc1ae12479650747e849709d6cea3bec84f3c5138f06cd5345c7b3a1a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb791fef4893a0c16383853dc594ec5bed3b9bb6c7da0372227a6c36b44beabe9993c0eb5dee39782d779996e9a804644843a1de88b33f761abeb39320ad1ccd08ac9fb005d8c443;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80ddc9fbc2cd38068c2815387d5be3e330ea99825b9f832a5ca61678ada222b5771f6bfe4a7e8663a7d10c151db206a39ce89db143b9bd07e5529381100c4f01c99d966c8f25692f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5281c75c1f23bd0bf795af37389ff08102feefbb516109d794dd365256a146ccfe62a9eef0a69053276359437b535808316af695cc6f9c916e1dbc664cbdfee2b9dce6ec06bca828;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h951bd44f666d61e7736a9ac12e4f832a72baa32bd779f52b4f0db446e0458b696812d65e02c10cf66b54d8335f7e2bc004aa73edf505acf0477578c63eb5dfdee1e62cd247f89f6c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9996193a076aabc1586d548d2ef4a3e11ef11e01e9f2c32debc6af39a23a9d49156eff1c0eaf8884044e335360c9915d01094bab65fcc0994ea44bfff3e04386aa2cb6d9b65fd0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ad96c11d418dd8a24ef7764b8274bd21bb80831bbe8719b617b3d443f57181d40b7ff319087c681e55ed7126a97cce1874888ddadbb17758da873545b50ace14e5aeedb83efbf00;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h360cee1ac511937094cf2ee7c73e3ab137c43a60d131f227d2bf33fd9d56802e9a56b0f162334d68a2e3b2a6ea423e8feb0919a36090ad80a4e74a6e9aa34feddf9cb71e038f5632;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67db8b868a613c57f7ff7bf52f5c4d1441cb68e905c818183321fe5d5f82e0d097fd51db7434f21bbfb3e6ae7ac3e99beb281837fbd9d8f6f0c64cfb2c2dd553d7028a72172bfdf4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h187b546b2ba2aa75c5dc902210c94653b0bb2d9fe3456a88980237c98738a151de7c35b1e34af19b0a7357d4d0ae358cab43ea1f94c40003623d4cc11b2a357681af1878dd92b05a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h825601ed8b3ad27a11e4ac4cf170ad5e637d925b060ffe6f27478478daf5acea6b17818c1af72518584f4ae93c79c51ad98ce6fba2eb695496804b935b97f140a57b96ed94c832c1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf99974ad71114f95977b450eb205972b84fe625bef17cb31c996d352aeb2ef5aa038ceb21c340f0d9c49b38f239fab831f565ce98873524f16950a8ff891e8d94fbaca214f735b72;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13fa848d2580ec64eb4ac20e076133c86a251522955c65c4e65f6ea67b65b7a16838bec530cedd1324ef64f31fce76f5a7ec035ddb194ef00cb0bd20b6851e8648c9d9ce0177d412;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc27349ed360177e378f9781df746920c214888e0f92645235416b1b83737ed1e27020096624f3e19c1f0bbfb01b62ba7d4421636ececf8f7b058ad5ba467a17a5f2f4e0eecba2920;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64b63803b5a43a128a16d5b075b5b8da9eb4f5e3f4c119cb5df7f83a0477313d4859cf82655b4a67b72b3a9b262289304f12b98c103524806896b24ae985181e5c2e74dc6393e8d4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ef53d7d830a12119cb07c9c899b750b69123dbf94eba5fff4e5ab283072996a19c58b175c6380ae467a3888048b9fb750d3716fa8c609279a68014935068a56e1b306eeaae9032f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5017c26458cf158cd1b5839eb09e4028fdb11def48d16126eb55324d3bd58f064f69dffa2f53ba7ff2b6fb31fbcb07d6a87b65a98d5ef09238b0ab532b6d33ba2e0c49325b9ba66;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b7115606a624001af2b56cfdc4e8bd5ef61e5c2622e6ac9334561c3599e609f59c4f8e8f3dc842b43ed00f24806c8719819f845310b160809a915e16acdbd371b714d638a4cd926;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h523d0450a46b5c592ac32c3649c034e891b7b23108e44d81474057c9fc5269c413a9ddddd210ee06be94314b730c5d1927e427ddbe1eb97a14704e7e7a31e84e7b9a2315b881e330;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf83e8d9ad85d8394e3431040c13fb4f4c91559257fba86f20832b80517f3ca8dfdd2bf13f5122ddc2c1079382069b1852d38b2fce7b510ffc6291edfef02cb5242da8c4d5ef1e5d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h919cb22c4773ea09c2fda46aaecdcc5bc5abc2d059452df7129ac2d6ba087c7cb408374dfde37ee22f6e507046d3661055f176775f063c4d3c541b3d4a439b8674975effdef6797b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae4737eb6efcf0c74d1ff79bc0df2c47f6e4448aa03e7fa816067ec57c784a93bb0c16f36d3eaef491320e820349d1b9e6229e7bf34d0854c482f7f686e87df6316b4d9cd86be558;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71eca8ba531b681c729dacdc24d9bc0a0ad9d89613109442011e0dc4d8a222c080a32bf75d49b0c1ce3a9ed79e612a6aacb1b2f4ad8c8975aa92e6ed843b3be5ffd05ef60091566e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c8bf3328bf484c856c06009334487fc4e4513fcc512777a3a077ef7f8fb2e6fc96a078b8379ad94b643540c60fafdeaa4a22ef3ac401660be96a6f936e8f2fd2a0b9cbbfc47cde8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26946cc446d55c5117d812a6157b7374b21d75e8ee7429e107186bdab2d535a45fe91eefa30dcd15a9ce63165c878aa6a73a5bf181a068a832d920d7aa9e4906ea75b085ca2e5e38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87ebf56845277873746c3ba5b47a82f667c671f0a431de355b461ad039fe0a74877ff5eaf4a5b88ddbc4888ef5310897e4de5933641c3d25d031f8c5b4e5b8eea4c07134e53030f8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffefeebc7e14a00d3430bca8812d13815478f6365acbf97326268982c752b409124b151386996ec4e0d515dda7596d263a0088b28a5653b159dbdc016a6eba389034b586c9ce230;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9bc34f641f8d47a5a48f7d73af35a55050d9a7b96bf92d650cf273fc93e8d48a6f4afdd78143ead1134ab57aea3bd96762de12e523434a9043105d95eb2dfa9d1aff1a6069f82a5e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52da2b1ea941ba85ae613053eaab1653d7c3b540a47c2f25cf5786f077d99d0314fb9b1789cc27109dd257cef46dbf3f347487944f9e8c842c1a619f886ec99def381d9c4d1694dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4dfd0bda3549d84676edd2b78b5306a5ce323593377c66c62d0b9f3dcdb08ca3142ca793093482bd42f9c9432f4147e3714dbf228623451816febada3bcc2f9dcc95542d92e25497;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c2e74bf46fdb2a043afe271762607bb582967ff10c6928cbc8f9c2944fd8c1fc69812580c828e083b2e379def9cf955a383edec13eb338d4879b1de249b4f9a72b3d9d6f8606c90;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74d1c6a64014893aac9ca4c7a09933a0343aeb83db0d3900d19009496a4e7c3d3e8d4327e6fa1cdacae7f551564ab3e5dca413049c7784bbed165054a0b4f5efb8d14d64017c79a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2256daa279f99e17d112751be30a44b081f467002506f522d0649ab3b80f546144082a76e28a4e15b21aa8959fb78b95a86bb4c023bad99f6d20b018e156d93eb8ff4f43ab99975b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1da40a9eb7d9861bb207d19f545595b40b8adfa008078d8a673ebaa915854e7e2b42f14200745b5d05c3f0cdf66077aa54ea2be86aeca18e1aa5230cdceb625f61de26ed65c8d7e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ca0f81c399a9fe5974170a93f3177726ebbd5761615568cbecee508fbaa082ddccae862bff698ee769b7db318fcf139e3c94eaee5c52ad5b6f6e706bde655bbbe6bbe527d949087;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b093119110774b5ec78f7123d09cdc9f2d5f89d08105bf84a927893285223ddb83b8f5e6057bac8aec89d0fa9708f1dd779067b2a1a3fb82635bebc238f105ce2dee0d8ca541a53;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66b73dea96c53f2f516262b732e5190ef860cb96acfdb3e875ceb165059ec5d55775ca05c9d1506f6c249bd66c0e6083eec40627a3729ad4816e8f7a29ee6680c901b8af59ff3797;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f385bdf0754e34bb5678cc0e72969fd62439771d471e82dd1bfaf35143a97da2d2831e615634cf8cbd56a43e62f9da19612e5f64ddbfc3e72045bb00ec2311b8fcd16217b6b5a81;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7a0949f6e3dfd954d170d490bcdbdc7f2aac9e95f1fc44154050e5e6b0fb446f725466dbf93f798a103911efae0c6a0c3e8e3455194c5482fb4e3af4cda5734a931e96e3de92a60;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e63bc0c2ab96241273dc47b8e22064476ad79aba97a7652877e76327ba43218b84c1e276b00445be3375585813359562686a96a4d783aa0213ea300798a5884aba1477d032668f9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35256ea1c75e47402ec094787b77352b0962d207014c5f8722a6e72e7571c6b7a00f23a43bc6d9ea51f5c1e64f93b666c99ca267e4c8144d915c448ff8c9868c221ed4374d1e4d49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd10c3a3ca9dbe040ba3dd6d6c662b37f423bb76405c5f31efdb347992949796c0883b1642cc197516fb7058472cb4facf907630a9c3bf8f06e8b794fc4b6785b9ab2f7b84f4f1f18;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h869805272d740ce30b8828f2aa8564bfaeeb496cc1bd1128a1cb1094112e170a822187692d01e26a540d170bb468c6dbea678d24c98e956dee955e979b9c17228dab889e493e8d06;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d7361d50e18936773676d8a0b80caf28a5acdbb5fb18672d07fd489d4083345b5cd2979b895e39a37cd151f66a9a31eba03ecaa0eaa1a40e5dbef90a6504cb239f8ba7527ed1f0d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbddda1a8caef88c137644d87a8ab9cb07398eb45300fce94f77be4b56cd1ef69706d64e4f2ffe8ed460d4ba223fcf724b6a0b097d12c5155fceec62c33c6f08d20b861d19a7ec4f9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3de23d0af188e1b7ac4654c2eeefcd61f0fd5515d1fb1af71803202b97a3524079be90640814a735f5512cc001087c9d854d523c63aed5e066b75c182c3cc0bacd7c3a84b33d126d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95db02df403481561140d57b9d77f4e5b3404d32d9e48ee6be1044f04fcd59a84a2406f6f5abe5f69d2848879cb06ad2d0567c2170c2c8556752967d7453e180148df88e84129b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38cc6a212e9b8fbc21d9483730711b9a22f64bb7d73c80b6191a0b438f25ede682d0515b68081024bf66a4edf64244ddb30ab38a88e3e34d3ed115869b38bc36df5c3baf9fe02cee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h307771d0cf7005e74a779796af19c4b8dcfb8897da5c04e376fa4757ab414540e677ac9fde7f1ba143893fb7777463da614f419d7dfebaf5f35cc558652b74ee884224903dd9eb0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdabe35481482d31fee533389ff01fd49cbd2ce4dfbeded19205cb447c6a2643ad3613427858457285de9750d027a8fc812b2eeea312ae85d5dc8cf611a8fc57ab2333d37a569414b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc632d5b0607ba7aaa3c47b1bbc939fdc24074934ec26634805d79d7cb1c0424930e97cfc8a698da692526d071ba78efe9795948b7e7bbf4cfc9094889eab1fa030dcdc2089cb28b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b0fe2f7e791f94b96e21f650ffb3a5daf38415198131678851fe0300a27085f56f5f8cfe2d1dbeba2f8b0f87349ea02b0cb26cde64b2d4acdb1d53eeb4324d93a453fb0507e19b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h895d2e766e918afd0f3ab643252c95006f4d1f90a76753231ceababf9f363f3bf9df3b82e31f76916f056e48ab6e8026859037c8172a4dff5bd430020f8fdd5a017979f6cf79cdf7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61da5aaeeffc90e259afffb08abad666c6f2eb0ae6468aa9539b7239e2a10cd967d6f6faccd2d713052042fc06074fbaaf60054731895ad7a4976da5f0d8e14352e2948166457b09;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h37cf83462e97661a6222f5c70cfc1ad7397c16d0617f3fdbd168cb9cae5ba23b9e42a9b79cb902d5ce39e40a7324537f4d69a2428eceba7efae19b7aa7546fe9a7574a2656bee0c3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heed575c52aebec61cac0481cc6d79c11b28a15fa77a27d8ea1d67a9f7f547453e12636b2cfeb409061d3342db2fefa44dfa81975d2c60c54310845d71998c32d701e3aa32587ddd5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7bb6f7fd5e39e58bedf094414e510781c7494f90c774ae4c30d7ff62c85891502f1ec8a2fe7e097cfe36574dc094b97ccaed4e9d6b8ef06868044d19d80fe8a535a6bb08a8761af;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9580a6d89f64912bc058eb0a668d876edf2415710e40293b16043f9c2f48f4afce5af798ce13312172a623bbfe6cdcc6dafa13c460d13196eb76d21f5530a3514ff4d1002167e035;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2d870f9a1bf9909fcb9afd7b30bdd52707993901e740a5bcc7ea8bf563b636357ec00937cb6cb2a3a2aedf75cd98b93788b9bbd9e3cecfc89814d1596222873f21657485c6cacae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2d3983b5f589539bfaa42e72d257a14dc1e06c863a6887f4376889c65b3c3b61274b97f97c1fd98e9c851b360b8688457e184b8be1619c22fb98ad93158b68651ba979b3c7b7863;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2fcd163086857dad6d7d3dd75a06f3484b65a72f70b19e90b3a8a59c52a2a0a99f150ba7f463db9cc30ec0a421d26f7beee4444086f54eeef069d7c2e56a3e7b8312ce721010f38e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda42d589bbf20bd1671cfebee1e5f3fb479089edc0702d3c78eb2178bc02383400059bcfc442946b9f2f53f6018ec98a7e46e234042178cd02ddbbfea7ab09c23635537d86f8025f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdcd15d18d915b823ef9d27f9fb305c5b308fe891c5e8ae6f96e924542fedab1e012a7fd22b79a5d5a2035e7314bab210751fca9f6c2abc25c65fec05b11792fc85f32de0c3a85c8e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92ba89db3f59d87b123a346044af89e47304d4085f753b2bbe68295f3fce491543f85218c0665136c5e342228e257b36a54314c15ee20626b7cdc6bd03b77eec925808b4370f248f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd49b8a52de7d63d35254b245a6c7cf815aa9ceee97c519735b04cbdae91306e168d765d841111f47cc765f01960f8d47a75d27f2fc38dd684c628771b1f288d27912a3d15f133043;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8626333f5edefbd1a26fa38ba159a1606139d84215b2474f0487c1953d52ab30d744b662440d48cb977e884f2d2f121fa690145bb5b443080539715ac6011ed62306d95ad509132e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h622983fd4a7ed16027fb8efad63e1f738eb09e562c5e2d776b98ec5d09306a3eedddfd6a5da3aa7b7663b134be2c44ecff98101f84b180f82a44e93988b3dbdfc35f861cbdfd434b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8a6a08843d237132c9ce4eb12127e08fb278048027c99db27bfad4e1f4a21dad6055b7ed252fbed6979ff4414e56c657166a27f59eb6636d0f190b590e867fba1f0c2f52467e667;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdddf97800cb223e39e7113fb784a6fec0a336de40a1b541af4de22c7283c5f9ea599903c5ff1c1128b602a8090b51c7f6a45e43fe5fd0795b911f6596112a841d3dcea6e0a835f3a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdb232961f67904d7fb998b73dc84505eb06c038c848a515296c2a99e5059e5c31cc05e193e858424635443f13905b798fffcfae64ec64c7a2f7776ae38b7979eadc37ad5acf7aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he027e6dfdf6a6f96b97ee5c24673bbccb80d5c78a4d76d899ac0f0104c2fd5c590e64814f38de945f070d2e6347b37417bd6d1d228064a8df2d371a5e9ecdffe401d9fe910f21191;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb63c42989c0b79230c77e58a25d27f5e24254cf8a1a2a4cea4ee4b9e4c3b3ecf6c9896639e04638e985852bb7a9e541aa6ef4159168abd4db03b78d1fa2a9baedc980bd727c926a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2cd1a78d28cbb3610520f896d1dfeeb5feb4dd62f54988041526b00fb0611f7716f11d42ba77518391c031edcd378411f6726443e924b7585251032df6f39b990304386e53aa53e6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h354c812bfee19cbf5798f5af1a2401c97b7f214f3aee56c61bc855f611da6de00711fc245ec51179319b17daffb8e0731eb3afc5171871ec9c931f63f8895657156cee27dba62638;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heecccb34e5a056dfba57021062393d91bec00a650e9543f53b9dc78d16b5c2cb9cecd785e31571e320b452ca071124de5af17e3f24ae7eeb979926fef7cc947ca4ba003c98af3e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c59f7ba47cdaae513f717ce3175f41e9b835e83a617e5a994c8923ff774dec4f4cc9aed0852c9c93d55025398a7ec81b3a1f946542595e3eefeef20c91fa1722cc93753f7f5493;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc0047e01a833a05de4e901449bf815e06969d7f877181eb73b5ed944bb03bb57e12268a261d016f82485f19b1f007bd9cb8030394b41abadee1478413a784c67ede85d3d38da4cd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27efbc2db51b60e886a9e51f9e6b8e917dff6b0ed6cb3d861851f1ec575be1d2cec05205c33c65f57ba9073eed0e7ab0c32c516c9d663a3c60ffcc094bf30daaada8ad539fbebe21;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbbee0bcc8e52b29d25b90ccba54511427576a3306453fb65a9740b65ec1251dadc16af5b9a2e5bdd7b3bec264d42b0285c7d7abf53a7bd1bf0fd53be3f985dcf992acd2c32434d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7faf244aea40a43372cb40a345c12f1175a47bbd66c2f085ff57d44522c3897d197d3ea0bdadc8169c72a1757da8168ca70cc553632b23197ad1341cf1e93ddc1c67eb99267fde2e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4be23fb5baf39877c8f72cb639b61b4818255796f237f863bf8c197d6917c008d27c6eb66d285152fe84b69c2845860db78adbb662ca839bca63bd8edb3088733d7e5cea9d4e5116;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8427ee3b1e82d63948c11424bef5f912eede6262d6760f21839605fb7ae27d931eab7b1b776fa39f74c97d6f6e428b33a6d319f462785c4e04f9d1f2827bacc956626fce7584f493;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5406235a6fcea64eb0ef8f82eea5af7698f39eb16615c33a4b57ca568d67628b2df1d34dc6cc2701ce98710a61961e1b33cbf0029f1ffcd4b7eab8a2e3b32df7e614ec5808ee6af9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0cd7977684ae6c01069c8a267c0df3caf767bdd5e74cd92c89fc3271ce4b489155681206e1eb2b487b3b6528f181589de8a4d12f78a14bbfb5445b46016c44ff24c0607d4bf92f4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h594c5547da1152861131b4554f0fbcc4c5f6cca8d7367d93ebc18b285a916b48d89f7d7ec0798789c95c0e741b24c08f6cd7584b633e940700b568abd2def8f6dabfa90d24277428;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26f509cffc4e32cbc3171d1c9a1c5c07ba71be1e57a2999c52b800ef035d624740b3a425f3d80a41eeacd8164a3f0db2c54d29fa2181763d9faf799e32b32e42d512c10a9b58d99b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d4e0d9e719aae218bf15b7b44d35c24eec53d33e640351836b809ed26022f88707f1ce25b55e3bb1f013ee1c7da1b40145624ff04413cf66576b581c3fc931558abf06741e6c07c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff470ba9d3109290baf03025722744f8f72ba2fdd2e4a2ba5614d30d652ae144951198ff62206d71ca8b73bac837c6f2497a71f68ae350fe805398d73256487eaa0a2c1d60bebf0e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb40f91e6d75496823f29bce58a7e6777810d80997b4fb4e309cbbd4d83b2211ccbf9d6f37d7ee562ec3f11b6693d4727a3efd7e4a9ef34e347830815f2891d1a5ed4d077602b17e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c6c27ef393a4d619aaab56e7382db11978f89db8c33daa2178fea303cf5f8eb7b4d955760603d4533fa3193f2c07c94294a7c42d81c1422407c488893bcefe955b142598f9cb308;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e326203a6aa83c8cb58a1136831d4cf2d48c50fbd66772b091f9b08ce5653f473fe4529e29c1f119b293e3f87eb2f2fe47ff4d8546af7adfdce6b8ff672b0b0908dabea5d711fb6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b85141e1813694c7af83a5ba619f23dbb30224aa140477a2508bdbb1a2b3b2b4778332bb3554ed0e6ccf49143845287c3a4f1b862cb6bac11c5e42b5adb06d00ce8a24c2591b5e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h200a9c1ada8f9dcf4d849e93fb0399902c85e6bbda8d44e7fb4d67a0f23e36527340de91e1d805ec64c794933617b242e07ad6dab2c9a4664503a11e00b6bddfb139eb0f7fc0d1d2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9aaf81317fa0a1edeb09a1c5d0da7d126889cb0ef3365b57162507cdf67525738b621dc116a89110e4f21876d99e7182744f847d55fd9c050c777fa6d66ed783dac91832df3b2e18;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c034fbe08a5753c6a7d1d532528f8dd6156d48b810989715ef11f966d12171bc96fc35c483a0040a0922a237439bbabb27a4e4af89f0afeac71102c3507c5fc064975a3ec5a8820;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95ecd21efb334ac6594b994ba9efaa5c3e7c67e523bb9a2b410e6199c61a9f99ed78b9a87cc9129a1456492c39e64241b0aa7af81024573e16cc031aebf21f998f0e85188be6e84;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f6fc240982fdddeae3fb8613274bd94e978835d2d771eb5d000f5094fac731816612411613be369920f49756ce1a4b4152396aec6907c50e9159e5bfcc4c239ff1e4078609a98fd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35a5702185cee159f12056b35ea6d14c22037075b9382305774164845df84986b19940f8fc1875a61b5030f654f00dc6a2011270a18892f1ee073d3d28b97fec9d7217ca78d62dba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he69b946cff8759cd8bb723e579c397b2eb917cadbec27723eff04d9f2a1f0c7b4af99c18bce80e53310dcb5e7c45a26c10b066703e8a099ca3d605ab9e8ce1ef4b4a81be0e98bc87;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf7196748e3ba4aa5b6dd5eaae482cc3f6f88d330661593488aaf69440305d0679545d466835e5ab4d951b3adfb6af98ac82bd7ceb7fbc6b32a582b38fd3fc9fdbe49e902edcd1fc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48a84e8d00e9990f7fd6bd3ce20b41d7b761005cef4d7cf77817e8122963a573e30437d14ab6f7ed2d07f64d351340d66c2a2cd360712bedd3f848bfd7291f87db4adc7e1a0c056b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd6b3102d6ed5dae12217be4770a97f3cadd718f4170c26ea2980e101d24b9f88175c10d4022efb1771ee40fcbb2ec8d24927f9c6a6f8c0ae2ea25bdaf7cd3e13877a88abb01aa6c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc7f9ec3d1957d273f4ed86cdb7f06127de1df89b0c84f2af3e029114a7b95ed011144cccdd28df8e0d1afc2f09d5699b87baaf1cbdc942175a76f33956cf91b32f953833bdd6e3e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb09f062d59797b85be79a26c1f29a57100cd40bd5af3966a2a96093d89ce23b7e24ee440363bcf1659b6a62b6ee8b185f10ec3d27bd1445b3ee4addcf7beaee12c10842fbfbae502;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7b9565d1a0cc437fb7d8c489050631206d5f94c007e1eb901c5027c5524c900d4ccbd01ca889d58fae82ab44e85eb1ff997aee41a3d56bbdbd3479eed957da59d485e4ebfd1da25;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h521d55e5e27b93db58ff9e8a9bed8e443ae76bd12caf53481a53e5ddbc976e759897cc01134f5ec85c62be27d9e4d5d5d12c58d9ed2c9b1527d7ce3f4a3db329f65046503f0925c3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h37e1700ab02339b65ba154aab58aea8d339df158a98a80797c9f570672b8fa527364f01adebe632cecb121871b084066bc798e278fa73ef2aef02ccce8fef9fd909763537b4c5d99;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4de07d36f95b909f7c5b924ea8cf1b7bab891a500246a87fd0e55ea6f7159a8a16adcd50b2ee40eb98597ec6f23d6fdae4b07625edfe568cebc4a4d6ae7f0bdef8a3ba94d5260957;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19a927e6f4b071990cb80287cf9a249d25dcf87e124b81830a261a318fe40bc81c4d4b77f8dbcd54ab2ada0f1fcc1ac60cefb3fb2ddae208a9db23c7bfd51ab22f65471d56c7911d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f4be4668a8a65d44d4ef1ad71ef272d9018d0cca5879d1637dd8efc1e7c141a9a17ab28e144e65c253666a32a2930ba7ad3f0358b856da05a0ad0fe0537b896159bf452cd3ba221;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb45a2657f642d1b2bc4262f4d8686c16654c6af9e8da267dda450df35792844993e41788606134ead79dea22bc9d70a5c714701c7c74ce8d2e04a324636b98457d0b3836f86c0a3a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h773b3df8352d552f0ca404a409b055f188de5cf60b9a9be86a5c43f66ccd8972b37f39e13946e2fbe6ad8217befe7d2e411d2b99dc7e1cf461fac5b0e2f0118c8c456c7a98155d1b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50d7f536fc9aaa20a3e375062275dea0af802852f3786dc3e711d22137b25e9e567d197ebc33f3aee2e3b0a856ebf78e5117a73d4e7019493e3a959f2fdd5b332dc4184be9e56036;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde327a410c95351a51d0a09c8389ba60d1080237c7cd9201f0ab078843335b100700851518c1f5617fc6d71afbbde7ff0caca9d927da010c93b7a311790e35afbbf57e178a74c010;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf008f0d4ce0ccf07ea49c93ee92657ed7f0714e53e21c86bd2ed144ae2f891354306f61e64f18c0e4a410c8946d8c371b0e48f7682435bbc8f02d71e67688a6fd1b11cf7afa03dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1212b6caf6160b0f1a5f67fb93a2ffefbb9c0fafb553231dfb8b479779471df7e0cb4097a9efebfec7d6c88a3737feb1e012624b8c6af69057940f0eccf8f014efb4de48f3644057;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1ffb44357a0f0215d5b78e21e214b215ae77ac9b05eef0a89e347820a9e21f440ecf60941b9733567f11cfcaae05731ee5dfac97a3328023309e1f1ff6b07a064ce917b3958cdfd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc1672bc214780f95d2aad641661bf8c2688fee085cf4b76df84a86bd7c160f0d78a802541b0a5650404443cd9b60af93ab9e07625f830961c8acb8257b54f8aa70003424edf99f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h597ab2f25f6e7fc7b7331477959c8fb4e7408c708c3caa2f3de2d3bdc821ae05fb50e1e9bbf17202c73c7ffb8c3e18530d0da43e4946377aa7e592c39f56ccbeb03922e45feeea9b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6d1b5ad8240d73a48c7c784cfb44796175471fcc80479c7c65b04d1774c919b9051ad50e2a26c954dcf6539f604fc5e296111a29a7682b04110937d08f271d9f5c26256f3b79f34;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18bbac6b705f98b1d66c48e1fe9e245d06013709905209c92bdd0239a5721a0c15c16a317ebd8e964cf9880e21d76ee1fd1e25990f7b2f1dd7616e92ff82f0e92ea38d882bc3349a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h171e5b2fb75f42202a48d63f7f1e6c415937570406f0d515b90e90f0f0d81032409c1935c14efebf6d9bdc88363d60a18e2620c3478e075c0213015e97fe4edbec690356398ceb07;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87f6847a647b28d4e2cf27b086d9e634beb21e0d962462cc675c1c439fbe36beb90ba5689443badc48196a695686a04d39e1c98a7d81eea3ab257e7753f1c5c6cbe76573f796f11f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha47f41a5676b004d87367144a81a49ca5a254d1339b745a250734dd887443c3b7077da0bb74e09c777d4968ae335052389249855dc86283f61c76d32d537d624dbbb72db8594fba3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49e1fe93cb454d7f7c8c594dec98c8d784688c3e73f3d9a8304fd7b72890af99d9cf05254bb1d6e6ab7d138600cade38f4566720d01ef05ef95557616fb0085736b5eb164105d08e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd8a3fea64e83e59e41ac521c8a4c8ac140b74c070397e48d11bb9fc346bbcec71982a5878b0184be16375981d14066ba72eb7de8d00eccb1b0f64896cda08b390617c0ac99717ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h442a675b2ac3156fc3acd0737a7c85d9f3ec038ec7f9f924a32e4d821b5bac2c9bbc0d7ba858e39f6810ab6129827c4163e2c15ed91c58e19a77637c9207c9587c6538701ab9a9b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c83ff771f494a5c3bf0d780587b78b289f6cf38211fdb077d90b1ef00a130024c5eeb306ae45859cc2318d821e5dac5e339a63c04a973c389100bf7f6894f5d52a3f54e1ebc9cee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1a29476d710f1312e3b22944dd87ed35023b3f8f0c4dc1838aa7a7e91294aeb032325e20a050adeddf352bb934b9f2d62035b3c788b81be6fc373c429832b4f7b06c208c2e9ed5b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h530800325aaafbb62d27d0f334dca12d91f8e9848971bbe83677f4c76cae419a6783632ace816b5d4a4abd12d9faf0c42992d492ff5872ba59f1807a9842b61b106011f7a469f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f8cc4d8e2348904f392a0d4857e1146fb0e222c35ffa4718bc0e7e605201db00137e4779e2cc11edd68f96394e2c23c9b877eb5d60fffe26cdcb5e07378387d66ce610e5e22b656;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92bd951c509dc4e7f94ea89ca820628e47eee9d1492bcb6f28d71bae202f0815e02bb84d4eafcaa7ed8df1e4c55446a70d18a7a177ea9b837e802e9eaf179b90e72f6bd94bd7fc0d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h126de6ed1a2ffdac04126d5754216748bcf5f75dd109c19a1ccfc2f41889788660cfbc106e8a29892b2c9d85d90ca723d39946b16119258963f3efa36962c22f33881e68b4097132;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h635d35f49e9dad4693587e0a246e19a2b3401b76601f38e36ecaf9edf0dc30de9e7a8efb5cf438c7ab96936a9aee806df6bc2e101e4739dcc4361f86bb8c5c46f5072ce0d09543cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h407212edf14e80208c2a92d8a7ed058a929b02ad9692266d763ef230c3aa9222fb6f4e55b0f2b636e2aebbb19379e75d0a3365227ec0f5893a32a853603e9502dc4359086556f2f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a1b78667b589309aed53a6071d57d64ecf2e3979b48215558d45e7f8be317fe7ebd2500b4fc64e5bd2b65227f8df8bb01bff256d6f4c11cd811ac4ef95c17cf3a0f2370eaf337b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4fe978482fbef932ec6564aaa3b7b693e6bcde2486fe8e90fad8f7fef8fbdea57a4c45b733e304845e7894dcf7b249283669403cfc4e9caa87e5dd595597b4f1cfb638d4d9851e7c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32c1efb963c0403e2e9af72472e255b212109fbe8fb1e16f5b6143150829db139cdc8a7d06cc7d90efaccf113f61bd7177c13421f921db20d9e1b5e6615e5aa6e4b41e8a016b1cda;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86db62ecbcd0c730d97d079e26cb14930c2a8b1558c1a46165b46c2ff538b0762f096e140e9af63e4bfc0f68d870d22894c22d5e8722fcf3eaf1667fb5e3b41841ab5ec44ff86f1d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0ef1655aed91ec947bf3691f2c8eb5ef0cbeac16085c7e21b351c211bee67e5972579b0d6f61b738a676aa9314a1c7cdc1ec98dec914334ec0080ba6173c0685f30fa10a99f93e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68635b5c1b5688f79c7fee1c6557ae2af0286da0d5c28b63c3cac4c1c51b43ea7669c9e7a9906c5fe8966ad2be49675f0bbbfa9e2087773453a9b56dff5a66f6bb5c61b1d931d65;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfef48efe5e96dc05d2a23ef865aaf41791f47f6fb21503ea905365bb0b11d0fe344d985f85b03f9c6ffd9adaccb70dcb6531c1bfca7605c0fb8d473f2f228ecb5bc2b0d650928a8c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4ca8cd67915833897835998166f185698e32a9b2ef535c5ad2992c592214e4204b4f068c651af20962d20acf39148fdfe6a18e348017fc774c5323670e451f134bd503f1fccfcd7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1bb84fa30743122c9f916c3fd5310ad2124dd767506ea704dc47b98f8d61410b8d384623d20d73453d6d80be230cf421a61c98e8acdc9410023d3d27e936439ebf3fd058c49e67a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a3742b5f224915f76d3a54b35764e66387b08c05b1f9b76bd3a1ea082a7ec8fe99a0c8108a988e4a7f82f9a8cc67fbc0ba78fd03604853d031e23d95ad4a466bfad90c5bc940550;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57378bb7f7d422955bbcc30b18ff22817018255e064dd525278e5ca1768f1dea7f076d1e020b732440a369526054cf873afa8e173d62f2e6297ca8f0e5f3e1ed1e56d94d6b00290c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf796f8fc4f4d0fddea35e6b1afc20b9a5c62421e6b21f6631075507b52f28bb78714f6f1a3ff42acf5e1f07f91de26886fcae540b5cb05d0767f8268742ddc7974c32c98d1976008;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h787a177c4eb664279f10b8473538ab7b202b24ebf3b30c5442d54d5f1a3f5998e22df741ead79da58b130624f9804fc5bb44660f1230bd0212c8fa7916041cfe8fd39d498c950ed5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf16d35f502c945678c525b70e142850760471f6dd60063c20559697bbf80667f6c0570c753d240f2682b8a5d18a4b43215098cfe35f04811a2046e237929a9b02fcf49a030609c1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b23a6acca71bf97ed08c3911d5ba7830c6ff4622aa216983d20625cd145335cf3abcf49d4bc6797c1da1c3aa0f23d5629aaf2aef9911ac5d3acdff150242929644e893333e04768;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2cc4cf14234c8626aa187dab7049803bd0a44329889edf4ed8980ce2431d69024d742ec031336b8bf1bae6afbcbabb832ac9e0e2f0bf8b748bb4dc7e26a6c576ac2cb2fdf7071d2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8e68b26290c1c5135ca4975096b1714d3c1d7b54d4923206efe5336bfee8d9bb2364ce1d6ef8664e973fbc64609bb22a578a2b444fca9ef0e81550ab3451e8bf80f4d3aa85bb317;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34eb5a1eeeba6950505572ac61a89e3d0033f1cb898a6a67d78e94c9b22722c6e641387ba8a6a6ccc457019d999129ca2bf4694a46945ebaaad30dac83fcc92967862271c3b55617;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h812bb5fdcb1dc869281e2aa8b01e681e232a9d6c6e5105e62f80dddff7e9b5cf22d3b6e71c83a19186997dfb993e7836b2b5abc564f2401ca892925ad221c132b6c864c8dbbde52d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55e5abf26b8ab01cfed3bf82ec0ba6b322f4b7704da5fbb05cd9e8282d34002ad1a4928ea3d93084b08796b3ef3eacc0e573cc6ef45ae1914ac48434dc06d62f42138b057f01ee0f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36d8c1e5ee39a1500cd921b683a6a3cf81611d779e00c915d109c051aa8469d6934aefbb4c679d0213a88b6b3f872be69e91c3eb7896a6b74633008ef829ce53301c1badeda926bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd329552cf64451361447c3a8b294631f1f54a870578657d8ee4a04e2f51a43cafdbcbfb1a635ab5afce6fb924d2da626d27de79a755449f1164474947480713d0f5d85fd98622fe2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b6ac8cbdfde0fe257dfa659da16171dbace64c751019d5a8ce3b622c1da5cbf3f28f088a41ae53dfb4a3c8604ae9445c7e01b9a4e72291fcef78c1e10697b1415a578342513dad5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3ee05b12fa61ddc5c88de31ea24defeefc795220caca245611cd4de90a53a2137c110ff4b044a4b694f1354dd12a046248ea44a3ceaa8108e26e6c69fcad48744b75f5a821a564;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7811addd04dff1eebe0d764c1df4ced6de69cdc4819b8e925007b0d9729d0916aab4f825dcfcd74162124c1d1af0a049bd95570870dd20713b2899f682da9ae9d9ce1ee8c4877e12;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf372aa051b3503aeb7a04b21a5e73d14ba1cf0ef3f60a1c1b667044877f2d22a776045a9f0b124a434782176a6cc514d13bf037f92aff4f2205067b9ac331258f40681efe494536;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf814c6725db9bd47383b1f9e012b5e9f52dbf6cc600ece598b341410412c5ad9536a9ce3eea9b5b0027ef1d49e3e484910306c69e7a32d8cd14cd6c8c42c7a9b7c53b38544fdc891;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5869641b1d942710f47b27f6cbad7dd9cbd4d70b629591b3fbe8dd59b282e483c9cacf30341ce637d8a68c7f10aa463cad6726c106e858d98dcac55221d8961d70e70a9a77607764;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9b04d9c6e51032f944bfec31caff983e487ff2aec2573be630d6f6c759e50cdc05851a934fb2a10a6f0d063584b8917af81f4d3401ab419796f7f40c027ab6b563f287ffd5ea9e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haaf7a5d2fb45a9be5d752bea53b42a91ce54548af3fa5b41dd10adaadfadd80412ed3e8d0c0c3703bbadd00bf3262716fdd61b33810528b51b775c6c6fc16169d6b4519e3f6c3f0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb289289694742f2579b5f23ffc20ddb2df8ff9543a72043b20f6fb2043bc0d808775bdf5ba306d0de419c5b9fa997a58b7559befbfbe94351ca7301b0be05798c31f5bbc8ddd78fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6c8b2060bd2057c79f711d79f87288af5a33d6e2891e384badb5de5bc9539c6b80a6e0869e80f27a09db28c015e9f6ad635ee20cee55b51e9cd283c278f206a4e463efff08c2120;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c13a2b59838f3cb88143ed14094ac62d9915fc9e50bd8f87ca8d1ef77ffd7cabced7af723ed0043f7504acc22eee929da16bd44d0305ae28af2176d398a731fae763573257befbb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd2d090617c699f3da887176f6ec155e78c74d392a85d0ccc6bd82ec83cc880d5323c279481a3751f6b795252a80aeb04cbef19fe538e07d94d4c38a37fa9d6169c70cd81b641328;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87e40be3c31543bcd32373a5b2194e441084a687b50af23624bcf64220ced602dbc1a1594f2eea685da728182ea50fb62dec02f0ef3b7cda5baddda903e60583b39c5fdd065cfa34;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ab156e8c76411c6cd0f5484e9910330164a005f5da680d4609b257339bcef32d5b00ed7a80fd913fb38fcfb5d031fa726137a71c3aa41909828544dbc5bf17d546560939b867695;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedea17ddb6008af8e1449b8d39438314db05e080992c4bae618f599957f431847e50c52771a9faeba04778dacc9d98f46ad79d744567a2dbf00ccb6e0fb7b74dd49a57a54bbce37c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75251831d292d7f46d290970e4172ee5fb1eb3d57f7d79efe1239bf01b189abc049978fc5685f0299d7027c4172036e7f4713824ec864a4f1bb8c04118436ef8867322ffb415d923;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9a0b42b467e0e545548a0c0f1f6b67f81cb6adb063a321bf2e6eb539f56d2a42efb740e885c5c5cce641ac0e001e39656ac368ac5fbae147cbc5035fae99459644610a6b8955a8e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1e2fdb2afd6ce6f28c750ead67ad290e8ad19127632994ad790654bf664da67d664c589297227b6e5bd53833536bd0298131c12e727d337a0fad9ac4d41e4da288913a9338bef69;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52e5115e29b81e2319ca3e194746ee7b233f47a696ab4f290c3ca2fdad2e67ae7afddf43d82716e03e8c3476efd57d311aeecfc96e66bfcd7738d12b94936ca90d1ddd22f46b49bc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a7255b4832761aa6e3bcd6cc286c03966bb6ba43947784ec63f6761c07b7944e64db5248d53533b2b133c0767b3f415e9bc6a085fc9897466846be22a4bd277d036a88c73026ed0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb7b953914532fae627f85faf81c6bf78401308c0083f22e5417f9015f53c712bc3cccebc42dea43187b28a9063a6f276cbeaab22b591f177a382ee9cd4008076617d4709ef42e00;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb810aa81c79b87dcd56ee4ce237d6ff8e66f9688e10b30d16b66298d2aa2ec55a4dfe47968084635cc97967077f3e7f827363317e32d8b30262666a42d8e885917baa73d9beb114;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3dd9b1147b6106d00dee35834af3e925b18c621ea6803cad9234fdcfb2d56db2ec55725799056791e0bf2acb15b7a12215f55661614e3e550141bfa7dfc8d2b78a482cdd433fb77e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3909056174bae6ad339a030e789c0d1f58c5ad04bc43c0860dcac2d91abf919014cad6fc3d030325f81f804f2c51600c5c6bddaddca0e0d09032c24f60501939bdcf7943144705af;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9916410082d750f9388d00767d90a3c18b43ab28e0115200bc2694afbf90b5da2fb09bdbf33d3e4f9d45b484b09f08e11f03da5fa1f4cd6d7cfc9a56d3126bf3aa718e587000d7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd1f0f85f7d5853705cd145e8a034755d70b545de26c073aaef32cf7fb87c3fda6e11067319f13297002f8073ec9608f5cbc234135d5378e80c8d327ffa4e7ace9d19a09ddb65088;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa0a59d140418c744ac1b6bd742601fe0170b33c93fdd6688cfcec8883eaa140184759c7eeb7cbc852ac96d3343e759906754432f09f631e7ceea892458518a94aed4907c3590ed1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a3ec4b043a5860e06077ccd37509107bc537f067675cb2aa65c7bfdebded15decef393f9400caeba10964a08b2d4ce162184d084bbeaaa006f055a52c19196686d0b3df24aafad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1fed12d6300e3183e74699f3a13e6051b903515f2b361a56200883a5e6ac98f7312bfd8a304718361f78640670906935b09f48913ba83446a9cc6a34e18d6a9f175cd01896336f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h512246d1fbaad45ea1c564c43f0a37c422532d438c7188b4bcc68debfe3ce77e38cca557db892dea671b513f9ac074f28169312c6a0e493ed0e1f2e9c09e8d69265284d6fe948c33;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2353b01337c36b6f6bd421c6453215177c86f66cf30666fcba592a5d88ca4a9ac7e3e43b853f5184be4793b433cdf5e75c96a3fe30e3454399f6b643e873dd4054ba0d82c3aa9e60;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36a33bc1e816e5e78eb046cb8f2c73f0443487e246220d46a2198fce8135d18800ae5c7e0290c21a2e9ad2b2ac7c4376e69b6b10f99a02b6519546f28f9a6e5de37d59433c647a02;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3722d2fe916b9307b78b92060334f21dda351a47b7c3b170417af1efad80c80a4cb015162b9750f46ab0f95c84e90dea8fcc7beff5d62be03d00d6d04cf972a5017a28353c44eb72;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47ad1def3cea10d80ef34d9e2ecba64fdbfb3094f169c557faca870cea08463cc20fd3793569012e40254874737fd4442838f22109530079bc908e2c0f867ee2625485c0ff572585;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdc50425d124fd99debfe013d035e0323a4e5319b3a0b0d4dd0b69d71d42591de57a91622469952e2b7bc1a533ef7929053f4a5e1856d0686deb7141f45b6f15490319a2af9adba9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef9c7ac19f1da04141625115f5e228af63427200d346e45089ced0267d2413dd9b13a0d91dd884c09f7c51286f92c42454d017fd385ca56b0e954a1e98f1de04871a9ec2691b1ba0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23af5566c131fecbf1a74e12923085d2ffa369c90a6a09459effa6c655539bbd2cd629a26714003b019581a9fff9c2c596b107e521b931995e20449ea158b490a6dfcf8b43029530;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6463c7dcc6ffc4d0c5d8ffb9550cce2ed1cb39bf589df0f933fb73e77f72015a3df18a2a9071573091e6f2271e8ad76f565ca4d24906a3fb620a12b775bbd8ac8bba06499d527891;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a0b983d92ff16f71c01daef37efe79adc381c6195dff405a7a7ea3f8ecbb8cd1cc907d07d7e2415c08fbb5e41188b70749c5c57573f4e5f23e1e10b5c113fb4d1dd7eb580f30aed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd848097f081e3bc3408b312f275f848d261cf19c5f1d3fd1f54e3f29c88cc503ea839c531e1789d7631a8a9163008b9d5b67cc468d902334f27e8d4e4137451548f2fcf381775e4d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3caa4fec6a4e6dece6bce23030e2895f9b18195452b40821007adbf6fa2955a6b66f3004896ff7c1ea076fd7c626cd541ed1dec6e77a9627fb5c41efae24157cc08896b49aac6789;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb6988c9776b17b73a643da66e497ec195f8de1540ea6752f03bee0cc65ff697f8007c436a7d850cda65681cb9a1e32c00280aaee61cf200eb780b7cd7190334cb23ef8df8e3ec62;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1aa308aa11fce6d639c8361adbe50970a5739a9dc1a083fbe9ffa1ad564cecec929e7f558674a87275c8eef4f99008689d787e8c82078990daace7f120fd3512c9e3d24a6db168ec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3aa761b6a75cb39200a0333a6297d107577704e2aff96430a36eb096923fce171bda7bcff89b66ce424a0421a85074372e05802a210587d4f17aff7dcc3f304f38c1e3f783f17d2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ad92d76472f1ec5619a20ec7cc3baf74701eaa73adde1dd109bb20a980bf5ecf6d798229769bcce683b17f880991bd3f9d0b643a1fd6b7693f5d86e5fdd7f1b080806c86389dc45;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb14aadd3e3061642b8c531b79386a152a6270c1779f1313e5931f7bc4d491fcf012cf9fd72db6b8fe77fd0dbdad910a299063e5ebd7e60f87380860bc531382c34f9deab995ae9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfde442222a7eb2b94d1a85911e82a4cde2db0220504e0df17c56cef4ae049e46993026c6c7adc0a4830a4eb9c9e7cbaebfb683854315b402290b5bffe5a1be994d3de7b35a4aa496;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h864d7a38201a43644bd08437a7bfd90475032a581ee05eebc041e8e9c1d169c8ccfdbac392002e4c01587bd3630e559944f5844d419381fa5d014db9c311e1eb1d6e647ed81b4315;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc32478a2b24b71203a080de2c48acb5b4b7ba295fdd93b8b1d9bf1743bf358cd0a1eb0a252d8cba007ddde93d39f4663835dd0e2debc60893b6eec5b015eb90fefff0279cf79ddd0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd16f68dd0b1bbe5209b78a2fefde5f62f7dbf6089a0fb21222ea37d3c83d77da83d531e95babc709d8dc1989bf7ae41f5151d7e286e4e428ae45a4be1ce38dfe4b075a3faf77cb1f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3a1a7cbbdee0a2e727e15872de6ea2147b5b37c080a842f21dd75715947bbbf23c0adbb40e6882e9b0912ee7dc92680796b2b8504d29f447c306a144241d7e0092571ba5d95c185;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h326717df6c249111b682e5605604d69f98da7d1dd78f1c66b1662255f3911a89c137e4e33de71a393fa89f1225f9a22ece94a44a549fa005857912d1b4ef4263c845e39a7b71d719;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbfc3145b37e521aab2355d21e8f94bfa6ac010c33c6a4ff0042ebff6e85a30b55190c1bf34a54b64d20485c1c79ff87bd31405d2b27f898a739e389fd95fca0ce7fbbddcf4cfbe1b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8660212b0f7896b8f3e63c7a8a351cea0b688431730b51e6bce98bbebfc10683e0bbe28599d1af8f096d6970932a5ef45d8bcf2fd27340e2424cb203aafc91715da1f5d0cf410fa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40898c6d318d4cfa68f270010146a262f8560ab7018327d15edbe49c7dc6aa4ce2f190537f5de332f60395640d4cdcf866fd25409b2d1a06c699c215ff9e9c9776a7e294f4a434bc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b728e8da64579df07a57fe8c9062fd629b466db1f112f14e3295f8e8ae22fb47bad2aca6ef309100ece3b06b6c3c19a01ff8589bec192ebc0ad8b1d8eb033bda9fe1ee5e58eaf64;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9764dfb2070126eb0416f3f94cc274aae08429ca67ab0a8016f5a52f7408b703da7267039c7e14cbb1b2ea44ab787b515234514f6b9c4d22dbce69ec8c9a4e02431cac3282841f2d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd2a5d757c3a728f91b3cd1d85dba2aaf35606f298fe8c0da80a2b93fed40c97b9dea36b6ec234798ee0dba768748464f746d49ef72c850365d17c850f2f90102119456c4e9a40d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a1f9f75027932fea11df56c0114035268206954381fed85e22acd2806ac4ad04af28daac589ce2374439b1b05ee98d20c0839baed786e58389277b38c49db737816c8c7019f2975;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21b1ed45e3be012be64f9f3fc835f87746d2a4da3b2a42c6d6fc8813e6a6bc279ea85640eff1c161748d9bd36d9c83f8bf4f2d40a5679603baa17496ef85a1fe3d49433036c0822e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd73a29d129e0b3f9002a5ccdfc6a8a845d9e18479a5914ddc44faf0c8115da7ea28a45ea74bf1f8940e0fdc6e3458fba10a676d677020995a8fc63e1f25f26f0d447742c96526f69;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6117a9f49cb67029acec9d045a2ce4292ee9adf8e2bbca60bed8e7f96b2e92699fc0016cc45713d171cd86e7ec4c09409e4b7c4b71caf5e4919921918a0d6fc3d7628f8b129373e6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7de348463f5221ed9058f5a4fe9580fd7ed54814de411d2b7ffc1f2e279d96173ea765c6fcc092a0faa8494c84c4cbe5da64d6d411d3bf84fefa970b52b261937306cdafa4775716;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ea364a4225e176ae6e7a5efce142c2c315d39a0bc7d29374b4b785b3eccdb002c16dcf4ca67d3b18ba4de8f35218e2eafb4aa591eb6f67af7da570c93c689f77b8d96c823e9520f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9f74d46d70292c394edf618e770f0b7a91e7f19cd06d3bcc36a227dc0937037a2a3c0a4a6eaf96896d53ad1d0c6b9e28ee34eab12675a247624a92eae8dd8b6c963333ac982bda1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h214ed216fa19169d39776e7ed28ea591be78ae34594ba92333a595bf2fd341e784c10b4da4554fbaf4c1271e5a6dca945131b832065c13553dd21c5b17483b7f9faa29d28eee8dc4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc17e43e2ada7e1f891bec8bddb72527b256f533b91ac76d3424ceda9679dff5cacf38122058d4894fe538c018d27068325fc390444caad46f8c8f5d1483468bbcdc06c0f1e10b4b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h859ba390646951fc4b0a6026a2be9801f87e08815ce1c20d9f57ffb2b90068cc1e7d50ff68717cc175d4c389101b4804b422217a45d79b4e608a73d6cb3f789bd65b18a01eeb7d82;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heaa5fab8998edebe2028b6c605d5b2c191fcc96500bd247bc296a3c5f632d8ccfd72b8d5aa26505c434fc6cccbd0d2142d53b45528216712efd7cde0bb34b66b081a603e990ad83;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a995167cc34ddc743ec334391474df5466743d1c71bca72502d5c47a057a6c27a2a2a983b34a40856cd0cbe2aab939189a8b6c7cda20f80de6395f8a8180aac81fff55c4b47559f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1c24aa44f31138f5d612c1a662cfb2f490d07f02c9c929430169baeb882d51da2e5f54d75fe345d57942c8da6f0a92c0d3e7ce3866db652d4735320ff300847ebc4c09d092a191a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8400fdfd8867e43a8439b5775455285d83570476b88cf47cd9beb80931c5d5e9045f6a4914f905d193e95a9157570dbbfce2a29e4e95c50a2a24304963672d70ff8d76e6142f48e9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ef4efdab6c35b96fdc3f432ed7b6326c3a6ba7848c29d3dcc3174e16864511b919aa087cb82846068921317dc399d2b6ac459bf5fb08052a57113721f9d9ebbc09a4ec35d742a40;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc4044254c2aee1fbf39e01faab92a82af530f24261758037bfe6da5e7ea1dcbe2583bd7cc190261317dbc79e0ff94ff06cf6361542315f7413b9c8b1c46222ca072194f3d067128;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hadd7e70d0d9fb849303439978c38e0042c05a39a907f5ee746aea5f9a9383de222a28846724e4025d579d411f17741e2211de7e72167a3742a76bd68ace0670fe8718f1ff97cdf62;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41251881566d29dc23c9b71204b8a6908dfe30fd3c955475bc5468fc59f4334495b0bd5f45a3ab952ff027cbca273cef1f11f83516b42a71210d79936191227ac781fb03e8fcc5b0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8df590a953618adc225a2e9eab8293b1df40e7318d32eec8763395d40be33323045e3bb359247799cf799e0cc3873fd84b67a13522f21d8bef7497d7a5983cb0fb9751e1bb53d55;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9d3394821a92390acdbf780c4c4292a3ed44e9223823584d2d4ded7b4f164943e49a533dbb22160ac8f9b8e3b846cb229eb4238e918c0a501cdbd04039d56e2921f25d8881cf483;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8c87b57850363df7b7eb5c2e41e4bd50b6ecbb072ff158c1fe574a0e5fe919b0c5862f23e917bb57eb109080870eaa9fbb80d93d80f343568cd53ccd5a1f021b19e3f53224f18dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92c8133004d0616933f621ff2259a5ee6de2fdd7495c130554b877fbb7e9e40d45f1538431e90136e08533a81b3b57e7761793d653e55fddf1456d4d0640e2962c76834ff890c61b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa1d1acbdb733ea444df69854d83420b8ac8499cfe065b0534aa867e68ca033a98a15bf332d411c9c3cf47120342ba1b50a932f8412db4c47a1a1e02cf839ced3286d49b95722f08;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc97c6e49ae528c771dee7571bf370657f63b466a2b6710ea388d5384b0cb218ac477149e79a6f5bcf0d8cc434f4ee9910bd24f989d1238549de0aec11125826b338876a0a4abf7d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60f259ac556335f5415c1b435acde4611b000c5d43a56d882d921fc433138f9d3e222e5f63eab901944dcbea6bde5651f1f61476674bda86cc4a57ca192dc555b14cb557d61fcaf5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8af4890f65c31cc0b5b9d3c0892ba8aad1edb00ab57e6c635701953b14e3d00c9aa011e3a511ef2a3abc0156db55a932b7b01432ea0da8af7d82824691f4cd9eb9c1ecfd6907fd89;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e269901935f342413491b41f922ab92cccb1d7bdc0c440a635ccf6551865f772bde61710e1ec0bf00a73fa54d8c0147896624d9aea9ff6c41fdabc16742d27e0f357ebd6f179428;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4fa6d582051dc08f21c51330b6bf3bc5685394fa93db0c9e75ca60f07ad5c52905265ecf5fddd11c0b2fc9ad5c2a40d5da40a15b1b46c4336c06fab24578f774ff6ba6214448b20b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hafd9f64a459b31aaf7041405f04b2a492de82ca02e7383b75168fbd66ee78b438a450b488c4c01bb51e710b70aee7ae4732b76b4cb3a0f34052200a80c62c16f2ae6b02a006d6f71;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb1bbb835bbfcc63060dd90cfdb86fc5a6242386601ba7e323232fbb57af5cf9859884f2dbe490e443ac01078ae0f5bee148654fb0d3301212c8906428c72999925d31a57e019c1d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h866c9e9aa9e3039b962607575da5621537bf802aa7584f6d8d0490d1887538509203101376bfbed98f78edef38b65e7c0922761e9d8c77803785d53e946664aaa1d427f7a833af0b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47415e65af7e00382dbbca43defdd6297144a0ded6dc756f1d840f7b0c37a46ab88dc1cc755a1e147f1141d62ce54a202810a22bfdad1aa9964ee28e54fdd7022d74ebcf006dc47;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b057708c373ff6e7411e6a1d105099a3a126853549cc375c88637387d07da3941f1c6ff64f4ff2311a6390457a638aec3c247fc670e165121be29a6efe2d0d7d412f767c086a936;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1f39d6c5902856b541b5cd53b4d9c89c04d784faefe29cc176954f7242353a1e6bc7f2446c31a968e7977629fed44e1695fda6057329c89b90395674b187a844d5b16eb9ea625ba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2517c313ecfdd40cea682f560bdaf2b446945d0d6c3db124d97c100dae05000c7818ec9d880a0a0f3c8a4938377b53b7a2218421a7ce17333e5e05399e1c3eff71833e1a92151ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45214a7c367cd6ebad530004ab97c84bd46c3f5df82bbf54bb6db25ef8f8c73558854fd1e14942b7a4314956a58d4da6c5a5fceb7878563dbef7ec80d46f049f5ddfad5380b79782;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5e3b990947139a4018a99049ccab9f06547b8f3499ef9520b6ab5518e75dc8737cc52b9e64b7824f6ad13df7d2570ff2149121f4564654112789e531be5e29f5f7de33a958811c0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cd521b08ba9f0f22fcded8c3df3028dc16b3097d311fc497b0f1082c14a2d3af637d3881bd9bf622d03717a30c98b734277839ad32b221e9a5392a79d3a1100bcfceb932c2f01cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haedaaa2793e4e2e97096a9bdf7d6cbfe41cfac9f5b6bbd89458cf897c7b9e1bc8e82d1f655d7d526845e794d53c2933f4e8ac3be6768c90f714128fad75338c7a684e18af96dd14;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12a66f9a3c8313b636fc0117c53f0f7a2ee9e7aba3bbdfaca4c37d9200408a1454c4f4d82d525dbcf54e091c6d7c536e2d04d70fee8fc21b11317b902b80245c1e65c13e3a153312;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55cf17e13d114d7caa54fb7658343b06efbe654622bcc56576b478d42bf2469942a7666d115d4eed7826e742b22499ea3b4024fcaadccbfa0b889d28716c8b7ad78445e8a4d09e28;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b50d21bc0d6f23baf5576dcd5edba5b854762b78cfdcdc61c6e3d8eb487e90c9ae3c34b3807a07a1137ad3d26c218761941e24f2f84ca99126d4af3a2cc5d19dde690ffea242b0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fb40c9abfcd717056500e152a65ef4428f67477d6189302ba69fa3e8e6e8fc6d7e9912b2401f75cf40fea98982200270b7adfe864a623a9cbdd354738ea232e64b718007a74db36;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha882995047b2e4c1470cdf6a18715dac7e5f9cda137a41be437ef0fbae90b650c527079fab5048e5a2491a0e9bf10141d4b1fc2e8f5e9e2c94d85a981bbbccf221c5f053ee9fa6fa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc9cd3949598a42176f0e9d7bade011885145b044a6c7a2a5c3f3e4426187366a651b9801fc50424ebdf7de120ad0c1c141843640e6daa3d5fd8b3632f1110b9bc074ea078ac94a2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h103765505f9381215da003b97fb03e9e9add33db67dca5beeda9c167b19cb6dbc46bbf6c0b1b9b80013d2d3f4dbd02a2a04cf39ae04763b882efab05ab0b1e30eafdc366cd2c98bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d68c87da2fc1777430ecca59d7349fab0c08c839b1934c459a473c905bdd8913cadbad8df3d9b0f5beed16d7446ead754d4e9aae5b5ded253f03e86af29d29ce0cad5d64f183e77;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f356aa9436eac78616e7acb66cd0943949a4a0564aee397831a095cebc23467a3b8ec907741e1545e6fa053313198639e591aa013a97e45cdeea89fd993dd1e2410574570df5a20;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd028868c0a1eb9280c39c0c650ccc873c2e87f0ddb8a23d7ed5ff304750b56813d79f693663ce589a9c370853641c8ed9bcacaaec910812ca999ec0d163af5c2018cb8918b00045;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf66eafcf3012ec079d292ff004b747abffc8ece2c069594b4410caf6e09260dfd6be1fb12f42d0ab30f1e3b6bfc90cb974e346d74a7769077c383dc7a986e25f777f731d2c688eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha662fe2ff87b617ca8bdae8154b863f098aeb2c04969b26a17f9f18053733132ef3fc9224b47c8f16627c853bc1ac4a17f9fbee338a4b3bc6086463d83ddaf5e94951a9e416cc7a8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdcc296a7259209cd6abc84c0c19578a805a1026852a5a81d4bbc9ae51acef2156eee61021bcd68ed3af3709f36777aa7b00e3905f739c65a31f554eb53ed7d6fad07d032c59c39ea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ab388e0c349ccc7be7eec1857b27fe74bf52ce7af335c2e14bf5ebf799f6ae86c6a592f85415f0f21e9f9dc594e5cec6478b4cb5303c12c743757139a570f05c6a2788cc6806c88;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b77cc0e038d42c39ed0397b7c74db2259e5c86167db7df5a3b3df5228881feb6390398c09b2d03a9cf78022170bc513c494af2396f15ff0c2a0ca518d9e00f10d84e078aa27da48;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7579546ca72a405231416bcd84f01b760e7afbd3b58e0f74647cf4a1d90af7e843febd3b2ef09836d92c5e94484a187d984db6e0adf44139605e9ec973f5115b361161943b09468d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb822ddbb746d078ee100b12c89562ea69a2cc19ddf8cf0d03365ebc4c9e4865370bf33277991f7e4fe30f69cdb0466e1983980ce0be80d7f43d5c6d1a84a2b319ede2ae417214642;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8621e2bd3c4ee2855a59adac8421691c1479c85a691f5e4ee9d08b8f46123eaae74d455181483f749ffe2de0a80fa40634e6faaebfa263d4643a533f683d7abe9823042894bc8110;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55e6d284bd17553a93044e1bab0efaa050f377d303c73ac359cb3084d73f9c663c0017a9d8982f56807f162c48d1b05bae99f3345ec488543c5c46192f3c8ba41fca1fd5987ead1c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0b386c8619e950b836e1cb52f7cd28640f13ad13b322ca3437a2ce1bfe88e7d94f2e269dfbd2106c4077ecd10fd0cbeb190fcb08ab4fa34f1fb49cbbaa971d252c13492b788a466;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa1cce449a3f8548062cc1f8612b6c03751adb2a636406c8feabf8c6ee31eede1f1bc79bb7a3a6da77b80cbf606f8ac294d188a554219bcc337b02c1835d7e2b2d85f22b5c09b241;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea0fbb477a59b9a4b9352b45c8db24fcd00f6e9218f34fdbaa4aa3c6fd9252a1af3e4ba74e97eb03d478109ab7e61c9e7eda1e3483b5b31a91b21045d8b74ce9eb21bf8c78fb844b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0df2b3c31949f524551dae167e61d95ee9a6a02a7a4bcbe20309c1fea573827a7890ca17a7af94463bcaff7bfd03d5269ba600305cdbba8882e3ee9b2f34ab8f062c6478330747b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc17bec6d38f5b932fb18c7742dbeb3b73ce77a9a8c8812a1c96e3e320c7f0ae972cdcd2eaec05f2bb146f0c305bc5dfab6362431b6a93375d4ebc3589c0f8424ac19937a8d9beaac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda3b18f9f858b44a4ea52f6d386a51e7af52bc90965f40d3d6e83246585d951fcae5347b0ffd5c783ad428adcd779bb0feec00c1d5f2dd1e28ca6a2c498f35d16396fd9f53ddc84d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41965948d8e4eea400b5fc99f8181915e1fca46e22d6e21507c0539d425706f670f7527e0ce5bc5d1fdbda5ab8c508a460e632bf837e6914cb44274518707369ef723560eb4e98c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b327ffa57e69b1a18496543501d22af0e62e83aab84569dd22903adfd28b70dc86fcccdeb2aadc1a6ce4f17b20161c7de5440abeface134051b723b1285478a4cc29f53aff16a00;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha39aee2b96addffab34b82e4bec69382c009b50fee978c967a07401585740f8d7f19bf9b18554b0e8824b71f496fc3538b95bfc72f287aa6689f52ba28c15f1b02bdf8616d04306f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb92f762eb2e5e239130209e8af0da84d38d4c79b98e53d436a54add9a084a846aa7d2dfc18812a5f2e3d9efa3e8a7bb2f7566543687b692d88d6a649f9bf3d065c9f156bc8a0f94;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1092eb5a5123cb05f81b25945dda6b1274e9ad320e31d5128de3e04e15cb9364b91c5fd197678e1ae88b92bca454bb6dd6956869bb5272a50f14a0f6eaa8d3161f1be73e65cd026;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93ceee1a6ff98b4eba9fa2ced4d9e95e9013648a6ac5e737f78bce8e84dbae11a81c4310ea98c5e4471020c1532846415880ffffd6a7067ccda611d6a3fbc643845fc89801b8b465;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa3ea3e4fd03fb4c98f9f2e11581478dc6aebe3d86a4f2ab686cad586c662ade3161a4e7cfbe4835efbf93cfba1779941405fbaeabe70b9551484f6f89b15d3f235218b239756bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42fa1d5a0e3f98b9cb2c832c47c9fcde2bb12a585c382252997486dd08e57db9d224d63c504a2e225e732e6f7a28e4193ecf679b007c827fd90cdd120272fb3e77e6eb83c7481d10;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d692174551ce31acc8a63d17f5f81d281582e798e8fc2f856e8726495e5961cde31a9cba843bc1447c650a152d7da7286c368ad271a58ec13bd8e7b6d05d08f9ac0dc26673dd899;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5678cf843d1e1ea5aedadcb12ebbdf6f8edf00b10ee5e89c5345dbaf58b4ec51e4f8e4b0fdb7626507166ba8bfe936d3e6312ebdcf4f640f2d6f11538ef8d0ca29f218f893385971;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he45e52edc7cd122ac808bea095c462f9290b97af9d65b9fdc3c709549d2f4abf4f02311411eebc6bcf8e1668bb9f1824ba247b36c300bb01d4cddb36b2a9f7afb423cb5a3665b29f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5291f690cf45e5cb0ac76e4b7cbd416e44f4309014d5ec2d30a27e9caee6cd05b2cdf1e90b21e6cfdd8d78eb873cc5421bc321f95c4201524ac379a229ccfe8bca004ea0dbc513e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h546daecc7917882878bbe74c35f24c502503e5635c28d04dc8c509f16deadb342c4fcef9f811c25391ef383579d5a90492f1da5c93307ad546654fb8692ded12f632a51afe45a4b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h841625877bf13621b42604738b8cd88a192c0680c57fcd642696012098039962be144d34ee5f404b1ff8a44c2bd68252acd21eef549c02b5d0dbe481fd36c7eca4702cec1c4fa4ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab00e40fe1ce11af7e17e74fc3cdc49b78def675673b1f880365e54612d7a60fa899d5e321fdec4f0e2bb43eacf2d65c2a8e9e642f5c57f6361af73c480c9d6e13661b608829d1b2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26a4697d2d235522e2f2ee85283fe4c7952442d8e26eb90a75477bfda81c26b48eff7a1cb73669280c430c07fa0c44a6c7c9a86a0697ad41e48a6ab58e3ec60dd29550226b1cd5e6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3024a6a0d1d72eabf5741874191d9a2498cfd9d1cc80fa8bda2d200082d20ac787c5cc63d72274b86afbeaad4031a2e2802e3e160ceedca1f1c8ca0bd2543bf15e4c43dd650854fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c27ff35916eb612546f5239067e20e947f987d29df1f371c14fa80bea23a522f89cc010b709e3a25bd9e92eda7c0471640a26a58a7d666b703bb6217df0e38520756b6bbd19b9c0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92bd0c9b38fc5fbd92ec5910bd9a4c245b374d53abba4b81da75bd76802a71480ed26682796f5de23d50eb42e7c9b81e211788b9bd8fc52b51a4e174017b414d0fe1aead5377fbc6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21512a1092f4407f1a5913d378458069e0325056b4e39469eeb52549032cbe291e8bac937af055d8ecd4cf31bf70c2b687fe536b7b9c0a19631142431424bc14fa26e6e3639e0b56;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90b71b38345a916fb25492092b3f7bc079d54ea7404b458b97a0d8e0a9499d416f71ccadb70d00dcebfd31635b3fbff40bd1f6491979229d5843c1bb9c0e5b74ebc37e4507f98877;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9467badbba62bb24bbf215fe1cd38331905df868b529937e669e101faf474c723a80dfdb12f923e1a8933e126e66c672a919168e14d9bb09fa128c0f6c9a9e7c04f4ff511537134a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ab6660a9f8743606d2f9300455ae8cc505103a4f15b4b214171ab6c01fcfb5201d05268760988c979c2a7f68ee5e172ed4cd543e8a84aff20938b507969e73e4ad3cf446160128e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2f6f7dc04f0c4e2f7d49897925d0ee167a5ec7dd59b80c6c27d5845fa3fb16a1a88ddf7abbad28d9ce3f96e0d1f3b3920225dc7fd09c39b5a377cacf89611b81c0010a341780da5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f2a4685fd9d57e17d11e24d628495e5611b728484c280ee9748d447e77232d14472b8a23a9fe1e499737a82eae85101c14dd6cb1c58f707389681493be51f6137377f2f3f0cf6a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h457a10f1c10ceb8948385156b0c020d734e824521735c2faf51b6309167cb903fe4cb64159317de1e4249894addf8453dde586a1504b390c5076b7c710654633039498b87f8b0c7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ffd61700102036d03dd545abf9b8e6c8013c9ee4bc58d70627a76a0955fd44f1c04e11373a5bf91825a9b0071c896b2e3a8994b42fd47a76688223e2cc00b74f89895e6fdca2701;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35b4932dbb4dd470592f4bd6a26fc6229df6d5839a6248bb3f4f0d35a0c3f81d12caa890570716ec47436124a4ce0c9574a5c0e1d6864b74c45af267522df38cb497d62f4dac4bc7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36563e0af2d95f4932745e3a4c50dcdd16de2be1c8b0a8195b85f2b92e18fb68b4372babeaf57b05c037da358788514a2844c88bafa3cdf8393e502f4ca59bcab99d16dc40e8c7d2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd7a6c38d6c1b5a17838fc0a23b41ca0d368015cda413370c34a91f5fe2030160558240e498817ee1bf490db2d3da8b0fe840f3b498c0ff801009576b571cac4562c164e1f663de7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ab1443db5e415fd3295e1b3178cc6221559f16d35c18f566181e91ceb0834703a87a609c2537e948e3d27b31bb2c6a6448e71d65bda1afb5ffd166d66feac1cf20a58a3153bcc7c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd376ce1c6e0d61414275abe8991e4740e375a83879eba7d3504b31192cae2a10d8040719910e27f4ed5c1144d9d9dc816432698b10b998d88430087a4ed1ee7193e37ee32daf45a2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99f7105b27ffe7f5e49f440b089309a71e0049e46b079120019d63b546d22fec534e75bd53dd476be06bc4fc2ac6a14fae9c47de257e4f1a77619bb0faa795048bcf7d17cd4dfad1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1661a26d02c5dd891c241dc49865c65cbe424db2d9607a1223fff87a600d14598a90cfdae57734da72ce55b87ffdf7c8e78a4621cee22e1e4a911debffdd074d5a79947c43d99996;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1041972284dfec47866b41a74e21a9bd26886507e01e54ad073f5f6fb80a05568e35a2d79a690eb97b58a19feda980134c3a80ea30cbd174a2fdf0c1d0b65f17d98ad83379204b64;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc29468afb68a47b66283a73bf5fd01e2de33ab9c4ce34b185ee3688c01b657bb3e125222bbddf2f374fe9336b1d446e3ea06de7eed8977407215ddd70edea33f36f1c06ad902eb81;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a23633ba4447627ee7c925f39003bacdf596b64d569db5d96825ab889953447b13f9dce2a26681cf7238a47ab950b930e7bde70056c5d30ec148c015b1aa64b23c098be6166d1ad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e0c53114717a8d0c0f1cbc857984c25f387b9bb6cb569e3425a700bf72ca81233519c2680f460445cbd0822e8e9eac698fbc05ac7291db9da7bfc9e010d5777ac448854ea0e5f1f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he556952a7611fdc00795397f21010f303edb1f5d7a1436663dc346618450cb2b5c87ed24b2aa95b0def844a468e0ca3bef6e57b210abb88d38f183dbdd8385d138264d57f7247d8d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31bff07982157ca00aebf619a0045d0703231f860ede8d26c415b11187d9594c9502ce708c30a011b6eec1e54368a029cfe253a22c68efc39806484436d08b1e5c578e6730989d03;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1ad7265113a5a66d8f33a5aecc6517e51390828ebeefd9b151d629eb140f9d9007361f69f13499e1ef8ad6166007b699d8d582957a5f0e119d6ae9168cec855544c6c5e769e24b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h369efdce77b254e2ddcde5930aa18b89b8873c69de58df8cf7afbf48fd91cf53a595e1bc6e9db544d941f9c14def390e504c177e7c4b30b23b85dffc4bd8aa29480b598f29d8dc4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he34fa98887b6b4cb61c2230219ba185b882ca43a8f449d3d6fe2515f582cda9ff98591636c44844f77d0a0dbd5f15a8ac2bf1ff09fb4dd67d2415ad0eda24801a05c4969843c7a65;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96636ea875a979ab3f435a9660b0efc81967de37690af4c5cdb46e5cdb6631c46a953a6d4dc66952795b5c10b2112ffa4752518d429e135d1a7c64af7b2841f2d6c3f6c0139d034e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he85c4548387383c2f3372143b86164d26290c6fab1c537200f5efc63488cca4ddb15f6d1bfc6d7a37d1d2f5f37a264bc8a6a9856012ee0f67f565eebc5cf2bdc4e8c217e63d773c0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3617ff8c6707c4c57a5dde2b3153d4eac856983db1904ffd122f2ff4c7499e393a6b9f95d171988a2dabaa672b2d27ce5d6f1617139d8a05a3ebf867af15db94852e9814e74bd6e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4abf4a612ead38a4c1e9110fc01dd43f4af7c2c1fa77c59ba8fbd4ade541576b021c037ed61224445564af177b8990f30a5721836288ce774e6c60983cdded4d2f7964f031680a6c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e01596001ccf88e0dabe9e98c9bc7844d643e1facbb7f7121add31967f71276e625d16efa4ab36944238223e241cd6399b552ea3b2ba72f62658853beab13cb028b4ef6c0b05f18;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcb989632a06f8898c8bd907d3131f8f8034b8affbb31362ff63949c49f6e7caaaef5420d7a6124a3a88285a9c531eba0ee0e3c92ebd608aa06cdda1d92153d7ee7e08f56dd6515f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c0493a0a44744673453320edf58eccb58c6313848c77407711736d198c19cee2c011fdd54715d163509daf0c2cd2e9a1193b7fbf7d96cc5098734210b8273138d063ddf72c5469e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3678d0a8107641a8bf4120f0b8997bb49346abf48fbf0978fbdc3a52fb7248142d419a471aa00274dd3e6327f729601e9be42efc0d8f801f1c9d8da043f5fac76648269df0c412d0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd4c4ce0481541e1aa5b16be6705e55e43cf75030f3d5901803b52fb7cac47dd0c17967310b241231b44063a37797998e87512c4b0ae4b71754013d047cb33da01d8ed5528739a5e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6554b7eede24e5ba8e37d53d5081faf4481057c2ea701e31a0ea5fb9e2f9b37bb34a0c9e5d678efe1ebdb4ba740fe7c8de59a61650e7fc653b866567594f7481c502f8411c49d476;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb64e94505c3ebb39838bbf489e7f86fcaf36e009b37864ac245865be19aa9aac4339ac96c699524d1521701331eff5333c523502c2242a3891a9795328b4db4b50df03c5028e94c0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97584fd2405c30e7d9d47d19c31170ad5582a35e1925bc72ac93cf7d72085ecf92dd01aed9729b226a6171762038c7aebd212666b7df7a4e6767f88da7eee48f180343abb2b005aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb27704e636d0d2460ec7b9d308bd35a1889a3fd272b22993c967871b9d2242d5f1614d22e1ff9f9696fcc6e502cd31df4163d91ad78af9f6b5d249ac7676ab1c4d039e8572780868;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88c22184e86566807c0c9a0cea3ad6e3a38b62fdae529c4b82866bbe4715d3cb6afa5b37c7e63f3844e68a34788af80efe439fd516f3394c08bc3c95552eac75b7eadc935b73dcce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haebc18b64ca7298a98a51892720140004729a4297fa43a0e8e0fef5d421c2bd06c99ad3bc0c25eb07f4967e69aecff9f8d893376f9d3945f3b47df7cdafc669c71728598e26cee11;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h190d8b074ed7a3b7d428a0f0d88b936de06cbc09587220f3e25747b183fd8d326c5dfbf223edc4425ca7f3b2dcac7def64ddb01ad79a219f02c26d0ab5ec728235a6d828068a9454;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb96a564fb202a39aa7df269acdec1c5ff524253713ecefe318e6f841c4079980f4dab5377069d70cc976ef9c6a118e82992d5e8c983af7240633e0a3b95ec13d288f5bf7c8894678;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8fe15a6eac1e506c84316e42e2051a33094252322321ac2c74cc81535866be224ce3dd01a2b5d1191e978b836a65241a00e726b0137558192a504a8c499e312055e5ac96e803f1db;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68e68bc66f09a963c8c41b90e19b6f5dd0bd7ac5471ba9845de83f160fb1995dda55b6614822bd78295ce33a11c160b0cb531c8dd98be0c35dc86b2db88c39ad5425965ba0086bef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he38567bd6197761378c41a0e2a952244fb71be3f446504c905483074ad12e1b13a5b2faa8d9a3e9a22cfa02e07cd5724c0678dfa48cebd2dae3302171875e1651c48b3a4561694a2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h769d85b32b898dc85bdf77f372482789c9ab9a6c6350ba7ba8de8b5b2c789aa81e5230485baf3d40cf7b370723c7e0848b1e4fb497699deade31b0bae056a2438ab7ef26095f5cff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93e5f5a20c4eda0d1c09c83bf7d24fbd06ac20df1be649d2a3f696b53e8e4afd7276a3edf05effd688dc248f64a1c4866a0bda0ba4c99cff5082a251840c371685342b33dd1f69b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca048f979b9cf24a2e843100f9dd50932838b08b0379e393eca25d34b840aacca28d06764c10bedee5a7e34f64a60ff429e1da106f2a8bde026bd5dfe94c269c2edfa6b6e37f5c73;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6219a85e950fe54d6f9109e1c8f1d4db5bd862d693a4d0d02fb97c3c195f353bca3e53a5bffaeac80a7273b7c345d2d8b714e44ee3a1f496ed8cdff6c97395e91bfae17b7c4700fd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49d645ffed9ff260f17423b42fe34c3ca18540b2b9fd2e75fffa93ff4fb6f0a20926ccb3410f91962846edea0d5875f2bd655e1093021091431f80c373af7a56d2d026a61745575c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3fb83c130a657b57b1d154ad1e487805447f86316177ec8ad426a0c879968f9ae7dfae580b2ce2615910efc933006e8083086aca15e74818390a463a1972e42bdb20b1bb16babbb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86284a2990e2992b8b6095f8669288e6866fe4af7e75214d0a4adb9f2343a4fe1d3bad7805453e8f5e20783560d86b5051f17626929abc9fc37b3b9411fde5fd570c58848bc4a0e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41d6180870b72857bee280c69e9ac09fe9e5447db7d00fc039d19eb56c8c67222e350c36475b43addb64e36a5760b63b900fbaddcdabf0bbcafb73c7789dc83ef33fbb299b5ddc43;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed3248d31916ee5bec770e3f5c2ea880aa8ffb0ae4dc398694ebcfeb583474dc0321b66dfd7a31ccdfc14d6f2814e81bba77ccc47f1cdaa0d99df8c87bb899849f140e88371e9792;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f15f17e4ec88b5245c677d2efb2fa75803a66a153127af270d97b286a6e94f9918ac62ef641a85af263485b2e5f78c0c2bce9ae25f63af3c2fc78eb13c197392d1d25300a5a795e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h615a39cdd8fc7222543ec2e04b3210988cdf86089e1d51e7abae035ea93d69200a22b00afcb692d4d05d3d77f9804882c4fbf3e00a120187c486e37e37bd74ff1b58d10f10f17887;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9bc642be3da193457e8b02fc89c693630650d0b2a824c8dfa6e404b9496109e57329bf7420c721cc4a11a7468c458fb9007bd0acb6ab645876c9cebb4f04112c93e9debdf5ee51b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h229bf41b9bb3ba67220c3450f4ef946fc1407c118ee7d0a262f15e58b8aa34a0631cd68cb80393b24c7a55863bcd13a99320ef11cade2d0dda0e248e02ec5472b492d0c54de8ccea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfae58dabff908655fbbd148e4a84a2d4f928e670c455b8e362e4da94a1d6e8f11a74cc6157793e95084ff01da4b0f7b1d2a92bf34f8e7ff8b54a13b29b1a84db131f076f7ecba80e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd297e6829a6b6508b3fdcca95093b69a12941e9584c98af7d76511bbc40372bb82ab17d39f418a5de637dcd24b08771bfb446c7c034ef4ac7841ee959ed19a0a91f19582db5ad7a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b241841eb61723e0e6b299b826f7405561faf997e8ad021ede8ec924298bb97237466166774c5a444f2781c2c939cfbdb182d8367dbaf64ca403d86975eebf5bcd6957705c91515;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36b3d6c461f1a5f1ef6e85daca5e0123d2a013847060f59e5dc79442ef926adc4d5a54191563239db2bd2eff8bf545a1cb1e172c13abb8de293b29e76cc9ff5266332f0e9db04816;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae9e5d5e58b0fd5231b546c71a85b53422cec80da674adc6428970d743d42cf857f7766b1c6018e8820070af5aa63800962585aa23416b2b61ea76a686442941697ef2591267ca35;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19eedce875d18240f2ad3b76fd1b355211713165e4905c6a76c565761e984826dcf1600c33b258bb3a52fc026be82b4df05022f6ea0015b0488422c78c1db65d3071b8d13d60ac56;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63aeff6d1fe330fb2551f9ee4f11764a7d76616a32f7b791f1aa75c5f0bea539d2567d5a78e15422fab523e81f7a82be9b4eaf2d46ff2c8b9331790d1bb4262378459971e62f7729;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53fbfcc41b643335b76c4df6bcea1af6600092646b25cf57a81827313e2abbd30159930920ed4a4df9c185b395034ac0ccbf8f0ee0a98a1435c29cd487d16529de9e2cadb6e2383a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae142de09f36c3ceea549507dd5e520220a2a9d3729bb61017b6b6cedcd34efcf21d8a18b41ce51699dc5e625b5d8383f5d4d6925a278c4c23191ba67c706e2ca51d31fa38672f9a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdb1cbe3eadfce2f8656ec50a4bfa29ad988ae70008c655e226ec399024b89d89884fcd41cd28545068fed2e894fcabf3401c867478bcd1b467f4173d163fe47ca15342103933167;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26eca782fe4fe39193a0573b7c1748cd45e1dee28b2d46b3171886c5efcb91cb7003809998229ccf8383de38a92e5f4c873fdd7413f1525f50d6cf41ef9d21b4d9d3fbc8510e327f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd74dd2c8a59b303188ee11ace414e98651162bf958d91a5ef17088b7c488d3b31ee5ac2a1601f12558f11b1a534bbe61a70cd97cb2a1548bbf8788e716cfc34f8c6ee0e1844711c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1541f0962d66baf7e2f00b74102e204abf3a5475f09df48d441bb2a2dba00c1f6296989998bda3038a6167ea9c286731321b73760fb4ea6cb4145ab36117a8bd31e3aef9df7c67;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d6260afef89368189e5a7e742d2c32c35515acbbcce4871bab881dc8443b6406b010defb5f22cdd1e9b8e791d59ae7435959233572b020e360ff7a412f7311a92f5bb571e9ce4fe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70284f95074293b6b15de2aac05fa446db3c824708738f36ebe3dd51070418dc82b02baa5d47273e310ac2e7eb818c1d745dde1f39fd6dabf08d52ad33fd4be3f861ae2a05d0ae76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a3e725872d1b4f79f4a8c29661e5b63ff044cb1347d6b302fa7af4362d6ec56703ec7b15a501f8aff75e448d171044d2a22eff377422753c777e7d5e2da6f96b7a70fe354996712;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc26f5fc6d85205c61af415a6b72e3ada8ea43584f9958961c95187106fc16e8096ea57d1973b403b8888fab19acce0deae455dd28551075b333b76fcbb95cb79a7c0d8b87b039ff6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75e03bcce68129d2e70f53101c1d76ba8454b04b80445cabb2a5eae3f4f7db22d9a859225c4fad5ae3b957008ce51ded45a9a5bb05d4a245fb9b5b0359bc2e91956077528d496faf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97bf0a981bccac49fd2695ed25d5e61fe221fd912cc7f1c4fecd03393e7b92e3b15b1a96bb8201d190648f449f04c7fa49158a4340a7771049c83877bf37ee6785c312d38d2ca74e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b77d0dc79984e13b338a36b8b569d5bf47925e152347058254c8d08b30e303f4d27e30f08d4b037c329b354f0754024a5f86e1710634b5eaf5057855130d039ba5f3af0f050363;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha95cd13082b3dd82766ed1f07eb706057d2c510db0dc69f96227ea32588937d81d1bc5038623bd7a06ff447b333da259fc132a5c702b547cce4ad6e48efa195b25416960ce9caf4a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b4a0d2f82324d6787536d0fee9956cec27102ce2c3793b8096af5affe957dc70f882259e7ab6eddef7b58e17382fb227328ebb747c7e0ae8ef980c4a38f7ec799e753c3ce5673e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35602c16c9f6c417d48077557946efaff721fc2534d56ed4c38eaf5e7a15ab8c0519fa8e7471e5fcff0444beef1109dbb3220814e2b88f92b34ef30e2a65aa850273cfdae4a0b47c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1a357daa0e314316fa6d609e9350d5646de06400fa2a5077b78fd7d4509462e3bc71af79e134b42ccd1775ef6522dec20d554616ca9eade5b05fcd96ae3e77dd3da030c3cf2e800;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc98d28524aed92da1138ed5659d28c8893c9e3010a467ea6e9b6e491c13b2921e0d5b8c3806d7b2c34862f343fd00e337cdef439c8ace2c874d2b68414637ab8bed7486ca61c0ab;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab0e59c9ffddb71c3187671e6fc69caab4a5d04b427178b33515d84ef98850618d883086704befc7bf8147b24f896815f523d7201dec82c152e85a2cbcf7d8e3dbc84630ddeb75e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6749de93cd930f57b4ae82a1af1a1949cb996d0d48f43d51dd79399629b29b7c1434e600529b41526712152c6cc04c5a7901331a1667b8af27ff75afe08769f65ebb9066e16c81c5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25eafbb8cf05715687a2ebc1981804ac20e78eeec1f89bda83b31130e92a93c89ae129977ef0bf92ca8a3296f5dc00508796034b75f8dd572d62c92c9abf8528d503a9a99f2cb9e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb028ba1a2e6064b73c2afd24180aa017a080cbf2056ede98d11877c022b1dbf6d3ddc0b7463b53445dc3427b664a1b866110018914f7525934b710f604c1ae546008e3f44d5ab4f8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h392878344ff7a3060499387fca58a85d124c48549f8d437266025c4a0fc77137026d290f161c1147ca1aee245a4eafb5f9d2e0da69408fcaedf86db07c176efb9c3b22c2296f0255;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h913ab9e537d7ceec32ab8692a67ff910450165be307287d42b78eb8b9dc9f6e6bb4bd006c5b6e785e9d9cb06067d8da65527c1dcfcb637ab635c8da0f2422ec4c3e8c47cda47d2d2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5352244d95eb3c069621c451dfb98ef0a05b0ea2230af21114792de8d4164ff9cb2ac79fd4b4f09a8e3c12c000754a8e4049b27dd97f32e205ca9c21dece4ad59f727fbee7a7ba43;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h641b830636b52b5433f0bb041516e11acd6ffd60037e35c11ddbbecf46f247d830838eec2797b4abb68a279a862412b50a2b9ae5ab8858409b9d6051c15b89d87b9d3033e45e9965;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3666ea2e344c74b7cf88efa14fb44240b2a629d8547149592970d372a15c91ca749d3c5f175da18ee96773bb6ab0eee50cead1dd0d3fc1b6997c10d4a8c91ee9c4cb02e16f49a30;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb82f4942003cccc83deb4a51dfb399ce35385a94cdb71d0289f56bddebd24172551b8b8a1c344f3a75978ccf9c8c0c94e242259978573e71f7894a3280469c27845d1b727d96f273;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ebf29f05b2c7b51610f732b78d57909fd042ac2a5fecfc20b80cfc2fed8356a9b22847688eb302d2c7d962e6a9595547362061c6166fdcafaa438148a7599e192247cad6cfe313f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc58bce1ee9c8b8e53252bb4712d0429f93845e7b2dd5ff6ce9a1efe986c150741bbf462959ec2aea810131cb54110d002e052185d7776a6a5e39aa5a3175e2760756f8365ae0a649;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha158db94f0b968db5fd7629e2edc00c82b9ed28790c2959cac643015d9875fe27754ba671f78da77be07fdd03f9f50fe30b19843574175267764d05f41f5e0cf7c5e4f9890d08d3b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had07798ea77673bba9dfd29d79466445143b1c63811edd1f4e363c1f0ed43fc3bd307797f6d7cd2b510bc64b30d9c0c0081efc52cf468c21b776421c24f21bce77c1eeacfecda0f3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h716e0a91147e3373aab98c1ed6c2dfbd7c9f10208ac18508097be048917c4cf10713345f59a9f587372353b1bac14e8a1c69bbe10e696ea54c2c60f956f10b4d45b175bab5bce3f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h357e53043dc825c1800b97bfdd5aeb06d9a2722210626c2b84745debff7771a6f9b804ffbf63eadeba57bf051bf43877a5528ef8f9bb482e32e1dc8821d87d58963163b1c61c0592;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2a63fba29ccfacc86dbe69d46228af028b0d640ac4d5598d9f1871d5412f9aff3c71ad8194d22b36127ff442f40eba0a40df0d5e78bc56524fe76db768a602a206abe5a33c2804c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa2f92f7ed31f8a4f813795a93083d78aeeb3ce840a23c4f24c3c347d8704f948517dccd26289b6616768c671c6cf35cb2b391ff60c5d73c17d4f711cf9ad319d2212ab918a30ed0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3322c21f21a8db65b8a88b921f3a3ae33948e89bcef600f9c64fb601dacd1c716b1d70bfac25ef886a1eca048558d69c47879668f234411dcf85b3a0cd52f28e86e0a4ceffa19afc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78803116c1717c3ab131aba678f33ead19be445d41a253818c381a31c26b7d933007d8164d582469e4688ea581fc7450bc96d22b78eee1d4ef358319d5ce4f3b55faedf3f15ef210;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0f1190103fd50ba9b2e3aedaab5380b532c8922d7fe8a07f989da41032f696de69dc1b15e2dd5c4e59ae67d6a65ba5dc1965d7641302c8f7a0663a7951c68ab0ec2ae9b45ab506;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h954419513e4577653eb4a099e6250f8a6309e6fa57345d85b625ce4f329aef003e44fd2a258d06963bd4811d0a698600776949220750850925943654d272ebebb04e7930ee9b70b0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h489b8419b16f9a86d8442075df69ef56086528095d8c3c454bfcfa4598e1572dedd017d172c5e91593b587ac1ceae316529efa90a00bdc02a9a4465226f41cd9bf5c6edb19ef202;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ae552b687080e682236e9c21607f0c0647ab17adff923487a2a6b6a8f444f6aa43ef96118b27cec792540d980af5565d23d605fecf90b66f8071982263fc81d4599176911c864c0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ffc545abb0ac9c398de5a1bc0d4012c10ee8244459a511fd028a970e8307bc9021a70ef3f882b66f346be6f694d9a6a19aa387d22e6eb611c1847f0e5c6f6179b5ec70d3dd8781a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habcb474c060bca21d84e6fc84d52d132c3246820b68337ec1bcafa45a7f1b90aa51a0ac8203ff6d0f73ecc75bf3789941ad49adba19cdc9007add3c2ad7743cdd22a1a8ad2229e20;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e689dd525c32620a14b1c7306c21604b6106aa835045e7928507a3831a4acca2c8f3a97a1bdd335b9e6a39115d105f458ab4429a4fea99672b70f25968581eedf5f4457b7b066dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h146c94bfa79bfc9bc0f7f9f3bc8b97442bcea27095d96beaab42689b481aaf2cf752bbff230fd33e56c1a94c80af7358503771f265f6c165ff9c8cde61272fd33bd88edb3c715960;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95774d8e1b6788a416fdbd9f3837f6053828ef3c877dc5061c2de592c7d8244b9c6241c303b4ff70fdab481895a8f277e9aed1e164a7e8c67483c04cb75841b69e984c5daa4f7f13;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cd6017b4a98214476b5aa0fb24aee9a1cd2c1b0c64b798f791c73daeade12e97587c0e568307f239947ec3cdb4d06632965c6cea14bb0666e7b6ebdeaee0a242bd87467a2fa9277;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb54bd1a8d9ad26d34ed85bbfe05f8c3ea03c3352ae2a0bf19a11855c618ae7dd898f54cfa7f8da7f0d41f7bfa76dc33f34b45b9d2d456d8862667fd3ac102f7d0144c16413d4d8ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c0c330551efde54aafe74f51ca923b84e418ad3c9e2757ca061ea5a904da1e2dd78d3009ef947563d488d3bce7063a95585806a1787ae4aebf7e6b412855909bd6fb122d9d5fa56;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fa29c339ab1c9a4e1fb723248208c9f966a2c2e018a137d3cee93d0ee8d2507e289be546498c9ff6179b62eb2f56c4f6e30bbd8cadd6f472c99613232dff9f2f0150e36a965dbbe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96363898130474663735814c214cbd9add28b3e0635a4aa7fcf0a65b358655603fa888601117aefadd92d58edbae675a652659a4132d91e4653d5b9eab1827cd80a0e151df689686;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3ad7a2418383c5c95ba4d01a431db042ca920dcd99129487ffeae62c278f0832af99561ec7370b311f8e8be04e620be310dd1d40f951e7ca58c553094504ac7b7fa91da638c1f53;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38b2045990aebfc334ba02e871507fb4a0eb33e6311d614b14b66e62548b62a7c2239d112dc891446b788ea45833ec4d03831bd3acaeeee874952c331542b8d250dd0b911a9ee29c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14723aa1a5e6e676132c9de1bd0b7daf0ab1c363046c13db70b1fab5b84efe6ec55252b816b064dbdd16a17f08958fd21b05b9daeff35fbda6edbec114f397e37c78dfb3f888a2c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha95ca1c79f3359dae81b9787db47ee3e2363894b6d7af1491d8cdb9c5c8a7a8887c5db0de6ecde4ca6599b99f0f8766a0a117b10582a3c6f1b60e6212e31ed28ba5c806afc51c7a2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h306f99a2f6afd23dcfed2bad5250e9d67bcbea91e39dad14ca0aded8362a3876d8a7efbc286be8ed6f20234f1a9233ac10a3a53c85504cbf4f5cc6179f29e7c716c1a89da9746d11;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0e345458ece6111db52bb79e3ce0b5adba5909a9e8ba8d0f3612535552a4de45cb8797af7afb479472ec0e9cc0b673fa95013f87c5f685bf6f5d1617fe90358c667ee50cad2e8c1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h700c67201df228f26ec271e88a2ebda70aed6a4ee95916c65ad987268f9ec3c81fdbb0fc7e9bc9cb4f91c5a8ce7305cdf0be996fed7b1fb8a5500b3a5c5d2be5cf2bb41d17c783ff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbcc56d2e0da1b7395428f42be5aa2144133361520a3a99e118eab61ebbb7c27619cb148ba3c45e70b61bb5db0e7e851faf2627956f3daab31f6208bdcb23b9e6ef97592fec023bd;
        #1
        $finish();
    end
endmodule
