module compressor2_1_128_16_shiftregister(input clk, input in_data0, input in_data1, input in_data2, input in_data3, input in_data4, input in_data5, input in_data6, input in_data7, input in_data8, input in_data9, input in_data10, input in_data11, input in_data12, input in_data13, input in_data14, input in_data15, input in_data16, input in_data17, input in_data18, input in_data19, input in_data20, input in_data21, input in_data22, input in_data23, input in_data24, input in_data25, input in_data26, input in_data27, input in_data28, input in_data29, input in_data30, input in_data31, input in_data32, input in_data33, input in_data34, input in_data35, input in_data36, input in_data37, input in_data38, input in_data39, input in_data40, input in_data41, input in_data42, input in_data43, input in_data44, input in_data45, input in_data46, input in_data47, input in_data48, input in_data49, input in_data50, input in_data51, input in_data52, input in_data53, input in_data54, input in_data55, input in_data56, input in_data57, input in_data58, input in_data59, input in_data60, input in_data61, input in_data62, input in_data63, input in_data64, input in_data65, input in_data66, input in_data67, input in_data68, input in_data69, input in_data70, input in_data71, input in_data72, input in_data73, input in_data74, input in_data75, input in_data76, input in_data77, input in_data78, input in_data79, input in_data80, input in_data81, input in_data82, input in_data83, input in_data84, input in_data85, input in_data86, input in_data87, input in_data88, input in_data89, input in_data90, input in_data91, input in_data92, input in_data93, input in_data94, input in_data95, input in_data96, input in_data97, input in_data98, input in_data99, input in_data100, input in_data101, input in_data102, input in_data103, input in_data104, input in_data105, input in_data106, input in_data107, input in_data108, input in_data109, input in_data110, input in_data111, input in_data112, input in_data113, input in_data114, input in_data115, input in_data116, input in_data117, input in_data118, input in_data119, input in_data120, input in_data121, input in_data122, input in_data123, input in_data124, input in_data125, input in_data126, input in_data127, output [22:0]dst);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    reg [15:0] src54;
    reg [15:0] src55;
    reg [15:0] src56;
    reg [15:0] src57;
    reg [15:0] src58;
    reg [15:0] src59;
    reg [15:0] src60;
    reg [15:0] src61;
    reg [15:0] src62;
    reg [15:0] src63;
    reg [15:0] src64;
    reg [15:0] src65;
    reg [15:0] src66;
    reg [15:0] src67;
    reg [15:0] src68;
    reg [15:0] src69;
    reg [15:0] src70;
    reg [15:0] src71;
    reg [15:0] src72;
    reg [15:0] src73;
    reg [15:0] src74;
    reg [15:0] src75;
    reg [15:0] src76;
    reg [15:0] src77;
    reg [15:0] src78;
    reg [15:0] src79;
    reg [15:0] src80;
    reg [15:0] src81;
    reg [15:0] src82;
    reg [15:0] src83;
    reg [15:0] src84;
    reg [15:0] src85;
    reg [15:0] src86;
    reg [15:0] src87;
    reg [15:0] src88;
    reg [15:0] src89;
    reg [15:0] src90;
    reg [15:0] src91;
    reg [15:0] src92;
    reg [15:0] src93;
    reg [15:0] src94;
    reg [15:0] src95;
    reg [15:0] src96;
    reg [15:0] src97;
    reg [15:0] src98;
    reg [15:0] src99;
    reg [15:0] src100;
    reg [15:0] src101;
    reg [15:0] src102;
    reg [15:0] src103;
    reg [15:0] src104;
    reg [15:0] src105;
    reg [15:0] src106;
    reg [15:0] src107;
    reg [15:0] src108;
    reg [15:0] src109;
    reg [15:0] src110;
    reg [15:0] src111;
    reg [15:0] src112;
    reg [15:0] src113;
    reg [15:0] src114;
    reg [15:0] src115;
    reg [15:0] src116;
    reg [15:0] src117;
    reg [15:0] src118;
    reg [15:0] src119;
    reg [15:0] src120;
    reg [15:0] src121;
    reg [15:0] src122;
    reg [15:0] src123;
    reg [15:0] src124;
    reg [15:0] src125;
    reg [15:0] src126;
    reg [15:0] src127;
    compressor2_1_128_16 compressor2_1_128_16(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .src26(src26), .src27(src27), .src28(src28), .src29(src29), .src30(src30), .src31(src31), .src32(src32), .src33(src33), .src34(src34), .src35(src35), .src36(src36), .src37(src37), .src38(src38), .src39(src39), .src40(src40), .src41(src41), .src42(src42), .src43(src43), .src44(src44), .src45(src45), .src46(src46), .src47(src47), .src48(src48), .src49(src49), .src50(src50), .src51(src51), .src52(src52), .src53(src53), .src54(src54), .src55(src55), .src56(src56), .src57(src57), .src58(src58), .src59(src59), .src60(src60), .src61(src61), .src62(src62), .src63(src63), .src64(src64), .src65(src65), .src66(src66), .src67(src67), .src68(src68), .src69(src69), .src70(src70), .src71(src71), .src72(src72), .src73(src73), .src74(src74), .src75(src75), .src76(src76), .src77(src77), .src78(src78), .src79(src79), .src80(src80), .src81(src81), .src82(src82), .src83(src83), .src84(src84), .src85(src85), .src86(src86), .src87(src87), .src88(src88), .src89(src89), .src90(src90), .src91(src91), .src92(src92), .src93(src93), .src94(src94), .src95(src95), .src96(src96), .src97(src97), .src98(src98), .src99(src99), .src100(src100), .src101(src101), .src102(src102), .src103(src103), .src104(src104), .src105(src105), .src106(src106), .src107(src107), .src108(src108), .src109(src109), .src110(src110), .src111(src111), .src112(src112), .src113(src113), .src114(src114), .src115(src115), .src116(src116), .src117(src117), .src118(src118), .src119(src119), .src120(src120), .src121(src121), .src122(src122), .src123(src123), .src124(src124), .src125(src125), .src126(src126), .src127(src127), .dst(dst));
    initial begin
        src0 <= 0;
        src1 <= 0;
        src2 <= 0;
        src3 <= 0;
        src4 <= 0;
        src5 <= 0;
        src6 <= 0;
        src7 <= 0;
        src8 <= 0;
        src9 <= 0;
        src10 <= 0;
        src11 <= 0;
        src12 <= 0;
        src13 <= 0;
        src14 <= 0;
        src15 <= 0;
        src16 <= 0;
        src17 <= 0;
        src18 <= 0;
        src19 <= 0;
        src20 <= 0;
        src21 <= 0;
        src22 <= 0;
        src23 <= 0;
        src24 <= 0;
        src25 <= 0;
        src26 <= 0;
        src27 <= 0;
        src28 <= 0;
        src29 <= 0;
        src30 <= 0;
        src31 <= 0;
        src32 <= 0;
        src33 <= 0;
        src34 <= 0;
        src35 <= 0;
        src36 <= 0;
        src37 <= 0;
        src38 <= 0;
        src39 <= 0;
        src40 <= 0;
        src41 <= 0;
        src42 <= 0;
        src43 <= 0;
        src44 <= 0;
        src45 <= 0;
        src46 <= 0;
        src47 <= 0;
        src48 <= 0;
        src49 <= 0;
        src50 <= 0;
        src51 <= 0;
        src52 <= 0;
        src53 <= 0;
        src54 <= 0;
        src55 <= 0;
        src56 <= 0;
        src57 <= 0;
        src58 <= 0;
        src59 <= 0;
        src60 <= 0;
        src61 <= 0;
        src62 <= 0;
        src63 <= 0;
        src64 <= 0;
        src65 <= 0;
        src66 <= 0;
        src67 <= 0;
        src68 <= 0;
        src69 <= 0;
        src70 <= 0;
        src71 <= 0;
        src72 <= 0;
        src73 <= 0;
        src74 <= 0;
        src75 <= 0;
        src76 <= 0;
        src77 <= 0;
        src78 <= 0;
        src79 <= 0;
        src80 <= 0;
        src81 <= 0;
        src82 <= 0;
        src83 <= 0;
        src84 <= 0;
        src85 <= 0;
        src86 <= 0;
        src87 <= 0;
        src88 <= 0;
        src89 <= 0;
        src90 <= 0;
        src91 <= 0;
        src92 <= 0;
        src93 <= 0;
        src94 <= 0;
        src95 <= 0;
        src96 <= 0;
        src97 <= 0;
        src98 <= 0;
        src99 <= 0;
        src100 <= 0;
        src101 <= 0;
        src102 <= 0;
        src103 <= 0;
        src104 <= 0;
        src105 <= 0;
        src106 <= 0;
        src107 <= 0;
        src108 <= 0;
        src109 <= 0;
        src110 <= 0;
        src111 <= 0;
        src112 <= 0;
        src113 <= 0;
        src114 <= 0;
        src115 <= 0;
        src116 <= 0;
        src117 <= 0;
        src118 <= 0;
        src119 <= 0;
        src120 <= 0;
        src121 <= 0;
        src122 <= 0;
        src123 <= 0;
        src124 <= 0;
        src125 <= 0;
        src126 <= 0;
        src127 <= 0;
    end
    always @(posedge clk) begin
        src0 <= {src0[14:0], in_data0};
        src1 <= {src1[14:0], in_data1};
        src2 <= {src2[14:0], in_data2};
        src3 <= {src3[14:0], in_data3};
        src4 <= {src4[14:0], in_data4};
        src5 <= {src5[14:0], in_data5};
        src6 <= {src6[14:0], in_data6};
        src7 <= {src7[14:0], in_data7};
        src8 <= {src8[14:0], in_data8};
        src9 <= {src9[14:0], in_data9};
        src10 <= {src10[14:0], in_data10};
        src11 <= {src11[14:0], in_data11};
        src12 <= {src12[14:0], in_data12};
        src13 <= {src13[14:0], in_data13};
        src14 <= {src14[14:0], in_data14};
        src15 <= {src15[14:0], in_data15};
        src16 <= {src16[14:0], in_data16};
        src17 <= {src17[14:0], in_data17};
        src18 <= {src18[14:0], in_data18};
        src19 <= {src19[14:0], in_data19};
        src20 <= {src20[14:0], in_data20};
        src21 <= {src21[14:0], in_data21};
        src22 <= {src22[14:0], in_data22};
        src23 <= {src23[14:0], in_data23};
        src24 <= {src24[14:0], in_data24};
        src25 <= {src25[14:0], in_data25};
        src26 <= {src26[14:0], in_data26};
        src27 <= {src27[14:0], in_data27};
        src28 <= {src28[14:0], in_data28};
        src29 <= {src29[14:0], in_data29};
        src30 <= {src30[14:0], in_data30};
        src31 <= {src31[14:0], in_data31};
        src32 <= {src32[14:0], in_data32};
        src33 <= {src33[14:0], in_data33};
        src34 <= {src34[14:0], in_data34};
        src35 <= {src35[14:0], in_data35};
        src36 <= {src36[14:0], in_data36};
        src37 <= {src37[14:0], in_data37};
        src38 <= {src38[14:0], in_data38};
        src39 <= {src39[14:0], in_data39};
        src40 <= {src40[14:0], in_data40};
        src41 <= {src41[14:0], in_data41};
        src42 <= {src42[14:0], in_data42};
        src43 <= {src43[14:0], in_data43};
        src44 <= {src44[14:0], in_data44};
        src45 <= {src45[14:0], in_data45};
        src46 <= {src46[14:0], in_data46};
        src47 <= {src47[14:0], in_data47};
        src48 <= {src48[14:0], in_data48};
        src49 <= {src49[14:0], in_data49};
        src50 <= {src50[14:0], in_data50};
        src51 <= {src51[14:0], in_data51};
        src52 <= {src52[14:0], in_data52};
        src53 <= {src53[14:0], in_data53};
        src54 <= {src54[14:0], in_data54};
        src55 <= {src55[14:0], in_data55};
        src56 <= {src56[14:0], in_data56};
        src57 <= {src57[14:0], in_data57};
        src58 <= {src58[14:0], in_data58};
        src59 <= {src59[14:0], in_data59};
        src60 <= {src60[14:0], in_data60};
        src61 <= {src61[14:0], in_data61};
        src62 <= {src62[14:0], in_data62};
        src63 <= {src63[14:0], in_data63};
        src64 <= {src64[14:0], in_data64};
        src65 <= {src65[14:0], in_data65};
        src66 <= {src66[14:0], in_data66};
        src67 <= {src67[14:0], in_data67};
        src68 <= {src68[14:0], in_data68};
        src69 <= {src69[14:0], in_data69};
        src70 <= {src70[14:0], in_data70};
        src71 <= {src71[14:0], in_data71};
        src72 <= {src72[14:0], in_data72};
        src73 <= {src73[14:0], in_data73};
        src74 <= {src74[14:0], in_data74};
        src75 <= {src75[14:0], in_data75};
        src76 <= {src76[14:0], in_data76};
        src77 <= {src77[14:0], in_data77};
        src78 <= {src78[14:0], in_data78};
        src79 <= {src79[14:0], in_data79};
        src80 <= {src80[14:0], in_data80};
        src81 <= {src81[14:0], in_data81};
        src82 <= {src82[14:0], in_data82};
        src83 <= {src83[14:0], in_data83};
        src84 <= {src84[14:0], in_data84};
        src85 <= {src85[14:0], in_data85};
        src86 <= {src86[14:0], in_data86};
        src87 <= {src87[14:0], in_data87};
        src88 <= {src88[14:0], in_data88};
        src89 <= {src89[14:0], in_data89};
        src90 <= {src90[14:0], in_data90};
        src91 <= {src91[14:0], in_data91};
        src92 <= {src92[14:0], in_data92};
        src93 <= {src93[14:0], in_data93};
        src94 <= {src94[14:0], in_data94};
        src95 <= {src95[14:0], in_data95};
        src96 <= {src96[14:0], in_data96};
        src97 <= {src97[14:0], in_data97};
        src98 <= {src98[14:0], in_data98};
        src99 <= {src99[14:0], in_data99};
        src100 <= {src100[14:0], in_data100};
        src101 <= {src101[14:0], in_data101};
        src102 <= {src102[14:0], in_data102};
        src103 <= {src103[14:0], in_data103};
        src104 <= {src104[14:0], in_data104};
        src105 <= {src105[14:0], in_data105};
        src106 <= {src106[14:0], in_data106};
        src107 <= {src107[14:0], in_data107};
        src108 <= {src108[14:0], in_data108};
        src109 <= {src109[14:0], in_data109};
        src110 <= {src110[14:0], in_data110};
        src111 <= {src111[14:0], in_data111};
        src112 <= {src112[14:0], in_data112};
        src113 <= {src113[14:0], in_data113};
        src114 <= {src114[14:0], in_data114};
        src115 <= {src115[14:0], in_data115};
        src116 <= {src116[14:0], in_data116};
        src117 <= {src117[14:0], in_data117};
        src118 <= {src118[14:0], in_data118};
        src119 <= {src119[14:0], in_data119};
        src120 <= {src120[14:0], in_data120};
        src121 <= {src121[14:0], in_data121};
        src122 <= {src122[14:0], in_data122};
        src123 <= {src123[14:0], in_data123};
        src124 <= {src124[14:0], in_data124};
        src125 <= {src125[14:0], in_data125};
        src126 <= {src126[14:0], in_data126};
        src127 <= {src127[14:0], in_data127};
    end
endmodule

module compressor2_1_128_16(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    input [15:0]src12,
    input [15:0]src13,
    input [15:0]src14,
    input [15:0]src15,
    input [15:0]src16,
    input [15:0]src17,
    input [15:0]src18,
    input [15:0]src19,
    input [15:0]src20,
    input [15:0]src21,
    input [15:0]src22,
    input [15:0]src23,
    input [15:0]src24,
    input [15:0]src25,
    input [15:0]src26,
    input [15:0]src27,
    input [15:0]src28,
    input [15:0]src29,
    input [15:0]src30,
    input [15:0]src31,
    input [15:0]src32,
    input [15:0]src33,
    input [15:0]src34,
    input [15:0]src35,
    input [15:0]src36,
    input [15:0]src37,
    input [15:0]src38,
    input [15:0]src39,
    input [15:0]src40,
    input [15:0]src41,
    input [15:0]src42,
    input [15:0]src43,
    input [15:0]src44,
    input [15:0]src45,
    input [15:0]src46,
    input [15:0]src47,
    input [15:0]src48,
    input [15:0]src49,
    input [15:0]src50,
    input [15:0]src51,
    input [15:0]src52,
    input [15:0]src53,
    input [15:0]src54,
    input [15:0]src55,
    input [15:0]src56,
    input [15:0]src57,
    input [15:0]src58,
    input [15:0]src59,
    input [15:0]src60,
    input [15:0]src61,
    input [15:0]src62,
    input [15:0]src63,
    input [15:0]src64,
    input [15:0]src65,
    input [15:0]src66,
    input [15:0]src67,
    input [15:0]src68,
    input [15:0]src69,
    input [15:0]src70,
    input [15:0]src71,
    input [15:0]src72,
    input [15:0]src73,
    input [15:0]src74,
    input [15:0]src75,
    input [15:0]src76,
    input [15:0]src77,
    input [15:0]src78,
    input [15:0]src79,
    input [15:0]src80,
    input [15:0]src81,
    input [15:0]src82,
    input [15:0]src83,
    input [15:0]src84,
    input [15:0]src85,
    input [15:0]src86,
    input [15:0]src87,
    input [15:0]src88,
    input [15:0]src89,
    input [15:0]src90,
    input [15:0]src91,
    input [15:0]src92,
    input [15:0]src93,
    input [15:0]src94,
    input [15:0]src95,
    input [15:0]src96,
    input [15:0]src97,
    input [15:0]src98,
    input [15:0]src99,
    input [15:0]src100,
    input [15:0]src101,
    input [15:0]src102,
    input [15:0]src103,
    input [15:0]src104,
    input [15:0]src105,
    input [15:0]src106,
    input [15:0]src107,
    input [15:0]src108,
    input [15:0]src109,
    input [15:0]src110,
    input [15:0]src111,
    input [15:0]src112,
    input [15:0]src113,
    input [15:0]src114,
    input [15:0]src115,
    input [15:0]src116,
    input [15:0]src117,
    input [15:0]src118,
    input [15:0]src119,
    input [15:0]src120,
    input [15:0]src121,
    input [15:0]src122,
    input [15:0]src123,
    input [15:0]src124,
    input [15:0]src125,
    input [15:0]src126,
    input [15:0]src127,
    output [22:0]dst);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [0:0] comp_out21;
    wire [0:0] comp_out22;
    wire [23:0] out;
    compressor compressor_inst(
        .src0({src127[0], src126[0], src125[0], src124[0], src123[0], src122[0], src121[0], src120[0], src119[0], src118[0], src117[0], src116[0], src115[0], src114[0], src113[0], src112[0], src111[0], src110[0], src109[0], src108[0], src107[0], src106[0], src105[0], src104[0], src103[0], src102[0], src101[0], src100[0], src99[0], src98[0], src97[0], src96[0], src95[0], src94[0], src93[0], src92[0], src91[0], src90[0], src89[0], src88[0], src87[0], src86[0], src85[0], src84[0], src83[0], src82[0], src81[0], src80[0], src79[0], src78[0], src77[0], src76[0], src75[0], src74[0], src73[0], src72[0], src71[0], src70[0], src69[0], src68[0], src67[0], src66[0], src65[0], src64[0], src63[0], src62[0], src61[0], src60[0], src59[0], src58[0], src57[0], src56[0], src55[0], src54[0], src53[0], src52[0], src51[0], src50[0], src49[0], src48[0], src47[0], src46[0], src45[0], src44[0], src43[0], src42[0], src41[0], src40[0], src39[0], src38[0], src37[0], src36[0], src35[0], src34[0], src33[0], src32[0], src31[0], src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}),
        .src1({src127[1], src126[1], src125[1], src124[1], src123[1], src122[1], src121[1], src120[1], src119[1], src118[1], src117[1], src116[1], src115[1], src114[1], src113[1], src112[1], src111[1], src110[1], src109[1], src108[1], src107[1], src106[1], src105[1], src104[1], src103[1], src102[1], src101[1], src100[1], src99[1], src98[1], src97[1], src96[1], src95[1], src94[1], src93[1], src92[1], src91[1], src90[1], src89[1], src88[1], src87[1], src86[1], src85[1], src84[1], src83[1], src82[1], src81[1], src80[1], src79[1], src78[1], src77[1], src76[1], src75[1], src74[1], src73[1], src72[1], src71[1], src70[1], src69[1], src68[1], src67[1], src66[1], src65[1], src64[1], src63[1], src62[1], src61[1], src60[1], src59[1], src58[1], src57[1], src56[1], src55[1], src54[1], src53[1], src52[1], src51[1], src50[1], src49[1], src48[1], src47[1], src46[1], src45[1], src44[1], src43[1], src42[1], src41[1], src40[1], src39[1], src38[1], src37[1], src36[1], src35[1], src34[1], src33[1], src32[1], src31[1], src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}),
        .src2({src127[2], src126[2], src125[2], src124[2], src123[2], src122[2], src121[2], src120[2], src119[2], src118[2], src117[2], src116[2], src115[2], src114[2], src113[2], src112[2], src111[2], src110[2], src109[2], src108[2], src107[2], src106[2], src105[2], src104[2], src103[2], src102[2], src101[2], src100[2], src99[2], src98[2], src97[2], src96[2], src95[2], src94[2], src93[2], src92[2], src91[2], src90[2], src89[2], src88[2], src87[2], src86[2], src85[2], src84[2], src83[2], src82[2], src81[2], src80[2], src79[2], src78[2], src77[2], src76[2], src75[2], src74[2], src73[2], src72[2], src71[2], src70[2], src69[2], src68[2], src67[2], src66[2], src65[2], src64[2], src63[2], src62[2], src61[2], src60[2], src59[2], src58[2], src57[2], src56[2], src55[2], src54[2], src53[2], src52[2], src51[2], src50[2], src49[2], src48[2], src47[2], src46[2], src45[2], src44[2], src43[2], src42[2], src41[2], src40[2], src39[2], src38[2], src37[2], src36[2], src35[2], src34[2], src33[2], src32[2], src31[2], src30[2], src29[2], src28[2], src27[2], src26[2], src25[2], src24[2], src23[2], src22[2], src21[2], src20[2], src19[2], src18[2], src17[2], src16[2], src15[2], src14[2], src13[2], src12[2], src11[2], src10[2], src9[2], src8[2], src7[2], src6[2], src5[2], src4[2], src3[2], src2[2], src1[2], src0[2]}),
        .src3({src127[3], src126[3], src125[3], src124[3], src123[3], src122[3], src121[3], src120[3], src119[3], src118[3], src117[3], src116[3], src115[3], src114[3], src113[3], src112[3], src111[3], src110[3], src109[3], src108[3], src107[3], src106[3], src105[3], src104[3], src103[3], src102[3], src101[3], src100[3], src99[3], src98[3], src97[3], src96[3], src95[3], src94[3], src93[3], src92[3], src91[3], src90[3], src89[3], src88[3], src87[3], src86[3], src85[3], src84[3], src83[3], src82[3], src81[3], src80[3], src79[3], src78[3], src77[3], src76[3], src75[3], src74[3], src73[3], src72[3], src71[3], src70[3], src69[3], src68[3], src67[3], src66[3], src65[3], src64[3], src63[3], src62[3], src61[3], src60[3], src59[3], src58[3], src57[3], src56[3], src55[3], src54[3], src53[3], src52[3], src51[3], src50[3], src49[3], src48[3], src47[3], src46[3], src45[3], src44[3], src43[3], src42[3], src41[3], src40[3], src39[3], src38[3], src37[3], src36[3], src35[3], src34[3], src33[3], src32[3], src31[3], src30[3], src29[3], src28[3], src27[3], src26[3], src25[3], src24[3], src23[3], src22[3], src21[3], src20[3], src19[3], src18[3], src17[3], src16[3], src15[3], src14[3], src13[3], src12[3], src11[3], src10[3], src9[3], src8[3], src7[3], src6[3], src5[3], src4[3], src3[3], src2[3], src1[3], src0[3]}),
        .src4({src127[4], src126[4], src125[4], src124[4], src123[4], src122[4], src121[4], src120[4], src119[4], src118[4], src117[4], src116[4], src115[4], src114[4], src113[4], src112[4], src111[4], src110[4], src109[4], src108[4], src107[4], src106[4], src105[4], src104[4], src103[4], src102[4], src101[4], src100[4], src99[4], src98[4], src97[4], src96[4], src95[4], src94[4], src93[4], src92[4], src91[4], src90[4], src89[4], src88[4], src87[4], src86[4], src85[4], src84[4], src83[4], src82[4], src81[4], src80[4], src79[4], src78[4], src77[4], src76[4], src75[4], src74[4], src73[4], src72[4], src71[4], src70[4], src69[4], src68[4], src67[4], src66[4], src65[4], src64[4], src63[4], src62[4], src61[4], src60[4], src59[4], src58[4], src57[4], src56[4], src55[4], src54[4], src53[4], src52[4], src51[4], src50[4], src49[4], src48[4], src47[4], src46[4], src45[4], src44[4], src43[4], src42[4], src41[4], src40[4], src39[4], src38[4], src37[4], src36[4], src35[4], src34[4], src33[4], src32[4], src31[4], src30[4], src29[4], src28[4], src27[4], src26[4], src25[4], src24[4], src23[4], src22[4], src21[4], src20[4], src19[4], src18[4], src17[4], src16[4], src15[4], src14[4], src13[4], src12[4], src11[4], src10[4], src9[4], src8[4], src7[4], src6[4], src5[4], src4[4], src3[4], src2[4], src1[4], src0[4]}),
        .src5({src127[5], src126[5], src125[5], src124[5], src123[5], src122[5], src121[5], src120[5], src119[5], src118[5], src117[5], src116[5], src115[5], src114[5], src113[5], src112[5], src111[5], src110[5], src109[5], src108[5], src107[5], src106[5], src105[5], src104[5], src103[5], src102[5], src101[5], src100[5], src99[5], src98[5], src97[5], src96[5], src95[5], src94[5], src93[5], src92[5], src91[5], src90[5], src89[5], src88[5], src87[5], src86[5], src85[5], src84[5], src83[5], src82[5], src81[5], src80[5], src79[5], src78[5], src77[5], src76[5], src75[5], src74[5], src73[5], src72[5], src71[5], src70[5], src69[5], src68[5], src67[5], src66[5], src65[5], src64[5], src63[5], src62[5], src61[5], src60[5], src59[5], src58[5], src57[5], src56[5], src55[5], src54[5], src53[5], src52[5], src51[5], src50[5], src49[5], src48[5], src47[5], src46[5], src45[5], src44[5], src43[5], src42[5], src41[5], src40[5], src39[5], src38[5], src37[5], src36[5], src35[5], src34[5], src33[5], src32[5], src31[5], src30[5], src29[5], src28[5], src27[5], src26[5], src25[5], src24[5], src23[5], src22[5], src21[5], src20[5], src19[5], src18[5], src17[5], src16[5], src15[5], src14[5], src13[5], src12[5], src11[5], src10[5], src9[5], src8[5], src7[5], src6[5], src5[5], src4[5], src3[5], src2[5], src1[5], src0[5]}),
        .src6({src127[6], src126[6], src125[6], src124[6], src123[6], src122[6], src121[6], src120[6], src119[6], src118[6], src117[6], src116[6], src115[6], src114[6], src113[6], src112[6], src111[6], src110[6], src109[6], src108[6], src107[6], src106[6], src105[6], src104[6], src103[6], src102[6], src101[6], src100[6], src99[6], src98[6], src97[6], src96[6], src95[6], src94[6], src93[6], src92[6], src91[6], src90[6], src89[6], src88[6], src87[6], src86[6], src85[6], src84[6], src83[6], src82[6], src81[6], src80[6], src79[6], src78[6], src77[6], src76[6], src75[6], src74[6], src73[6], src72[6], src71[6], src70[6], src69[6], src68[6], src67[6], src66[6], src65[6], src64[6], src63[6], src62[6], src61[6], src60[6], src59[6], src58[6], src57[6], src56[6], src55[6], src54[6], src53[6], src52[6], src51[6], src50[6], src49[6], src48[6], src47[6], src46[6], src45[6], src44[6], src43[6], src42[6], src41[6], src40[6], src39[6], src38[6], src37[6], src36[6], src35[6], src34[6], src33[6], src32[6], src31[6], src30[6], src29[6], src28[6], src27[6], src26[6], src25[6], src24[6], src23[6], src22[6], src21[6], src20[6], src19[6], src18[6], src17[6], src16[6], src15[6], src14[6], src13[6], src12[6], src11[6], src10[6], src9[6], src8[6], src7[6], src6[6], src5[6], src4[6], src3[6], src2[6], src1[6], src0[6]}),
        .src7({src127[7], src126[7], src125[7], src124[7], src123[7], src122[7], src121[7], src120[7], src119[7], src118[7], src117[7], src116[7], src115[7], src114[7], src113[7], src112[7], src111[7], src110[7], src109[7], src108[7], src107[7], src106[7], src105[7], src104[7], src103[7], src102[7], src101[7], src100[7], src99[7], src98[7], src97[7], src96[7], src95[7], src94[7], src93[7], src92[7], src91[7], src90[7], src89[7], src88[7], src87[7], src86[7], src85[7], src84[7], src83[7], src82[7], src81[7], src80[7], src79[7], src78[7], src77[7], src76[7], src75[7], src74[7], src73[7], src72[7], src71[7], src70[7], src69[7], src68[7], src67[7], src66[7], src65[7], src64[7], src63[7], src62[7], src61[7], src60[7], src59[7], src58[7], src57[7], src56[7], src55[7], src54[7], src53[7], src52[7], src51[7], src50[7], src49[7], src48[7], src47[7], src46[7], src45[7], src44[7], src43[7], src42[7], src41[7], src40[7], src39[7], src38[7], src37[7], src36[7], src35[7], src34[7], src33[7], src32[7], src31[7], src30[7], src29[7], src28[7], src27[7], src26[7], src25[7], src24[7], src23[7], src22[7], src21[7], src20[7], src19[7], src18[7], src17[7], src16[7], src15[7], src14[7], src13[7], src12[7], src11[7], src10[7], src9[7], src8[7], src7[7], src6[7], src5[7], src4[7], src3[7], src2[7], src1[7], src0[7]}),
        .src8({src127[8], src126[8], src125[8], src124[8], src123[8], src122[8], src121[8], src120[8], src119[8], src118[8], src117[8], src116[8], src115[8], src114[8], src113[8], src112[8], src111[8], src110[8], src109[8], src108[8], src107[8], src106[8], src105[8], src104[8], src103[8], src102[8], src101[8], src100[8], src99[8], src98[8], src97[8], src96[8], src95[8], src94[8], src93[8], src92[8], src91[8], src90[8], src89[8], src88[8], src87[8], src86[8], src85[8], src84[8], src83[8], src82[8], src81[8], src80[8], src79[8], src78[8], src77[8], src76[8], src75[8], src74[8], src73[8], src72[8], src71[8], src70[8], src69[8], src68[8], src67[8], src66[8], src65[8], src64[8], src63[8], src62[8], src61[8], src60[8], src59[8], src58[8], src57[8], src56[8], src55[8], src54[8], src53[8], src52[8], src51[8], src50[8], src49[8], src48[8], src47[8], src46[8], src45[8], src44[8], src43[8], src42[8], src41[8], src40[8], src39[8], src38[8], src37[8], src36[8], src35[8], src34[8], src33[8], src32[8], src31[8], src30[8], src29[8], src28[8], src27[8], src26[8], src25[8], src24[8], src23[8], src22[8], src21[8], src20[8], src19[8], src18[8], src17[8], src16[8], src15[8], src14[8], src13[8], src12[8], src11[8], src10[8], src9[8], src8[8], src7[8], src6[8], src5[8], src4[8], src3[8], src2[8], src1[8], src0[8]}),
        .src9({src127[9], src126[9], src125[9], src124[9], src123[9], src122[9], src121[9], src120[9], src119[9], src118[9], src117[9], src116[9], src115[9], src114[9], src113[9], src112[9], src111[9], src110[9], src109[9], src108[9], src107[9], src106[9], src105[9], src104[9], src103[9], src102[9], src101[9], src100[9], src99[9], src98[9], src97[9], src96[9], src95[9], src94[9], src93[9], src92[9], src91[9], src90[9], src89[9], src88[9], src87[9], src86[9], src85[9], src84[9], src83[9], src82[9], src81[9], src80[9], src79[9], src78[9], src77[9], src76[9], src75[9], src74[9], src73[9], src72[9], src71[9], src70[9], src69[9], src68[9], src67[9], src66[9], src65[9], src64[9], src63[9], src62[9], src61[9], src60[9], src59[9], src58[9], src57[9], src56[9], src55[9], src54[9], src53[9], src52[9], src51[9], src50[9], src49[9], src48[9], src47[9], src46[9], src45[9], src44[9], src43[9], src42[9], src41[9], src40[9], src39[9], src38[9], src37[9], src36[9], src35[9], src34[9], src33[9], src32[9], src31[9], src30[9], src29[9], src28[9], src27[9], src26[9], src25[9], src24[9], src23[9], src22[9], src21[9], src20[9], src19[9], src18[9], src17[9], src16[9], src15[9], src14[9], src13[9], src12[9], src11[9], src10[9], src9[9], src8[9], src7[9], src6[9], src5[9], src4[9], src3[9], src2[9], src1[9], src0[9]}),
        .src10({src127[10], src126[10], src125[10], src124[10], src123[10], src122[10], src121[10], src120[10], src119[10], src118[10], src117[10], src116[10], src115[10], src114[10], src113[10], src112[10], src111[10], src110[10], src109[10], src108[10], src107[10], src106[10], src105[10], src104[10], src103[10], src102[10], src101[10], src100[10], src99[10], src98[10], src97[10], src96[10], src95[10], src94[10], src93[10], src92[10], src91[10], src90[10], src89[10], src88[10], src87[10], src86[10], src85[10], src84[10], src83[10], src82[10], src81[10], src80[10], src79[10], src78[10], src77[10], src76[10], src75[10], src74[10], src73[10], src72[10], src71[10], src70[10], src69[10], src68[10], src67[10], src66[10], src65[10], src64[10], src63[10], src62[10], src61[10], src60[10], src59[10], src58[10], src57[10], src56[10], src55[10], src54[10], src53[10], src52[10], src51[10], src50[10], src49[10], src48[10], src47[10], src46[10], src45[10], src44[10], src43[10], src42[10], src41[10], src40[10], src39[10], src38[10], src37[10], src36[10], src35[10], src34[10], src33[10], src32[10], src31[10], src30[10], src29[10], src28[10], src27[10], src26[10], src25[10], src24[10], src23[10], src22[10], src21[10], src20[10], src19[10], src18[10], src17[10], src16[10], src15[10], src14[10], src13[10], src12[10], src11[10], src10[10], src9[10], src8[10], src7[10], src6[10], src5[10], src4[10], src3[10], src2[10], src1[10], src0[10]}),
        .src11({src127[11], src126[11], src125[11], src124[11], src123[11], src122[11], src121[11], src120[11], src119[11], src118[11], src117[11], src116[11], src115[11], src114[11], src113[11], src112[11], src111[11], src110[11], src109[11], src108[11], src107[11], src106[11], src105[11], src104[11], src103[11], src102[11], src101[11], src100[11], src99[11], src98[11], src97[11], src96[11], src95[11], src94[11], src93[11], src92[11], src91[11], src90[11], src89[11], src88[11], src87[11], src86[11], src85[11], src84[11], src83[11], src82[11], src81[11], src80[11], src79[11], src78[11], src77[11], src76[11], src75[11], src74[11], src73[11], src72[11], src71[11], src70[11], src69[11], src68[11], src67[11], src66[11], src65[11], src64[11], src63[11], src62[11], src61[11], src60[11], src59[11], src58[11], src57[11], src56[11], src55[11], src54[11], src53[11], src52[11], src51[11], src50[11], src49[11], src48[11], src47[11], src46[11], src45[11], src44[11], src43[11], src42[11], src41[11], src40[11], src39[11], src38[11], src37[11], src36[11], src35[11], src34[11], src33[11], src32[11], src31[11], src30[11], src29[11], src28[11], src27[11], src26[11], src25[11], src24[11], src23[11], src22[11], src21[11], src20[11], src19[11], src18[11], src17[11], src16[11], src15[11], src14[11], src13[11], src12[11], src11[11], src10[11], src9[11], src8[11], src7[11], src6[11], src5[11], src4[11], src3[11], src2[11], src1[11], src0[11]}),
        .src12({src127[12], src126[12], src125[12], src124[12], src123[12], src122[12], src121[12], src120[12], src119[12], src118[12], src117[12], src116[12], src115[12], src114[12], src113[12], src112[12], src111[12], src110[12], src109[12], src108[12], src107[12], src106[12], src105[12], src104[12], src103[12], src102[12], src101[12], src100[12], src99[12], src98[12], src97[12], src96[12], src95[12], src94[12], src93[12], src92[12], src91[12], src90[12], src89[12], src88[12], src87[12], src86[12], src85[12], src84[12], src83[12], src82[12], src81[12], src80[12], src79[12], src78[12], src77[12], src76[12], src75[12], src74[12], src73[12], src72[12], src71[12], src70[12], src69[12], src68[12], src67[12], src66[12], src65[12], src64[12], src63[12], src62[12], src61[12], src60[12], src59[12], src58[12], src57[12], src56[12], src55[12], src54[12], src53[12], src52[12], src51[12], src50[12], src49[12], src48[12], src47[12], src46[12], src45[12], src44[12], src43[12], src42[12], src41[12], src40[12], src39[12], src38[12], src37[12], src36[12], src35[12], src34[12], src33[12], src32[12], src31[12], src30[12], src29[12], src28[12], src27[12], src26[12], src25[12], src24[12], src23[12], src22[12], src21[12], src20[12], src19[12], src18[12], src17[12], src16[12], src15[12], src14[12], src13[12], src12[12], src11[12], src10[12], src9[12], src8[12], src7[12], src6[12], src5[12], src4[12], src3[12], src2[12], src1[12], src0[12]}),
        .src13({src127[13], src126[13], src125[13], src124[13], src123[13], src122[13], src121[13], src120[13], src119[13], src118[13], src117[13], src116[13], src115[13], src114[13], src113[13], src112[13], src111[13], src110[13], src109[13], src108[13], src107[13], src106[13], src105[13], src104[13], src103[13], src102[13], src101[13], src100[13], src99[13], src98[13], src97[13], src96[13], src95[13], src94[13], src93[13], src92[13], src91[13], src90[13], src89[13], src88[13], src87[13], src86[13], src85[13], src84[13], src83[13], src82[13], src81[13], src80[13], src79[13], src78[13], src77[13], src76[13], src75[13], src74[13], src73[13], src72[13], src71[13], src70[13], src69[13], src68[13], src67[13], src66[13], src65[13], src64[13], src63[13], src62[13], src61[13], src60[13], src59[13], src58[13], src57[13], src56[13], src55[13], src54[13], src53[13], src52[13], src51[13], src50[13], src49[13], src48[13], src47[13], src46[13], src45[13], src44[13], src43[13], src42[13], src41[13], src40[13], src39[13], src38[13], src37[13], src36[13], src35[13], src34[13], src33[13], src32[13], src31[13], src30[13], src29[13], src28[13], src27[13], src26[13], src25[13], src24[13], src23[13], src22[13], src21[13], src20[13], src19[13], src18[13], src17[13], src16[13], src15[13], src14[13], src13[13], src12[13], src11[13], src10[13], src9[13], src8[13], src7[13], src6[13], src5[13], src4[13], src3[13], src2[13], src1[13], src0[13]}),
        .src14({src127[14], src126[14], src125[14], src124[14], src123[14], src122[14], src121[14], src120[14], src119[14], src118[14], src117[14], src116[14], src115[14], src114[14], src113[14], src112[14], src111[14], src110[14], src109[14], src108[14], src107[14], src106[14], src105[14], src104[14], src103[14], src102[14], src101[14], src100[14], src99[14], src98[14], src97[14], src96[14], src95[14], src94[14], src93[14], src92[14], src91[14], src90[14], src89[14], src88[14], src87[14], src86[14], src85[14], src84[14], src83[14], src82[14], src81[14], src80[14], src79[14], src78[14], src77[14], src76[14], src75[14], src74[14], src73[14], src72[14], src71[14], src70[14], src69[14], src68[14], src67[14], src66[14], src65[14], src64[14], src63[14], src62[14], src61[14], src60[14], src59[14], src58[14], src57[14], src56[14], src55[14], src54[14], src53[14], src52[14], src51[14], src50[14], src49[14], src48[14], src47[14], src46[14], src45[14], src44[14], src43[14], src42[14], src41[14], src40[14], src39[14], src38[14], src37[14], src36[14], src35[14], src34[14], src33[14], src32[14], src31[14], src30[14], src29[14], src28[14], src27[14], src26[14], src25[14], src24[14], src23[14], src22[14], src21[14], src20[14], src19[14], src18[14], src17[14], src16[14], src15[14], src14[14], src13[14], src12[14], src11[14], src10[14], src9[14], src8[14], src7[14], src6[14], src5[14], src4[14], src3[14], src2[14], src1[14], src0[14]}),
        .src15({src127[15], src126[15], src125[15], src124[15], src123[15], src122[15], src121[15], src120[15], src119[15], src118[15], src117[15], src116[15], src115[15], src114[15], src113[15], src112[15], src111[15], src110[15], src109[15], src108[15], src107[15], src106[15], src105[15], src104[15], src103[15], src102[15], src101[15], src100[15], src99[15], src98[15], src97[15], src96[15], src95[15], src94[15], src93[15], src92[15], src91[15], src90[15], src89[15], src88[15], src87[15], src86[15], src85[15], src84[15], src83[15], src82[15], src81[15], src80[15], src79[15], src78[15], src77[15], src76[15], src75[15], src74[15], src73[15], src72[15], src71[15], src70[15], src69[15], src68[15], src67[15], src66[15], src65[15], src64[15], src63[15], src62[15], src61[15], src60[15], src59[15], src58[15], src57[15], src56[15], src55[15], src54[15], src53[15], src52[15], src51[15], src50[15], src49[15], src48[15], src47[15], src46[15], src45[15], src44[15], src43[15], src42[15], src41[15], src40[15], src39[15], src38[15], src37[15], src36[15], src35[15], src34[15], src33[15], src32[15], src31[15], src30[15], src29[15], src28[15], src27[15], src26[15], src25[15], src24[15], src23[15], src22[15], src21[15], src20[15], src19[15], src18[15], src17[15], src16[15], src15[15], src14[15], src13[15], src12[15], src11[15], src10[15], src9[15], src8[15], src7[15], src6[15], src5[15], src4[15], src3[15], src2[15], src1[15], src0[15]}),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22)
    );
    rowadder2_1_23 rowadder2_1inst(
        .src0({comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0(out)
    );
    assign dst = out[22:0];
endmodule
module compressor (
      input wire [127:0] src0,
      input wire [127:0] src1,
      input wire [127:0] src2,
      input wire [127:0] src3,
      input wire [127:0] src4,
      input wire [127:0] src5,
      input wire [127:0] src6,
      input wire [127:0] src7,
      input wire [127:0] src8,
      input wire [127:0] src9,
      input wire [127:0] src10,
      input wire [127:0] src11,
      input wire [127:0] src12,
      input wire [127:0] src13,
      input wire [127:0] src14,
      input wire [127:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [0:0] dst21,
      output wire [0:0] dst22);

   wire [127:0] stage0_0;
   wire [127:0] stage0_1;
   wire [127:0] stage0_2;
   wire [127:0] stage0_3;
   wire [127:0] stage0_4;
   wire [127:0] stage0_5;
   wire [127:0] stage0_6;
   wire [127:0] stage0_7;
   wire [127:0] stage0_8;
   wire [127:0] stage0_9;
   wire [127:0] stage0_10;
   wire [127:0] stage0_11;
   wire [127:0] stage0_12;
   wire [127:0] stage0_13;
   wire [127:0] stage0_14;
   wire [127:0] stage0_15;
   wire [45:0] stage1_0;
   wire [63:0] stage1_1;
   wire [38:0] stage1_2;
   wire [48:0] stage1_3;
   wire [59:0] stage1_4;
   wire [56:0] stage1_5;
   wire [47:0] stage1_6;
   wire [64:0] stage1_7;
   wire [55:0] stage1_8;
   wire [57:0] stage1_9;
   wire [53:0] stage1_10;
   wire [51:0] stage1_11;
   wire [56:0] stage1_12;
   wire [71:0] stage1_13;
   wire [70:0] stage1_14;
   wire [37:0] stage1_15;
   wire [35:0] stage1_16;
   wire [20:0] stage1_17;
   wire [14:0] stage2_0;
   wire [13:0] stage2_1;
   wire [19:0] stage2_2;
   wire [19:0] stage2_3;
   wire [27:0] stage2_4;
   wire [27:0] stage2_5;
   wire [16:0] stage2_6;
   wire [30:0] stage2_7;
   wire [28:0] stage2_8;
   wire [20:0] stage2_9;
   wire [17:0] stage2_10;
   wire [37:0] stage2_11;
   wire [28:0] stage2_12;
   wire [18:0] stage2_13;
   wire [34:0] stage2_14;
   wire [26:0] stage2_15;
   wire [19:0] stage2_16;
   wire [19:0] stage2_17;
   wire [6:0] stage2_18;
   wire [1:0] stage2_19;
   wire [14:0] stage3_0;
   wire [8:0] stage3_1;
   wire [12:0] stage3_2;
   wire [10:0] stage3_3;
   wire [8:0] stage3_4;
   wire [9:0] stage3_5;
   wire [10:0] stage3_6;
   wire [8:0] stage3_7;
   wire [13:0] stage3_8;
   wire [12:0] stage3_9;
   wire [7:0] stage3_10;
   wire [16:0] stage3_11;
   wire [13:0] stage3_12;
   wire [11:0] stage3_13;
   wire [15:0] stage3_14;
   wire [10:0] stage3_15;
   wire [19:0] stage3_16;
   wire [6:0] stage3_17;
   wire [5:0] stage3_18;
   wire [5:0] stage3_19;
   wire [0:0] stage3_20;
   wire [5:0] stage4_0;
   wire [9:0] stage4_1;
   wire [2:0] stage4_2;
   wire [10:0] stage4_3;
   wire [5:0] stage4_4;
   wire [4:0] stage4_5;
   wire [3:0] stage4_6;
   wire [4:0] stage4_7;
   wire [4:0] stage4_8;
   wire [6:0] stage4_9;
   wire [5:0] stage4_10;
   wire [3:0] stage4_11;
   wire [5:0] stage4_12;
   wire [5:0] stage4_13;
   wire [5:0] stage4_14;
   wire [7:0] stage4_15;
   wire [6:0] stage4_16;
   wire [5:0] stage4_17;
   wire [3:0] stage4_18;
   wire [1:0] stage4_19;
   wire [2:0] stage4_20;
   wire [0:0] stage4_21;
   wire [1:0] stage5_0;
   wire [3:0] stage5_1;
   wire [2:0] stage5_2;
   wire [6:0] stage5_3;
   wire [2:0] stage5_4;
   wire [5:0] stage5_5;
   wire [0:0] stage5_6;
   wire [4:0] stage5_7;
   wire [1:0] stage5_8;
   wire [6:0] stage5_9;
   wire [0:0] stage5_10;
   wire [4:0] stage5_11;
   wire [1:0] stage5_12;
   wire [6:0] stage5_13;
   wire [0:0] stage5_14;
   wire [4:0] stage5_15;
   wire [5:0] stage5_16;
   wire [5:0] stage5_17;
   wire [2:0] stage5_18;
   wire [0:0] stage5_19;
   wire [0:0] stage5_20;
   wire [0:0] stage5_21;
   wire [0:0] stage5_22;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [0:0] stage6_21;
   wire [0:0] stage6_22;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6]},
      {stage1_5[0],stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17]}
   );
   gpc606_5 gpc18 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[1],stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18]}
   );
   gpc606_5 gpc19 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18]},
      {stage1_5[2],stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19]}
   );
   gpc606_5 gpc20 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24]},
      {stage1_5[3],stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20]}
   );
   gpc606_5 gpc21 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30]},
      {stage1_5[4],stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21]}
   );
   gpc606_5 gpc22 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36]},
      {stage1_5[5],stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22]}
   );
   gpc606_5 gpc23 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42]},
      {stage1_5[6],stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23]}
   );
   gpc606_5 gpc24 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48]},
      {stage1_5[7],stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24]}
   );
   gpc606_5 gpc25 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage1_5[8],stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25]}
   );
   gpc606_5 gpc26 (
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60]},
      {stage1_5[9],stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26]}
   );
   gpc606_5 gpc27 (
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66]},
      {stage1_5[10],stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72]},
      {stage1_5[11],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78]},
      {stage1_5[12],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84]},
      {stage1_5[13],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90]},
      {stage1_5[14],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[15],stage1_4[32],stage1_3[32],stage1_2[32]}
   );
   gpc606_5 gpc33 (
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[16],stage1_4[33],stage1_3[33],stage1_2[33]}
   );
   gpc606_5 gpc34 (
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[17],stage1_4[34],stage1_3[34],stage1_2[34]}
   );
   gpc606_5 gpc35 (
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[18],stage1_4[35],stage1_3[35],stage1_2[35]}
   );
   gpc615_5 gpc36 (
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125]},
      {stage0_3[91]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[19],stage1_4[36],stage1_3[36],stage1_2[36]}
   );
   gpc615_5 gpc37 (
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage0_4[30]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[5],stage1_5[20],stage1_4[37],stage1_3[37]}
   );
   gpc615_5 gpc38 (
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101]},
      {stage0_4[31]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[6],stage1_5[21],stage1_4[38],stage1_3[38]}
   );
   gpc615_5 gpc39 (
      {stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage0_4[32]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[7],stage1_5[22],stage1_4[39],stage1_3[39]}
   );
   gpc615_5 gpc40 (
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage0_4[33]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[8],stage1_5[23],stage1_4[40],stage1_3[40]}
   );
   gpc615_5 gpc41 (
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage0_4[34]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[9],stage1_5[24],stage1_4[41],stage1_3[41]}
   );
   gpc615_5 gpc42 (
      {stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121]},
      {stage0_4[35]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[10],stage1_5[25],stage1_4[42],stage1_3[42]}
   );
   gpc606_5 gpc43 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[6],stage1_6[11],stage1_5[26],stage1_4[43]}
   );
   gpc606_5 gpc44 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[7],stage1_6[12],stage1_5[27],stage1_4[44]}
   );
   gpc606_5 gpc45 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[8],stage1_6[13],stage1_5[28],stage1_4[45]}
   );
   gpc606_5 gpc46 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[9],stage1_6[14],stage1_5[29],stage1_4[46]}
   );
   gpc606_5 gpc47 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[10],stage1_6[15],stage1_5[30],stage1_4[47]}
   );
   gpc606_5 gpc48 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[11],stage1_6[16],stage1_5[31],stage1_4[48]}
   );
   gpc606_5 gpc49 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[12],stage1_6[17],stage1_5[32],stage1_4[49]}
   );
   gpc606_5 gpc50 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[13],stage1_6[18],stage1_5[33],stage1_4[50]}
   );
   gpc606_5 gpc51 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[14],stage1_6[19],stage1_5[34],stage1_4[51]}
   );
   gpc606_5 gpc52 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[15],stage1_6[20],stage1_5[35],stage1_4[52]}
   );
   gpc606_5 gpc53 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[16],stage1_6[21],stage1_5[36],stage1_4[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[17],stage1_6[22],stage1_5[37],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[18],stage1_6[23],stage1_5[38],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[19],stage1_6[24],stage1_5[39],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[20],stage1_6[25],stage1_5[40],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[15],stage1_7[21],stage1_6[26],stage1_5[41]}
   );
   gpc606_5 gpc59 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[16],stage1_7[22],stage1_6[27],stage1_5[42]}
   );
   gpc606_5 gpc60 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[17],stage1_7[23],stage1_6[28],stage1_5[43]}
   );
   gpc606_5 gpc61 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[18],stage1_7[24],stage1_6[29],stage1_5[44]}
   );
   gpc606_5 gpc62 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[19],stage1_7[25],stage1_6[30],stage1_5[45]}
   );
   gpc606_5 gpc63 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[20],stage1_7[26],stage1_6[31],stage1_5[46]}
   );
   gpc606_5 gpc64 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[21],stage1_7[27],stage1_6[32],stage1_5[47]}
   );
   gpc606_5 gpc65 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[22],stage1_7[28],stage1_6[33],stage1_5[48]}
   );
   gpc606_5 gpc66 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[23],stage1_7[29],stage1_6[34],stage1_5[49]}
   );
   gpc606_5 gpc67 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[24],stage1_7[30],stage1_6[35],stage1_5[50]}
   );
   gpc606_5 gpc68 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[25],stage1_7[31],stage1_6[36],stage1_5[51]}
   );
   gpc606_5 gpc69 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[26],stage1_7[32],stage1_6[37],stage1_5[52]}
   );
   gpc615_5 gpc70 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112]},
      {stage0_6[90]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[27],stage1_7[33],stage1_6[38],stage1_5[53]}
   );
   gpc615_5 gpc71 (
      {stage0_5[113], stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117]},
      {stage0_6[91]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[28],stage1_7[34],stage1_6[39],stage1_5[54]}
   );
   gpc615_5 gpc72 (
      {stage0_5[118], stage0_5[119], stage0_5[120], stage0_5[121], stage0_5[122]},
      {stage0_6[92]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[29],stage1_7[35],stage1_6[40],stage1_5[55]}
   );
   gpc615_5 gpc73 (
      {stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126], stage0_5[127]},
      {stage0_6[93]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[30],stage1_7[36],stage1_6[41],stage1_5[56]}
   );
   gpc606_5 gpc74 (
      {stage0_6[94], stage0_6[95], stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[16],stage1_8[31],stage1_7[37],stage1_6[42]}
   );
   gpc606_5 gpc75 (
      {stage0_6[100], stage0_6[101], stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[17],stage1_8[32],stage1_7[38],stage1_6[43]}
   );
   gpc606_5 gpc76 (
      {stage0_6[106], stage0_6[107], stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[18],stage1_8[33],stage1_7[39],stage1_6[44]}
   );
   gpc606_5 gpc77 (
      {stage0_6[112], stage0_6[113], stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[19],stage1_8[34],stage1_7[40],stage1_6[45]}
   );
   gpc615_5 gpc78 (
      {stage0_6[118], stage0_6[119], stage0_6[120], stage0_6[121], stage0_6[122]},
      {stage0_7[96]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[20],stage1_8[35],stage1_7[41],stage1_6[46]}
   );
   gpc615_5 gpc79 (
      {stage0_6[123], stage0_6[124], stage0_6[125], stage0_6[126], stage0_6[127]},
      {stage0_7[97]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[21],stage1_8[36],stage1_7[42],stage1_6[47]}
   );
   gpc615_5 gpc80 (
      {stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101], stage0_7[102]},
      {stage0_8[36]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[6],stage1_9[22],stage1_8[37],stage1_7[43]}
   );
   gpc615_5 gpc81 (
      {stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage0_8[37]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[7],stage1_9[23],stage1_8[38],stage1_7[44]}
   );
   gpc606_5 gpc82 (
      {stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[2],stage1_10[8],stage1_9[24],stage1_8[39]}
   );
   gpc606_5 gpc83 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48], stage0_8[49]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[3],stage1_10[9],stage1_9[25],stage1_8[40]}
   );
   gpc606_5 gpc84 (
      {stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53], stage0_8[54], stage0_8[55]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[4],stage1_10[10],stage1_9[26],stage1_8[41]}
   );
   gpc606_5 gpc85 (
      {stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[5],stage1_10[11],stage1_9[27],stage1_8[42]}
   );
   gpc606_5 gpc86 (
      {stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66], stage0_8[67]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[6],stage1_10[12],stage1_9[28],stage1_8[43]}
   );
   gpc606_5 gpc87 (
      {stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72], stage0_8[73]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[7],stage1_10[13],stage1_9[29],stage1_8[44]}
   );
   gpc606_5 gpc88 (
      {stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77], stage0_8[78], stage0_8[79]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[8],stage1_10[14],stage1_9[30],stage1_8[45]}
   );
   gpc606_5 gpc89 (
      {stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83], stage0_8[84], stage0_8[85]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[9],stage1_10[15],stage1_9[31],stage1_8[46]}
   );
   gpc606_5 gpc90 (
      {stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[10],stage1_10[16],stage1_9[32],stage1_8[47]}
   );
   gpc606_5 gpc91 (
      {stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[11],stage1_10[17],stage1_9[33],stage1_8[48]}
   );
   gpc606_5 gpc92 (
      {stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[12],stage1_10[18],stage1_9[34],stage1_8[49]}
   );
   gpc606_5 gpc93 (
      {stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[13],stage1_10[19],stage1_9[35],stage1_8[50]}
   );
   gpc606_5 gpc94 (
      {stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[14],stage1_10[20],stage1_9[36],stage1_8[51]}
   );
   gpc615_5 gpc95 (
      {stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120]},
      {stage0_9[12]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[15],stage1_10[21],stage1_9[37],stage1_8[52]}
   );
   gpc615_5 gpc96 (
      {stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_9[13]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[16],stage1_10[22],stage1_9[38],stage1_8[53]}
   );
   gpc606_5 gpc97 (
      {stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[15],stage1_11[17],stage1_10[23],stage1_9[39]}
   );
   gpc606_5 gpc98 (
      {stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[16],stage1_11[18],stage1_10[24],stage1_9[40]}
   );
   gpc606_5 gpc99 (
      {stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[17],stage1_11[19],stage1_10[25],stage1_9[41]}
   );
   gpc606_5 gpc100 (
      {stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[18],stage1_11[20],stage1_10[26],stage1_9[42]}
   );
   gpc606_5 gpc101 (
      {stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[19],stage1_11[21],stage1_10[27],stage1_9[43]}
   );
   gpc606_5 gpc102 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[20],stage1_11[22],stage1_10[28],stage1_9[44]}
   );
   gpc606_5 gpc103 (
      {stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[21],stage1_11[23],stage1_10[29],stage1_9[45]}
   );
   gpc606_5 gpc104 (
      {stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[22],stage1_11[24],stage1_10[30],stage1_9[46]}
   );
   gpc606_5 gpc105 (
      {stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[23],stage1_11[25],stage1_10[31],stage1_9[47]}
   );
   gpc606_5 gpc106 (
      {stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[24],stage1_11[26],stage1_10[32],stage1_9[48]}
   );
   gpc606_5 gpc107 (
      {stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[25],stage1_11[27],stage1_10[33],stage1_9[49]}
   );
   gpc606_5 gpc108 (
      {stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[26],stage1_11[28],stage1_10[34],stage1_9[50]}
   );
   gpc606_5 gpc109 (
      {stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[27],stage1_11[29],stage1_10[35],stage1_9[51]}
   );
   gpc606_5 gpc110 (
      {stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[28],stage1_11[30],stage1_10[36],stage1_9[52]}
   );
   gpc606_5 gpc111 (
      {stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[29],stage1_11[31],stage1_10[37],stage1_9[53]}
   );
   gpc606_5 gpc112 (
      {stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[30],stage1_11[32],stage1_10[38],stage1_9[54]}
   );
   gpc606_5 gpc113 (
      {stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[31],stage1_11[33],stage1_10[39],stage1_9[55]}
   );
   gpc606_5 gpc114 (
      {stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[32],stage1_11[34],stage1_10[40],stage1_9[56]}
   );
   gpc606_5 gpc115 (
      {stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126], stage0_9[127]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[33],stage1_11[35],stage1_10[41],stage1_9[57]}
   );
   gpc606_5 gpc116 (
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[19],stage1_12[34],stage1_11[36],stage1_10[42]}
   );
   gpc606_5 gpc117 (
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[20],stage1_12[35],stage1_11[37],stage1_10[43]}
   );
   gpc615_5 gpc118 (
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106]},
      {stage0_11[114]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[21],stage1_12[36],stage1_11[38],stage1_10[44]}
   );
   gpc615_5 gpc119 (
      {stage0_10[107], stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111]},
      {stage0_11[115]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[22],stage1_12[37],stage1_11[39],stage1_10[45]}
   );
   gpc615_5 gpc120 (
      {stage0_10[112], stage0_10[113], stage0_10[114], stage0_10[115], stage0_10[116]},
      {stage0_11[116]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[23],stage1_12[38],stage1_11[40],stage1_10[46]}
   );
   gpc615_5 gpc121 (
      {stage0_10[117], stage0_10[118], stage0_10[119], stage0_10[120], stage0_10[121]},
      {stage0_11[117]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[24],stage1_12[39],stage1_11[41],stage1_10[47]}
   );
   gpc606_5 gpc122 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[0],stage1_14[6],stage1_13[25],stage1_12[40]}
   );
   gpc606_5 gpc123 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[1],stage1_14[7],stage1_13[26],stage1_12[41]}
   );
   gpc606_5 gpc124 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[2],stage1_14[8],stage1_13[27],stage1_12[42]}
   );
   gpc606_5 gpc125 (
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[3],stage1_14[9],stage1_13[28],stage1_12[43]}
   );
   gpc606_5 gpc126 (
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[4],stage1_14[10],stage1_13[29],stage1_12[44]}
   );
   gpc606_5 gpc127 (
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[5],stage1_14[11],stage1_13[30],stage1_12[45]}
   );
   gpc606_5 gpc128 (
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[6],stage1_14[12],stage1_13[31],stage1_12[46]}
   );
   gpc606_5 gpc129 (
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[7],stage1_14[13],stage1_13[32],stage1_12[47]}
   );
   gpc606_5 gpc130 (
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[8],stage1_14[14],stage1_13[33],stage1_12[48]}
   );
   gpc606_5 gpc131 (
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[9],stage1_14[15],stage1_13[34],stage1_12[49]}
   );
   gpc606_5 gpc132 (
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[10],stage1_14[16],stage1_13[35],stage1_12[50]}
   );
   gpc606_5 gpc133 (
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[11],stage1_14[17],stage1_13[36],stage1_12[51]}
   );
   gpc606_5 gpc134 (
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[12],stage1_14[18],stage1_13[37],stage1_12[52]}
   );
   gpc606_5 gpc135 (
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[13],stage1_14[19],stage1_13[38],stage1_12[53]}
   );
   gpc606_5 gpc136 (
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[14],stage1_14[20],stage1_13[39],stage1_12[54]}
   );
   gpc606_5 gpc137 (
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[15],stage1_15[15],stage1_14[21],stage1_13[40]}
   );
   gpc606_5 gpc138 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[16],stage1_15[16],stage1_14[22],stage1_13[41]}
   );
   gpc606_5 gpc139 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[17],stage1_15[17],stage1_14[23],stage1_13[42]}
   );
   gpc606_5 gpc140 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[18],stage1_15[18],stage1_14[24],stage1_13[43]}
   );
   gpc606_5 gpc141 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[19],stage1_15[19],stage1_14[25],stage1_13[44]}
   );
   gpc606_5 gpc142 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[20],stage1_15[20],stage1_14[26],stage1_13[45]}
   );
   gpc606_5 gpc143 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[21],stage1_15[21],stage1_14[27],stage1_13[46]}
   );
   gpc606_5 gpc144 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[22],stage1_15[22],stage1_14[28],stage1_13[47]}
   );
   gpc606_5 gpc145 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[23],stage1_15[23],stage1_14[29],stage1_13[48]}
   );
   gpc606_5 gpc146 (
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[24],stage1_15[24],stage1_14[30],stage1_13[49]}
   );
   gpc606_5 gpc147 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[25],stage1_15[25],stage1_14[31],stage1_13[50]}
   );
   gpc606_5 gpc148 (
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[26],stage1_15[26],stage1_14[32],stage1_13[51]}
   );
   gpc615_5 gpc149 (
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76]},
      {stage0_14[90]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[27],stage1_15[27],stage1_14[33],stage1_13[52]}
   );
   gpc615_5 gpc150 (
      {stage0_13[77], stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81]},
      {stage0_14[91]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[28],stage1_15[28],stage1_14[34],stage1_13[53]}
   );
   gpc615_5 gpc151 (
      {stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85], stage0_13[86]},
      {stage0_14[92]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[29],stage1_15[29],stage1_14[35],stage1_13[54]}
   );
   gpc615_5 gpc152 (
      {stage0_13[87], stage0_13[88], stage0_13[89], stage0_13[90], stage0_13[91]},
      {stage0_14[93]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[30],stage1_15[30],stage1_14[36],stage1_13[55]}
   );
   gpc615_5 gpc153 (
      {stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95], stage0_13[96]},
      {stage0_14[94]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[31],stage1_15[31],stage1_14[37],stage1_13[56]}
   );
   gpc615_5 gpc154 (
      {stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage0_14[95]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[32],stage1_15[32],stage1_14[38],stage1_13[57]}
   );
   gpc615_5 gpc155 (
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106]},
      {stage0_14[96]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[33],stage1_15[33],stage1_14[39],stage1_13[58]}
   );
   gpc615_5 gpc156 (
      {stage0_13[107], stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111]},
      {stage0_14[97]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[34],stage1_15[34],stage1_14[40],stage1_13[59]}
   );
   gpc615_5 gpc157 (
      {stage0_13[112], stage0_13[113], stage0_13[114], stage0_13[115], stage0_13[116]},
      {stage0_14[98]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[35],stage1_15[35],stage1_14[41],stage1_13[60]}
   );
   gpc1_1 gpc158 (
      {stage0_0[99]},
      {stage1_0[17]}
   );
   gpc1_1 gpc159 (
      {stage0_0[100]},
      {stage1_0[18]}
   );
   gpc1_1 gpc160 (
      {stage0_0[101]},
      {stage1_0[19]}
   );
   gpc1_1 gpc161 (
      {stage0_0[102]},
      {stage1_0[20]}
   );
   gpc1_1 gpc162 (
      {stage0_0[103]},
      {stage1_0[21]}
   );
   gpc1_1 gpc163 (
      {stage0_0[104]},
      {stage1_0[22]}
   );
   gpc1_1 gpc164 (
      {stage0_0[105]},
      {stage1_0[23]}
   );
   gpc1_1 gpc165 (
      {stage0_0[106]},
      {stage1_0[24]}
   );
   gpc1_1 gpc166 (
      {stage0_0[107]},
      {stage1_0[25]}
   );
   gpc1_1 gpc167 (
      {stage0_0[108]},
      {stage1_0[26]}
   );
   gpc1_1 gpc168 (
      {stage0_0[109]},
      {stage1_0[27]}
   );
   gpc1_1 gpc169 (
      {stage0_0[110]},
      {stage1_0[28]}
   );
   gpc1_1 gpc170 (
      {stage0_0[111]},
      {stage1_0[29]}
   );
   gpc1_1 gpc171 (
      {stage0_0[112]},
      {stage1_0[30]}
   );
   gpc1_1 gpc172 (
      {stage0_0[113]},
      {stage1_0[31]}
   );
   gpc1_1 gpc173 (
      {stage0_0[114]},
      {stage1_0[32]}
   );
   gpc1_1 gpc174 (
      {stage0_0[115]},
      {stage1_0[33]}
   );
   gpc1_1 gpc175 (
      {stage0_0[116]},
      {stage1_0[34]}
   );
   gpc1_1 gpc176 (
      {stage0_0[117]},
      {stage1_0[35]}
   );
   gpc1_1 gpc177 (
      {stage0_0[118]},
      {stage1_0[36]}
   );
   gpc1_1 gpc178 (
      {stage0_0[119]},
      {stage1_0[37]}
   );
   gpc1_1 gpc179 (
      {stage0_0[120]},
      {stage1_0[38]}
   );
   gpc1_1 gpc180 (
      {stage0_0[121]},
      {stage1_0[39]}
   );
   gpc1_1 gpc181 (
      {stage0_0[122]},
      {stage1_0[40]}
   );
   gpc1_1 gpc182 (
      {stage0_0[123]},
      {stage1_0[41]}
   );
   gpc1_1 gpc183 (
      {stage0_0[124]},
      {stage1_0[42]}
   );
   gpc1_1 gpc184 (
      {stage0_0[125]},
      {stage1_0[43]}
   );
   gpc1_1 gpc185 (
      {stage0_0[126]},
      {stage1_0[44]}
   );
   gpc1_1 gpc186 (
      {stage0_0[127]},
      {stage1_0[45]}
   );
   gpc1_1 gpc187 (
      {stage0_1[96]},
      {stage1_1[32]}
   );
   gpc1_1 gpc188 (
      {stage0_1[97]},
      {stage1_1[33]}
   );
   gpc1_1 gpc189 (
      {stage0_1[98]},
      {stage1_1[34]}
   );
   gpc1_1 gpc190 (
      {stage0_1[99]},
      {stage1_1[35]}
   );
   gpc1_1 gpc191 (
      {stage0_1[100]},
      {stage1_1[36]}
   );
   gpc1_1 gpc192 (
      {stage0_1[101]},
      {stage1_1[37]}
   );
   gpc1_1 gpc193 (
      {stage0_1[102]},
      {stage1_1[38]}
   );
   gpc1_1 gpc194 (
      {stage0_1[103]},
      {stage1_1[39]}
   );
   gpc1_1 gpc195 (
      {stage0_1[104]},
      {stage1_1[40]}
   );
   gpc1_1 gpc196 (
      {stage0_1[105]},
      {stage1_1[41]}
   );
   gpc1_1 gpc197 (
      {stage0_1[106]},
      {stage1_1[42]}
   );
   gpc1_1 gpc198 (
      {stage0_1[107]},
      {stage1_1[43]}
   );
   gpc1_1 gpc199 (
      {stage0_1[108]},
      {stage1_1[44]}
   );
   gpc1_1 gpc200 (
      {stage0_1[109]},
      {stage1_1[45]}
   );
   gpc1_1 gpc201 (
      {stage0_1[110]},
      {stage1_1[46]}
   );
   gpc1_1 gpc202 (
      {stage0_1[111]},
      {stage1_1[47]}
   );
   gpc1_1 gpc203 (
      {stage0_1[112]},
      {stage1_1[48]}
   );
   gpc1_1 gpc204 (
      {stage0_1[113]},
      {stage1_1[49]}
   );
   gpc1_1 gpc205 (
      {stage0_1[114]},
      {stage1_1[50]}
   );
   gpc1_1 gpc206 (
      {stage0_1[115]},
      {stage1_1[51]}
   );
   gpc1_1 gpc207 (
      {stage0_1[116]},
      {stage1_1[52]}
   );
   gpc1_1 gpc208 (
      {stage0_1[117]},
      {stage1_1[53]}
   );
   gpc1_1 gpc209 (
      {stage0_1[118]},
      {stage1_1[54]}
   );
   gpc1_1 gpc210 (
      {stage0_1[119]},
      {stage1_1[55]}
   );
   gpc1_1 gpc211 (
      {stage0_1[120]},
      {stage1_1[56]}
   );
   gpc1_1 gpc212 (
      {stage0_1[121]},
      {stage1_1[57]}
   );
   gpc1_1 gpc213 (
      {stage0_1[122]},
      {stage1_1[58]}
   );
   gpc1_1 gpc214 (
      {stage0_1[123]},
      {stage1_1[59]}
   );
   gpc1_1 gpc215 (
      {stage0_1[124]},
      {stage1_1[60]}
   );
   gpc1_1 gpc216 (
      {stage0_1[125]},
      {stage1_1[61]}
   );
   gpc1_1 gpc217 (
      {stage0_1[126]},
      {stage1_1[62]}
   );
   gpc1_1 gpc218 (
      {stage0_1[127]},
      {stage1_1[63]}
   );
   gpc1_1 gpc219 (
      {stage0_2[126]},
      {stage1_2[37]}
   );
   gpc1_1 gpc220 (
      {stage0_2[127]},
      {stage1_2[38]}
   );
   gpc1_1 gpc221 (
      {stage0_3[122]},
      {stage1_3[43]}
   );
   gpc1_1 gpc222 (
      {stage0_3[123]},
      {stage1_3[44]}
   );
   gpc1_1 gpc223 (
      {stage0_3[124]},
      {stage1_3[45]}
   );
   gpc1_1 gpc224 (
      {stage0_3[125]},
      {stage1_3[46]}
   );
   gpc1_1 gpc225 (
      {stage0_3[126]},
      {stage1_3[47]}
   );
   gpc1_1 gpc226 (
      {stage0_3[127]},
      {stage1_3[48]}
   );
   gpc1_1 gpc227 (
      {stage0_4[126]},
      {stage1_4[58]}
   );
   gpc1_1 gpc228 (
      {stage0_4[127]},
      {stage1_4[59]}
   );
   gpc1_1 gpc229 (
      {stage0_7[108]},
      {stage1_7[45]}
   );
   gpc1_1 gpc230 (
      {stage0_7[109]},
      {stage1_7[46]}
   );
   gpc1_1 gpc231 (
      {stage0_7[110]},
      {stage1_7[47]}
   );
   gpc1_1 gpc232 (
      {stage0_7[111]},
      {stage1_7[48]}
   );
   gpc1_1 gpc233 (
      {stage0_7[112]},
      {stage1_7[49]}
   );
   gpc1_1 gpc234 (
      {stage0_7[113]},
      {stage1_7[50]}
   );
   gpc1_1 gpc235 (
      {stage0_7[114]},
      {stage1_7[51]}
   );
   gpc1_1 gpc236 (
      {stage0_7[115]},
      {stage1_7[52]}
   );
   gpc1_1 gpc237 (
      {stage0_7[116]},
      {stage1_7[53]}
   );
   gpc1_1 gpc238 (
      {stage0_7[117]},
      {stage1_7[54]}
   );
   gpc1_1 gpc239 (
      {stage0_7[118]},
      {stage1_7[55]}
   );
   gpc1_1 gpc240 (
      {stage0_7[119]},
      {stage1_7[56]}
   );
   gpc1_1 gpc241 (
      {stage0_7[120]},
      {stage1_7[57]}
   );
   gpc1_1 gpc242 (
      {stage0_7[121]},
      {stage1_7[58]}
   );
   gpc1_1 gpc243 (
      {stage0_7[122]},
      {stage1_7[59]}
   );
   gpc1_1 gpc244 (
      {stage0_7[123]},
      {stage1_7[60]}
   );
   gpc1_1 gpc245 (
      {stage0_7[124]},
      {stage1_7[61]}
   );
   gpc1_1 gpc246 (
      {stage0_7[125]},
      {stage1_7[62]}
   );
   gpc1_1 gpc247 (
      {stage0_7[126]},
      {stage1_7[63]}
   );
   gpc1_1 gpc248 (
      {stage0_7[127]},
      {stage1_7[64]}
   );
   gpc1_1 gpc249 (
      {stage0_8[126]},
      {stage1_8[54]}
   );
   gpc1_1 gpc250 (
      {stage0_8[127]},
      {stage1_8[55]}
   );
   gpc1_1 gpc251 (
      {stage0_10[122]},
      {stage1_10[48]}
   );
   gpc1_1 gpc252 (
      {stage0_10[123]},
      {stage1_10[49]}
   );
   gpc1_1 gpc253 (
      {stage0_10[124]},
      {stage1_10[50]}
   );
   gpc1_1 gpc254 (
      {stage0_10[125]},
      {stage1_10[51]}
   );
   gpc1_1 gpc255 (
      {stage0_10[126]},
      {stage1_10[52]}
   );
   gpc1_1 gpc256 (
      {stage0_10[127]},
      {stage1_10[53]}
   );
   gpc1_1 gpc257 (
      {stage0_11[118]},
      {stage1_11[42]}
   );
   gpc1_1 gpc258 (
      {stage0_11[119]},
      {stage1_11[43]}
   );
   gpc1_1 gpc259 (
      {stage0_11[120]},
      {stage1_11[44]}
   );
   gpc1_1 gpc260 (
      {stage0_11[121]},
      {stage1_11[45]}
   );
   gpc1_1 gpc261 (
      {stage0_11[122]},
      {stage1_11[46]}
   );
   gpc1_1 gpc262 (
      {stage0_11[123]},
      {stage1_11[47]}
   );
   gpc1_1 gpc263 (
      {stage0_11[124]},
      {stage1_11[48]}
   );
   gpc1_1 gpc264 (
      {stage0_11[125]},
      {stage1_11[49]}
   );
   gpc1_1 gpc265 (
      {stage0_11[126]},
      {stage1_11[50]}
   );
   gpc1_1 gpc266 (
      {stage0_11[127]},
      {stage1_11[51]}
   );
   gpc1_1 gpc267 (
      {stage0_12[126]},
      {stage1_12[55]}
   );
   gpc1_1 gpc268 (
      {stage0_12[127]},
      {stage1_12[56]}
   );
   gpc1_1 gpc269 (
      {stage0_13[117]},
      {stage1_13[61]}
   );
   gpc1_1 gpc270 (
      {stage0_13[118]},
      {stage1_13[62]}
   );
   gpc1_1 gpc271 (
      {stage0_13[119]},
      {stage1_13[63]}
   );
   gpc1_1 gpc272 (
      {stage0_13[120]},
      {stage1_13[64]}
   );
   gpc1_1 gpc273 (
      {stage0_13[121]},
      {stage1_13[65]}
   );
   gpc1_1 gpc274 (
      {stage0_13[122]},
      {stage1_13[66]}
   );
   gpc1_1 gpc275 (
      {stage0_13[123]},
      {stage1_13[67]}
   );
   gpc1_1 gpc276 (
      {stage0_13[124]},
      {stage1_13[68]}
   );
   gpc1_1 gpc277 (
      {stage0_13[125]},
      {stage1_13[69]}
   );
   gpc1_1 gpc278 (
      {stage0_13[126]},
      {stage1_13[70]}
   );
   gpc1_1 gpc279 (
      {stage0_13[127]},
      {stage1_13[71]}
   );
   gpc1_1 gpc280 (
      {stage0_14[99]},
      {stage1_14[42]}
   );
   gpc1_1 gpc281 (
      {stage0_14[100]},
      {stage1_14[43]}
   );
   gpc1_1 gpc282 (
      {stage0_14[101]},
      {stage1_14[44]}
   );
   gpc1_1 gpc283 (
      {stage0_14[102]},
      {stage1_14[45]}
   );
   gpc1_1 gpc284 (
      {stage0_14[103]},
      {stage1_14[46]}
   );
   gpc1_1 gpc285 (
      {stage0_14[104]},
      {stage1_14[47]}
   );
   gpc1_1 gpc286 (
      {stage0_14[105]},
      {stage1_14[48]}
   );
   gpc1_1 gpc287 (
      {stage0_14[106]},
      {stage1_14[49]}
   );
   gpc1_1 gpc288 (
      {stage0_14[107]},
      {stage1_14[50]}
   );
   gpc1_1 gpc289 (
      {stage0_14[108]},
      {stage1_14[51]}
   );
   gpc1_1 gpc290 (
      {stage0_14[109]},
      {stage1_14[52]}
   );
   gpc1_1 gpc291 (
      {stage0_14[110]},
      {stage1_14[53]}
   );
   gpc1_1 gpc292 (
      {stage0_14[111]},
      {stage1_14[54]}
   );
   gpc1_1 gpc293 (
      {stage0_14[112]},
      {stage1_14[55]}
   );
   gpc1_1 gpc294 (
      {stage0_14[113]},
      {stage1_14[56]}
   );
   gpc1_1 gpc295 (
      {stage0_14[114]},
      {stage1_14[57]}
   );
   gpc1_1 gpc296 (
      {stage0_14[115]},
      {stage1_14[58]}
   );
   gpc1_1 gpc297 (
      {stage0_14[116]},
      {stage1_14[59]}
   );
   gpc1_1 gpc298 (
      {stage0_14[117]},
      {stage1_14[60]}
   );
   gpc1_1 gpc299 (
      {stage0_14[118]},
      {stage1_14[61]}
   );
   gpc1_1 gpc300 (
      {stage0_14[119]},
      {stage1_14[62]}
   );
   gpc1_1 gpc301 (
      {stage0_14[120]},
      {stage1_14[63]}
   );
   gpc1_1 gpc302 (
      {stage0_14[121]},
      {stage1_14[64]}
   );
   gpc1_1 gpc303 (
      {stage0_14[122]},
      {stage1_14[65]}
   );
   gpc1_1 gpc304 (
      {stage0_14[123]},
      {stage1_14[66]}
   );
   gpc1_1 gpc305 (
      {stage0_14[124]},
      {stage1_14[67]}
   );
   gpc1_1 gpc306 (
      {stage0_14[125]},
      {stage1_14[68]}
   );
   gpc1_1 gpc307 (
      {stage0_14[126]},
      {stage1_14[69]}
   );
   gpc1_1 gpc308 (
      {stage0_14[127]},
      {stage1_14[70]}
   );
   gpc1_1 gpc309 (
      {stage0_15[126]},
      {stage1_15[36]}
   );
   gpc1_1 gpc310 (
      {stage0_15[127]},
      {stage1_15[37]}
   );
   gpc1163_5 gpc311 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc312 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc313 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc314 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc315 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc316 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc317 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc318 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc606_5 gpc319 (
      {stage1_0[24], stage1_0[25], stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc606_5 gpc320 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc606_5 gpc321 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1406_5 gpc322 (
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage1_4[0]},
      {stage2_5[0],stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11]}
   );
   gpc615_5 gpc323 (
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58]},
      {stage1_2[26]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[1],stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12]}
   );
   gpc615_5 gpc324 (
      {stage1_1[59], stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63]},
      {stage1_2[27]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[2],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc325 (
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage2_6[0],stage2_5[3],stage2_4[14],stage2_3[14],stage2_2[14]}
   );
   gpc615_5 gpc326 (
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28]},
      {stage1_4[7]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[1],stage2_5[4],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc327 (
      {stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage1_4[8]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[2],stage2_5[5],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc328 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38]},
      {stage1_4[9]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[3],stage2_5[6],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc329 (
      {stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage1_4[10]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[4],stage2_5[7],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc330 (
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48]},
      {stage1_4[11]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[5],stage2_5[8],stage2_4[19],stage2_3[19]}
   );
   gpc606_5 gpc331 (
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[5],stage2_6[6],stage2_5[9],stage2_4[20]}
   );
   gpc606_5 gpc332 (
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[6],stage2_6[7],stage2_5[10],stage2_4[21]}
   );
   gpc606_5 gpc333 (
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[7],stage2_6[8],stage2_5[11],stage2_4[22]}
   );
   gpc606_5 gpc334 (
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[8],stage2_6[9],stage2_5[12],stage2_4[23]}
   );
   gpc606_5 gpc335 (
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[9],stage2_6[10],stage2_5[13],stage2_4[24]}
   );
   gpc606_5 gpc336 (
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[10],stage2_6[11],stage2_5[14],stage2_4[25]}
   );
   gpc606_5 gpc337 (
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[11],stage2_6[12],stage2_5[15],stage2_4[26]}
   );
   gpc606_5 gpc338 (
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[12],stage2_6[13],stage2_5[16],stage2_4[27]}
   );
   gpc207_4 gpc339 (
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36]},
      {stage1_7[0], stage1_7[1]},
      {stage2_8[8],stage2_7[13],stage2_6[14],stage2_5[17]}
   );
   gpc606_5 gpc340 (
      {stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41], stage1_5[42]},
      {stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7]},
      {stage2_9[0],stage2_8[9],stage2_7[14],stage2_6[15],stage2_5[18]}
   );
   gpc606_5 gpc341 (
      {stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47], stage1_5[48]},
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13]},
      {stage2_9[1],stage2_8[10],stage2_7[15],stage2_6[16],stage2_5[19]}
   );
   gpc615_5 gpc342 (
      {stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[2],stage2_8[11],stage2_7[16]}
   );
   gpc615_5 gpc343 (
      {stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage1_8[1]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[1],stage2_9[3],stage2_8[12],stage2_7[17]}
   );
   gpc615_5 gpc344 (
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28]},
      {stage1_8[2]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[2],stage2_9[4],stage2_8[13],stage2_7[18]}
   );
   gpc615_5 gpc345 (
      {stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33]},
      {stage1_8[3]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[3],stage2_9[5],stage2_8[14],stage2_7[19]}
   );
   gpc615_5 gpc346 (
      {stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37], stage1_7[38]},
      {stage1_8[4]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[4],stage2_9[6],stage2_8[15],stage2_7[20]}
   );
   gpc615_5 gpc347 (
      {stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage1_8[5]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[5],stage2_9[7],stage2_8[16],stage2_7[21]}
   );
   gpc615_5 gpc348 (
      {stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage1_8[6]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[6],stage2_9[8],stage2_8[17],stage2_7[22]}
   );
   gpc615_5 gpc349 (
      {stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage1_8[7]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[7],stage2_9[9],stage2_8[18],stage2_7[23]}
   );
   gpc615_5 gpc350 (
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58]},
      {stage1_8[8]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[8],stage2_9[10],stage2_8[19],stage2_7[24]}
   );
   gpc606_5 gpc351 (
      {stage1_8[9], stage1_8[10], stage1_8[11], stage1_8[12], stage1_8[13], stage1_8[14]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[9],stage2_10[9],stage2_9[11],stage2_8[20]}
   );
   gpc606_5 gpc352 (
      {stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19], stage1_8[20]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[10],stage2_10[10],stage2_9[12],stage2_8[21]}
   );
   gpc606_5 gpc353 (
      {stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[11],stage2_10[11],stage2_9[13],stage2_8[22]}
   );
   gpc606_5 gpc354 (
      {stage1_8[27], stage1_8[28], stage1_8[29], stage1_8[30], stage1_8[31], stage1_8[32]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[12],stage2_10[12],stage2_9[14],stage2_8[23]}
   );
   gpc606_5 gpc355 (
      {stage1_8[33], stage1_8[34], stage1_8[35], stage1_8[36], stage1_8[37], stage1_8[38]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[13],stage2_10[13],stage2_9[15],stage2_8[24]}
   );
   gpc606_5 gpc356 (
      {stage1_8[39], stage1_8[40], stage1_8[41], stage1_8[42], stage1_8[43], stage1_8[44]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[14],stage2_10[14],stage2_9[16],stage2_8[25]}
   );
   gpc615_5 gpc357 (
      {stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48], stage1_8[49]},
      {stage1_9[54]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[15],stage2_10[15],stage2_9[17],stage2_8[26]}
   );
   gpc615_5 gpc358 (
      {stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53], stage1_8[54]},
      {stage1_9[55]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[16],stage2_10[16],stage2_9[18],stage2_8[27]}
   );
   gpc606_5 gpc359 (
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[0],stage2_12[8],stage2_11[17],stage2_10[17]}
   );
   gpc615_5 gpc360 (
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[1],stage2_13[1],stage2_12[9],stage2_11[18]}
   );
   gpc615_5 gpc361 (
      {stage1_11[5], stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9]},
      {stage1_12[7]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[2],stage2_13[2],stage2_12[10],stage2_11[19]}
   );
   gpc615_5 gpc362 (
      {stage1_11[10], stage1_11[11], stage1_11[12], stage1_11[13], stage1_11[14]},
      {stage1_12[8]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[3],stage2_13[3],stage2_12[11],stage2_11[20]}
   );
   gpc615_5 gpc363 (
      {stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18], stage1_11[19]},
      {stage1_12[9]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[4],stage2_13[4],stage2_12[12],stage2_11[21]}
   );
   gpc615_5 gpc364 (
      {stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage1_12[10]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[5],stage2_13[5],stage2_12[13],stage2_11[22]}
   );
   gpc615_5 gpc365 (
      {stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage1_12[11]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[6],stage2_13[6],stage2_12[14],stage2_11[23]}
   );
   gpc615_5 gpc366 (
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34]},
      {stage1_12[12]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[7],stage2_13[7],stage2_12[15],stage2_11[24]}
   );
   gpc615_5 gpc367 (
      {stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39]},
      {stage1_12[13]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[8],stage2_13[8],stage2_12[16],stage2_11[25]}
   );
   gpc207_4 gpc368 (
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19], stage1_12[20]},
      {stage1_14[0], stage1_14[1]},
      {stage2_15[8],stage2_14[9],stage2_13[9],stage2_12[17]}
   );
   gpc606_5 gpc369 (
      {stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25], stage1_12[26]},
      {stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6], stage1_14[7]},
      {stage2_16[0],stage2_15[9],stage2_14[10],stage2_13[10],stage2_12[18]}
   );
   gpc606_5 gpc370 (
      {stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30], stage1_12[31], stage1_12[32]},
      {stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12], stage1_14[13]},
      {stage2_16[1],stage2_15[10],stage2_14[11],stage2_13[11],stage2_12[19]}
   );
   gpc606_5 gpc371 (
      {stage1_12[33], stage1_12[34], stage1_12[35], stage1_12[36], stage1_12[37], stage1_12[38]},
      {stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18], stage1_14[19]},
      {stage2_16[2],stage2_15[11],stage2_14[12],stage2_13[12],stage2_12[20]}
   );
   gpc606_5 gpc372 (
      {stage1_12[39], stage1_12[40], stage1_12[41], stage1_12[42], stage1_12[43], stage1_12[44]},
      {stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25]},
      {stage2_16[3],stage2_15[12],stage2_14[13],stage2_13[13],stage2_12[21]}
   );
   gpc606_5 gpc373 (
      {stage1_12[45], stage1_12[46], stage1_12[47], stage1_12[48], stage1_12[49], stage1_12[50]},
      {stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31]},
      {stage2_16[4],stage2_15[13],stage2_14[14],stage2_13[14],stage2_12[22]}
   );
   gpc606_5 gpc374 (
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[5],stage2_15[14],stage2_14[15],stage2_13[15]}
   );
   gpc606_5 gpc375 (
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[6],stage2_15[15],stage2_14[16],stage2_13[16]}
   );
   gpc606_5 gpc376 (
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[7],stage2_15[16],stage2_14[17],stage2_13[17]}
   );
   gpc606_5 gpc377 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[8],stage2_15[17],stage2_14[18],stage2_13[18]}
   );
   gpc606_5 gpc378 (
      {stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36], stage1_14[37]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[4],stage2_16[9],stage2_15[18],stage2_14[19]}
   );
   gpc606_5 gpc379 (
      {stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42], stage1_14[43]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[5],stage2_16[10],stage2_15[19],stage2_14[20]}
   );
   gpc606_5 gpc380 (
      {stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47], stage1_14[48], stage1_14[49]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[6],stage2_16[11],stage2_15[20],stage2_14[21]}
   );
   gpc615_5 gpc381 (
      {stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53], stage1_14[54]},
      {stage1_15[24]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[7],stage2_16[12],stage2_15[21],stage2_14[22]}
   );
   gpc615_5 gpc382 (
      {stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage1_15[25]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[8],stage2_16[13],stage2_15[22],stage2_14[23]}
   );
   gpc615_5 gpc383 (
      {stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29], stage1_15[30]},
      {stage1_16[30]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[5],stage2_17[9],stage2_16[14],stage2_15[23]}
   );
   gpc615_5 gpc384 (
      {stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage1_16[31]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[6],stage2_17[10],stage2_16[15],stage2_15[24]}
   );
   gpc1_1 gpc385 (
      {stage1_0[42]},
      {stage2_0[11]}
   );
   gpc1_1 gpc386 (
      {stage1_0[43]},
      {stage2_0[12]}
   );
   gpc1_1 gpc387 (
      {stage1_0[44]},
      {stage2_0[13]}
   );
   gpc1_1 gpc388 (
      {stage1_0[45]},
      {stage2_0[14]}
   );
   gpc1_1 gpc389 (
      {stage1_2[34]},
      {stage2_2[15]}
   );
   gpc1_1 gpc390 (
      {stage1_2[35]},
      {stage2_2[16]}
   );
   gpc1_1 gpc391 (
      {stage1_2[36]},
      {stage2_2[17]}
   );
   gpc1_1 gpc392 (
      {stage1_2[37]},
      {stage2_2[18]}
   );
   gpc1_1 gpc393 (
      {stage1_2[38]},
      {stage2_2[19]}
   );
   gpc1_1 gpc394 (
      {stage1_5[49]},
      {stage2_5[20]}
   );
   gpc1_1 gpc395 (
      {stage1_5[50]},
      {stage2_5[21]}
   );
   gpc1_1 gpc396 (
      {stage1_5[51]},
      {stage2_5[22]}
   );
   gpc1_1 gpc397 (
      {stage1_5[52]},
      {stage2_5[23]}
   );
   gpc1_1 gpc398 (
      {stage1_5[53]},
      {stage2_5[24]}
   );
   gpc1_1 gpc399 (
      {stage1_5[54]},
      {stage2_5[25]}
   );
   gpc1_1 gpc400 (
      {stage1_5[55]},
      {stage2_5[26]}
   );
   gpc1_1 gpc401 (
      {stage1_5[56]},
      {stage2_5[27]}
   );
   gpc1_1 gpc402 (
      {stage1_7[59]},
      {stage2_7[25]}
   );
   gpc1_1 gpc403 (
      {stage1_7[60]},
      {stage2_7[26]}
   );
   gpc1_1 gpc404 (
      {stage1_7[61]},
      {stage2_7[27]}
   );
   gpc1_1 gpc405 (
      {stage1_7[62]},
      {stage2_7[28]}
   );
   gpc1_1 gpc406 (
      {stage1_7[63]},
      {stage2_7[29]}
   );
   gpc1_1 gpc407 (
      {stage1_7[64]},
      {stage2_7[30]}
   );
   gpc1_1 gpc408 (
      {stage1_8[55]},
      {stage2_8[28]}
   );
   gpc1_1 gpc409 (
      {stage1_9[56]},
      {stage2_9[19]}
   );
   gpc1_1 gpc410 (
      {stage1_9[57]},
      {stage2_9[20]}
   );
   gpc1_1 gpc411 (
      {stage1_11[40]},
      {stage2_11[26]}
   );
   gpc1_1 gpc412 (
      {stage1_11[41]},
      {stage2_11[27]}
   );
   gpc1_1 gpc413 (
      {stage1_11[42]},
      {stage2_11[28]}
   );
   gpc1_1 gpc414 (
      {stage1_11[43]},
      {stage2_11[29]}
   );
   gpc1_1 gpc415 (
      {stage1_11[44]},
      {stage2_11[30]}
   );
   gpc1_1 gpc416 (
      {stage1_11[45]},
      {stage2_11[31]}
   );
   gpc1_1 gpc417 (
      {stage1_11[46]},
      {stage2_11[32]}
   );
   gpc1_1 gpc418 (
      {stage1_11[47]},
      {stage2_11[33]}
   );
   gpc1_1 gpc419 (
      {stage1_11[48]},
      {stage2_11[34]}
   );
   gpc1_1 gpc420 (
      {stage1_11[49]},
      {stage2_11[35]}
   );
   gpc1_1 gpc421 (
      {stage1_11[50]},
      {stage2_11[36]}
   );
   gpc1_1 gpc422 (
      {stage1_11[51]},
      {stage2_11[37]}
   );
   gpc1_1 gpc423 (
      {stage1_12[51]},
      {stage2_12[23]}
   );
   gpc1_1 gpc424 (
      {stage1_12[52]},
      {stage2_12[24]}
   );
   gpc1_1 gpc425 (
      {stage1_12[53]},
      {stage2_12[25]}
   );
   gpc1_1 gpc426 (
      {stage1_12[54]},
      {stage2_12[26]}
   );
   gpc1_1 gpc427 (
      {stage1_12[55]},
      {stage2_12[27]}
   );
   gpc1_1 gpc428 (
      {stage1_12[56]},
      {stage2_12[28]}
   );
   gpc1_1 gpc429 (
      {stage1_14[60]},
      {stage2_14[24]}
   );
   gpc1_1 gpc430 (
      {stage1_14[61]},
      {stage2_14[25]}
   );
   gpc1_1 gpc431 (
      {stage1_14[62]},
      {stage2_14[26]}
   );
   gpc1_1 gpc432 (
      {stage1_14[63]},
      {stage2_14[27]}
   );
   gpc1_1 gpc433 (
      {stage1_14[64]},
      {stage2_14[28]}
   );
   gpc1_1 gpc434 (
      {stage1_14[65]},
      {stage2_14[29]}
   );
   gpc1_1 gpc435 (
      {stage1_14[66]},
      {stage2_14[30]}
   );
   gpc1_1 gpc436 (
      {stage1_14[67]},
      {stage2_14[31]}
   );
   gpc1_1 gpc437 (
      {stage1_14[68]},
      {stage2_14[32]}
   );
   gpc1_1 gpc438 (
      {stage1_14[69]},
      {stage2_14[33]}
   );
   gpc1_1 gpc439 (
      {stage1_14[70]},
      {stage2_14[34]}
   );
   gpc1_1 gpc440 (
      {stage1_15[36]},
      {stage2_15[25]}
   );
   gpc1_1 gpc441 (
      {stage1_15[37]},
      {stage2_15[26]}
   );
   gpc1_1 gpc442 (
      {stage1_16[32]},
      {stage2_16[16]}
   );
   gpc1_1 gpc443 (
      {stage1_16[33]},
      {stage2_16[17]}
   );
   gpc1_1 gpc444 (
      {stage1_16[34]},
      {stage2_16[18]}
   );
   gpc1_1 gpc445 (
      {stage1_16[35]},
      {stage2_16[19]}
   );
   gpc1_1 gpc446 (
      {stage1_17[12]},
      {stage2_17[11]}
   );
   gpc1_1 gpc447 (
      {stage1_17[13]},
      {stage2_17[12]}
   );
   gpc1_1 gpc448 (
      {stage1_17[14]},
      {stage2_17[13]}
   );
   gpc1_1 gpc449 (
      {stage1_17[15]},
      {stage2_17[14]}
   );
   gpc1_1 gpc450 (
      {stage1_17[16]},
      {stage2_17[15]}
   );
   gpc1_1 gpc451 (
      {stage1_17[17]},
      {stage2_17[16]}
   );
   gpc1_1 gpc452 (
      {stage1_17[18]},
      {stage2_17[17]}
   );
   gpc1_1 gpc453 (
      {stage1_17[19]},
      {stage2_17[18]}
   );
   gpc1_1 gpc454 (
      {stage1_17[20]},
      {stage2_17[19]}
   );
   gpc606_5 gpc455 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc615_5 gpc456 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4]},
      {stage2_3[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc615_5 gpc457 (
      {stage2_2[5], stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9]},
      {stage2_3[7]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[2],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc1163_5 gpc458 (
      {stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage2_5[0]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[2],stage3_5[3],stage3_4[3],stage3_3[3]}
   );
   gpc1163_5 gpc459 (
      {stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage2_5[1]},
      {stage2_6[1]},
      {stage3_7[1],stage3_6[3],stage3_5[4],stage3_4[4],stage3_3[4]}
   );
   gpc606_5 gpc460 (
      {stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[0],stage3_7[2],stage3_6[4],stage3_5[5]}
   );
   gpc615_5 gpc461 (
      {stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12]},
      {stage2_6[2]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[1],stage3_7[3],stage3_6[5],stage3_5[6]}
   );
   gpc615_5 gpc462 (
      {stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage2_6[3]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[2],stage3_7[4],stage3_6[6],stage3_5[7]}
   );
   gpc615_5 gpc463 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22]},
      {stage2_6[4]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[3],stage3_7[5],stage3_6[7],stage3_5[8]}
   );
   gpc615_5 gpc464 (
      {stage2_5[23], stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27]},
      {stage2_6[5]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[4],stage3_7[6],stage3_6[8],stage3_5[9]}
   );
   gpc606_5 gpc465 (
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[5],stage3_8[5],stage3_7[7],stage3_6[9]}
   );
   gpc615_5 gpc466 (
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16]},
      {stage2_7[30]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[6],stage3_8[6],stage3_7[8],stage3_6[10]}
   );
   gpc606_5 gpc467 (
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[2],stage3_9[7],stage3_8[7]}
   );
   gpc606_5 gpc468 (
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[1],stage3_10[3],stage3_9[8],stage3_8[8]}
   );
   gpc1163_5 gpc469 (
      {stage2_9[0], stage2_9[1], stage2_9[2]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage2_11[0]},
      {stage2_12[0]},
      {stage3_13[0],stage3_12[2],stage3_11[2],stage3_10[4],stage3_9[9]}
   );
   gpc606_5 gpc470 (
      {stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6], stage2_9[7], stage2_9[8]},
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage3_13[1],stage3_12[3],stage3_11[3],stage3_10[5],stage3_9[10]}
   );
   gpc606_5 gpc471 (
      {stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12], stage2_9[13], stage2_9[14]},
      {stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11], stage2_11[12]},
      {stage3_13[2],stage3_12[4],stage3_11[4],stage3_10[6],stage3_9[11]}
   );
   gpc606_5 gpc472 (
      {stage2_9[15], stage2_9[16], stage2_9[17], stage2_9[18], stage2_9[19], stage2_9[20]},
      {stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18]},
      {stage3_13[3],stage3_12[5],stage3_11[5],stage3_10[7],stage3_9[12]}
   );
   gpc615_5 gpc473 (
      {stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage2_12[1]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[4],stage3_12[6],stage3_11[6]}
   );
   gpc615_5 gpc474 (
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28]},
      {stage2_12[2]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[5],stage3_12[7],stage3_11[7]}
   );
   gpc606_5 gpc475 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[2],stage3_14[2],stage3_13[6],stage3_12[8]}
   );
   gpc606_5 gpc476 (
      {stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[3],stage3_14[3],stage3_13[7],stage3_12[9]}
   );
   gpc606_5 gpc477 (
      {stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18], stage2_12[19], stage2_12[20]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[4],stage3_14[4],stage3_13[8],stage3_12[10]}
   );
   gpc606_5 gpc478 (
      {stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25], stage2_12[26]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[5],stage3_14[5],stage3_13[9],stage3_12[11]}
   );
   gpc606_5 gpc479 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[6],stage3_14[6],stage3_13[10]}
   );
   gpc1163_5 gpc480 (
      {stage2_14[24], stage2_14[25], stage2_14[26]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage2_16[0]},
      {stage2_17[0]},
      {stage3_18[0],stage3_17[1],stage3_16[5],stage3_15[7],stage3_14[7]}
   );
   gpc615_5 gpc481 (
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16]},
      {stage2_16[1]},
      {stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6]},
      {stage3_19[0],stage3_18[1],stage3_17[2],stage3_16[6],stage3_15[8]}
   );
   gpc615_5 gpc482 (
      {stage2_15[17], stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21]},
      {stage2_16[2]},
      {stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12]},
      {stage3_19[1],stage3_18[2],stage3_17[3],stage3_16[7],stage3_15[9]}
   );
   gpc615_5 gpc483 (
      {stage2_15[22], stage2_15[23], stage2_15[24], stage2_15[25], stage2_15[26]},
      {stage2_16[3]},
      {stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17], stage2_17[18]},
      {stage3_19[2],stage3_18[3],stage3_17[4],stage3_16[8],stage3_15[10]}
   );
   gpc606_5 gpc484 (
      {stage2_16[4], stage2_16[5], stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[3],stage3_18[4],stage3_17[5],stage3_16[9]}
   );
   gpc1_1 gpc485 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc486 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc487 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc488 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc489 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc490 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc491 (
      {stage2_0[6]},
      {stage3_0[6]}
   );
   gpc1_1 gpc492 (
      {stage2_0[7]},
      {stage3_0[7]}
   );
   gpc1_1 gpc493 (
      {stage2_0[8]},
      {stage3_0[8]}
   );
   gpc1_1 gpc494 (
      {stage2_0[9]},
      {stage3_0[9]}
   );
   gpc1_1 gpc495 (
      {stage2_0[10]},
      {stage3_0[10]}
   );
   gpc1_1 gpc496 (
      {stage2_0[11]},
      {stage3_0[11]}
   );
   gpc1_1 gpc497 (
      {stage2_0[12]},
      {stage3_0[12]}
   );
   gpc1_1 gpc498 (
      {stage2_0[13]},
      {stage3_0[13]}
   );
   gpc1_1 gpc499 (
      {stage2_0[14]},
      {stage3_0[14]}
   );
   gpc1_1 gpc500 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc501 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc502 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc503 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc504 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc505 (
      {stage2_1[11]},
      {stage3_1[6]}
   );
   gpc1_1 gpc506 (
      {stage2_1[12]},
      {stage3_1[7]}
   );
   gpc1_1 gpc507 (
      {stage2_1[13]},
      {stage3_1[8]}
   );
   gpc1_1 gpc508 (
      {stage2_2[10]},
      {stage3_2[3]}
   );
   gpc1_1 gpc509 (
      {stage2_2[11]},
      {stage3_2[4]}
   );
   gpc1_1 gpc510 (
      {stage2_2[12]},
      {stage3_2[5]}
   );
   gpc1_1 gpc511 (
      {stage2_2[13]},
      {stage3_2[6]}
   );
   gpc1_1 gpc512 (
      {stage2_2[14]},
      {stage3_2[7]}
   );
   gpc1_1 gpc513 (
      {stage2_2[15]},
      {stage3_2[8]}
   );
   gpc1_1 gpc514 (
      {stage2_2[16]},
      {stage3_2[9]}
   );
   gpc1_1 gpc515 (
      {stage2_2[17]},
      {stage3_2[10]}
   );
   gpc1_1 gpc516 (
      {stage2_2[18]},
      {stage3_2[11]}
   );
   gpc1_1 gpc517 (
      {stage2_2[19]},
      {stage3_2[12]}
   );
   gpc1_1 gpc518 (
      {stage2_3[14]},
      {stage3_3[5]}
   );
   gpc1_1 gpc519 (
      {stage2_3[15]},
      {stage3_3[6]}
   );
   gpc1_1 gpc520 (
      {stage2_3[16]},
      {stage3_3[7]}
   );
   gpc1_1 gpc521 (
      {stage2_3[17]},
      {stage3_3[8]}
   );
   gpc1_1 gpc522 (
      {stage2_3[18]},
      {stage3_3[9]}
   );
   gpc1_1 gpc523 (
      {stage2_3[19]},
      {stage3_3[10]}
   );
   gpc1_1 gpc524 (
      {stage2_4[24]},
      {stage3_4[5]}
   );
   gpc1_1 gpc525 (
      {stage2_4[25]},
      {stage3_4[6]}
   );
   gpc1_1 gpc526 (
      {stage2_4[26]},
      {stage3_4[7]}
   );
   gpc1_1 gpc527 (
      {stage2_4[27]},
      {stage3_4[8]}
   );
   gpc1_1 gpc528 (
      {stage2_8[24]},
      {stage3_8[9]}
   );
   gpc1_1 gpc529 (
      {stage2_8[25]},
      {stage3_8[10]}
   );
   gpc1_1 gpc530 (
      {stage2_8[26]},
      {stage3_8[11]}
   );
   gpc1_1 gpc531 (
      {stage2_8[27]},
      {stage3_8[12]}
   );
   gpc1_1 gpc532 (
      {stage2_8[28]},
      {stage3_8[13]}
   );
   gpc1_1 gpc533 (
      {stage2_11[29]},
      {stage3_11[8]}
   );
   gpc1_1 gpc534 (
      {stage2_11[30]},
      {stage3_11[9]}
   );
   gpc1_1 gpc535 (
      {stage2_11[31]},
      {stage3_11[10]}
   );
   gpc1_1 gpc536 (
      {stage2_11[32]},
      {stage3_11[11]}
   );
   gpc1_1 gpc537 (
      {stage2_11[33]},
      {stage3_11[12]}
   );
   gpc1_1 gpc538 (
      {stage2_11[34]},
      {stage3_11[13]}
   );
   gpc1_1 gpc539 (
      {stage2_11[35]},
      {stage3_11[14]}
   );
   gpc1_1 gpc540 (
      {stage2_11[36]},
      {stage3_11[15]}
   );
   gpc1_1 gpc541 (
      {stage2_11[37]},
      {stage3_11[16]}
   );
   gpc1_1 gpc542 (
      {stage2_12[27]},
      {stage3_12[12]}
   );
   gpc1_1 gpc543 (
      {stage2_12[28]},
      {stage3_12[13]}
   );
   gpc1_1 gpc544 (
      {stage2_13[18]},
      {stage3_13[11]}
   );
   gpc1_1 gpc545 (
      {stage2_14[27]},
      {stage3_14[8]}
   );
   gpc1_1 gpc546 (
      {stage2_14[28]},
      {stage3_14[9]}
   );
   gpc1_1 gpc547 (
      {stage2_14[29]},
      {stage3_14[10]}
   );
   gpc1_1 gpc548 (
      {stage2_14[30]},
      {stage3_14[11]}
   );
   gpc1_1 gpc549 (
      {stage2_14[31]},
      {stage3_14[12]}
   );
   gpc1_1 gpc550 (
      {stage2_14[32]},
      {stage3_14[13]}
   );
   gpc1_1 gpc551 (
      {stage2_14[33]},
      {stage3_14[14]}
   );
   gpc1_1 gpc552 (
      {stage2_14[34]},
      {stage3_14[15]}
   );
   gpc1_1 gpc553 (
      {stage2_16[10]},
      {stage3_16[10]}
   );
   gpc1_1 gpc554 (
      {stage2_16[11]},
      {stage3_16[11]}
   );
   gpc1_1 gpc555 (
      {stage2_16[12]},
      {stage3_16[12]}
   );
   gpc1_1 gpc556 (
      {stage2_16[13]},
      {stage3_16[13]}
   );
   gpc1_1 gpc557 (
      {stage2_16[14]},
      {stage3_16[14]}
   );
   gpc1_1 gpc558 (
      {stage2_16[15]},
      {stage3_16[15]}
   );
   gpc1_1 gpc559 (
      {stage2_16[16]},
      {stage3_16[16]}
   );
   gpc1_1 gpc560 (
      {stage2_16[17]},
      {stage3_16[17]}
   );
   gpc1_1 gpc561 (
      {stage2_16[18]},
      {stage3_16[18]}
   );
   gpc1_1 gpc562 (
      {stage2_16[19]},
      {stage3_16[19]}
   );
   gpc1_1 gpc563 (
      {stage2_17[19]},
      {stage3_17[6]}
   );
   gpc1_1 gpc564 (
      {stage2_18[6]},
      {stage3_18[5]}
   );
   gpc1_1 gpc565 (
      {stage2_19[0]},
      {stage3_19[4]}
   );
   gpc1_1 gpc566 (
      {stage2_19[1]},
      {stage3_19[5]}
   );
   gpc606_5 gpc567 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc568 (
      {stage3_0[6], stage3_0[7], stage3_0[8], stage3_0[9], stage3_0[10]},
      {stage3_1[0]},
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1],stage4_0[1]}
   );
   gpc1163_5 gpc569 (
      {stage3_3[0], stage3_3[1], stage3_3[2]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_5[0]},
      {stage3_6[0]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[2],stage4_3[2]}
   );
   gpc606_5 gpc570 (
      {stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1]}
   );
   gpc615_5 gpc571 (
      {stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage3_7[6]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[2],stage4_6[2]}
   );
   gpc615_5 gpc572 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[7]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[2],stage4_8[2],stage4_7[3],stage4_6[3]}
   );
   gpc606_5 gpc573 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[2],stage4_9[3]}
   );
   gpc615_5 gpc574 (
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10]},
      {stage3_10[0]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[1],stage4_10[3],stage4_9[4]}
   );
   gpc606_5 gpc575 (
      {stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[2],stage4_12[2],stage4_11[2],stage4_10[4]}
   );
   gpc615_5 gpc576 (
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16]},
      {stage3_12[6]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[1],stage4_13[3],stage4_12[3],stage4_11[3]}
   );
   gpc606_5 gpc577 (
      {stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11], stage3_12[12]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[2],stage4_13[4],stage4_12[4]}
   );
   gpc606_5 gpc578 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[3],stage4_13[5]}
   );
   gpc615_5 gpc579 (
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10]},
      {stage3_15[6]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[1],stage4_16[2],stage4_15[3],stage4_14[4]}
   );
   gpc615_5 gpc580 (
      {stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15]},
      {stage3_15[7]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[2],stage4_16[3],stage4_15[4],stage4_14[5]}
   );
   gpc606_5 gpc581 (
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[2],stage4_17[3],stage4_16[4]}
   );
   gpc606_5 gpc582 (
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[1],stage4_19[1],stage4_18[3],stage4_17[4]}
   );
   gpc1_1 gpc583 (
      {stage3_0[11]},
      {stage4_0[2]}
   );
   gpc1_1 gpc584 (
      {stage3_0[12]},
      {stage4_0[3]}
   );
   gpc1_1 gpc585 (
      {stage3_0[13]},
      {stage4_0[4]}
   );
   gpc1_1 gpc586 (
      {stage3_0[14]},
      {stage4_0[5]}
   );
   gpc1_1 gpc587 (
      {stage3_1[1]},
      {stage4_1[2]}
   );
   gpc1_1 gpc588 (
      {stage3_1[2]},
      {stage4_1[3]}
   );
   gpc1_1 gpc589 (
      {stage3_1[3]},
      {stage4_1[4]}
   );
   gpc1_1 gpc590 (
      {stage3_1[4]},
      {stage4_1[5]}
   );
   gpc1_1 gpc591 (
      {stage3_1[5]},
      {stage4_1[6]}
   );
   gpc1_1 gpc592 (
      {stage3_1[6]},
      {stage4_1[7]}
   );
   gpc1_1 gpc593 (
      {stage3_1[7]},
      {stage4_1[8]}
   );
   gpc1_1 gpc594 (
      {stage3_1[8]},
      {stage4_1[9]}
   );
   gpc1_1 gpc595 (
      {stage3_2[12]},
      {stage4_2[2]}
   );
   gpc1_1 gpc596 (
      {stage3_3[3]},
      {stage4_3[3]}
   );
   gpc1_1 gpc597 (
      {stage3_3[4]},
      {stage4_3[4]}
   );
   gpc1_1 gpc598 (
      {stage3_3[5]},
      {stage4_3[5]}
   );
   gpc1_1 gpc599 (
      {stage3_3[6]},
      {stage4_3[6]}
   );
   gpc1_1 gpc600 (
      {stage3_3[7]},
      {stage4_3[7]}
   );
   gpc1_1 gpc601 (
      {stage3_3[8]},
      {stage4_3[8]}
   );
   gpc1_1 gpc602 (
      {stage3_3[9]},
      {stage4_3[9]}
   );
   gpc1_1 gpc603 (
      {stage3_3[10]},
      {stage4_3[10]}
   );
   gpc1_1 gpc604 (
      {stage3_4[6]},
      {stage4_4[3]}
   );
   gpc1_1 gpc605 (
      {stage3_4[7]},
      {stage4_4[4]}
   );
   gpc1_1 gpc606 (
      {stage3_4[8]},
      {stage4_4[5]}
   );
   gpc1_1 gpc607 (
      {stage3_5[7]},
      {stage4_5[2]}
   );
   gpc1_1 gpc608 (
      {stage3_5[8]},
      {stage4_5[3]}
   );
   gpc1_1 gpc609 (
      {stage3_5[9]},
      {stage4_5[4]}
   );
   gpc1_1 gpc610 (
      {stage3_7[8]},
      {stage4_7[4]}
   );
   gpc1_1 gpc611 (
      {stage3_8[12]},
      {stage4_8[3]}
   );
   gpc1_1 gpc612 (
      {stage3_8[13]},
      {stage4_8[4]}
   );
   gpc1_1 gpc613 (
      {stage3_9[11]},
      {stage4_9[5]}
   );
   gpc1_1 gpc614 (
      {stage3_9[12]},
      {stage4_9[6]}
   );
   gpc1_1 gpc615 (
      {stage3_10[7]},
      {stage4_10[5]}
   );
   gpc1_1 gpc616 (
      {stage3_12[13]},
      {stage4_12[5]}
   );
   gpc1_1 gpc617 (
      {stage3_15[8]},
      {stage4_15[5]}
   );
   gpc1_1 gpc618 (
      {stage3_15[9]},
      {stage4_15[6]}
   );
   gpc1_1 gpc619 (
      {stage3_15[10]},
      {stage4_15[7]}
   );
   gpc1_1 gpc620 (
      {stage3_16[18]},
      {stage4_16[5]}
   );
   gpc1_1 gpc621 (
      {stage3_16[19]},
      {stage4_16[6]}
   );
   gpc1_1 gpc622 (
      {stage3_17[6]},
      {stage4_17[5]}
   );
   gpc1_1 gpc623 (
      {stage3_20[0]},
      {stage4_20[2]}
   );
   gpc2135_5 gpc624 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4]},
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0]},
      {stage4_3[0], stage4_3[1]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc1415_5 gpc625 (
      {stage4_1[3], stage4_1[4], stage4_1[5], stage4_1[6], stage4_1[7]},
      {stage4_2[1]},
      {stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage4_4[0]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc1415_5 gpc626 (
      {stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_5[0]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3]},
      {stage4_7[0]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[1],stage5_4[2]}
   );
   gpc615_5 gpc627 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[0]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[0],stage5_8[1]}
   );
   gpc606_5 gpc628 (
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[0],stage5_12[1]}
   );
   gpc135_4 gpc629 (
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4]},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[1]}
   );
   gpc1343_5 gpc630 (
      {stage4_18[0], stage4_18[1], stage4_18[2]},
      {stage4_19[0], stage4_19[1], 1'b0, 1'b0},
      {stage4_20[0], stage4_20[1], stage4_20[2]},
      {stage4_21[0]},
      {stage5_22[0],stage5_21[0],stage5_20[0],stage5_19[0],stage5_18[1]}
   );
   gpc1_1 gpc631 (
      {stage4_0[5]},
      {stage5_0[1]}
   );
   gpc1_1 gpc632 (
      {stage4_1[8]},
      {stage5_1[2]}
   );
   gpc1_1 gpc633 (
      {stage4_1[9]},
      {stage5_1[3]}
   );
   gpc1_1 gpc634 (
      {stage4_2[2]},
      {stage5_2[2]}
   );
   gpc1_1 gpc635 (
      {stage4_3[6]},
      {stage5_3[2]}
   );
   gpc1_1 gpc636 (
      {stage4_3[7]},
      {stage5_3[3]}
   );
   gpc1_1 gpc637 (
      {stage4_3[8]},
      {stage5_3[4]}
   );
   gpc1_1 gpc638 (
      {stage4_3[9]},
      {stage5_3[5]}
   );
   gpc1_1 gpc639 (
      {stage4_3[10]},
      {stage5_3[6]}
   );
   gpc1_1 gpc640 (
      {stage4_5[1]},
      {stage5_5[2]}
   );
   gpc1_1 gpc641 (
      {stage4_5[2]},
      {stage5_5[3]}
   );
   gpc1_1 gpc642 (
      {stage4_5[3]},
      {stage5_5[4]}
   );
   gpc1_1 gpc643 (
      {stage4_5[4]},
      {stage5_5[5]}
   );
   gpc1_1 gpc644 (
      {stage4_7[1]},
      {stage5_7[1]}
   );
   gpc1_1 gpc645 (
      {stage4_7[2]},
      {stage5_7[2]}
   );
   gpc1_1 gpc646 (
      {stage4_7[3]},
      {stage5_7[3]}
   );
   gpc1_1 gpc647 (
      {stage4_7[4]},
      {stage5_7[4]}
   );
   gpc1_1 gpc648 (
      {stage4_9[1]},
      {stage5_9[1]}
   );
   gpc1_1 gpc649 (
      {stage4_9[2]},
      {stage5_9[2]}
   );
   gpc1_1 gpc650 (
      {stage4_9[3]},
      {stage5_9[3]}
   );
   gpc1_1 gpc651 (
      {stage4_9[4]},
      {stage5_9[4]}
   );
   gpc1_1 gpc652 (
      {stage4_9[5]},
      {stage5_9[5]}
   );
   gpc1_1 gpc653 (
      {stage4_9[6]},
      {stage5_9[6]}
   );
   gpc1_1 gpc654 (
      {stage4_11[0]},
      {stage5_11[1]}
   );
   gpc1_1 gpc655 (
      {stage4_11[1]},
      {stage5_11[2]}
   );
   gpc1_1 gpc656 (
      {stage4_11[2]},
      {stage5_11[3]}
   );
   gpc1_1 gpc657 (
      {stage4_11[3]},
      {stage5_11[4]}
   );
   gpc1_1 gpc658 (
      {stage4_13[0]},
      {stage5_13[1]}
   );
   gpc1_1 gpc659 (
      {stage4_13[1]},
      {stage5_13[2]}
   );
   gpc1_1 gpc660 (
      {stage4_13[2]},
      {stage5_13[3]}
   );
   gpc1_1 gpc661 (
      {stage4_13[3]},
      {stage5_13[4]}
   );
   gpc1_1 gpc662 (
      {stage4_13[4]},
      {stage5_13[5]}
   );
   gpc1_1 gpc663 (
      {stage4_13[5]},
      {stage5_13[6]}
   );
   gpc1_1 gpc664 (
      {stage4_15[5]},
      {stage5_15[2]}
   );
   gpc1_1 gpc665 (
      {stage4_15[6]},
      {stage5_15[3]}
   );
   gpc1_1 gpc666 (
      {stage4_15[7]},
      {stage5_15[4]}
   );
   gpc1_1 gpc667 (
      {stage4_16[3]},
      {stage5_16[2]}
   );
   gpc1_1 gpc668 (
      {stage4_16[4]},
      {stage5_16[3]}
   );
   gpc1_1 gpc669 (
      {stage4_16[5]},
      {stage5_16[4]}
   );
   gpc1_1 gpc670 (
      {stage4_16[6]},
      {stage5_16[5]}
   );
   gpc1_1 gpc671 (
      {stage4_17[1]},
      {stage5_17[1]}
   );
   gpc1_1 gpc672 (
      {stage4_17[2]},
      {stage5_17[2]}
   );
   gpc1_1 gpc673 (
      {stage4_17[3]},
      {stage5_17[3]}
   );
   gpc1_1 gpc674 (
      {stage4_17[4]},
      {stage5_17[4]}
   );
   gpc1_1 gpc675 (
      {stage4_17[5]},
      {stage5_17[5]}
   );
   gpc1_1 gpc676 (
      {stage4_18[3]},
      {stage5_18[2]}
   );
   gpc2223_5 gpc677 (
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0], stage5_2[1]},
      {stage5_3[0], stage5_3[1]},
      {stage5_4[0], stage5_4[1]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0]}
   );
   gpc615_5 gpc678 (
      {stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5], stage5_3[6]},
      {stage5_4[2]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc615_5 gpc679 (
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4]},
      {stage5_8[0]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[1]}
   );
   gpc615_5 gpc680 (
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4]},
      {stage5_12[0]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[0],stage6_11[1]}
   );
   gpc615_5 gpc681 (
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4]},
      {stage5_16[0]},
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage6_19[0],stage6_18[0],stage6_17[0],stage6_16[0],stage6_15[1]}
   );
   gpc1415_5 gpc682 (
      {stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5]},
      {1'b0},
      {stage5_18[0], stage5_18[1], stage5_18[2], 1'b0},
      {stage5_19[0]},
      {stage6_20[0],stage6_19[1],stage6_18[1],stage6_17[1],stage6_16[1]}
   );
   gpc1_1 gpc683 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc684 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc685 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc686 (
      {stage5_2[2]},
      {stage6_2[1]}
   );
   gpc1_1 gpc687 (
      {stage5_6[0]},
      {stage6_6[1]}
   );
   gpc1_1 gpc688 (
      {stage5_8[1]},
      {stage6_8[1]}
   );
   gpc1_1 gpc689 (
      {stage5_9[6]},
      {stage6_9[1]}
   );
   gpc1_1 gpc690 (
      {stage5_10[0]},
      {stage6_10[1]}
   );
   gpc1_1 gpc691 (
      {stage5_12[1]},
      {stage6_12[1]}
   );
   gpc1_1 gpc692 (
      {stage5_13[6]},
      {stage6_13[1]}
   );
   gpc1_1 gpc693 (
      {stage5_14[0]},
      {stage6_14[1]}
   );
   gpc1_1 gpc694 (
      {stage5_20[0]},
      {stage6_20[1]}
   );
   gpc1_1 gpc695 (
      {stage5_21[0]},
      {stage6_21[0]}
   );
   gpc1_1 gpc696 (
      {stage5_22[0]},
      {stage6_22[0]}
   );
endmodule
module rowadder2_1_23(input [22:0] src0, input [22:0] src1, output [23:0] dst0);
    wire [22:0] gene;
    wire [22:0] prop;
    wire [23:0] out;
    wire [23:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI({1'h0, gene[22:20]}),
        .S({1'h0, prop[22:20]})
    );
    assign dst0 = {carryout[22], out[22:0]};
endmodule


module comp2_1test_128_16();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    reg [15:0] src54;
    reg [15:0] src55;
    reg [15:0] src56;
    reg [15:0] src57;
    reg [15:0] src58;
    reg [15:0] src59;
    reg [15:0] src60;
    reg [15:0] src61;
    reg [15:0] src62;
    reg [15:0] src63;
    reg [15:0] src64;
    reg [15:0] src65;
    reg [15:0] src66;
    reg [15:0] src67;
    reg [15:0] src68;
    reg [15:0] src69;
    reg [15:0] src70;
    reg [15:0] src71;
    reg [15:0] src72;
    reg [15:0] src73;
    reg [15:0] src74;
    reg [15:0] src75;
    reg [15:0] src76;
    reg [15:0] src77;
    reg [15:0] src78;
    reg [15:0] src79;
    reg [15:0] src80;
    reg [15:0] src81;
    reg [15:0] src82;
    reg [15:0] src83;
    reg [15:0] src84;
    reg [15:0] src85;
    reg [15:0] src86;
    reg [15:0] src87;
    reg [15:0] src88;
    reg [15:0] src89;
    reg [15:0] src90;
    reg [15:0] src91;
    reg [15:0] src92;
    reg [15:0] src93;
    reg [15:0] src94;
    reg [15:0] src95;
    reg [15:0] src96;
    reg [15:0] src97;
    reg [15:0] src98;
    reg [15:0] src99;
    reg [15:0] src100;
    reg [15:0] src101;
    reg [15:0] src102;
    reg [15:0] src103;
    reg [15:0] src104;
    reg [15:0] src105;
    reg [15:0] src106;
    reg [15:0] src107;
    reg [15:0] src108;
    reg [15:0] src109;
    reg [15:0] src110;
    reg [15:0] src111;
    reg [15:0] src112;
    reg [15:0] src113;
    reg [15:0] src114;
    reg [15:0] src115;
    reg [15:0] src116;
    reg [15:0] src117;
    reg [15:0] src118;
    reg [15:0] src119;
    reg [15:0] src120;
    reg [15:0] src121;
    reg [15:0] src122;
    reg [15:0] src123;
    reg [15:0] src124;
    reg [15:0] src125;
    reg [15:0] src126;
    reg [15:0] src127;
    reg [22:0] exp;
    wire [22:0] dst;
    assign test = dst == exp;
    compressor2_1_128_16 compressor2_1_128_16_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .src64(src64),
        .src65(src65),
        .src66(src66),
        .src67(src67),
        .src68(src68),
        .src69(src69),
        .src70(src70),
        .src71(src71),
        .src72(src72),
        .src73(src73),
        .src74(src74),
        .src75(src75),
        .src76(src76),
        .src77(src77),
        .src78(src78),
        .src79(src79),
        .src80(src80),
        .src81(src81),
        .src82(src82),
        .src83(src83),
        .src84(src84),
        .src85(src85),
        .src86(src86),
        .src87(src87),
        .src88(src88),
        .src89(src89),
        .src90(src90),
        .src91(src91),
        .src92(src92),
        .src93(src93),
        .src94(src94),
        .src95(src95),
        .src96(src96),
        .src97(src97),
        .src98(src98),
        .src99(src99),
        .src100(src100),
        .src101(src101),
        .src102(src102),
        .src103(src103),
        .src104(src104),
        .src105(src105),
        .src106(src106),
        .src107(src107),
        .src108(src108),
        .src109(src109),
        .src110(src110),
        .src111(src111),
        .src112(src112),
        .src113(src113),
        .src114(src114),
        .src115(src115),
        .src116(src116),
        .src117(src117),
        .src118(src118),
        .src119(src119),
        .src120(src120),
        .src121(src121),
        .src122(src122),
        .src123(src123),
        .src124(src124),
        .src125(src125),
        .src126(src126),
        .src127(src127),
        .dst(dst)
    );
    initial begin
        $monitor("0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x %x", src0, src1, src2, src3, src4, src5, src6, src7, src8, src9, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, src32, src33, src34, src35, src36, src37, src38, src39, src40, src41, src42, src43, src44, src45, src46, src47, src48, src49, src50, src51, src52, src53, src54, src55, src56, src57, src58, src59, src60, src61, src62, src63, src64, src65, src66, src67, src68, src69, src70, src71, src72, src73, src74, src75, src76, src77, src78, src79, src80, src81, src82, src83, src84, src85, src86, src87, src88, src89, src90, src91, src92, src93, src94, src95, src96, src97, src98, src99, src100, src101, src102, src103, src104, src105, src106, src107, src108, src109, src110, src111, src112, src113, src114, src115, src116, src117, src118, src119, src120, src121, src122, src123, src124, src125, src126, src127, dst, exp, test);
        src0 <= 16'hd1c0;
        src1 <= 16'h340e;
        src2 <= 16'h6f87;
        src3 <= 16'h4506;
        src4 <= 16'h672;
        src5 <= 16'he3ba;
        src6 <= 16'h6f1f;
        src7 <= 16'h93d4;
        src8 <= 16'h364e;
        src9 <= 16'ha17e;
        src10 <= 16'hbdcc;
        src11 <= 16'hc501;
        src12 <= 16'h826c;
        src13 <= 16'h42ef;
        src14 <= 16'h1a86;
        src15 <= 16'h8528;
        src16 <= 16'ha344;
        src17 <= 16'ha358;
        src18 <= 16'h757e;
        src19 <= 16'h87b0;
        src20 <= 16'h28f3;
        src21 <= 16'hd191;
        src22 <= 16'h4e22;
        src23 <= 16'h76c3;
        src24 <= 16'h7e2a;
        src25 <= 16'he9c7;
        src26 <= 16'h6eb1;
        src27 <= 16'hd8e2;
        src28 <= 16'hc5f;
        src29 <= 16'h1af6;
        src30 <= 16'h4bd3;
        src31 <= 16'h48b4;
        src32 <= 16'h75a8;
        src33 <= 16'h382e;
        src34 <= 16'he17e;
        src35 <= 16'h81bb;
        src36 <= 16'hffd4;
        src37 <= 16'h908a;
        src38 <= 16'h998d;
        src39 <= 16'hbd3d;
        src40 <= 16'hebf9;
        src41 <= 16'h3704;
        src42 <= 16'h1a02;
        src43 <= 16'h8151;
        src44 <= 16'hca6c;
        src45 <= 16'h583c;
        src46 <= 16'h19f0;
        src47 <= 16'h5477;
        src48 <= 16'h9fae;
        src49 <= 16'hed51;
        src50 <= 16'h58d7;
        src51 <= 16'h3f66;
        src52 <= 16'he814;
        src53 <= 16'hdbe7;
        src54 <= 16'haaaa;
        src55 <= 16'hf179;
        src56 <= 16'h3c3;
        src57 <= 16'h7ffc;
        src58 <= 16'h1571;
        src59 <= 16'h2f93;
        src60 <= 16'hacfe;
        src61 <= 16'h9e57;
        src62 <= 16'h7f78;
        src63 <= 16'hb72d;
        src64 <= 16'he5bd;
        src65 <= 16'h9f02;
        src66 <= 16'h8157;
        src67 <= 16'hd6e;
        src68 <= 16'h12fe;
        src69 <= 16'h22be;
        src70 <= 16'ha1e8;
        src71 <= 16'h96a2;
        src72 <= 16'h4c07;
        src73 <= 16'h2db3;
        src74 <= 16'hd269;
        src75 <= 16'haafa;
        src76 <= 16'h6537;
        src77 <= 16'h7287;
        src78 <= 16'h5292;
        src79 <= 16'h17cc;
        src80 <= 16'ha559;
        src81 <= 16'h6c50;
        src82 <= 16'hf804;
        src83 <= 16'h8fdc;
        src84 <= 16'h128e;
        src85 <= 16'ha838;
        src86 <= 16'h1e7e;
        src87 <= 16'hc533;
        src88 <= 16'h94d6;
        src89 <= 16'hcaec;
        src90 <= 16'hd28b;
        src91 <= 16'h5d7a;
        src92 <= 16'h9f35;
        src93 <= 16'hae3f;
        src94 <= 16'h7b;
        src95 <= 16'h9dad;
        src96 <= 16'h4f66;
        src97 <= 16'h28f1;
        src98 <= 16'h3a29;
        src99 <= 16'h9a02;
        src100 <= 16'h3df8;
        src101 <= 16'h7f93;
        src102 <= 16'h22c6;
        src103 <= 16'h97e2;
        src104 <= 16'he2a4;
        src105 <= 16'hf880;
        src106 <= 16'hf085;
        src107 <= 16'hfdb1;
        src108 <= 16'hf92b;
        src109 <= 16'hedab;
        src110 <= 16'h43d7;
        src111 <= 16'ha9c2;
        src112 <= 16'ha68e;
        src113 <= 16'h1ed4;
        src114 <= 16'h5bf8;
        src115 <= 16'hafec;
        src116 <= 16'h3bf8;
        src117 <= 16'h1f64;
        src118 <= 16'ha516;
        src119 <= 16'hac3d;
        src120 <= 16'h59fa;
        src121 <= 16'h36ee;
        src122 <= 16'h68af;
        src123 <= 16'h7cae;
        src124 <= 16'hbd98;
        src125 <= 16'h9af9;
        src126 <= 16'h8bf4;
        src127 <= 16'hc88;
        exp <= 23'h3fa387;
        #1
        src0 <= 16'hc660;
        src1 <= 16'h96ee;
        src2 <= 16'ha586;
        src3 <= 16'h1c2c;
        src4 <= 16'he10;
        src5 <= 16'hb0b9;
        src6 <= 16'hea9e;
        src7 <= 16'h552e;
        src8 <= 16'h5e1e;
        src9 <= 16'h8dcd;
        src10 <= 16'h3231;
        src11 <= 16'h4dd9;
        src12 <= 16'h18bc;
        src13 <= 16'h1896;
        src14 <= 16'hdf78;
        src15 <= 16'hc4bd;
        src16 <= 16'h89f3;
        src17 <= 16'h4452;
        src18 <= 16'h5029;
        src19 <= 16'h739;
        src20 <= 16'h8d0b;
        src21 <= 16'h8c27;
        src22 <= 16'hc6da;
        src23 <= 16'h6d37;
        src24 <= 16'ha4f6;
        src25 <= 16'h81d8;
        src26 <= 16'hae2;
        src27 <= 16'h81b2;
        src28 <= 16'h4153;
        src29 <= 16'h1b0c;
        src30 <= 16'hfd44;
        src31 <= 16'hcb91;
        src32 <= 16'h9c8b;
        src33 <= 16'he484;
        src34 <= 16'h4b99;
        src35 <= 16'h9fe6;
        src36 <= 16'h72a2;
        src37 <= 16'hd9ea;
        src38 <= 16'hd47f;
        src39 <= 16'he758;
        src40 <= 16'h62b2;
        src41 <= 16'he508;
        src42 <= 16'hd43f;
        src43 <= 16'hf200;
        src44 <= 16'h20ad;
        src45 <= 16'he76e;
        src46 <= 16'hc179;
        src47 <= 16'h8bc;
        src48 <= 16'h1d08;
        src49 <= 16'h462c;
        src50 <= 16'h72be;
        src51 <= 16'hd9b2;
        src52 <= 16'ha6bf;
        src53 <= 16'h9e03;
        src54 <= 16'hb892;
        src55 <= 16'h67cb;
        src56 <= 16'h2a90;
        src57 <= 16'hded8;
        src58 <= 16'h44f;
        src59 <= 16'h243f;
        src60 <= 16'h7ea9;
        src61 <= 16'h9a31;
        src62 <= 16'h3fe8;
        src63 <= 16'h2ffc;
        src64 <= 16'hfead;
        src65 <= 16'hb229;
        src66 <= 16'h8e27;
        src67 <= 16'h4331;
        src68 <= 16'h864a;
        src69 <= 16'he32f;
        src70 <= 16'h57c5;
        src71 <= 16'hde01;
        src72 <= 16'hbdb5;
        src73 <= 16'h738e;
        src74 <= 16'h9b64;
        src75 <= 16'h93ab;
        src76 <= 16'h798c;
        src77 <= 16'h1399;
        src78 <= 16'h5c3f;
        src79 <= 16'hb88f;
        src80 <= 16'h9b06;
        src81 <= 16'hea68;
        src82 <= 16'hd7b6;
        src83 <= 16'hb0d2;
        src84 <= 16'hbdd2;
        src85 <= 16'hde50;
        src86 <= 16'h7c4b;
        src87 <= 16'hc34;
        src88 <= 16'h78e1;
        src89 <= 16'h8f62;
        src90 <= 16'h9461;
        src91 <= 16'h1671;
        src92 <= 16'h4831;
        src93 <= 16'h6b43;
        src94 <= 16'hc2b6;
        src95 <= 16'hba05;
        src96 <= 16'hd4e7;
        src97 <= 16'h6eaa;
        src98 <= 16'hbcf8;
        src99 <= 16'h3c59;
        src100 <= 16'h92ea;
        src101 <= 16'hb154;
        src102 <= 16'h7295;
        src103 <= 16'h7308;
        src104 <= 16'hdd44;
        src105 <= 16'hc925;
        src106 <= 16'hd2b3;
        src107 <= 16'hc029;
        src108 <= 16'hc882;
        src109 <= 16'h2ed0;
        src110 <= 16'h7df9;
        src111 <= 16'h929d;
        src112 <= 16'h5a63;
        src113 <= 16'hb008;
        src114 <= 16'hcac;
        src115 <= 16'h77;
        src116 <= 16'h4585;
        src117 <= 16'h72ad;
        src118 <= 16'h8878;
        src119 <= 16'ha57;
        src120 <= 16'h65ae;
        src121 <= 16'hb00f;
        src122 <= 16'h9d57;
        src123 <= 16'hcbab;
        src124 <= 16'h7ffa;
        src125 <= 16'h5137;
        src126 <= 16'ha149;
        src127 <= 16'h8274;
        exp <= 23'h4286f5;
        #1
        src0 <= 16'hf5dc;
        src1 <= 16'h44a9;
        src2 <= 16'hec14;
        src3 <= 16'h892f;
        src4 <= 16'h3881;
        src5 <= 16'h626f;
        src6 <= 16'h53f7;
        src7 <= 16'h16af;
        src8 <= 16'h6a03;
        src9 <= 16'h721b;
        src10 <= 16'haa55;
        src11 <= 16'h775;
        src12 <= 16'hea1c;
        src13 <= 16'h2f20;
        src14 <= 16'hc670;
        src15 <= 16'h7f1;
        src16 <= 16'hc71d;
        src17 <= 16'h494c;
        src18 <= 16'hc5da;
        src19 <= 16'h1541;
        src20 <= 16'h96c6;
        src21 <= 16'ha893;
        src22 <= 16'hbb96;
        src23 <= 16'ha470;
        src24 <= 16'h7bcc;
        src25 <= 16'hf6af;
        src26 <= 16'hfdf;
        src27 <= 16'hc7c1;
        src28 <= 16'h39c0;
        src29 <= 16'h3a8d;
        src30 <= 16'h5e0f;
        src31 <= 16'h87fe;
        src32 <= 16'hd2e2;
        src33 <= 16'h2590;
        src34 <= 16'h3e66;
        src35 <= 16'h112c;
        src36 <= 16'hc276;
        src37 <= 16'hb526;
        src38 <= 16'hf413;
        src39 <= 16'h5add;
        src40 <= 16'hd392;
        src41 <= 16'h2b57;
        src42 <= 16'h246;
        src43 <= 16'hcda5;
        src44 <= 16'hfce3;
        src45 <= 16'hd7ac;
        src46 <= 16'h2afa;
        src47 <= 16'hb15f;
        src48 <= 16'ha465;
        src49 <= 16'h8a1e;
        src50 <= 16'h1101;
        src51 <= 16'hd77c;
        src52 <= 16'h6737;
        src53 <= 16'hc54;
        src54 <= 16'ha964;
        src55 <= 16'h8888;
        src56 <= 16'hefdd;
        src57 <= 16'hc8a5;
        src58 <= 16'h3a8a;
        src59 <= 16'ha64d;
        src60 <= 16'hda74;
        src61 <= 16'hd605;
        src62 <= 16'ha12c;
        src63 <= 16'h9238;
        src64 <= 16'h94d1;
        src65 <= 16'hed1e;
        src66 <= 16'he47d;
        src67 <= 16'h1d4f;
        src68 <= 16'hbc01;
        src69 <= 16'he508;
        src70 <= 16'h6e9c;
        src71 <= 16'hddb4;
        src72 <= 16'h8787;
        src73 <= 16'hfdfa;
        src74 <= 16'hf458;
        src75 <= 16'h63ad;
        src76 <= 16'h6908;
        src77 <= 16'hf594;
        src78 <= 16'ha4dc;
        src79 <= 16'h2a6f;
        src80 <= 16'ha7ca;
        src81 <= 16'he16f;
        src82 <= 16'h92e4;
        src83 <= 16'hd10;
        src84 <= 16'hcee7;
        src85 <= 16'hcec9;
        src86 <= 16'hb5a0;
        src87 <= 16'h385f;
        src88 <= 16'h8a23;
        src89 <= 16'hba41;
        src90 <= 16'he243;
        src91 <= 16'hb854;
        src92 <= 16'hb8fd;
        src93 <= 16'h2a26;
        src94 <= 16'hf3af;
        src95 <= 16'h6559;
        src96 <= 16'h32f5;
        src97 <= 16'h832e;
        src98 <= 16'h65ca;
        src99 <= 16'h8810;
        src100 <= 16'h2bed;
        src101 <= 16'h5bec;
        src102 <= 16'hac26;
        src103 <= 16'hdf02;
        src104 <= 16'h292d;
        src105 <= 16'hf168;
        src106 <= 16'h786;
        src107 <= 16'h9749;
        src108 <= 16'h3362;
        src109 <= 16'ha479;
        src110 <= 16'hc056;
        src111 <= 16'h3a7b;
        src112 <= 16'ha8a8;
        src113 <= 16'h5100;
        src114 <= 16'h382;
        src115 <= 16'h8717;
        src116 <= 16'h583f;
        src117 <= 16'h36b7;
        src118 <= 16'h82de;
        src119 <= 16'h96c;
        src120 <= 16'hae7;
        src121 <= 16'hd629;
        src122 <= 16'h864b;
        src123 <= 16'hf7aa;
        src124 <= 16'h6a09;
        src125 <= 16'h4462;
        src126 <= 16'h619d;
        src127 <= 16'hee8f;
        exp <= 23'h43aee2;
        #1
        src0 <= 16'h67b0;
        src1 <= 16'hc837;
        src2 <= 16'hc153;
        src3 <= 16'h606a;
        src4 <= 16'hdeb0;
        src5 <= 16'h2903;
        src6 <= 16'h2a3c;
        src7 <= 16'hb0bd;
        src8 <= 16'h6a5c;
        src9 <= 16'h8155;
        src10 <= 16'hb23f;
        src11 <= 16'h569e;
        src12 <= 16'hd90a;
        src13 <= 16'h5feb;
        src14 <= 16'hdee2;
        src15 <= 16'hec0c;
        src16 <= 16'h60a9;
        src17 <= 16'h1a02;
        src18 <= 16'h4596;
        src19 <= 16'hd406;
        src20 <= 16'ha9ac;
        src21 <= 16'hd327;
        src22 <= 16'hc472;
        src23 <= 16'h113d;
        src24 <= 16'h5367;
        src25 <= 16'h342f;
        src26 <= 16'he083;
        src27 <= 16'h868c;
        src28 <= 16'h9b92;
        src29 <= 16'ha2eb;
        src30 <= 16'ha506;
        src31 <= 16'h91c;
        src32 <= 16'h519a;
        src33 <= 16'h46a1;
        src34 <= 16'hbaec;
        src35 <= 16'h7c71;
        src36 <= 16'hf30a;
        src37 <= 16'h5b4b;
        src38 <= 16'h70dd;
        src39 <= 16'h56a;
        src40 <= 16'h1703;
        src41 <= 16'hca86;
        src42 <= 16'h3256;
        src43 <= 16'h4e9c;
        src44 <= 16'h219d;
        src45 <= 16'haa2b;
        src46 <= 16'hf048;
        src47 <= 16'h11ca;
        src48 <= 16'h575f;
        src49 <= 16'h2bcf;
        src50 <= 16'hcef1;
        src51 <= 16'hb926;
        src52 <= 16'hb940;
        src53 <= 16'h1869;
        src54 <= 16'hb53b;
        src55 <= 16'h2faf;
        src56 <= 16'hd7e5;
        src57 <= 16'h695;
        src58 <= 16'h9ede;
        src59 <= 16'h6e51;
        src60 <= 16'hfdc3;
        src61 <= 16'ha7e4;
        src62 <= 16'he2fb;
        src63 <= 16'h1702;
        src64 <= 16'hda2d;
        src65 <= 16'h55ae;
        src66 <= 16'h1a2;
        src67 <= 16'hcdff;
        src68 <= 16'h1f97;
        src69 <= 16'heda6;
        src70 <= 16'hd70d;
        src71 <= 16'hb2ca;
        src72 <= 16'ha48c;
        src73 <= 16'h4c46;
        src74 <= 16'hdf2e;
        src75 <= 16'h3c73;
        src76 <= 16'h1303;
        src77 <= 16'hf4f4;
        src78 <= 16'h2070;
        src79 <= 16'hc137;
        src80 <= 16'h2d7a;
        src81 <= 16'h498f;
        src82 <= 16'h30aa;
        src83 <= 16'hb8e5;
        src84 <= 16'h5f85;
        src85 <= 16'h8dc;
        src86 <= 16'hfbe9;
        src87 <= 16'ha3ae;
        src88 <= 16'h95f8;
        src89 <= 16'h2ac6;
        src90 <= 16'h436a;
        src91 <= 16'h5bbf;
        src92 <= 16'h6ae7;
        src93 <= 16'hfe12;
        src94 <= 16'h77a2;
        src95 <= 16'he707;
        src96 <= 16'h53ed;
        src97 <= 16'h820c;
        src98 <= 16'h82d6;
        src99 <= 16'hf502;
        src100 <= 16'hbfaf;
        src101 <= 16'h4188;
        src102 <= 16'h274b;
        src103 <= 16'hc5b7;
        src104 <= 16'he6fe;
        src105 <= 16'h786b;
        src106 <= 16'hc090;
        src107 <= 16'he45d;
        src108 <= 16'h4d3b;
        src109 <= 16'hd980;
        src110 <= 16'h773a;
        src111 <= 16'hd40c;
        src112 <= 16'hf4ff;
        src113 <= 16'ha832;
        src114 <= 16'h972f;
        src115 <= 16'h1c48;
        src116 <= 16'h2c97;
        src117 <= 16'h854c;
        src118 <= 16'hd01d;
        src119 <= 16'hce1c;
        src120 <= 16'hf90e;
        src121 <= 16'hb762;
        src122 <= 16'h72b2;
        src123 <= 16'h6da1;
        src124 <= 16'h7f97;
        src125 <= 16'h78e0;
        src126 <= 16'h1ef9;
        src127 <= 16'hf3bf;
        exp <= 23'h430c4d;
        #1
        src0 <= 16'h5ee;
        src1 <= 16'h9cb1;
        src2 <= 16'h3ebc;
        src3 <= 16'h552a;
        src4 <= 16'h420a;
        src5 <= 16'hfb74;
        src6 <= 16'ha939;
        src7 <= 16'h3878;
        src8 <= 16'hcd73;
        src9 <= 16'h51b7;
        src10 <= 16'hca03;
        src11 <= 16'h92ca;
        src12 <= 16'h8332;
        src13 <= 16'hb07e;
        src14 <= 16'h5689;
        src15 <= 16'h386f;
        src16 <= 16'he856;
        src17 <= 16'h2454;
        src18 <= 16'h98d1;
        src19 <= 16'he79d;
        src20 <= 16'he1c1;
        src21 <= 16'h3884;
        src22 <= 16'hf1a5;
        src23 <= 16'hbe1d;
        src24 <= 16'h361a;
        src25 <= 16'h324c;
        src26 <= 16'h14e3;
        src27 <= 16'h1b47;
        src28 <= 16'h61b4;
        src29 <= 16'hcc4e;
        src30 <= 16'h2a25;
        src31 <= 16'h6cc1;
        src32 <= 16'h111;
        src33 <= 16'ha43a;
        src34 <= 16'h963e;
        src35 <= 16'h804d;
        src36 <= 16'hcfda;
        src37 <= 16'h28fe;
        src38 <= 16'h9e99;
        src39 <= 16'h3ca0;
        src40 <= 16'h2995;
        src41 <= 16'hd56f;
        src42 <= 16'had19;
        src43 <= 16'h86dd;
        src44 <= 16'h24a8;
        src45 <= 16'h4c07;
        src46 <= 16'h996;
        src47 <= 16'he0a9;
        src48 <= 16'hd883;
        src49 <= 16'ha2ae;
        src50 <= 16'hd2c9;
        src51 <= 16'h225b;
        src52 <= 16'h4154;
        src53 <= 16'heb6d;
        src54 <= 16'h3ef1;
        src55 <= 16'hdd41;
        src56 <= 16'h8b0;
        src57 <= 16'h7a0b;
        src58 <= 16'hb7b5;
        src59 <= 16'h4dbe;
        src60 <= 16'h1923;
        src61 <= 16'h6d94;
        src62 <= 16'h91d4;
        src63 <= 16'hb4e2;
        src64 <= 16'hbff8;
        src65 <= 16'hb75f;
        src66 <= 16'h1597;
        src67 <= 16'h69f9;
        src68 <= 16'h56ae;
        src69 <= 16'he1c7;
        src70 <= 16'h597a;
        src71 <= 16'h6560;
        src72 <= 16'ha6e0;
        src73 <= 16'hab80;
        src74 <= 16'h35a0;
        src75 <= 16'hbfac;
        src76 <= 16'hd6b1;
        src77 <= 16'hf14f;
        src78 <= 16'h781e;
        src79 <= 16'h4700;
        src80 <= 16'h8547;
        src81 <= 16'hc92f;
        src82 <= 16'h83c1;
        src83 <= 16'hfd57;
        src84 <= 16'hc644;
        src85 <= 16'ha887;
        src86 <= 16'h5756;
        src87 <= 16'hc2ac;
        src88 <= 16'hbfb3;
        src89 <= 16'h82d5;
        src90 <= 16'hf316;
        src91 <= 16'h780;
        src92 <= 16'hdf23;
        src93 <= 16'h4a68;
        src94 <= 16'h11ef;
        src95 <= 16'h4719;
        src96 <= 16'h2750;
        src97 <= 16'he3c5;
        src98 <= 16'he5c6;
        src99 <= 16'h578b;
        src100 <= 16'h64b9;
        src101 <= 16'h81c;
        src102 <= 16'h460e;
        src103 <= 16'h9a7f;
        src104 <= 16'h1245;
        src105 <= 16'h83ef;
        src106 <= 16'h7a6a;
        src107 <= 16'ha9ea;
        src108 <= 16'hbd29;
        src109 <= 16'hcaf9;
        src110 <= 16'h5158;
        src111 <= 16'hfffd;
        src112 <= 16'h63d8;
        src113 <= 16'hdaab;
        src114 <= 16'h8b77;
        src115 <= 16'h22ac;
        src116 <= 16'h8b9e;
        src117 <= 16'hc5e4;
        src118 <= 16'ha295;
        src119 <= 16'h49c6;
        src120 <= 16'h7edb;
        src121 <= 16'hdb22;
        src122 <= 16'h7ca8;
        src123 <= 16'ha5c2;
        src124 <= 16'h2c84;
        src125 <= 16'ha2e5;
        src126 <= 16'hef26;
        src127 <= 16'haa5c;
        exp <= 23'h418444;
        #1
        src0 <= 16'h249c;
        src1 <= 16'h36c6;
        src2 <= 16'h1ed8;
        src3 <= 16'hf77b;
        src4 <= 16'h5ddd;
        src5 <= 16'h9f32;
        src6 <= 16'h9a41;
        src7 <= 16'h8481;
        src8 <= 16'hd540;
        src9 <= 16'ha4e6;
        src10 <= 16'h5b30;
        src11 <= 16'hb2d;
        src12 <= 16'h57b2;
        src13 <= 16'h5b17;
        src14 <= 16'h4c7a;
        src15 <= 16'hec6d;
        src16 <= 16'h1528;
        src17 <= 16'hc976;
        src18 <= 16'h25f4;
        src19 <= 16'h8861;
        src20 <= 16'hd274;
        src21 <= 16'hf29;
        src22 <= 16'h1fa3;
        src23 <= 16'hec46;
        src24 <= 16'hcc70;
        src25 <= 16'hafe5;
        src26 <= 16'h1c3f;
        src27 <= 16'h2d13;
        src28 <= 16'h8513;
        src29 <= 16'h6c36;
        src30 <= 16'h4977;
        src31 <= 16'hce86;
        src32 <= 16'hbc04;
        src33 <= 16'hc7be;
        src34 <= 16'hf748;
        src35 <= 16'hd0d6;
        src36 <= 16'hc125;
        src37 <= 16'hccf9;
        src38 <= 16'h71c7;
        src39 <= 16'h2fb5;
        src40 <= 16'he0c4;
        src41 <= 16'h382d;
        src42 <= 16'hb266;
        src43 <= 16'h8f94;
        src44 <= 16'hb87;
        src45 <= 16'h64d2;
        src46 <= 16'h6577;
        src47 <= 16'h59b6;
        src48 <= 16'h9527;
        src49 <= 16'h5e46;
        src50 <= 16'h3c67;
        src51 <= 16'hbbea;
        src52 <= 16'hf6;
        src53 <= 16'he563;
        src54 <= 16'hf2a8;
        src55 <= 16'h6bcf;
        src56 <= 16'hc5e9;
        src57 <= 16'hb106;
        src58 <= 16'h7de3;
        src59 <= 16'h4c7c;
        src60 <= 16'h4239;
        src61 <= 16'h3286;
        src62 <= 16'h9d6a;
        src63 <= 16'haee8;
        src64 <= 16'h4fd0;
        src65 <= 16'h16e7;
        src66 <= 16'h69bf;
        src67 <= 16'hdd5a;
        src68 <= 16'h143a;
        src69 <= 16'hd529;
        src70 <= 16'h1beb;
        src71 <= 16'ha5db;
        src72 <= 16'he209;
        src73 <= 16'h1dc9;
        src74 <= 16'hba08;
        src75 <= 16'h7a95;
        src76 <= 16'h23eb;
        src77 <= 16'h9dff;
        src78 <= 16'h93ab;
        src79 <= 16'h43a5;
        src80 <= 16'h899e;
        src81 <= 16'h4628;
        src82 <= 16'h31b6;
        src83 <= 16'h89ca;
        src84 <= 16'h1747;
        src85 <= 16'hb547;
        src86 <= 16'ha40;
        src87 <= 16'hba53;
        src88 <= 16'ha07e;
        src89 <= 16'h8dc1;
        src90 <= 16'h4356;
        src91 <= 16'h2bcd;
        src92 <= 16'h20ad;
        src93 <= 16'h8152;
        src94 <= 16'he68a;
        src95 <= 16'h2345;
        src96 <= 16'ha073;
        src97 <= 16'h8ff8;
        src98 <= 16'hee30;
        src99 <= 16'he8b5;
        src100 <= 16'h2667;
        src101 <= 16'h8d1a;
        src102 <= 16'hd790;
        src103 <= 16'h8995;
        src104 <= 16'h9217;
        src105 <= 16'ha7c0;
        src106 <= 16'h887e;
        src107 <= 16'h76b0;
        src108 <= 16'hcd36;
        src109 <= 16'h5126;
        src110 <= 16'hffb;
        src111 <= 16'hf8f8;
        src112 <= 16'hfdaa;
        src113 <= 16'h115c;
        src114 <= 16'hb360;
        src115 <= 16'h3259;
        src116 <= 16'h9638;
        src117 <= 16'hd9aa;
        src118 <= 16'hf3a3;
        src119 <= 16'h90de;
        src120 <= 16'he0b0;
        src121 <= 16'hdd17;
        src122 <= 16'hd89b;
        src123 <= 16'hf78b;
        src124 <= 16'h8c86;
        src125 <= 16'ha455;
        src126 <= 16'h6dc4;
        src127 <= 16'hdea1;
        exp <= 23'h41d8c9;
        #1
        src0 <= 16'h54e8;
        src1 <= 16'h6301;
        src2 <= 16'had7b;
        src3 <= 16'h5252;
        src4 <= 16'h9b16;
        src5 <= 16'h96fe;
        src6 <= 16'hf37;
        src7 <= 16'h1617;
        src8 <= 16'h4002;
        src9 <= 16'hf522;
        src10 <= 16'hedd3;
        src11 <= 16'hb3a9;
        src12 <= 16'hcae6;
        src13 <= 16'had66;
        src14 <= 16'h8a38;
        src15 <= 16'h3e38;
        src16 <= 16'h5b32;
        src17 <= 16'ha892;
        src18 <= 16'hebac;
        src19 <= 16'h5fb1;
        src20 <= 16'h9e27;
        src21 <= 16'h8677;
        src22 <= 16'hb0b9;
        src23 <= 16'h92e0;
        src24 <= 16'h673;
        src25 <= 16'ha9ef;
        src26 <= 16'h30ce;
        src27 <= 16'h7852;
        src28 <= 16'hb6eb;
        src29 <= 16'h2916;
        src30 <= 16'ha165;
        src31 <= 16'h38d9;
        src32 <= 16'h448d;
        src33 <= 16'h2255;
        src34 <= 16'h58f8;
        src35 <= 16'hf90c;
        src36 <= 16'hf422;
        src37 <= 16'hc07;
        src38 <= 16'h51e4;
        src39 <= 16'h3f94;
        src40 <= 16'h915b;
        src41 <= 16'h74c0;
        src42 <= 16'hcfa;
        src43 <= 16'hdd30;
        src44 <= 16'hd13d;
        src45 <= 16'he160;
        src46 <= 16'h2039;
        src47 <= 16'h37f3;
        src48 <= 16'he661;
        src49 <= 16'h625d;
        src50 <= 16'h8409;
        src51 <= 16'h7601;
        src52 <= 16'h5265;
        src53 <= 16'had0c;
        src54 <= 16'h1c;
        src55 <= 16'h7f3f;
        src56 <= 16'h7f1b;
        src57 <= 16'hac46;
        src58 <= 16'h5f23;
        src59 <= 16'hf400;
        src60 <= 16'ha42f;
        src61 <= 16'h83c5;
        src62 <= 16'h2c32;
        src63 <= 16'h2d0f;
        src64 <= 16'h6831;
        src65 <= 16'hd2f6;
        src66 <= 16'hd107;
        src67 <= 16'h5c6d;
        src68 <= 16'h988a;
        src69 <= 16'h2395;
        src70 <= 16'h4d29;
        src71 <= 16'h1440;
        src72 <= 16'hc6fc;
        src73 <= 16'hf772;
        src74 <= 16'h6cb;
        src75 <= 16'h2bcb;
        src76 <= 16'h9871;
        src77 <= 16'h7678;
        src78 <= 16'hc5f9;
        src79 <= 16'h881;
        src80 <= 16'h74a4;
        src81 <= 16'h3d13;
        src82 <= 16'h4c2e;
        src83 <= 16'habd;
        src84 <= 16'h68c1;
        src85 <= 16'h2533;
        src86 <= 16'h959c;
        src87 <= 16'hfe94;
        src88 <= 16'hc137;
        src89 <= 16'h7f65;
        src90 <= 16'h1710;
        src91 <= 16'hbecb;
        src92 <= 16'h4913;
        src93 <= 16'hdfa3;
        src94 <= 16'h499d;
        src95 <= 16'he845;
        src96 <= 16'h42e5;
        src97 <= 16'h6411;
        src98 <= 16'h4f50;
        src99 <= 16'hbaeb;
        src100 <= 16'h3607;
        src101 <= 16'h630c;
        src102 <= 16'hdefd;
        src103 <= 16'h38c9;
        src104 <= 16'hd30;
        src105 <= 16'h5eae;
        src106 <= 16'hcc3f;
        src107 <= 16'h84e6;
        src108 <= 16'h2a5c;
        src109 <= 16'h94c8;
        src110 <= 16'h1122;
        src111 <= 16'hf6b2;
        src112 <= 16'h3b01;
        src113 <= 16'h99af;
        src114 <= 16'h88f8;
        src115 <= 16'ha0f5;
        src116 <= 16'h5969;
        src117 <= 16'hb64d;
        src118 <= 16'h5d2;
        src119 <= 16'h9931;
        src120 <= 16'hafbc;
        src121 <= 16'h5c56;
        src122 <= 16'hf6ad;
        src123 <= 16'h56f1;
        src124 <= 16'hb78;
        src125 <= 16'h8682;
        src126 <= 16'h4feb;
        src127 <= 16'h9224;
        exp <= 23'h3c49e2;
        #1
        src0 <= 16'he644;
        src1 <= 16'h33ed;
        src2 <= 16'hb7c1;
        src3 <= 16'h3700;
        src4 <= 16'h574;
        src5 <= 16'h27a4;
        src6 <= 16'ha4fb;
        src7 <= 16'hdd41;
        src8 <= 16'h5355;
        src9 <= 16'he62;
        src10 <= 16'h204;
        src11 <= 16'h72c1;
        src12 <= 16'h680c;
        src13 <= 16'h55a9;
        src14 <= 16'he926;
        src15 <= 16'h7009;
        src16 <= 16'h92b9;
        src17 <= 16'h98ed;
        src18 <= 16'hd39b;
        src19 <= 16'he50c;
        src20 <= 16'h93d4;
        src21 <= 16'h45e1;
        src22 <= 16'h663c;
        src23 <= 16'hc96f;
        src24 <= 16'hb3a;
        src25 <= 16'hed45;
        src26 <= 16'hf186;
        src27 <= 16'h59b0;
        src28 <= 16'hf72f;
        src29 <= 16'h259d;
        src30 <= 16'ha7c8;
        src31 <= 16'h4951;
        src32 <= 16'hca0;
        src33 <= 16'h174a;
        src34 <= 16'h49f1;
        src35 <= 16'h3e73;
        src36 <= 16'h3098;
        src37 <= 16'h8e03;
        src38 <= 16'hb6a0;
        src39 <= 16'hd8b6;
        src40 <= 16'h73fb;
        src41 <= 16'h142e;
        src42 <= 16'h4f65;
        src43 <= 16'hba9a;
        src44 <= 16'h1997;
        src45 <= 16'h3760;
        src46 <= 16'hb31;
        src47 <= 16'h68b9;
        src48 <= 16'h7e2a;
        src49 <= 16'hb3c2;
        src50 <= 16'h960d;
        src51 <= 16'h4c05;
        src52 <= 16'h24cc;
        src53 <= 16'ha09e;
        src54 <= 16'h3c88;
        src55 <= 16'he4f8;
        src56 <= 16'h649c;
        src57 <= 16'h427d;
        src58 <= 16'hbda1;
        src59 <= 16'h1c0e;
        src60 <= 16'h77f2;
        src61 <= 16'hceed;
        src62 <= 16'ha717;
        src63 <= 16'hc6c8;
        src64 <= 16'h69bb;
        src65 <= 16'hd9b5;
        src66 <= 16'h3059;
        src67 <= 16'h17b;
        src68 <= 16'h5b5d;
        src69 <= 16'h3c6b;
        src70 <= 16'he952;
        src71 <= 16'hace9;
        src72 <= 16'h2249;
        src73 <= 16'h12a2;
        src74 <= 16'hc0c5;
        src75 <= 16'hc80;
        src76 <= 16'h7a19;
        src77 <= 16'hbbaa;
        src78 <= 16'h29d5;
        src79 <= 16'hc4fa;
        src80 <= 16'h53c;
        src81 <= 16'hdfb6;
        src82 <= 16'h97dc;
        src83 <= 16'h1b34;
        src84 <= 16'h4855;
        src85 <= 16'h4c91;
        src86 <= 16'h7586;
        src87 <= 16'h3284;
        src88 <= 16'h35b0;
        src89 <= 16'h7484;
        src90 <= 16'h283a;
        src91 <= 16'hde59;
        src92 <= 16'h46e3;
        src93 <= 16'hcb80;
        src94 <= 16'ha632;
        src95 <= 16'h8413;
        src96 <= 16'hb4fa;
        src97 <= 16'hf4cd;
        src98 <= 16'hd1d7;
        src99 <= 16'h60f3;
        src100 <= 16'h21b0;
        src101 <= 16'h7736;
        src102 <= 16'he8e6;
        src103 <= 16'h2496;
        src104 <= 16'ha18b;
        src105 <= 16'h9894;
        src106 <= 16'ha31;
        src107 <= 16'hf0a9;
        src108 <= 16'h8f15;
        src109 <= 16'h3f3c;
        src110 <= 16'he6c2;
        src111 <= 16'h8066;
        src112 <= 16'haa39;
        src113 <= 16'h70c1;
        src114 <= 16'h1979;
        src115 <= 16'hd79d;
        src116 <= 16'h9a6e;
        src117 <= 16'h771a;
        src118 <= 16'h6cb;
        src119 <= 16'h65c0;
        src120 <= 16'h936d;
        src121 <= 16'h277c;
        src122 <= 16'h187c;
        src123 <= 16'hae69;
        src124 <= 16'h981a;
        src125 <= 16'h6e69;
        src126 <= 16'h677d;
        src127 <= 16'hffe;
        exp <= 23'h3a6a61;
        #1
        src0 <= 16'he0ee;
        src1 <= 16'h2672;
        src2 <= 16'h8826;
        src3 <= 16'h3c52;
        src4 <= 16'h928a;
        src5 <= 16'h4ddc;
        src6 <= 16'hccf2;
        src7 <= 16'h8ece;
        src8 <= 16'h76af;
        src9 <= 16'h3812;
        src10 <= 16'hbbc5;
        src11 <= 16'h7186;
        src12 <= 16'hb66a;
        src13 <= 16'h80b4;
        src14 <= 16'h9e73;
        src15 <= 16'h5039;
        src16 <= 16'hbc33;
        src17 <= 16'haa1b;
        src18 <= 16'h851;
        src19 <= 16'h7354;
        src20 <= 16'hd193;
        src21 <= 16'hdd4b;
        src22 <= 16'hf68c;
        src23 <= 16'h5676;
        src24 <= 16'h4828;
        src25 <= 16'hcb6a;
        src26 <= 16'h855a;
        src27 <= 16'hf953;
        src28 <= 16'hf3d0;
        src29 <= 16'h5d28;
        src30 <= 16'h712b;
        src31 <= 16'hec02;
        src32 <= 16'h31ec;
        src33 <= 16'h308;
        src34 <= 16'h9329;
        src35 <= 16'hf983;
        src36 <= 16'hab98;
        src37 <= 16'hc49c;
        src38 <= 16'h2bf1;
        src39 <= 16'h4daf;
        src40 <= 16'h8969;
        src41 <= 16'h3522;
        src42 <= 16'hd4ac;
        src43 <= 16'he610;
        src44 <= 16'h2985;
        src45 <= 16'hed24;
        src46 <= 16'hf052;
        src47 <= 16'h399;
        src48 <= 16'he851;
        src49 <= 16'ha5cb;
        src50 <= 16'he3af;
        src51 <= 16'hbda0;
        src52 <= 16'he285;
        src53 <= 16'h5345;
        src54 <= 16'hc25d;
        src55 <= 16'h958;
        src56 <= 16'hb435;
        src57 <= 16'h4c3c;
        src58 <= 16'h1a21;
        src59 <= 16'h37ab;
        src60 <= 16'h5db0;
        src61 <= 16'h493a;
        src62 <= 16'h3bfa;
        src63 <= 16'h33aa;
        src64 <= 16'hd855;
        src65 <= 16'hcca0;
        src66 <= 16'h391a;
        src67 <= 16'h2357;
        src68 <= 16'hef39;
        src69 <= 16'h1988;
        src70 <= 16'h9e5;
        src71 <= 16'hc31d;
        src72 <= 16'hdc05;
        src73 <= 16'h6c3a;
        src74 <= 16'h70b8;
        src75 <= 16'h879d;
        src76 <= 16'hea0f;
        src77 <= 16'h48f1;
        src78 <= 16'h2398;
        src79 <= 16'h620e;
        src80 <= 16'h2468;
        src81 <= 16'hb054;
        src82 <= 16'h63dd;
        src83 <= 16'ha686;
        src84 <= 16'hb199;
        src85 <= 16'h4567;
        src86 <= 16'hd5ab;
        src87 <= 16'h883;
        src88 <= 16'h8ff6;
        src89 <= 16'h527e;
        src90 <= 16'h6ae0;
        src91 <= 16'hf2bb;
        src92 <= 16'hcde1;
        src93 <= 16'he30d;
        src94 <= 16'h67ee;
        src95 <= 16'h1790;
        src96 <= 16'h8214;
        src97 <= 16'he3b4;
        src98 <= 16'h190d;
        src99 <= 16'h78b7;
        src100 <= 16'h4c6b;
        src101 <= 16'hf9b0;
        src102 <= 16'h4ef3;
        src103 <= 16'ha7da;
        src104 <= 16'h244c;
        src105 <= 16'hfdcc;
        src106 <= 16'h7914;
        src107 <= 16'h58ff;
        src108 <= 16'he11f;
        src109 <= 16'h6735;
        src110 <= 16'hc698;
        src111 <= 16'h2fc7;
        src112 <= 16'he9e6;
        src113 <= 16'he9a3;
        src114 <= 16'hafa5;
        src115 <= 16'hb159;
        src116 <= 16'h17da;
        src117 <= 16'hca3c;
        src118 <= 16'hc357;
        src119 <= 16'h919c;
        src120 <= 16'he557;
        src121 <= 16'hf9a6;
        src122 <= 16'ha376;
        src123 <= 16'h121c;
        src124 <= 16'hf0e0;
        src125 <= 16'hc1cc;
        src126 <= 16'hba8a;
        src127 <= 16'heef0;
        exp <= 23'h45a9d1;
        #1
        src0 <= 16'hc023;
        src1 <= 16'h448a;
        src2 <= 16'h50c9;
        src3 <= 16'hd4cc;
        src4 <= 16'h1063;
        src5 <= 16'h2f82;
        src6 <= 16'h425a;
        src7 <= 16'hd7c3;
        src8 <= 16'h1269;
        src9 <= 16'hce08;
        src10 <= 16'h9b14;
        src11 <= 16'h4e30;
        src12 <= 16'hce36;
        src13 <= 16'h7778;
        src14 <= 16'hd48e;
        src15 <= 16'h72a1;
        src16 <= 16'hfed0;
        src17 <= 16'h84e2;
        src18 <= 16'hd22e;
        src19 <= 16'h5817;
        src20 <= 16'h3af4;
        src21 <= 16'hcf94;
        src22 <= 16'h2e75;
        src23 <= 16'hbbfc;
        src24 <= 16'hbe38;
        src25 <= 16'h3bac;
        src26 <= 16'hb08a;
        src27 <= 16'had7b;
        src28 <= 16'hef30;
        src29 <= 16'h6dbb;
        src30 <= 16'h4f93;
        src31 <= 16'h17c5;
        src32 <= 16'ha3a;
        src33 <= 16'h15fe;
        src34 <= 16'h13de;
        src35 <= 16'h1216;
        src36 <= 16'h32e6;
        src37 <= 16'ha3e4;
        src38 <= 16'h7af3;
        src39 <= 16'hbbb4;
        src40 <= 16'h8a16;
        src41 <= 16'hf399;
        src42 <= 16'h722f;
        src43 <= 16'hb9b9;
        src44 <= 16'hed30;
        src45 <= 16'hcb9d;
        src46 <= 16'hb317;
        src47 <= 16'h7c2e;
        src48 <= 16'h2cac;
        src49 <= 16'hed66;
        src50 <= 16'hd565;
        src51 <= 16'h54d9;
        src52 <= 16'h55c;
        src53 <= 16'h8cf9;
        src54 <= 16'h151a;
        src55 <= 16'h520a;
        src56 <= 16'ha183;
        src57 <= 16'ha129;
        src58 <= 16'h93b;
        src59 <= 16'h2d3b;
        src60 <= 16'he0c8;
        src61 <= 16'h65a1;
        src62 <= 16'h18c0;
        src63 <= 16'h7823;
        src64 <= 16'hfd3b;
        src65 <= 16'h846a;
        src66 <= 16'hab55;
        src67 <= 16'ha222;
        src68 <= 16'hf67c;
        src69 <= 16'ha4d5;
        src70 <= 16'hab7b;
        src71 <= 16'hf563;
        src72 <= 16'hceec;
        src73 <= 16'ha989;
        src74 <= 16'hc872;
        src75 <= 16'hfb85;
        src76 <= 16'h5704;
        src77 <= 16'h46e6;
        src78 <= 16'h382f;
        src79 <= 16'h85c2;
        src80 <= 16'hae05;
        src81 <= 16'h6b86;
        src82 <= 16'h9351;
        src83 <= 16'hf014;
        src84 <= 16'h2d9;
        src85 <= 16'hc2c3;
        src86 <= 16'h9295;
        src87 <= 16'h46b0;
        src88 <= 16'hfe40;
        src89 <= 16'he89f;
        src90 <= 16'h1706;
        src91 <= 16'h5d07;
        src92 <= 16'h9439;
        src93 <= 16'h2c4a;
        src94 <= 16'he028;
        src95 <= 16'h64e4;
        src96 <= 16'h6cff;
        src97 <= 16'h93f0;
        src98 <= 16'h213d;
        src99 <= 16'he26e;
        src100 <= 16'h5b25;
        src101 <= 16'h3c25;
        src102 <= 16'h6c53;
        src103 <= 16'hc2a9;
        src104 <= 16'h3ce3;
        src105 <= 16'h4101;
        src106 <= 16'h8433;
        src107 <= 16'h5099;
        src108 <= 16'hf227;
        src109 <= 16'hdbbd;
        src110 <= 16'h370a;
        src111 <= 16'h6ac5;
        src112 <= 16'hfef6;
        src113 <= 16'hcc58;
        src114 <= 16'h6d21;
        src115 <= 16'h382e;
        src116 <= 16'hddb0;
        src117 <= 16'h6982;
        src118 <= 16'hceb0;
        src119 <= 16'h9c8c;
        src120 <= 16'he001;
        src121 <= 16'h9afa;
        src122 <= 16'hebc;
        src123 <= 16'h8bbb;
        src124 <= 16'h6525;
        src125 <= 16'hab93;
        src126 <= 16'hbc7b;
        src127 <= 16'h8363;
        exp <= 23'h4363a3;
        #1
        src0 <= 16'h766b;
        src1 <= 16'he522;
        src2 <= 16'h7980;
        src3 <= 16'h4ac8;
        src4 <= 16'h819a;
        src5 <= 16'hddbf;
        src6 <= 16'he593;
        src7 <= 16'hab81;
        src8 <= 16'h7003;
        src9 <= 16'h21fa;
        src10 <= 16'hf545;
        src11 <= 16'hf87b;
        src12 <= 16'h2476;
        src13 <= 16'h6dc1;
        src14 <= 16'hec6;
        src15 <= 16'h368d;
        src16 <= 16'h27f8;
        src17 <= 16'h7a40;
        src18 <= 16'hfc2;
        src19 <= 16'h2a31;
        src20 <= 16'h8e7e;
        src21 <= 16'hb105;
        src22 <= 16'h3ea4;
        src23 <= 16'hc2c1;
        src24 <= 16'hf315;
        src25 <= 16'h77e9;
        src26 <= 16'ha918;
        src27 <= 16'he5c2;
        src28 <= 16'he47c;
        src29 <= 16'h1ecd;
        src30 <= 16'hfa12;
        src31 <= 16'h38ae;
        src32 <= 16'h5a66;
        src33 <= 16'h9c3b;
        src34 <= 16'h2a1;
        src35 <= 16'h5939;
        src36 <= 16'h3075;
        src37 <= 16'hd1ea;
        src38 <= 16'h483c;
        src39 <= 16'h2077;
        src40 <= 16'heaf4;
        src41 <= 16'had8f;
        src42 <= 16'hb06e;
        src43 <= 16'hda4e;
        src44 <= 16'h4b02;
        src45 <= 16'ha769;
        src46 <= 16'hecb0;
        src47 <= 16'h565d;
        src48 <= 16'hca40;
        src49 <= 16'hc9de;
        src50 <= 16'h3308;
        src51 <= 16'h7807;
        src52 <= 16'h1df4;
        src53 <= 16'h7570;
        src54 <= 16'hc84;
        src55 <= 16'hb958;
        src56 <= 16'hdc93;
        src57 <= 16'h4f6e;
        src58 <= 16'h48c0;
        src59 <= 16'h6986;
        src60 <= 16'hfc5b;
        src61 <= 16'h28d4;
        src62 <= 16'hc932;
        src63 <= 16'h3504;
        src64 <= 16'hf3ed;
        src65 <= 16'h14b3;
        src66 <= 16'h36b8;
        src67 <= 16'hff93;
        src68 <= 16'hd47d;
        src69 <= 16'haa7b;
        src70 <= 16'hf8c8;
        src71 <= 16'h218b;
        src72 <= 16'hb272;
        src73 <= 16'h50b6;
        src74 <= 16'h8fa0;
        src75 <= 16'hf7c8;
        src76 <= 16'hcc37;
        src77 <= 16'h1189;
        src78 <= 16'h7109;
        src79 <= 16'h2564;
        src80 <= 16'hb5ea;
        src81 <= 16'h165c;
        src82 <= 16'hedfd;
        src83 <= 16'h23a4;
        src84 <= 16'h5613;
        src85 <= 16'h7e21;
        src86 <= 16'ha280;
        src87 <= 16'h7eff;
        src88 <= 16'h4925;
        src89 <= 16'h2ac3;
        src90 <= 16'h9376;
        src91 <= 16'h16bb;
        src92 <= 16'hbfe2;
        src93 <= 16'he9cd;
        src94 <= 16'h3e88;
        src95 <= 16'h5d35;
        src96 <= 16'he1ad;
        src97 <= 16'hdf8e;
        src98 <= 16'h6365;
        src99 <= 16'he71b;
        src100 <= 16'h24de;
        src101 <= 16'hca38;
        src102 <= 16'h12cb;
        src103 <= 16'h75c8;
        src104 <= 16'he116;
        src105 <= 16'h5577;
        src106 <= 16'h6e2b;
        src107 <= 16'h835d;
        src108 <= 16'h3098;
        src109 <= 16'hb6d4;
        src110 <= 16'hde0f;
        src111 <= 16'h6e36;
        src112 <= 16'h3580;
        src113 <= 16'hfd3a;
        src114 <= 16'h2119;
        src115 <= 16'head2;
        src116 <= 16'h2448;
        src117 <= 16'h2871;
        src118 <= 16'h3c19;
        src119 <= 16'hac33;
        src120 <= 16'hf42f;
        src121 <= 16'h28e6;
        src122 <= 16'hb984;
        src123 <= 16'h4db4;
        src124 <= 16'hfcb2;
        src125 <= 16'h45f3;
        src126 <= 16'he768;
        src127 <= 16'hd2b3;
        exp <= 23'h41e6cd;
        #1
        src0 <= 16'h30cf;
        src1 <= 16'h778e;
        src2 <= 16'heeac;
        src3 <= 16'h84b3;
        src4 <= 16'h3e03;
        src5 <= 16'h6c0;
        src6 <= 16'hf7b5;
        src7 <= 16'hd91c;
        src8 <= 16'h54a8;
        src9 <= 16'hb899;
        src10 <= 16'h5488;
        src11 <= 16'he335;
        src12 <= 16'h2341;
        src13 <= 16'h9103;
        src14 <= 16'ha373;
        src15 <= 16'hd687;
        src16 <= 16'h8d92;
        src17 <= 16'haca;
        src18 <= 16'h17c9;
        src19 <= 16'h9bad;
        src20 <= 16'hc46b;
        src21 <= 16'h409c;
        src22 <= 16'h78ea;
        src23 <= 16'hfc4d;
        src24 <= 16'h7dea;
        src25 <= 16'h9aa0;
        src26 <= 16'h1e29;
        src27 <= 16'h34ae;
        src28 <= 16'h543c;
        src29 <= 16'h9062;
        src30 <= 16'hfb74;
        src31 <= 16'hdd28;
        src32 <= 16'h474c;
        src33 <= 16'hea41;
        src34 <= 16'hc2ed;
        src35 <= 16'h3b5a;
        src36 <= 16'h6a05;
        src37 <= 16'h3e6d;
        src38 <= 16'h10cf;
        src39 <= 16'h784;
        src40 <= 16'hb694;
        src41 <= 16'h4253;
        src42 <= 16'he455;
        src43 <= 16'h9905;
        src44 <= 16'hb8a3;
        src45 <= 16'hbb4b;
        src46 <= 16'h9e3d;
        src47 <= 16'hda08;
        src48 <= 16'h96a6;
        src49 <= 16'h31c2;
        src50 <= 16'h6827;
        src51 <= 16'hcfd1;
        src52 <= 16'h70d2;
        src53 <= 16'hb5d3;
        src54 <= 16'hde73;
        src55 <= 16'ha30b;
        src56 <= 16'h39d3;
        src57 <= 16'hb05;
        src58 <= 16'h9336;
        src59 <= 16'h2d5d;
        src60 <= 16'h650f;
        src61 <= 16'hfa15;
        src62 <= 16'h8079;
        src63 <= 16'h5a05;
        src64 <= 16'h9109;
        src65 <= 16'hd31d;
        src66 <= 16'hee05;
        src67 <= 16'ha0b1;
        src68 <= 16'hffb9;
        src69 <= 16'heb54;
        src70 <= 16'h8a7d;
        src71 <= 16'h3a30;
        src72 <= 16'h740c;
        src73 <= 16'h25b6;
        src74 <= 16'h9a58;
        src75 <= 16'h1497;
        src76 <= 16'ha2d1;
        src77 <= 16'h4a2b;
        src78 <= 16'h11e4;
        src79 <= 16'h645f;
        src80 <= 16'h538c;
        src81 <= 16'h66e2;
        src82 <= 16'h4f38;
        src83 <= 16'h26fa;
        src84 <= 16'hbccb;
        src85 <= 16'hce8;
        src86 <= 16'hb846;
        src87 <= 16'h8903;
        src88 <= 16'hbdf6;
        src89 <= 16'hd235;
        src90 <= 16'h23a5;
        src91 <= 16'h2e8c;
        src92 <= 16'h68f2;
        src93 <= 16'h321c;
        src94 <= 16'h2d88;
        src95 <= 16'ha804;
        src96 <= 16'hce92;
        src97 <= 16'hb7e8;
        src98 <= 16'h6ca8;
        src99 <= 16'hd295;
        src100 <= 16'h7f6c;
        src101 <= 16'h5bf7;
        src102 <= 16'h8e2c;
        src103 <= 16'h6473;
        src104 <= 16'h22f6;
        src105 <= 16'ha575;
        src106 <= 16'had27;
        src107 <= 16'hf77c;
        src108 <= 16'hd17b;
        src109 <= 16'h13ae;
        src110 <= 16'hffb1;
        src111 <= 16'hb8e4;
        src112 <= 16'h2c4;
        src113 <= 16'h10ca;
        src114 <= 16'hc322;
        src115 <= 16'h972b;
        src116 <= 16'h2302;
        src117 <= 16'hb3ac;
        src118 <= 16'hca75;
        src119 <= 16'h32af;
        src120 <= 16'ha5d3;
        src121 <= 16'h913e;
        src122 <= 16'h142c;
        src123 <= 16'h9b7e;
        src124 <= 16'he801;
        src125 <= 16'h867c;
        src126 <= 16'he242;
        src127 <= 16'h6231;
        exp <= 23'h4124c9;
        #1
        src0 <= 16'hee43;
        src1 <= 16'h72e1;
        src2 <= 16'h7fe5;
        src3 <= 16'h41bf;
        src4 <= 16'hef53;
        src5 <= 16'h7784;
        src6 <= 16'hda4f;
        src7 <= 16'heba4;
        src8 <= 16'h7ef;
        src9 <= 16'hdb58;
        src10 <= 16'h3265;
        src11 <= 16'ha0b2;
        src12 <= 16'h2a93;
        src13 <= 16'hb44e;
        src14 <= 16'hf0b9;
        src15 <= 16'h6840;
        src16 <= 16'h359f;
        src17 <= 16'h1b17;
        src18 <= 16'h94f2;
        src19 <= 16'h8408;
        src20 <= 16'hd835;
        src21 <= 16'hf88c;
        src22 <= 16'h830b;
        src23 <= 16'hb269;
        src24 <= 16'hf784;
        src25 <= 16'hfac8;
        src26 <= 16'h2db3;
        src27 <= 16'he112;
        src28 <= 16'hde29;
        src29 <= 16'h3eb2;
        src30 <= 16'h63;
        src31 <= 16'h1e04;
        src32 <= 16'hbe27;
        src33 <= 16'hce81;
        src34 <= 16'hecf8;
        src35 <= 16'h5bc7;
        src36 <= 16'h5237;
        src37 <= 16'hdfe1;
        src38 <= 16'hbff0;
        src39 <= 16'h3011;
        src40 <= 16'h119f;
        src41 <= 16'h8353;
        src42 <= 16'h449f;
        src43 <= 16'h2450;
        src44 <= 16'h6049;
        src45 <= 16'hc166;
        src46 <= 16'h3ada;
        src47 <= 16'h899a;
        src48 <= 16'hff0;
        src49 <= 16'ha131;
        src50 <= 16'h13ec;
        src51 <= 16'h2678;
        src52 <= 16'hdaa9;
        src53 <= 16'hedb5;
        src54 <= 16'h179e;
        src55 <= 16'hef21;
        src56 <= 16'hadce;
        src57 <= 16'h5c22;
        src58 <= 16'hd33e;
        src59 <= 16'h6584;
        src60 <= 16'h5023;
        src61 <= 16'h23f5;
        src62 <= 16'he03b;
        src63 <= 16'h63ec;
        src64 <= 16'h6195;
        src65 <= 16'hd6b3;
        src66 <= 16'h944f;
        src67 <= 16'h34d;
        src68 <= 16'h98e3;
        src69 <= 16'h10af;
        src70 <= 16'h2cc2;
        src71 <= 16'h8bdc;
        src72 <= 16'h707d;
        src73 <= 16'h11e1;
        src74 <= 16'h72e7;
        src75 <= 16'hfa85;
        src76 <= 16'hb127;
        src77 <= 16'hcc71;
        src78 <= 16'ha6b8;
        src79 <= 16'h50d0;
        src80 <= 16'h29df;
        src81 <= 16'h83c;
        src82 <= 16'h7b;
        src83 <= 16'h934e;
        src84 <= 16'h5d6;
        src85 <= 16'h4e3a;
        src86 <= 16'h586e;
        src87 <= 16'h378f;
        src88 <= 16'h5420;
        src89 <= 16'h6048;
        src90 <= 16'h45b0;
        src91 <= 16'h4f28;
        src92 <= 16'h12f2;
        src93 <= 16'h3cbe;
        src94 <= 16'h90fa;
        src95 <= 16'hfad6;
        src96 <= 16'hbc2b;
        src97 <= 16'hc632;
        src98 <= 16'hdd4f;
        src99 <= 16'h2be3;
        src100 <= 16'h4cb9;
        src101 <= 16'h99c0;
        src102 <= 16'h78fd;
        src103 <= 16'hd925;
        src104 <= 16'hbcc7;
        src105 <= 16'h1b85;
        src106 <= 16'h22b9;
        src107 <= 16'h2a19;
        src108 <= 16'h7add;
        src109 <= 16'h18b6;
        src110 <= 16'he2e9;
        src111 <= 16'h5b0;
        src112 <= 16'h11d6;
        src113 <= 16'hd48a;
        src114 <= 16'h9e8b;
        src115 <= 16'h40d4;
        src116 <= 16'h8cef;
        src117 <= 16'h457f;
        src118 <= 16'hb0b7;
        src119 <= 16'hdfc4;
        src120 <= 16'h7f8a;
        src121 <= 16'h97cb;
        src122 <= 16'ha76b;
        src123 <= 16'h680e;
        src124 <= 16'hc3e5;
        src125 <= 16'he034;
        src126 <= 16'ha04d;
        src127 <= 16'h69af;
        exp <= 23'h3e43c7;
        #1
        src0 <= 16'haff5;
        src1 <= 16'he47b;
        src2 <= 16'h507;
        src3 <= 16'hc382;
        src4 <= 16'hca09;
        src5 <= 16'hd0f7;
        src6 <= 16'ha3b3;
        src7 <= 16'h7905;
        src8 <= 16'he675;
        src9 <= 16'h7e0f;
        src10 <= 16'hfeed;
        src11 <= 16'hd26c;
        src12 <= 16'hd68c;
        src13 <= 16'h979b;
        src14 <= 16'hc932;
        src15 <= 16'h8155;
        src16 <= 16'h1344;
        src17 <= 16'h4e24;
        src18 <= 16'h9ad9;
        src19 <= 16'h85a;
        src20 <= 16'h93d7;
        src21 <= 16'h41da;
        src22 <= 16'h641;
        src23 <= 16'h392c;
        src24 <= 16'h6f3b;
        src25 <= 16'h82ed;
        src26 <= 16'h148d;
        src27 <= 16'hfe2a;
        src28 <= 16'hf891;
        src29 <= 16'h9066;
        src30 <= 16'h3255;
        src31 <= 16'h7b17;
        src32 <= 16'h59dc;
        src33 <= 16'h990e;
        src34 <= 16'h1716;
        src35 <= 16'hc722;
        src36 <= 16'h8bfa;
        src37 <= 16'h5d14;
        src38 <= 16'hc3e1;
        src39 <= 16'hc066;
        src40 <= 16'h5053;
        src41 <= 16'h782;
        src42 <= 16'hd9c5;
        src43 <= 16'ha168;
        src44 <= 16'h463f;
        src45 <= 16'hbeb3;
        src46 <= 16'h7f24;
        src47 <= 16'h25bf;
        src48 <= 16'hdc15;
        src49 <= 16'hfb49;
        src50 <= 16'h77e4;
        src51 <= 16'h619a;
        src52 <= 16'ha4b;
        src53 <= 16'h1ea3;
        src54 <= 16'h4ad4;
        src55 <= 16'h140c;
        src56 <= 16'h2c09;
        src57 <= 16'h1faa;
        src58 <= 16'h387;
        src59 <= 16'h4deb;
        src60 <= 16'ha6ac;
        src61 <= 16'h5686;
        src62 <= 16'h6fa9;
        src63 <= 16'h2324;
        src64 <= 16'h6e4;
        src65 <= 16'h798e;
        src66 <= 16'h5179;
        src67 <= 16'hffe;
        src68 <= 16'h2b2;
        src69 <= 16'h44ef;
        src70 <= 16'h79f2;
        src71 <= 16'h1ea;
        src72 <= 16'h51de;
        src73 <= 16'h264f;
        src74 <= 16'hac25;
        src75 <= 16'hf693;
        src76 <= 16'h4824;
        src77 <= 16'h3349;
        src78 <= 16'hfffc;
        src79 <= 16'h12e4;
        src80 <= 16'h6971;
        src81 <= 16'hfbba;
        src82 <= 16'hb76b;
        src83 <= 16'h393e;
        src84 <= 16'h21a4;
        src85 <= 16'h9942;
        src86 <= 16'h4aba;
        src87 <= 16'h8bd;
        src88 <= 16'hb9ac;
        src89 <= 16'h68ab;
        src90 <= 16'hd980;
        src91 <= 16'h906a;
        src92 <= 16'h54cf;
        src93 <= 16'hf60f;
        src94 <= 16'h29c6;
        src95 <= 16'h78fd;
        src96 <= 16'hba82;
        src97 <= 16'hfc6a;
        src98 <= 16'hc53b;
        src99 <= 16'h50de;
        src100 <= 16'h3dc;
        src101 <= 16'h592f;
        src102 <= 16'h2a39;
        src103 <= 16'h55f2;
        src104 <= 16'ha798;
        src105 <= 16'hd253;
        src106 <= 16'he6b1;
        src107 <= 16'h1b28;
        src108 <= 16'hc716;
        src109 <= 16'h34b8;
        src110 <= 16'h5817;
        src111 <= 16'h4d14;
        src112 <= 16'h9a9e;
        src113 <= 16'h6cb3;
        src114 <= 16'hb465;
        src115 <= 16'h248a;
        src116 <= 16'hc75b;
        src117 <= 16'hd0cc;
        src118 <= 16'h9915;
        src119 <= 16'h2612;
        src120 <= 16'h2813;
        src121 <= 16'h56a0;
        src122 <= 16'hd947;
        src123 <= 16'h508a;
        src124 <= 16'ha1d9;
        src125 <= 16'h259;
        src126 <= 16'hacbc;
        src127 <= 16'he7f3;
        exp <= 23'h3b85e9;
        #1
        src0 <= 16'h5dd0;
        src1 <= 16'h1c66;
        src2 <= 16'he049;
        src3 <= 16'h81b9;
        src4 <= 16'hf6b2;
        src5 <= 16'hff52;
        src6 <= 16'h4510;
        src7 <= 16'hbcc0;
        src8 <= 16'h3d4f;
        src9 <= 16'hce0a;
        src10 <= 16'h91fb;
        src11 <= 16'h70a5;
        src12 <= 16'hd505;
        src13 <= 16'hd7d4;
        src14 <= 16'hed33;
        src15 <= 16'hb5ff;
        src16 <= 16'h2a;
        src17 <= 16'h1a9a;
        src18 <= 16'hd967;
        src19 <= 16'ha570;
        src20 <= 16'hb4bf;
        src21 <= 16'hc67a;
        src22 <= 16'hbe9b;
        src23 <= 16'h4152;
        src24 <= 16'h5fc6;
        src25 <= 16'h7e92;
        src26 <= 16'he842;
        src27 <= 16'h741f;
        src28 <= 16'ha697;
        src29 <= 16'hf8ff;
        src30 <= 16'h3fe7;
        src31 <= 16'h7a68;
        src32 <= 16'hb6f1;
        src33 <= 16'h3efd;
        src34 <= 16'h428d;
        src35 <= 16'hda0e;
        src36 <= 16'h4146;
        src37 <= 16'h423;
        src38 <= 16'h9739;
        src39 <= 16'h11ec;
        src40 <= 16'hf894;
        src41 <= 16'h3dc4;
        src42 <= 16'h9bee;
        src43 <= 16'h4aab;
        src44 <= 16'h5d7f;
        src45 <= 16'h7613;
        src46 <= 16'h8698;
        src47 <= 16'h9f37;
        src48 <= 16'hff07;
        src49 <= 16'h5571;
        src50 <= 16'h771a;
        src51 <= 16'h32d1;
        src52 <= 16'hbf3d;
        src53 <= 16'h1125;
        src54 <= 16'h6ff3;
        src55 <= 16'hfe0d;
        src56 <= 16'h3167;
        src57 <= 16'h3e7b;
        src58 <= 16'h89af;
        src59 <= 16'h162d;
        src60 <= 16'h56ae;
        src61 <= 16'h7c02;
        src62 <= 16'h1805;
        src63 <= 16'ha6e7;
        src64 <= 16'h6409;
        src65 <= 16'hc0da;
        src66 <= 16'hebcb;
        src67 <= 16'h2f39;
        src68 <= 16'h77bb;
        src69 <= 16'hb432;
        src70 <= 16'hdbc2;
        src71 <= 16'h59b6;
        src72 <= 16'h60bb;
        src73 <= 16'h13e4;
        src74 <= 16'h5808;
        src75 <= 16'h6de2;
        src76 <= 16'h8e20;
        src77 <= 16'had6f;
        src78 <= 16'hc4d5;
        src79 <= 16'h362b;
        src80 <= 16'he2f8;
        src81 <= 16'h651e;
        src82 <= 16'h4389;
        src83 <= 16'h88d;
        src84 <= 16'h7097;
        src85 <= 16'h4107;
        src86 <= 16'hb8ce;
        src87 <= 16'hcd16;
        src88 <= 16'h5374;
        src89 <= 16'h11a;
        src90 <= 16'hab7d;
        src91 <= 16'h30e4;
        src92 <= 16'h3cc3;
        src93 <= 16'h2c1e;
        src94 <= 16'hbc8a;
        src95 <= 16'hd120;
        src96 <= 16'h223b;
        src97 <= 16'h1573;
        src98 <= 16'hc506;
        src99 <= 16'h2175;
        src100 <= 16'h3726;
        src101 <= 16'hb49a;
        src102 <= 16'h1e3b;
        src103 <= 16'h14a3;
        src104 <= 16'hef7;
        src105 <= 16'hae54;
        src106 <= 16'h6674;
        src107 <= 16'hc209;
        src108 <= 16'h8d2a;
        src109 <= 16'hfe95;
        src110 <= 16'h1c7a;
        src111 <= 16'hc4b1;
        src112 <= 16'h9501;
        src113 <= 16'h5ea5;
        src114 <= 16'h4368;
        src115 <= 16'hab65;
        src116 <= 16'h7b;
        src117 <= 16'h9c71;
        src118 <= 16'h16ac;
        src119 <= 16'h1f8d;
        src120 <= 16'hc37;
        src121 <= 16'hcf18;
        src122 <= 16'ha41d;
        src123 <= 16'h80f;
        src124 <= 16'h6387;
        src125 <= 16'hba7a;
        src126 <= 16'ha935;
        src127 <= 16'h36e0;
        exp <= 23'h3ca125;
        #1
        src0 <= 16'h777e;
        src1 <= 16'h2a64;
        src2 <= 16'h7e1f;
        src3 <= 16'h4e7a;
        src4 <= 16'h96;
        src5 <= 16'h957c;
        src6 <= 16'h2e37;
        src7 <= 16'h27cb;
        src8 <= 16'hb54a;
        src9 <= 16'h4e66;
        src10 <= 16'h5e00;
        src11 <= 16'h9e7e;
        src12 <= 16'hb872;
        src13 <= 16'haba8;
        src14 <= 16'haa96;
        src15 <= 16'h4013;
        src16 <= 16'hef97;
        src17 <= 16'h9764;
        src18 <= 16'h3e51;
        src19 <= 16'h97b9;
        src20 <= 16'h99c0;
        src21 <= 16'h2e75;
        src22 <= 16'h17b;
        src23 <= 16'hdf50;
        src24 <= 16'h421a;
        src25 <= 16'h4eca;
        src26 <= 16'habb5;
        src27 <= 16'h3e1c;
        src28 <= 16'hf0e4;
        src29 <= 16'h3018;
        src30 <= 16'hfb54;
        src31 <= 16'hfe0;
        src32 <= 16'h47e2;
        src33 <= 16'h789d;
        src34 <= 16'ha908;
        src35 <= 16'hf5c3;
        src36 <= 16'hc436;
        src37 <= 16'h4259;
        src38 <= 16'h5b38;
        src39 <= 16'h1ea1;
        src40 <= 16'hcbd1;
        src41 <= 16'hd9ef;
        src42 <= 16'h4830;
        src43 <= 16'h14dc;
        src44 <= 16'h83df;
        src45 <= 16'h52e7;
        src46 <= 16'h8a6c;
        src47 <= 16'he2ae;
        src48 <= 16'hf284;
        src49 <= 16'h3d2e;
        src50 <= 16'hc1a8;
        src51 <= 16'h8739;
        src52 <= 16'hf4f0;
        src53 <= 16'h9827;
        src54 <= 16'h6aea;
        src55 <= 16'h527;
        src56 <= 16'h8c92;
        src57 <= 16'h2604;
        src58 <= 16'h1931;
        src59 <= 16'h1726;
        src60 <= 16'h6ce3;
        src61 <= 16'hd360;
        src62 <= 16'hd4a5;
        src63 <= 16'h4960;
        src64 <= 16'h4a4b;
        src65 <= 16'h923;
        src66 <= 16'h8f9d;
        src67 <= 16'hf51d;
        src68 <= 16'h4258;
        src69 <= 16'had80;
        src70 <= 16'h8af9;
        src71 <= 16'he418;
        src72 <= 16'h4a55;
        src73 <= 16'hd56a;
        src74 <= 16'h178a;
        src75 <= 16'h98c5;
        src76 <= 16'hfa99;
        src77 <= 16'hf814;
        src78 <= 16'hf858;
        src79 <= 16'h6e0c;
        src80 <= 16'hab98;
        src81 <= 16'h25a5;
        src82 <= 16'h542b;
        src83 <= 16'hb715;
        src84 <= 16'h3251;
        src85 <= 16'h6d3a;
        src86 <= 16'h809e;
        src87 <= 16'h499d;
        src88 <= 16'h1a20;
        src89 <= 16'ha609;
        src90 <= 16'h819b;
        src91 <= 16'hea7a;
        src92 <= 16'hbfba;
        src93 <= 16'h2e1;
        src94 <= 16'h608d;
        src95 <= 16'h5e82;
        src96 <= 16'h6ea9;
        src97 <= 16'h1bbd;
        src98 <= 16'h5963;
        src99 <= 16'hacf7;
        src100 <= 16'hcdaa;
        src101 <= 16'h589a;
        src102 <= 16'h857e;
        src103 <= 16'h179b;
        src104 <= 16'h1617;
        src105 <= 16'hf1d2;
        src106 <= 16'hb963;
        src107 <= 16'ha4b2;
        src108 <= 16'hacab;
        src109 <= 16'he41a;
        src110 <= 16'hcc8e;
        src111 <= 16'hd78e;
        src112 <= 16'h3c55;
        src113 <= 16'h6a1d;
        src114 <= 16'hed76;
        src115 <= 16'ha4e6;
        src116 <= 16'h6eaa;
        src117 <= 16'h2e55;
        src118 <= 16'h2704;
        src119 <= 16'hf1ce;
        src120 <= 16'h872d;
        src121 <= 16'h18ae;
        src122 <= 16'h3010;
        src123 <= 16'hcf47;
        src124 <= 16'hda7b;
        src125 <= 16'h83ee;
        src126 <= 16'h334d;
        src127 <= 16'h914f;
        exp <= 23'h3f27e5;
        #1
        src0 <= 16'hc262;
        src1 <= 16'h6cd3;
        src2 <= 16'h1de;
        src3 <= 16'h44fc;
        src4 <= 16'hdde1;
        src5 <= 16'hdf6c;
        src6 <= 16'ha2d9;
        src7 <= 16'h296d;
        src8 <= 16'h5609;
        src9 <= 16'h2ca3;
        src10 <= 16'heb0a;
        src11 <= 16'h21a3;
        src12 <= 16'h3ef5;
        src13 <= 16'h1168;
        src14 <= 16'ha025;
        src15 <= 16'h1adc;
        src16 <= 16'h541;
        src17 <= 16'ha633;
        src18 <= 16'hd86e;
        src19 <= 16'hb7a;
        src20 <= 16'ha0a3;
        src21 <= 16'h9316;
        src22 <= 16'hb21c;
        src23 <= 16'hf10a;
        src24 <= 16'hb35f;
        src25 <= 16'hf0c6;
        src26 <= 16'h7bd9;
        src27 <= 16'h439f;
        src28 <= 16'h9ae6;
        src29 <= 16'h9687;
        src30 <= 16'hb59f;
        src31 <= 16'h1180;
        src32 <= 16'h40cf;
        src33 <= 16'h6d82;
        src34 <= 16'hd6f1;
        src35 <= 16'hb3f;
        src36 <= 16'h8a63;
        src37 <= 16'h3682;
        src38 <= 16'hbf2c;
        src39 <= 16'h77c9;
        src40 <= 16'h7510;
        src41 <= 16'h643b;
        src42 <= 16'h5a89;
        src43 <= 16'h3b39;
        src44 <= 16'h892;
        src45 <= 16'h7994;
        src46 <= 16'hc378;
        src47 <= 16'h185a;
        src48 <= 16'h12ee;
        src49 <= 16'h642c;
        src50 <= 16'h59d;
        src51 <= 16'h98fb;
        src52 <= 16'hd13b;
        src53 <= 16'h6f58;
        src54 <= 16'h9624;
        src55 <= 16'h46c9;
        src56 <= 16'hb9a5;
        src57 <= 16'hbe3d;
        src58 <= 16'h6df1;
        src59 <= 16'h67bc;
        src60 <= 16'he5f6;
        src61 <= 16'h6848;
        src62 <= 16'h2a7d;
        src63 <= 16'h8593;
        src64 <= 16'h6311;
        src65 <= 16'hb736;
        src66 <= 16'h3dd3;
        src67 <= 16'hf713;
        src68 <= 16'h16ac;
        src69 <= 16'h9297;
        src70 <= 16'hf9e9;
        src71 <= 16'h9b33;
        src72 <= 16'h142e;
        src73 <= 16'hcc22;
        src74 <= 16'h96ff;
        src75 <= 16'hbb80;
        src76 <= 16'h26db;
        src77 <= 16'h8c6;
        src78 <= 16'hc085;
        src79 <= 16'hfb4;
        src80 <= 16'h5a28;
        src81 <= 16'ha054;
        src82 <= 16'hd8c0;
        src83 <= 16'h12d0;
        src84 <= 16'h3a06;
        src85 <= 16'h49a3;
        src86 <= 16'h8411;
        src87 <= 16'h9e24;
        src88 <= 16'h7a5a;
        src89 <= 16'he343;
        src90 <= 16'he294;
        src91 <= 16'hb61d;
        src92 <= 16'h28ff;
        src93 <= 16'ha385;
        src94 <= 16'h5296;
        src95 <= 16'hcedc;
        src96 <= 16'h72e8;
        src97 <= 16'h9b1c;
        src98 <= 16'h37ae;
        src99 <= 16'h45cb;
        src100 <= 16'h71e8;
        src101 <= 16'hd751;
        src102 <= 16'h22ab;
        src103 <= 16'hda1e;
        src104 <= 16'hba88;
        src105 <= 16'hcf16;
        src106 <= 16'ha510;
        src107 <= 16'hf19b;
        src108 <= 16'h7937;
        src109 <= 16'he62a;
        src110 <= 16'h278b;
        src111 <= 16'hecd7;
        src112 <= 16'h1945;
        src113 <= 16'h9b2;
        src114 <= 16'hf841;
        src115 <= 16'hd687;
        src116 <= 16'h897;
        src117 <= 16'hd861;
        src118 <= 16'h95da;
        src119 <= 16'h6a8f;
        src120 <= 16'hfda2;
        src121 <= 16'h8db4;
        src122 <= 16'h53c1;
        src123 <= 16'haa1d;
        src124 <= 16'h9989;
        src125 <= 16'h8bcb;
        src126 <= 16'he601;
        src127 <= 16'hce26;
        exp <= 23'h3ffce9;
        #1
        src0 <= 16'h488d;
        src1 <= 16'h1ab7;
        src2 <= 16'h53a4;
        src3 <= 16'h711e;
        src4 <= 16'hd26b;
        src5 <= 16'h8bdb;
        src6 <= 16'hcb51;
        src7 <= 16'hda18;
        src8 <= 16'h3e9;
        src9 <= 16'h3dab;
        src10 <= 16'h3e76;
        src11 <= 16'hccfc;
        src12 <= 16'h8342;
        src13 <= 16'ha8e8;
        src14 <= 16'ha53a;
        src15 <= 16'he19b;
        src16 <= 16'h438a;
        src17 <= 16'h82d6;
        src18 <= 16'h47a7;
        src19 <= 16'he542;
        src20 <= 16'hdc22;
        src21 <= 16'h3f80;
        src22 <= 16'h2e98;
        src23 <= 16'h6092;
        src24 <= 16'h610f;
        src25 <= 16'h2164;
        src26 <= 16'hab10;
        src27 <= 16'h9eaf;
        src28 <= 16'h6e6e;
        src29 <= 16'h9d97;
        src30 <= 16'h25d4;
        src31 <= 16'hadfc;
        src32 <= 16'h2fd9;
        src33 <= 16'hb60b;
        src34 <= 16'h2feb;
        src35 <= 16'hf3a6;
        src36 <= 16'h8ca3;
        src37 <= 16'h59d0;
        src38 <= 16'hc5de;
        src39 <= 16'hdbe5;
        src40 <= 16'h687a;
        src41 <= 16'hb2d0;
        src42 <= 16'h6457;
        src43 <= 16'h76de;
        src44 <= 16'h66d;
        src45 <= 16'h17c;
        src46 <= 16'h564b;
        src47 <= 16'h2ac;
        src48 <= 16'h7b85;
        src49 <= 16'h2be7;
        src50 <= 16'h332e;
        src51 <= 16'hbbf7;
        src52 <= 16'hec94;
        src53 <= 16'hfd4;
        src54 <= 16'ha0c0;
        src55 <= 16'h6717;
        src56 <= 16'hfe87;
        src57 <= 16'hfc17;
        src58 <= 16'hc7f1;
        src59 <= 16'h34b0;
        src60 <= 16'ha64f;
        src61 <= 16'hfc5f;
        src62 <= 16'h41d9;
        src63 <= 16'h64b8;
        src64 <= 16'h5028;
        src65 <= 16'h9362;
        src66 <= 16'hd7a2;
        src67 <= 16'hf703;
        src68 <= 16'h970;
        src69 <= 16'h71a4;
        src70 <= 16'h3454;
        src71 <= 16'hf222;
        src72 <= 16'h555;
        src73 <= 16'h8597;
        src74 <= 16'h118c;
        src75 <= 16'ha4f7;
        src76 <= 16'h44fc;
        src77 <= 16'hde42;
        src78 <= 16'h6bde;
        src79 <= 16'hd375;
        src80 <= 16'he5b0;
        src81 <= 16'h231d;
        src82 <= 16'h4883;
        src83 <= 16'h51d2;
        src84 <= 16'h325c;
        src85 <= 16'hc3cf;
        src86 <= 16'hab41;
        src87 <= 16'h30d6;
        src88 <= 16'hc7f;
        src89 <= 16'hbdf8;
        src90 <= 16'h4519;
        src91 <= 16'hae12;
        src92 <= 16'h796c;
        src93 <= 16'h2023;
        src94 <= 16'hb5ac;
        src95 <= 16'h7f4d;
        src96 <= 16'hf662;
        src97 <= 16'he13b;
        src98 <= 16'h826c;
        src99 <= 16'hbd2e;
        src100 <= 16'h21e1;
        src101 <= 16'h441f;
        src102 <= 16'h3904;
        src103 <= 16'h8da7;
        src104 <= 16'hc86;
        src105 <= 16'h7092;
        src106 <= 16'hca66;
        src107 <= 16'h7263;
        src108 <= 16'h3e8f;
        src109 <= 16'hee6d;
        src110 <= 16'h6371;
        src111 <= 16'haf72;
        src112 <= 16'h9ddd;
        src113 <= 16'h22e;
        src114 <= 16'h6196;
        src115 <= 16'h9964;
        src116 <= 16'hb1c9;
        src117 <= 16'hb6e0;
        src118 <= 16'h572d;
        src119 <= 16'h3731;
        src120 <= 16'h3306;
        src121 <= 16'h24f4;
        src122 <= 16'h59eb;
        src123 <= 16'hbba5;
        src124 <= 16'h6003;
        src125 <= 16'ha025;
        src126 <= 16'hacd0;
        src127 <= 16'h151e;
        exp <= 23'h3d32c3;
        #1
        src0 <= 16'hc7fd;
        src1 <= 16'he376;
        src2 <= 16'haf7a;
        src3 <= 16'hf276;
        src4 <= 16'h4015;
        src5 <= 16'h9c5d;
        src6 <= 16'h225b;
        src7 <= 16'h2810;
        src8 <= 16'h24a0;
        src9 <= 16'h7b3f;
        src10 <= 16'hf95a;
        src11 <= 16'hba70;
        src12 <= 16'h6e56;
        src13 <= 16'hb614;
        src14 <= 16'h8f86;
        src15 <= 16'h50da;
        src16 <= 16'hd7a2;
        src17 <= 16'ha24d;
        src18 <= 16'h6896;
        src19 <= 16'hbbf5;
        src20 <= 16'h8e7b;
        src21 <= 16'hf3dc;
        src22 <= 16'h3678;
        src23 <= 16'hbfa9;
        src24 <= 16'hde4f;
        src25 <= 16'hbb6e;
        src26 <= 16'h9e2a;
        src27 <= 16'he63;
        src28 <= 16'h48;
        src29 <= 16'h9eef;
        src30 <= 16'hf82f;
        src31 <= 16'h1178;
        src32 <= 16'h9ee6;
        src33 <= 16'h54e9;
        src34 <= 16'h746;
        src35 <= 16'hb80;
        src36 <= 16'h9e2b;
        src37 <= 16'hc5a7;
        src38 <= 16'h4041;
        src39 <= 16'hf880;
        src40 <= 16'h33d7;
        src41 <= 16'h96fc;
        src42 <= 16'h7fd;
        src43 <= 16'h5dbf;
        src44 <= 16'h2566;
        src45 <= 16'ha9b8;
        src46 <= 16'h6275;
        src47 <= 16'hac4d;
        src48 <= 16'hd562;
        src49 <= 16'h467c;
        src50 <= 16'h81dd;
        src51 <= 16'h7a86;
        src52 <= 16'hb3db;
        src53 <= 16'h87af;
        src54 <= 16'he3ce;
        src55 <= 16'h8613;
        src56 <= 16'h3a26;
        src57 <= 16'h3175;
        src58 <= 16'h2258;
        src59 <= 16'h5da0;
        src60 <= 16'h7383;
        src61 <= 16'h2708;
        src62 <= 16'h4333;
        src63 <= 16'hb143;
        src64 <= 16'h1714;
        src65 <= 16'h98af;
        src66 <= 16'h2693;
        src67 <= 16'h2f7b;
        src68 <= 16'hd95b;
        src69 <= 16'h830c;
        src70 <= 16'hd269;
        src71 <= 16'h6b5c;
        src72 <= 16'h4a43;
        src73 <= 16'hc0d1;
        src74 <= 16'hf746;
        src75 <= 16'hcfb1;
        src76 <= 16'h7ad4;
        src77 <= 16'haa8b;
        src78 <= 16'h95dd;
        src79 <= 16'hb42f;
        src80 <= 16'h5b67;
        src81 <= 16'hd14;
        src82 <= 16'hc892;
        src83 <= 16'h945c;
        src84 <= 16'h3096;
        src85 <= 16'h2636;
        src86 <= 16'h2bc4;
        src87 <= 16'h8a6a;
        src88 <= 16'hc523;
        src89 <= 16'hc113;
        src90 <= 16'hcca1;
        src91 <= 16'h3759;
        src92 <= 16'hfe17;
        src93 <= 16'hd310;
        src94 <= 16'hb2c9;
        src95 <= 16'hb840;
        src96 <= 16'h77e8;
        src97 <= 16'hcc7;
        src98 <= 16'h3049;
        src99 <= 16'h50d8;
        src100 <= 16'ha652;
        src101 <= 16'h2db;
        src102 <= 16'haf5f;
        src103 <= 16'h8d7c;
        src104 <= 16'hde92;
        src105 <= 16'h7c40;
        src106 <= 16'hb51;
        src107 <= 16'hab2b;
        src108 <= 16'h3f70;
        src109 <= 16'h6026;
        src110 <= 16'ha1b6;
        src111 <= 16'h4e;
        src112 <= 16'h61fb;
        src113 <= 16'h5d6e;
        src114 <= 16'h6031;
        src115 <= 16'hc176;
        src116 <= 16'h87c4;
        src117 <= 16'h57ad;
        src118 <= 16'h5246;
        src119 <= 16'h7197;
        src120 <= 16'hcdde;
        src121 <= 16'h3a6;
        src122 <= 16'hda06;
        src123 <= 16'h85e0;
        src124 <= 16'h9093;
        src125 <= 16'h1b8;
        src126 <= 16'hcf75;
        src127 <= 16'h957d;
        exp <= 23'h3f229f;
        #1
        src0 <= 16'h8ffe;
        src1 <= 16'hf0c9;
        src2 <= 16'hc87d;
        src3 <= 16'hf72b;
        src4 <= 16'h7387;
        src5 <= 16'he1c8;
        src6 <= 16'ha122;
        src7 <= 16'haad1;
        src8 <= 16'hb1f8;
        src9 <= 16'ha1dc;
        src10 <= 16'hf7bb;
        src11 <= 16'he43e;
        src12 <= 16'h4a9c;
        src13 <= 16'h643d;
        src14 <= 16'ha278;
        src15 <= 16'h7df5;
        src16 <= 16'h5aa8;
        src17 <= 16'hd98f;
        src18 <= 16'hb3a5;
        src19 <= 16'hd8be;
        src20 <= 16'h7ae6;
        src21 <= 16'h6101;
        src22 <= 16'hd505;
        src23 <= 16'h70ee;
        src24 <= 16'h626c;
        src25 <= 16'h43af;
        src26 <= 16'h33c2;
        src27 <= 16'ha634;
        src28 <= 16'h5a2a;
        src29 <= 16'h71ae;
        src30 <= 16'h74fe;
        src31 <= 16'haa49;
        src32 <= 16'h6ec0;
        src33 <= 16'h43d6;
        src34 <= 16'h5cba;
        src35 <= 16'hdba4;
        src36 <= 16'hddb7;
        src37 <= 16'h232c;
        src38 <= 16'ha1b0;
        src39 <= 16'h3501;
        src40 <= 16'h3a88;
        src41 <= 16'h6d05;
        src42 <= 16'h584d;
        src43 <= 16'h41c8;
        src44 <= 16'hde90;
        src45 <= 16'hf58;
        src46 <= 16'heb85;
        src47 <= 16'h562c;
        src48 <= 16'h16ce;
        src49 <= 16'he6ec;
        src50 <= 16'h19dc;
        src51 <= 16'h3666;
        src52 <= 16'h77a0;
        src53 <= 16'h44f8;
        src54 <= 16'h35a2;
        src55 <= 16'h7b8c;
        src56 <= 16'h2ebe;
        src57 <= 16'ha892;
        src58 <= 16'hd8dc;
        src59 <= 16'h6acd;
        src60 <= 16'hb462;
        src61 <= 16'h1f54;
        src62 <= 16'h8e03;
        src63 <= 16'h542e;
        src64 <= 16'he4c3;
        src65 <= 16'h7b7d;
        src66 <= 16'hff1a;
        src67 <= 16'h99a1;
        src68 <= 16'h6cd4;
        src69 <= 16'h7953;
        src70 <= 16'h398a;
        src71 <= 16'hfcb3;
        src72 <= 16'hb10b;
        src73 <= 16'hfda6;
        src74 <= 16'hcf2;
        src75 <= 16'he06b;
        src76 <= 16'hf5a;
        src77 <= 16'h5ce4;
        src78 <= 16'h9993;
        src79 <= 16'hd241;
        src80 <= 16'hb05e;
        src81 <= 16'h4997;
        src82 <= 16'hfaee;
        src83 <= 16'ha775;
        src84 <= 16'h547;
        src85 <= 16'h2b6f;
        src86 <= 16'he369;
        src87 <= 16'hc6b4;
        src88 <= 16'he3d7;
        src89 <= 16'hf492;
        src90 <= 16'h8ff2;
        src91 <= 16'h6aa;
        src92 <= 16'hfd80;
        src93 <= 16'hd46;
        src94 <= 16'heb13;
        src95 <= 16'h4cf7;
        src96 <= 16'hf6cc;
        src97 <= 16'he918;
        src98 <= 16'h8b64;
        src99 <= 16'h9f6e;
        src100 <= 16'h634b;
        src101 <= 16'h21d0;
        src102 <= 16'hc612;
        src103 <= 16'h9168;
        src104 <= 16'hf8ad;
        src105 <= 16'hf8a4;
        src106 <= 16'hb176;
        src107 <= 16'h5289;
        src108 <= 16'hd0d8;
        src109 <= 16'h2a19;
        src110 <= 16'h3edb;
        src111 <= 16'h4b1f;
        src112 <= 16'h9672;
        src113 <= 16'h753e;
        src114 <= 16'h41c1;
        src115 <= 16'h2e3c;
        src116 <= 16'hccf0;
        src117 <= 16'ha3c4;
        src118 <= 16'h7b98;
        src119 <= 16'hb1c0;
        src120 <= 16'h9873;
        src121 <= 16'h4429;
        src122 <= 16'h593e;
        src123 <= 16'h155;
        src124 <= 16'h181b;
        src125 <= 16'hdb6a;
        src126 <= 16'hbe95;
        src127 <= 16'h5bb6;
        exp <= 23'h44618a;
        #1
        src0 <= 16'h27b0;
        src1 <= 16'he959;
        src2 <= 16'h2324;
        src3 <= 16'hcb10;
        src4 <= 16'h350f;
        src5 <= 16'hb22b;
        src6 <= 16'h8c34;
        src7 <= 16'hd4af;
        src8 <= 16'h2746;
        src9 <= 16'hd087;
        src10 <= 16'h957d;
        src11 <= 16'heb6a;
        src12 <= 16'h776b;
        src13 <= 16'hcaf2;
        src14 <= 16'h929d;
        src15 <= 16'hc72a;
        src16 <= 16'h9265;
        src17 <= 16'h5ed;
        src18 <= 16'h844b;
        src19 <= 16'h335c;
        src20 <= 16'h31a0;
        src21 <= 16'he813;
        src22 <= 16'he704;
        src23 <= 16'h283b;
        src24 <= 16'h9a8e;
        src25 <= 16'h4bec;
        src26 <= 16'h2aa4;
        src27 <= 16'h4924;
        src28 <= 16'h7c6;
        src29 <= 16'h7391;
        src30 <= 16'h4a5b;
        src31 <= 16'he484;
        src32 <= 16'h175;
        src33 <= 16'hcee3;
        src34 <= 16'hf413;
        src35 <= 16'hd7f8;
        src36 <= 16'hf5b0;
        src37 <= 16'h7e95;
        src38 <= 16'hb622;
        src39 <= 16'hd44e;
        src40 <= 16'hed63;
        src41 <= 16'h2f7d;
        src42 <= 16'he2a;
        src43 <= 16'hdd1b;
        src44 <= 16'hede7;
        src45 <= 16'he171;
        src46 <= 16'hef1a;
        src47 <= 16'hb3ce;
        src48 <= 16'hfed1;
        src49 <= 16'h618;
        src50 <= 16'hd91;
        src51 <= 16'h8dac;
        src52 <= 16'h1b5c;
        src53 <= 16'hbd4d;
        src54 <= 16'h156d;
        src55 <= 16'h53f4;
        src56 <= 16'hc0c7;
        src57 <= 16'hef3b;
        src58 <= 16'hc8a4;
        src59 <= 16'hf35f;
        src60 <= 16'hebe9;
        src61 <= 16'h2c39;
        src62 <= 16'h350a;
        src63 <= 16'hebfd;
        src64 <= 16'hd0e3;
        src65 <= 16'h61cf;
        src66 <= 16'ha500;
        src67 <= 16'h7524;
        src68 <= 16'h8feb;
        src69 <= 16'h87c4;
        src70 <= 16'hc033;
        src71 <= 16'hc142;
        src72 <= 16'hfbab;
        src73 <= 16'h93aa;
        src74 <= 16'h86b5;
        src75 <= 16'h6bf2;
        src76 <= 16'h2a17;
        src77 <= 16'h5f51;
        src78 <= 16'h7018;
        src79 <= 16'h1579;
        src80 <= 16'h3d0a;
        src81 <= 16'hfdb0;
        src82 <= 16'he147;
        src83 <= 16'he222;
        src84 <= 16'h8e39;
        src85 <= 16'h2b8d;
        src86 <= 16'h6021;
        src87 <= 16'h2007;
        src88 <= 16'h8707;
        src89 <= 16'ha70a;
        src90 <= 16'hf2a3;
        src91 <= 16'hf6b8;
        src92 <= 16'h903c;
        src93 <= 16'hcfca;
        src94 <= 16'h57a6;
        src95 <= 16'hfc33;
        src96 <= 16'h642b;
        src97 <= 16'h9e5d;
        src98 <= 16'hbfb2;
        src99 <= 16'h599c;
        src100 <= 16'h4408;
        src101 <= 16'hcd76;
        src102 <= 16'h9b65;
        src103 <= 16'h3106;
        src104 <= 16'h12ad;
        src105 <= 16'h25ee;
        src106 <= 16'hf030;
        src107 <= 16'h83c9;
        src108 <= 16'h2ed;
        src109 <= 16'h4401;
        src110 <= 16'h9663;
        src111 <= 16'h2c1e;
        src112 <= 16'h9765;
        src113 <= 16'h51e9;
        src114 <= 16'h11a3;
        src115 <= 16'hfc39;
        src116 <= 16'heb4;
        src117 <= 16'h60dd;
        src118 <= 16'h6bc;
        src119 <= 16'he83b;
        src120 <= 16'ha73a;
        src121 <= 16'hb4b0;
        src122 <= 16'h50ef;
        src123 <= 16'h9720;
        src124 <= 16'h8d1a;
        src125 <= 16'hf401;
        src126 <= 16'hbca2;
        src127 <= 16'hacbf;
        exp <= 23'h4524a4;
        #1
        src0 <= 16'hb1e8;
        src1 <= 16'hc2c2;
        src2 <= 16'h322a;
        src3 <= 16'h8ca;
        src4 <= 16'hd196;
        src5 <= 16'h3f78;
        src6 <= 16'hb63e;
        src7 <= 16'hc7db;
        src8 <= 16'hb62a;
        src9 <= 16'ha952;
        src10 <= 16'haf73;
        src11 <= 16'h77ba;
        src12 <= 16'hc5f3;
        src13 <= 16'h1e4a;
        src14 <= 16'h6e10;
        src15 <= 16'h5090;
        src16 <= 16'h9380;
        src17 <= 16'he6c7;
        src18 <= 16'h1c05;
        src19 <= 16'h79fa;
        src20 <= 16'h2bcd;
        src21 <= 16'h8f19;
        src22 <= 16'hd65a;
        src23 <= 16'h4c65;
        src24 <= 16'h7fee;
        src25 <= 16'hbeb2;
        src26 <= 16'h3208;
        src27 <= 16'hbbc;
        src28 <= 16'hd11f;
        src29 <= 16'hc4e9;
        src30 <= 16'he06f;
        src31 <= 16'h9668;
        src32 <= 16'h27ed;
        src33 <= 16'hf1e7;
        src34 <= 16'hec2d;
        src35 <= 16'h7c06;
        src36 <= 16'h28ed;
        src37 <= 16'hcb9;
        src38 <= 16'h6ddf;
        src39 <= 16'h124b;
        src40 <= 16'h59fe;
        src41 <= 16'h537b;
        src42 <= 16'hc817;
        src43 <= 16'h8ef7;
        src44 <= 16'h909e;
        src45 <= 16'heb98;
        src46 <= 16'hf509;
        src47 <= 16'h7f91;
        src48 <= 16'h9d6;
        src49 <= 16'he876;
        src50 <= 16'h4530;
        src51 <= 16'hd077;
        src52 <= 16'h46c0;
        src53 <= 16'hbe82;
        src54 <= 16'he3f9;
        src55 <= 16'h63bc;
        src56 <= 16'hdaec;
        src57 <= 16'h4cba;
        src58 <= 16'hf8c2;
        src59 <= 16'hb36;
        src60 <= 16'hea90;
        src61 <= 16'h6f08;
        src62 <= 16'h4be5;
        src63 <= 16'h387b;
        src64 <= 16'h702;
        src65 <= 16'h57db;
        src66 <= 16'h3feb;
        src67 <= 16'hb009;
        src68 <= 16'he209;
        src69 <= 16'h3549;
        src70 <= 16'h78e2;
        src71 <= 16'hb269;
        src72 <= 16'h1db6;
        src73 <= 16'h1efd;
        src74 <= 16'h4c26;
        src75 <= 16'ha265;
        src76 <= 16'h8c6f;
        src77 <= 16'h730;
        src78 <= 16'h9d1f;
        src79 <= 16'hb5b7;
        src80 <= 16'h6c50;
        src81 <= 16'h2cf0;
        src82 <= 16'ha0cd;
        src83 <= 16'h8eb9;
        src84 <= 16'heea7;
        src85 <= 16'hd68f;
        src86 <= 16'h648b;
        src87 <= 16'hd673;
        src88 <= 16'h3cc3;
        src89 <= 16'h7c4c;
        src90 <= 16'h7e76;
        src91 <= 16'h2a1c;
        src92 <= 16'hc580;
        src93 <= 16'ha9dd;
        src94 <= 16'hfbff;
        src95 <= 16'hbae8;
        src96 <= 16'h4e97;
        src97 <= 16'h857d;
        src98 <= 16'ha359;
        src99 <= 16'h7adc;
        src100 <= 16'hd877;
        src101 <= 16'h1e07;
        src102 <= 16'h6b3c;
        src103 <= 16'hd07d;
        src104 <= 16'he3b5;
        src105 <= 16'hf44c;
        src106 <= 16'h4ef6;
        src107 <= 16'h257b;
        src108 <= 16'h5d41;
        src109 <= 16'h9fa9;
        src110 <= 16'h14c2;
        src111 <= 16'hbdcc;
        src112 <= 16'h950;
        src113 <= 16'hac5a;
        src114 <= 16'h1673;
        src115 <= 16'h1c18;
        src116 <= 16'h611f;
        src117 <= 16'hf72b;
        src118 <= 16'hc12f;
        src119 <= 16'h1922;
        src120 <= 16'h6f12;
        src121 <= 16'h7501;
        src122 <= 16'ha8c9;
        src123 <= 16'h40ea;
        src124 <= 16'h2cec;
        src125 <= 16'ha030;
        src126 <= 16'h2594;
        src127 <= 16'hbddd;
        exp <= 23'h4038b4;
        #1
        src0 <= 16'h5688;
        src1 <= 16'h9989;
        src2 <= 16'h8fa;
        src3 <= 16'h4c41;
        src4 <= 16'hc2b0;
        src5 <= 16'h1674;
        src6 <= 16'h6369;
        src7 <= 16'h95a0;
        src8 <= 16'h8b86;
        src9 <= 16'hf9c2;
        src10 <= 16'h64e0;
        src11 <= 16'h3c3;
        src12 <= 16'ha3f7;
        src13 <= 16'h95dc;
        src14 <= 16'hb263;
        src15 <= 16'h6e5f;
        src16 <= 16'h2c18;
        src17 <= 16'hec9e;
        src18 <= 16'haf78;
        src19 <= 16'h1ee4;
        src20 <= 16'h74e5;
        src21 <= 16'hd734;
        src22 <= 16'he1fc;
        src23 <= 16'hde07;
        src24 <= 16'h22c;
        src25 <= 16'h39af;
        src26 <= 16'hdc73;
        src27 <= 16'h243e;
        src28 <= 16'h1309;
        src29 <= 16'he09d;
        src30 <= 16'h8ebb;
        src31 <= 16'h3849;
        src32 <= 16'h7928;
        src33 <= 16'hb3cb;
        src34 <= 16'hb3a8;
        src35 <= 16'h2688;
        src36 <= 16'hd07e;
        src37 <= 16'heecd;
        src38 <= 16'hcd57;
        src39 <= 16'h7812;
        src40 <= 16'h4e64;
        src41 <= 16'he83;
        src42 <= 16'hb38e;
        src43 <= 16'hd998;
        src44 <= 16'h4c38;
        src45 <= 16'h435;
        src46 <= 16'hc8d6;
        src47 <= 16'h1958;
        src48 <= 16'hded2;
        src49 <= 16'h841b;
        src50 <= 16'h94b5;
        src51 <= 16'h8b26;
        src52 <= 16'h559e;
        src53 <= 16'h4b7e;
        src54 <= 16'hcc88;
        src55 <= 16'h935;
        src56 <= 16'h6063;
        src57 <= 16'h6789;
        src58 <= 16'ha87e;
        src59 <= 16'h5eab;
        src60 <= 16'hf293;
        src61 <= 16'hde39;
        src62 <= 16'h8a82;
        src63 <= 16'h72f;
        src64 <= 16'h7914;
        src65 <= 16'h421e;
        src66 <= 16'h4514;
        src67 <= 16'hd95f;
        src68 <= 16'h5ada;
        src69 <= 16'h4fb3;
        src70 <= 16'h7aa7;
        src71 <= 16'hf10a;
        src72 <= 16'he974;
        src73 <= 16'h9bf4;
        src74 <= 16'heba1;
        src75 <= 16'hcfad;
        src76 <= 16'h18c;
        src77 <= 16'h6d45;
        src78 <= 16'hd329;
        src79 <= 16'h5a95;
        src80 <= 16'h51c8;
        src81 <= 16'hbea4;
        src82 <= 16'h7979;
        src83 <= 16'h12ce;
        src84 <= 16'he08f;
        src85 <= 16'h2792;
        src86 <= 16'h7abc;
        src87 <= 16'h911e;
        src88 <= 16'h1459;
        src89 <= 16'h34f3;
        src90 <= 16'hfc2f;
        src91 <= 16'h80c0;
        src92 <= 16'hc76f;
        src93 <= 16'h63aa;
        src94 <= 16'h96e4;
        src95 <= 16'hbb75;
        src96 <= 16'h3bb7;
        src97 <= 16'h154d;
        src98 <= 16'h24f6;
        src99 <= 16'h40d;
        src100 <= 16'h138c;
        src101 <= 16'h2c72;
        src102 <= 16'h317a;
        src103 <= 16'h2312;
        src104 <= 16'hcb42;
        src105 <= 16'hc69f;
        src106 <= 16'h74fc;
        src107 <= 16'h3db8;
        src108 <= 16'h155f;
        src109 <= 16'hfe1b;
        src110 <= 16'h7ed0;
        src111 <= 16'h5036;
        src112 <= 16'h8832;
        src113 <= 16'h8bb4;
        src114 <= 16'h502f;
        src115 <= 16'h7b14;
        src116 <= 16'h5bc;
        src117 <= 16'he95;
        src118 <= 16'h892a;
        src119 <= 16'hbd33;
        src120 <= 16'h83c1;
        src121 <= 16'h620b;
        src122 <= 16'h94b1;
        src123 <= 16'hd848;
        src124 <= 16'h44f2;
        src125 <= 16'hcac0;
        src126 <= 16'hfbd5;
        src127 <= 16'hdbf9;
        exp <= 23'h3e0954;
        #1
        src0 <= 16'hede3;
        src1 <= 16'h60ae;
        src2 <= 16'ha215;
        src3 <= 16'he621;
        src4 <= 16'hee31;
        src5 <= 16'hee03;
        src6 <= 16'hd995;
        src7 <= 16'h8638;
        src8 <= 16'h5b84;
        src9 <= 16'hdf2;
        src10 <= 16'hebf1;
        src11 <= 16'h4495;
        src12 <= 16'h7d3b;
        src13 <= 16'h26b6;
        src14 <= 16'h24f9;
        src15 <= 16'h379c;
        src16 <= 16'hb9a2;
        src17 <= 16'h75b6;
        src18 <= 16'h366c;
        src19 <= 16'h3bba;
        src20 <= 16'h329e;
        src21 <= 16'ha1cf;
        src22 <= 16'hcefe;
        src23 <= 16'hb5cd;
        src24 <= 16'h10f8;
        src25 <= 16'h5907;
        src26 <= 16'h5cfd;
        src27 <= 16'h6bae;
        src28 <= 16'h393c;
        src29 <= 16'ha8db;
        src30 <= 16'h68a3;
        src31 <= 16'h480a;
        src32 <= 16'h6f86;
        src33 <= 16'h2c25;
        src34 <= 16'hff4d;
        src35 <= 16'h5fe1;
        src36 <= 16'h6911;
        src37 <= 16'hbd82;
        src38 <= 16'he64;
        src39 <= 16'h3271;
        src40 <= 16'h1631;
        src41 <= 16'h2a5c;
        src42 <= 16'h7240;
        src43 <= 16'h2f38;
        src44 <= 16'h5016;
        src45 <= 16'hf704;
        src46 <= 16'ha9e8;
        src47 <= 16'haaae;
        src48 <= 16'hee6c;
        src49 <= 16'h2fad;
        src50 <= 16'h626f;
        src51 <= 16'h2b74;
        src52 <= 16'h54cc;
        src53 <= 16'hc77b;
        src54 <= 16'h3eb7;
        src55 <= 16'hfabb;
        src56 <= 16'hd3a;
        src57 <= 16'h9f91;
        src58 <= 16'he9fd;
        src59 <= 16'hef29;
        src60 <= 16'h4bb3;
        src61 <= 16'hec5a;
        src62 <= 16'h3ad2;
        src63 <= 16'h115;
        src64 <= 16'he5d6;
        src65 <= 16'hd1eb;
        src66 <= 16'he23c;
        src67 <= 16'h7811;
        src68 <= 16'h6faf;
        src69 <= 16'h7658;
        src70 <= 16'h52a;
        src71 <= 16'hca0e;
        src72 <= 16'heb46;
        src73 <= 16'hcbf3;
        src74 <= 16'h5167;
        src75 <= 16'he16b;
        src76 <= 16'hc795;
        src77 <= 16'hfbfe;
        src78 <= 16'h3cf5;
        src79 <= 16'hfecc;
        src80 <= 16'h9c41;
        src81 <= 16'h5e08;
        src82 <= 16'h9f7a;
        src83 <= 16'h9f29;
        src84 <= 16'h1c46;
        src85 <= 16'hff4;
        src86 <= 16'h3a0d;
        src87 <= 16'h5802;
        src88 <= 16'hbf28;
        src89 <= 16'h127b;
        src90 <= 16'he119;
        src91 <= 16'h555e;
        src92 <= 16'he74d;
        src93 <= 16'h362d;
        src94 <= 16'hd9fc;
        src95 <= 16'h3874;
        src96 <= 16'hf713;
        src97 <= 16'h3bcb;
        src98 <= 16'h880e;
        src99 <= 16'hffe3;
        src100 <= 16'h15e2;
        src101 <= 16'h71cf;
        src102 <= 16'hf9cc;
        src103 <= 16'ha1a8;
        src104 <= 16'h6f7d;
        src105 <= 16'h10ac;
        src106 <= 16'h54a8;
        src107 <= 16'h2a1;
        src108 <= 16'h8830;
        src109 <= 16'h6e96;
        src110 <= 16'h69b1;
        src111 <= 16'h3461;
        src112 <= 16'h78ea;
        src113 <= 16'he9ff;
        src114 <= 16'h9978;
        src115 <= 16'hf19;
        src116 <= 16'h8001;
        src117 <= 16'h34a3;
        src118 <= 16'h5a06;
        src119 <= 16'hcb57;
        src120 <= 16'hb9f0;
        src121 <= 16'hf271;
        src122 <= 16'he0b;
        src123 <= 16'hf660;
        src124 <= 16'he8cc;
        src125 <= 16'h5002;
        src126 <= 16'h2dfa;
        src127 <= 16'h9365;
        exp <= 23'h400395;
        #1
        src0 <= 16'h4e60;
        src1 <= 16'h6084;
        src2 <= 16'h6d8e;
        src3 <= 16'hf86e;
        src4 <= 16'h93d;
        src5 <= 16'h772d;
        src6 <= 16'h774a;
        src7 <= 16'h21c5;
        src8 <= 16'h5206;
        src9 <= 16'hc67b;
        src10 <= 16'h33d6;
        src11 <= 16'h48e4;
        src12 <= 16'hf21c;
        src13 <= 16'h3845;
        src14 <= 16'hcc8c;
        src15 <= 16'h4f82;
        src16 <= 16'hfca5;
        src17 <= 16'heb16;
        src18 <= 16'h3803;
        src19 <= 16'h1f12;
        src20 <= 16'h1102;
        src21 <= 16'h5d11;
        src22 <= 16'h553c;
        src23 <= 16'hb05e;
        src24 <= 16'ha7d2;
        src25 <= 16'h3a4d;
        src26 <= 16'he947;
        src27 <= 16'hd512;
        src28 <= 16'hdb12;
        src29 <= 16'h861a;
        src30 <= 16'h7ccc;
        src31 <= 16'h6934;
        src32 <= 16'h9710;
        src33 <= 16'h9fba;
        src34 <= 16'he49d;
        src35 <= 16'h715d;
        src36 <= 16'hed3e;
        src37 <= 16'hf348;
        src38 <= 16'h366d;
        src39 <= 16'h1967;
        src40 <= 16'h99c3;
        src41 <= 16'h7257;
        src42 <= 16'h3918;
        src43 <= 16'h577a;
        src44 <= 16'h9e4c;
        src45 <= 16'hec35;
        src46 <= 16'h7663;
        src47 <= 16'hdba8;
        src48 <= 16'h44d3;
        src49 <= 16'h77a9;
        src50 <= 16'h353b;
        src51 <= 16'h791a;
        src52 <= 16'h4efb;
        src53 <= 16'hd83a;
        src54 <= 16'h83dc;
        src55 <= 16'hf8b7;
        src56 <= 16'h4225;
        src57 <= 16'haa2e;
        src58 <= 16'hd94;
        src59 <= 16'h527f;
        src60 <= 16'hbb0d;
        src61 <= 16'h5a5a;
        src62 <= 16'ha8c4;
        src63 <= 16'h1d79;
        src64 <= 16'h2c3a;
        src65 <= 16'hc9d2;
        src66 <= 16'h5081;
        src67 <= 16'ha7b6;
        src68 <= 16'h8c04;
        src69 <= 16'h20ad;
        src70 <= 16'h2893;
        src71 <= 16'h2633;
        src72 <= 16'hd592;
        src73 <= 16'h755;
        src74 <= 16'hcdac;
        src75 <= 16'had3f;
        src76 <= 16'h6250;
        src77 <= 16'h76f4;
        src78 <= 16'h807b;
        src79 <= 16'h46a1;
        src80 <= 16'h44f8;
        src81 <= 16'hc931;
        src82 <= 16'h69fc;
        src83 <= 16'h9cf9;
        src84 <= 16'h3851;
        src85 <= 16'h86f7;
        src86 <= 16'h7d96;
        src87 <= 16'h221f;
        src88 <= 16'h42a3;
        src89 <= 16'hd5d9;
        src90 <= 16'h66c8;
        src91 <= 16'hdfa7;
        src92 <= 16'h9f8c;
        src93 <= 16'h98c1;
        src94 <= 16'ha63c;
        src95 <= 16'h9e88;
        src96 <= 16'haac9;
        src97 <= 16'h9f70;
        src98 <= 16'h40d9;
        src99 <= 16'hf2cf;
        src100 <= 16'haec1;
        src101 <= 16'hb540;
        src102 <= 16'hf6d8;
        src103 <= 16'hcdda;
        src104 <= 16'hb18a;
        src105 <= 16'h964;
        src106 <= 16'h9cb3;
        src107 <= 16'h1304;
        src108 <= 16'hf9ea;
        src109 <= 16'hf4fd;
        src110 <= 16'hbc61;
        src111 <= 16'h39dc;
        src112 <= 16'h86d;
        src113 <= 16'h27a0;
        src114 <= 16'hdcf3;
        src115 <= 16'h63fc;
        src116 <= 16'h7d66;
        src117 <= 16'hcfc1;
        src118 <= 16'h1554;
        src119 <= 16'haf81;
        src120 <= 16'h29fb;
        src121 <= 16'h20d5;
        src122 <= 16'h91f0;
        src123 <= 16'hb791;
        src124 <= 16'h229a;
        src125 <= 16'hae1c;
        src126 <= 16'h7105;
        src127 <= 16'h2066;
        exp <= 23'h3fb2e7;
        #1
        src0 <= 16'h523a;
        src1 <= 16'h7f41;
        src2 <= 16'h19f3;
        src3 <= 16'hde75;
        src4 <= 16'hc2e3;
        src5 <= 16'hfd07;
        src6 <= 16'hb9d7;
        src7 <= 16'hcdb2;
        src8 <= 16'hb495;
        src9 <= 16'h2bd7;
        src10 <= 16'h64a;
        src11 <= 16'hee2f;
        src12 <= 16'h98c2;
        src13 <= 16'h1fe6;
        src14 <= 16'hb428;
        src15 <= 16'hd274;
        src16 <= 16'h159e;
        src17 <= 16'ha817;
        src18 <= 16'h1442;
        src19 <= 16'h1f95;
        src20 <= 16'hdd59;
        src21 <= 16'h56c3;
        src22 <= 16'h8ae0;
        src23 <= 16'ha6f2;
        src24 <= 16'he65b;
        src25 <= 16'h2c6d;
        src26 <= 16'hbe94;
        src27 <= 16'h31d2;
        src28 <= 16'hccb5;
        src29 <= 16'h9df;
        src30 <= 16'h335c;
        src31 <= 16'h50ba;
        src32 <= 16'hf4c7;
        src33 <= 16'h6b30;
        src34 <= 16'h5975;
        src35 <= 16'h59b;
        src36 <= 16'h789f;
        src37 <= 16'h4fbd;
        src38 <= 16'h6dd;
        src39 <= 16'h3422;
        src40 <= 16'h854e;
        src41 <= 16'h7ad4;
        src42 <= 16'h7afe;
        src43 <= 16'h7bb8;
        src44 <= 16'he586;
        src45 <= 16'h3f9c;
        src46 <= 16'h9e54;
        src47 <= 16'h5f47;
        src48 <= 16'hda9e;
        src49 <= 16'hf5dd;
        src50 <= 16'hcf01;
        src51 <= 16'h2305;
        src52 <= 16'he445;
        src53 <= 16'h1a40;
        src54 <= 16'h8f5a;
        src55 <= 16'h8dd9;
        src56 <= 16'hdc6e;
        src57 <= 16'hf005;
        src58 <= 16'hdf7d;
        src59 <= 16'hbb88;
        src60 <= 16'h3c74;
        src61 <= 16'h744a;
        src62 <= 16'h2efc;
        src63 <= 16'h3251;
        src64 <= 16'hd6f6;
        src65 <= 16'h3fed;
        src66 <= 16'h369c;
        src67 <= 16'he2d;
        src68 <= 16'h9e4;
        src69 <= 16'he7c1;
        src70 <= 16'h6375;
        src71 <= 16'h80b2;
        src72 <= 16'hdc97;
        src73 <= 16'h3ff4;
        src74 <= 16'hd6b2;
        src75 <= 16'h5419;
        src76 <= 16'h5149;
        src77 <= 16'h687e;
        src78 <= 16'h3a76;
        src79 <= 16'h1f24;
        src80 <= 16'h60d;
        src81 <= 16'h5193;
        src82 <= 16'h8465;
        src83 <= 16'hd79;
        src84 <= 16'hd0ae;
        src85 <= 16'he6b1;
        src86 <= 16'h5c6c;
        src87 <= 16'h7212;
        src88 <= 16'h7721;
        src89 <= 16'h273d;
        src90 <= 16'h951e;
        src91 <= 16'h85f2;
        src92 <= 16'h6a4d;
        src93 <= 16'h93a7;
        src94 <= 16'heafb;
        src95 <= 16'hbb54;
        src96 <= 16'h2215;
        src97 <= 16'h3eba;
        src98 <= 16'hb3a2;
        src99 <= 16'hbf86;
        src100 <= 16'h4d77;
        src101 <= 16'h6c17;
        src102 <= 16'h8d65;
        src103 <= 16'h548b;
        src104 <= 16'he836;
        src105 <= 16'h9762;
        src106 <= 16'hfa53;
        src107 <= 16'h37a0;
        src108 <= 16'h9c4d;
        src109 <= 16'hf433;
        src110 <= 16'h6021;
        src111 <= 16'h13b3;
        src112 <= 16'hc8bc;
        src113 <= 16'hf5d;
        src114 <= 16'hc787;
        src115 <= 16'hef9e;
        src116 <= 16'had53;
        src117 <= 16'h4d12;
        src118 <= 16'he25b;
        src119 <= 16'h6a70;
        src120 <= 16'h20ec;
        src121 <= 16'h24d0;
        src122 <= 16'h2f48;
        src123 <= 16'ha7d9;
        src124 <= 16'h6fea;
        src125 <= 16'h5845;
        src126 <= 16'hc7b6;
        src127 <= 16'h1515;
        exp <= 23'h3e2558;
        #1
        src0 <= 16'h59cb;
        src1 <= 16'h2d3f;
        src2 <= 16'h5beb;
        src3 <= 16'hb8f7;
        src4 <= 16'h44d7;
        src5 <= 16'h6398;
        src6 <= 16'hf57f;
        src7 <= 16'h588e;
        src8 <= 16'h5fa8;
        src9 <= 16'h9ca2;
        src10 <= 16'h7666;
        src11 <= 16'h318d;
        src12 <= 16'h9fb2;
        src13 <= 16'h9872;
        src14 <= 16'he26c;
        src15 <= 16'h10e;
        src16 <= 16'h45b0;
        src17 <= 16'h5fa7;
        src18 <= 16'hd704;
        src19 <= 16'h109d;
        src20 <= 16'h8b1c;
        src21 <= 16'h2a40;
        src22 <= 16'h6acb;
        src23 <= 16'hf481;
        src24 <= 16'h313e;
        src25 <= 16'h931c;
        src26 <= 16'ha3f4;
        src27 <= 16'h3df6;
        src28 <= 16'h210d;
        src29 <= 16'hf9ca;
        src30 <= 16'h6fba;
        src31 <= 16'hd4ee;
        src32 <= 16'h7232;
        src33 <= 16'ha76b;
        src34 <= 16'hb18a;
        src35 <= 16'hb08e;
        src36 <= 16'h76f8;
        src37 <= 16'h8df3;
        src38 <= 16'h1555;
        src39 <= 16'hff9d;
        src40 <= 16'h68ff;
        src41 <= 16'hc542;
        src42 <= 16'h3eb;
        src43 <= 16'hb0f3;
        src44 <= 16'hf1b;
        src45 <= 16'hdd41;
        src46 <= 16'h38d8;
        src47 <= 16'hdd35;
        src48 <= 16'h5906;
        src49 <= 16'h6ba7;
        src50 <= 16'h7bfa;
        src51 <= 16'h6eef;
        src52 <= 16'hbefc;
        src53 <= 16'h3b8f;
        src54 <= 16'h616a;
        src55 <= 16'h7d65;
        src56 <= 16'h6ab0;
        src57 <= 16'h257b;
        src58 <= 16'h229f;
        src59 <= 16'h34e6;
        src60 <= 16'hb0a5;
        src61 <= 16'ha5a2;
        src62 <= 16'hfd7;
        src63 <= 16'heee7;
        src64 <= 16'h7037;
        src65 <= 16'he62;
        src66 <= 16'h49f8;
        src67 <= 16'hd573;
        src68 <= 16'he1f0;
        src69 <= 16'h7b99;
        src70 <= 16'h3853;
        src71 <= 16'hd93e;
        src72 <= 16'h3c08;
        src73 <= 16'hdbb3;
        src74 <= 16'h1c19;
        src75 <= 16'h715c;
        src76 <= 16'h5047;
        src77 <= 16'h7e81;
        src78 <= 16'hf044;
        src79 <= 16'h653b;
        src80 <= 16'h15c4;
        src81 <= 16'hc4df;
        src82 <= 16'h212f;
        src83 <= 16'had9b;
        src84 <= 16'h1107;
        src85 <= 16'hd1f;
        src86 <= 16'h2fc7;
        src87 <= 16'hb379;
        src88 <= 16'h53da;
        src89 <= 16'hfa6d;
        src90 <= 16'h723a;
        src91 <= 16'h8b8f;
        src92 <= 16'h9013;
        src93 <= 16'hc910;
        src94 <= 16'h9597;
        src95 <= 16'hfeb8;
        src96 <= 16'hb88e;
        src97 <= 16'h80dc;
        src98 <= 16'hdbf9;
        src99 <= 16'h4acd;
        src100 <= 16'hee1c;
        src101 <= 16'h9fff;
        src102 <= 16'hdaaf;
        src103 <= 16'h18ac;
        src104 <= 16'ha130;
        src105 <= 16'h2751;
        src106 <= 16'h306c;
        src107 <= 16'h9c94;
        src108 <= 16'h89db;
        src109 <= 16'hcbc6;
        src110 <= 16'h3693;
        src111 <= 16'h9c63;
        src112 <= 16'h5c3c;
        src113 <= 16'h92cf;
        src114 <= 16'h9940;
        src115 <= 16'h24ff;
        src116 <= 16'hd380;
        src117 <= 16'h53c1;
        src118 <= 16'ha051;
        src119 <= 16'hff55;
        src120 <= 16'hca78;
        src121 <= 16'hffe6;
        src122 <= 16'h9e30;
        src123 <= 16'hc20b;
        src124 <= 16'hb20b;
        src125 <= 16'h27c0;
        src126 <= 16'h5bfa;
        src127 <= 16'h12fb;
        exp <= 23'h3f7c97;
        #1
        src0 <= 16'hefa1;
        src1 <= 16'hc08f;
        src2 <= 16'h8177;
        src3 <= 16'h5996;
        src4 <= 16'h815f;
        src5 <= 16'hbb62;
        src6 <= 16'h3d51;
        src7 <= 16'h7ba7;
        src8 <= 16'hf99c;
        src9 <= 16'h252b;
        src10 <= 16'hcebb;
        src11 <= 16'h8eb8;
        src12 <= 16'h193c;
        src13 <= 16'hb6d5;
        src14 <= 16'h407c;
        src15 <= 16'h24ad;
        src16 <= 16'hb89f;
        src17 <= 16'h9214;
        src18 <= 16'h7ee;
        src19 <= 16'h4180;
        src20 <= 16'h9580;
        src21 <= 16'h1712;
        src22 <= 16'hf4f8;
        src23 <= 16'hbc78;
        src24 <= 16'h4b00;
        src25 <= 16'hbc06;
        src26 <= 16'h691d;
        src27 <= 16'h7aae;
        src28 <= 16'hd638;
        src29 <= 16'h7544;
        src30 <= 16'h5959;
        src31 <= 16'hd744;
        src32 <= 16'h588c;
        src33 <= 16'hc2fe;
        src34 <= 16'h257e;
        src35 <= 16'h8fbe;
        src36 <= 16'h7c8c;
        src37 <= 16'hda4e;
        src38 <= 16'hcf71;
        src39 <= 16'h2223;
        src40 <= 16'haffb;
        src41 <= 16'h73d2;
        src42 <= 16'he7d7;
        src43 <= 16'h411e;
        src44 <= 16'hbc73;
        src45 <= 16'hcfd6;
        src46 <= 16'h42f9;
        src47 <= 16'hf42b;
        src48 <= 16'hed64;
        src49 <= 16'hd713;
        src50 <= 16'h8ca6;
        src51 <= 16'hb7b4;
        src52 <= 16'h97b2;
        src53 <= 16'h4401;
        src54 <= 16'h4fc9;
        src55 <= 16'h5a08;
        src56 <= 16'hd7f5;
        src57 <= 16'hb4c2;
        src58 <= 16'h8089;
        src59 <= 16'h70bd;
        src60 <= 16'hbf01;
        src61 <= 16'hce04;
        src62 <= 16'h2714;
        src63 <= 16'h4d3d;
        src64 <= 16'h90cb;
        src65 <= 16'h105;
        src66 <= 16'h1768;
        src67 <= 16'he685;
        src68 <= 16'haac9;
        src69 <= 16'hecae;
        src70 <= 16'he71f;
        src71 <= 16'h8c83;
        src72 <= 16'headd;
        src73 <= 16'h6697;
        src74 <= 16'h6dac;
        src75 <= 16'h399a;
        src76 <= 16'hba25;
        src77 <= 16'h5e33;
        src78 <= 16'h295a;
        src79 <= 16'hed40;
        src80 <= 16'h6597;
        src81 <= 16'h4c9e;
        src82 <= 16'hb60a;
        src83 <= 16'hd7cc;
        src84 <= 16'h77f2;
        src85 <= 16'h8ae5;
        src86 <= 16'ha0fb;
        src87 <= 16'h9c63;
        src88 <= 16'hc908;
        src89 <= 16'hb0c1;
        src90 <= 16'hc6d1;
        src91 <= 16'haa2c;
        src92 <= 16'h7083;
        src93 <= 16'h98e7;
        src94 <= 16'hed35;
        src95 <= 16'hb665;
        src96 <= 16'hd9f8;
        src97 <= 16'h10b1;
        src98 <= 16'hb53e;
        src99 <= 16'h3078;
        src100 <= 16'h6457;
        src101 <= 16'hc5a;
        src102 <= 16'hb29e;
        src103 <= 16'ha507;
        src104 <= 16'h3aff;
        src105 <= 16'h1c3c;
        src106 <= 16'hbf8a;
        src107 <= 16'hf069;
        src108 <= 16'h5c51;
        src109 <= 16'hc2a5;
        src110 <= 16'hf1fe;
        src111 <= 16'h9809;
        src112 <= 16'hd6aa;
        src113 <= 16'ha30f;
        src114 <= 16'h6e96;
        src115 <= 16'h31a1;
        src116 <= 16'h99c1;
        src117 <= 16'ha310;
        src118 <= 16'h5dd0;
        src119 <= 16'h1660;
        src120 <= 16'he9e;
        src121 <= 16'h3c8c;
        src122 <= 16'hc690;
        src123 <= 16'h44c6;
        src124 <= 16'hc756;
        src125 <= 16'hdc6b;
        src126 <= 16'he192;
        src127 <= 16'haec5;
        exp <= 23'h463b77;
        #1
        src0 <= 16'h3012;
        src1 <= 16'he919;
        src2 <= 16'h7977;
        src3 <= 16'h645;
        src4 <= 16'h3fff;
        src5 <= 16'h70a3;
        src6 <= 16'h4abb;
        src7 <= 16'hd5f4;
        src8 <= 16'h70f1;
        src9 <= 16'hf8b6;
        src10 <= 16'h1387;
        src11 <= 16'h115;
        src12 <= 16'haee6;
        src13 <= 16'h6b2;
        src14 <= 16'h8609;
        src15 <= 16'h10ca;
        src16 <= 16'h3bab;
        src17 <= 16'hd7b4;
        src18 <= 16'h2b9;
        src19 <= 16'ha044;
        src20 <= 16'h8ba0;
        src21 <= 16'hf9f2;
        src22 <= 16'h1e4f;
        src23 <= 16'h8b96;
        src24 <= 16'hd929;
        src25 <= 16'h818f;
        src26 <= 16'h2282;
        src27 <= 16'he602;
        src28 <= 16'h756a;
        src29 <= 16'h1922;
        src30 <= 16'h2ea2;
        src31 <= 16'h7ce1;
        src32 <= 16'h2e24;
        src33 <= 16'h52a7;
        src34 <= 16'hd1a3;
        src35 <= 16'h48fd;
        src36 <= 16'h245c;
        src37 <= 16'heebd;
        src38 <= 16'h61b5;
        src39 <= 16'h3c51;
        src40 <= 16'h9f5e;
        src41 <= 16'h188f;
        src42 <= 16'h5ae9;
        src43 <= 16'h1bef;
        src44 <= 16'h97db;
        src45 <= 16'hd850;
        src46 <= 16'h51e1;
        src47 <= 16'h89be;
        src48 <= 16'hd66d;
        src49 <= 16'h9128;
        src50 <= 16'h80f;
        src51 <= 16'ha050;
        src52 <= 16'h31ac;
        src53 <= 16'heaed;
        src54 <= 16'h7c49;
        src55 <= 16'h9008;
        src56 <= 16'h52af;
        src57 <= 16'h169;
        src58 <= 16'h9d75;
        src59 <= 16'h1d8b;
        src60 <= 16'hee3d;
        src61 <= 16'habb4;
        src62 <= 16'h29eb;
        src63 <= 16'hc205;
        src64 <= 16'h6d5c;
        src65 <= 16'hef6d;
        src66 <= 16'h4d77;
        src67 <= 16'he43b;
        src68 <= 16'h4f2a;
        src69 <= 16'hfe63;
        src70 <= 16'hc36e;
        src71 <= 16'ha060;
        src72 <= 16'h2b68;
        src73 <= 16'h7af8;
        src74 <= 16'h3b30;
        src75 <= 16'hb3ab;
        src76 <= 16'h8435;
        src77 <= 16'h96c9;
        src78 <= 16'hcf00;
        src79 <= 16'h8a1e;
        src80 <= 16'h1a09;
        src81 <= 16'hd13c;
        src82 <= 16'h2dd;
        src83 <= 16'hcd95;
        src84 <= 16'h7e36;
        src85 <= 16'h775a;
        src86 <= 16'hf6da;
        src87 <= 16'h3c2f;
        src88 <= 16'h85dc;
        src89 <= 16'hea6e;
        src90 <= 16'h479b;
        src91 <= 16'h475b;
        src92 <= 16'he3da;
        src93 <= 16'h7d6c;
        src94 <= 16'h50f5;
        src95 <= 16'h32f5;
        src96 <= 16'h943a;
        src97 <= 16'h7ccf;
        src98 <= 16'h6a8c;
        src99 <= 16'h80cc;
        src100 <= 16'h7030;
        src101 <= 16'h4cc3;
        src102 <= 16'h5ff;
        src103 <= 16'ha296;
        src104 <= 16'h5695;
        src105 <= 16'h9d22;
        src106 <= 16'h1d80;
        src107 <= 16'hc87a;
        src108 <= 16'h26e1;
        src109 <= 16'he86c;
        src110 <= 16'hd2c5;
        src111 <= 16'h4413;
        src112 <= 16'h17d0;
        src113 <= 16'h6966;
        src114 <= 16'habfc;
        src115 <= 16'hf820;
        src116 <= 16'hda97;
        src117 <= 16'h8f7c;
        src118 <= 16'h66fa;
        src119 <= 16'h5f38;
        src120 <= 16'h2bee;
        src121 <= 16'h60a;
        src122 <= 16'h1695;
        src123 <= 16'h4304;
        src124 <= 16'h27b0;
        src125 <= 16'h18f9;
        src126 <= 16'h675a;
        src127 <= 16'hecc6;
        exp <= 23'h3b3691;
        #1
        src0 <= 16'h2de;
        src1 <= 16'h4988;
        src2 <= 16'he531;
        src3 <= 16'hbe4f;
        src4 <= 16'h7def;
        src5 <= 16'h1371;
        src6 <= 16'hccdc;
        src7 <= 16'h910;
        src8 <= 16'hb14f;
        src9 <= 16'h1ee2;
        src10 <= 16'h14cf;
        src11 <= 16'ha67;
        src12 <= 16'h5017;
        src13 <= 16'h9923;
        src14 <= 16'hb592;
        src15 <= 16'hfd90;
        src16 <= 16'hf4e0;
        src17 <= 16'h5617;
        src18 <= 16'h281e;
        src19 <= 16'h55cb;
        src20 <= 16'hfe52;
        src21 <= 16'hab70;
        src22 <= 16'h5792;
        src23 <= 16'h3be0;
        src24 <= 16'hdac2;
        src25 <= 16'h90a3;
        src26 <= 16'h29b7;
        src27 <= 16'hc832;
        src28 <= 16'h2465;
        src29 <= 16'h5f0b;
        src30 <= 16'hb53;
        src31 <= 16'hf858;
        src32 <= 16'h1601;
        src33 <= 16'h2866;
        src34 <= 16'ha8d7;
        src35 <= 16'h40f7;
        src36 <= 16'h39d6;
        src37 <= 16'hce3b;
        src38 <= 16'h2ff9;
        src39 <= 16'h308d;
        src40 <= 16'hb9dd;
        src41 <= 16'h2ab5;
        src42 <= 16'h4214;
        src43 <= 16'h180;
        src44 <= 16'hbe1;
        src45 <= 16'hecec;
        src46 <= 16'h308;
        src47 <= 16'h5fcf;
        src48 <= 16'hb40b;
        src49 <= 16'h7bdf;
        src50 <= 16'h764b;
        src51 <= 16'h1ca7;
        src52 <= 16'hbfa8;
        src53 <= 16'h8e30;
        src54 <= 16'h95c2;
        src55 <= 16'h459a;
        src56 <= 16'ha612;
        src57 <= 16'hc28f;
        src58 <= 16'h3ebc;
        src59 <= 16'h7a71;
        src60 <= 16'hca1b;
        src61 <= 16'hc898;
        src62 <= 16'h6698;
        src63 <= 16'h7ec9;
        src64 <= 16'h4c1d;
        src65 <= 16'h7f19;
        src66 <= 16'hab7c;
        src67 <= 16'h659a;
        src68 <= 16'he629;
        src69 <= 16'h304c;
        src70 <= 16'hcca8;
        src71 <= 16'h700b;
        src72 <= 16'h1dfe;
        src73 <= 16'h4496;
        src74 <= 16'hff02;
        src75 <= 16'hd48c;
        src76 <= 16'hefba;
        src77 <= 16'h6789;
        src78 <= 16'h63cb;
        src79 <= 16'hce84;
        src80 <= 16'h1987;
        src81 <= 16'h50c;
        src82 <= 16'h311e;
        src83 <= 16'haec4;
        src84 <= 16'h479;
        src85 <= 16'hca62;
        src86 <= 16'hd4f0;
        src87 <= 16'hca6c;
        src88 <= 16'hda2b;
        src89 <= 16'hf99b;
        src90 <= 16'hcf24;
        src91 <= 16'hea8f;
        src92 <= 16'h22f0;
        src93 <= 16'h1196;
        src94 <= 16'h483f;
        src95 <= 16'h2862;
        src96 <= 16'h74dd;
        src97 <= 16'h86da;
        src98 <= 16'heaa2;
        src99 <= 16'hd516;
        src100 <= 16'hc301;
        src101 <= 16'h583b;
        src102 <= 16'hf93f;
        src103 <= 16'he3a;
        src104 <= 16'h74eb;
        src105 <= 16'hf68d;
        src106 <= 16'hc960;
        src107 <= 16'hbd60;
        src108 <= 16'hb7c1;
        src109 <= 16'h91b;
        src110 <= 16'h2cbd;
        src111 <= 16'hb1f6;
        src112 <= 16'h92c9;
        src113 <= 16'h1cf;
        src114 <= 16'h20d6;
        src115 <= 16'h6a6;
        src116 <= 16'h3f30;
        src117 <= 16'h6c32;
        src118 <= 16'h41f7;
        src119 <= 16'hed1b;
        src120 <= 16'h6792;
        src121 <= 16'hd9bd;
        src122 <= 16'h97df;
        src123 <= 16'h6b3;
        src124 <= 16'h777f;
        src125 <= 16'h7b8a;
        src126 <= 16'hb7ec;
        src127 <= 16'h3d4b;
        exp <= 23'h3cc502;
        #1
        src0 <= 16'hcffa;
        src1 <= 16'h5939;
        src2 <= 16'hf1c7;
        src3 <= 16'hfcae;
        src4 <= 16'h12aa;
        src5 <= 16'ha297;
        src6 <= 16'heed3;
        src7 <= 16'hd5b;
        src8 <= 16'h194e;
        src9 <= 16'h5497;
        src10 <= 16'h4bf3;
        src11 <= 16'hfcc4;
        src12 <= 16'hdeea;
        src13 <= 16'h557;
        src14 <= 16'h20e;
        src15 <= 16'h5fd;
        src16 <= 16'h2084;
        src17 <= 16'hb741;
        src18 <= 16'h4f87;
        src19 <= 16'h9f6e;
        src20 <= 16'h339d;
        src21 <= 16'h40c8;
        src22 <= 16'h6c8;
        src23 <= 16'h8d13;
        src24 <= 16'h864b;
        src25 <= 16'h944c;
        src26 <= 16'h3746;
        src27 <= 16'h6b84;
        src28 <= 16'he99d;
        src29 <= 16'he7b5;
        src30 <= 16'h9acf;
        src31 <= 16'hb6e4;
        src32 <= 16'hcf50;
        src33 <= 16'hccd9;
        src34 <= 16'h75f3;
        src35 <= 16'hdcd;
        src36 <= 16'hdb74;
        src37 <= 16'h1f9a;
        src38 <= 16'hcdeb;
        src39 <= 16'h4a88;
        src40 <= 16'hd6e1;
        src41 <= 16'he35d;
        src42 <= 16'h88d8;
        src43 <= 16'h6382;
        src44 <= 16'h1eab;
        src45 <= 16'h5d23;
        src46 <= 16'h7cd7;
        src47 <= 16'hdac1;
        src48 <= 16'h240b;
        src49 <= 16'haf5c;
        src50 <= 16'h5bd6;
        src51 <= 16'hf35c;
        src52 <= 16'h2f5b;
        src53 <= 16'h8936;
        src54 <= 16'h4b1f;
        src55 <= 16'hd8f5;
        src56 <= 16'h5bb5;
        src57 <= 16'hbf;
        src58 <= 16'h50a1;
        src59 <= 16'ha11d;
        src60 <= 16'h719f;
        src61 <= 16'h403f;
        src62 <= 16'hb517;
        src63 <= 16'hd954;
        src64 <= 16'h3076;
        src65 <= 16'h3ed0;
        src66 <= 16'h304c;
        src67 <= 16'hddf;
        src68 <= 16'h8546;
        src69 <= 16'h615f;
        src70 <= 16'h9bfb;
        src71 <= 16'h5ed7;
        src72 <= 16'hc156;
        src73 <= 16'h7aa4;
        src74 <= 16'hf64a;
        src75 <= 16'h2d58;
        src76 <= 16'hff22;
        src77 <= 16'hbf19;
        src78 <= 16'h2d77;
        src79 <= 16'h9024;
        src80 <= 16'h9004;
        src81 <= 16'ha671;
        src82 <= 16'h2a01;
        src83 <= 16'hc0e2;
        src84 <= 16'hcdb3;
        src85 <= 16'h292b;
        src86 <= 16'h2d65;
        src87 <= 16'ha93;
        src88 <= 16'hbf36;
        src89 <= 16'h178c;
        src90 <= 16'hb58b;
        src91 <= 16'hb7a9;
        src92 <= 16'h261a;
        src93 <= 16'ha08e;
        src94 <= 16'h9136;
        src95 <= 16'hc4a2;
        src96 <= 16'h7cfe;
        src97 <= 16'hea09;
        src98 <= 16'h830a;
        src99 <= 16'h54e0;
        src100 <= 16'h5d6e;
        src101 <= 16'hc914;
        src102 <= 16'h4242;
        src103 <= 16'hcd02;
        src104 <= 16'h57c9;
        src105 <= 16'h4b30;
        src106 <= 16'hc9bc;
        src107 <= 16'hc3fb;
        src108 <= 16'haaeb;
        src109 <= 16'h47b8;
        src110 <= 16'hec52;
        src111 <= 16'h7932;
        src112 <= 16'h2a8f;
        src113 <= 16'he447;
        src114 <= 16'hafd3;
        src115 <= 16'h4369;
        src116 <= 16'h8d8d;
        src117 <= 16'h7d1c;
        src118 <= 16'h270b;
        src119 <= 16'h760f;
        src120 <= 16'h839d;
        src121 <= 16'h4e31;
        src122 <= 16'h148c;
        src123 <= 16'hddc0;
        src124 <= 16'h76b5;
        src125 <= 16'he82c;
        src126 <= 16'h2181;
        src127 <= 16'ha3b3;
        exp <= 23'h3f0110;
        #1
        src0 <= 16'h932e;
        src1 <= 16'hc6be;
        src2 <= 16'h2d78;
        src3 <= 16'h181a;
        src4 <= 16'hc695;
        src5 <= 16'hde8d;
        src6 <= 16'h1396;
        src7 <= 16'h59d3;
        src8 <= 16'hf94;
        src9 <= 16'h2b55;
        src10 <= 16'h249c;
        src11 <= 16'h15fa;
        src12 <= 16'h3f7b;
        src13 <= 16'h3923;
        src14 <= 16'h3898;
        src15 <= 16'h796f;
        src16 <= 16'h3b32;
        src17 <= 16'he5b6;
        src18 <= 16'h486e;
        src19 <= 16'ha0bc;
        src20 <= 16'h47fb;
        src21 <= 16'h5d45;
        src22 <= 16'hfb7c;
        src23 <= 16'h38fa;
        src24 <= 16'hfe44;
        src25 <= 16'h4744;
        src26 <= 16'h10f;
        src27 <= 16'hd198;
        src28 <= 16'h2902;
        src29 <= 16'h679a;
        src30 <= 16'h526e;
        src31 <= 16'h2bc8;
        src32 <= 16'h7fd4;
        src33 <= 16'hb8b7;
        src34 <= 16'h30a7;
        src35 <= 16'h3211;
        src36 <= 16'h7e57;
        src37 <= 16'ha850;
        src38 <= 16'h144c;
        src39 <= 16'h987f;
        src40 <= 16'hd9d9;
        src41 <= 16'h1b89;
        src42 <= 16'hcc27;
        src43 <= 16'h3608;
        src44 <= 16'h686c;
        src45 <= 16'h308;
        src46 <= 16'hb191;
        src47 <= 16'hacaf;
        src48 <= 16'h2b10;
        src49 <= 16'hb11b;
        src50 <= 16'h70fd;
        src51 <= 16'h95d7;
        src52 <= 16'h1528;
        src53 <= 16'h6138;
        src54 <= 16'head7;
        src55 <= 16'hebcc;
        src56 <= 16'h4034;
        src57 <= 16'ha20a;
        src58 <= 16'h29a9;
        src59 <= 16'hf518;
        src60 <= 16'hb552;
        src61 <= 16'ha0d7;
        src62 <= 16'hef29;
        src63 <= 16'h1a3b;
        src64 <= 16'h1c66;
        src65 <= 16'h84d;
        src66 <= 16'h616;
        src67 <= 16'h39c0;
        src68 <= 16'h2fc4;
        src69 <= 16'h774;
        src70 <= 16'h6ad4;
        src71 <= 16'ha7e9;
        src72 <= 16'h87ed;
        src73 <= 16'h57a2;
        src74 <= 16'hbc9;
        src75 <= 16'ha17b;
        src76 <= 16'h372d;
        src77 <= 16'hafed;
        src78 <= 16'hc3e1;
        src79 <= 16'h982f;
        src80 <= 16'h1779;
        src81 <= 16'hb766;
        src82 <= 16'h97a8;
        src83 <= 16'h6a5f;
        src84 <= 16'he82f;
        src85 <= 16'h3258;
        src86 <= 16'hd3;
        src87 <= 16'hfc6c;
        src88 <= 16'hf17e;
        src89 <= 16'hd3d2;
        src90 <= 16'hfa75;
        src91 <= 16'h2d7f;
        src92 <= 16'h2306;
        src93 <= 16'hb171;
        src94 <= 16'hb8ae;
        src95 <= 16'hec64;
        src96 <= 16'h5a59;
        src97 <= 16'hf51d;
        src98 <= 16'hf255;
        src99 <= 16'ha985;
        src100 <= 16'h828b;
        src101 <= 16'h5dc2;
        src102 <= 16'h3daf;
        src103 <= 16'h68ea;
        src104 <= 16'h45f1;
        src105 <= 16'h24f4;
        src106 <= 16'h4378;
        src107 <= 16'hcc98;
        src108 <= 16'h77d1;
        src109 <= 16'ha806;
        src110 <= 16'h7db6;
        src111 <= 16'hcef8;
        src112 <= 16'hd750;
        src113 <= 16'h93d6;
        src114 <= 16'hec1d;
        src115 <= 16'h8ecf;
        src116 <= 16'hc141;
        src117 <= 16'h355c;
        src118 <= 16'hb301;
        src119 <= 16'haccb;
        src120 <= 16'h8a72;
        src121 <= 16'h1649;
        src122 <= 16'hcc30;
        src123 <= 16'haa67;
        src124 <= 16'h4057;
        src125 <= 16'h9496;
        src126 <= 16'hfacd;
        src127 <= 16'h99c5;
        exp <= 23'h3d026e;
        #1
        src0 <= 16'h4686;
        src1 <= 16'hbd27;
        src2 <= 16'h1597;
        src3 <= 16'h8cd8;
        src4 <= 16'h956d;
        src5 <= 16'h56ad;
        src6 <= 16'hac16;
        src7 <= 16'hf5f3;
        src8 <= 16'hfc47;
        src9 <= 16'h1b20;
        src10 <= 16'h73e2;
        src11 <= 16'hed6d;
        src12 <= 16'hc408;
        src13 <= 16'hd099;
        src14 <= 16'ha7e2;
        src15 <= 16'hf8c3;
        src16 <= 16'h4b57;
        src17 <= 16'h12b;
        src18 <= 16'h6e7e;
        src19 <= 16'hb0d1;
        src20 <= 16'h347e;
        src21 <= 16'hc373;
        src22 <= 16'h3a21;
        src23 <= 16'h7b12;
        src24 <= 16'he97;
        src25 <= 16'he23f;
        src26 <= 16'h86af;
        src27 <= 16'h71f9;
        src28 <= 16'h550d;
        src29 <= 16'ha21b;
        src30 <= 16'he1ec;
        src31 <= 16'h9269;
        src32 <= 16'hf466;
        src33 <= 16'h4126;
        src34 <= 16'h7659;
        src35 <= 16'h71d7;
        src36 <= 16'h1265;
        src37 <= 16'h62c9;
        src38 <= 16'h4944;
        src39 <= 16'he3b2;
        src40 <= 16'hf365;
        src41 <= 16'ha130;
        src42 <= 16'hf304;
        src43 <= 16'h4e18;
        src44 <= 16'h5252;
        src45 <= 16'h634;
        src46 <= 16'h2b6;
        src47 <= 16'h391c;
        src48 <= 16'hd7c1;
        src49 <= 16'h2c6a;
        src50 <= 16'h88ff;
        src51 <= 16'hbbd3;
        src52 <= 16'h5c28;
        src53 <= 16'hf6f0;
        src54 <= 16'h79df;
        src55 <= 16'hc4c;
        src56 <= 16'h3867;
        src57 <= 16'hfc99;
        src58 <= 16'hf762;
        src59 <= 16'h677b;
        src60 <= 16'h439e;
        src61 <= 16'haee0;
        src62 <= 16'h1ad9;
        src63 <= 16'hc65c;
        src64 <= 16'hb005;
        src65 <= 16'h619b;
        src66 <= 16'hd08f;
        src67 <= 16'hf7ab;
        src68 <= 16'hfcc4;
        src69 <= 16'h6d17;
        src70 <= 16'hf29b;
        src71 <= 16'h8ed0;
        src72 <= 16'h2730;
        src73 <= 16'h7046;
        src74 <= 16'h433d;
        src75 <= 16'h96b9;
        src76 <= 16'h4637;
        src77 <= 16'h7021;
        src78 <= 16'h46fc;
        src79 <= 16'h309;
        src80 <= 16'hcf4e;
        src81 <= 16'habed;
        src82 <= 16'hbce2;
        src83 <= 16'h255e;
        src84 <= 16'he247;
        src85 <= 16'h315d;
        src86 <= 16'hdde0;
        src87 <= 16'h1188;
        src88 <= 16'h947c;
        src89 <= 16'hf303;
        src90 <= 16'h1030;
        src91 <= 16'hbb49;
        src92 <= 16'hbc57;
        src93 <= 16'hcb0;
        src94 <= 16'h599f;
        src95 <= 16'ha5f1;
        src96 <= 16'hef3c;
        src97 <= 16'h2a59;
        src98 <= 16'h6cec;
        src99 <= 16'hd4d6;
        src100 <= 16'h9ab7;
        src101 <= 16'hc0eb;
        src102 <= 16'h4e89;
        src103 <= 16'hb808;
        src104 <= 16'h2735;
        src105 <= 16'hf9b2;
        src106 <= 16'haf1b;
        src107 <= 16'hb489;
        src108 <= 16'ha762;
        src109 <= 16'hba86;
        src110 <= 16'h1f12;
        src111 <= 16'hce6a;
        src112 <= 16'hd483;
        src113 <= 16'h59f8;
        src114 <= 16'h1fa9;
        src115 <= 16'h140;
        src116 <= 16'h5b0c;
        src117 <= 16'h27d6;
        src118 <= 16'h47ab;
        src119 <= 16'h17d4;
        src120 <= 16'h70c4;
        src121 <= 16'h2ab6;
        src122 <= 16'h75b7;
        src123 <= 16'h358d;
        src124 <= 16'h332f;
        src125 <= 16'h5a4;
        src126 <= 16'h4af0;
        src127 <= 16'h9233;
        exp <= 23'h3fd6d5;
        #1
        src0 <= 16'h5ff0;
        src1 <= 16'hd3ac;
        src2 <= 16'hbd73;
        src3 <= 16'h888e;
        src4 <= 16'h8f9e;
        src5 <= 16'h5b2d;
        src6 <= 16'h13da;
        src7 <= 16'hefa5;
        src8 <= 16'hc1bb;
        src9 <= 16'h9f98;
        src10 <= 16'h9853;
        src11 <= 16'h7b07;
        src12 <= 16'hc882;
        src13 <= 16'h5a30;
        src14 <= 16'h30ed;
        src15 <= 16'hed25;
        src16 <= 16'hd789;
        src17 <= 16'hf990;
        src18 <= 16'h276;
        src19 <= 16'he99e;
        src20 <= 16'h88d2;
        src21 <= 16'hd8b3;
        src22 <= 16'ha1ad;
        src23 <= 16'h3fde;
        src24 <= 16'h9a5b;
        src25 <= 16'h2768;
        src26 <= 16'he893;
        src27 <= 16'h8492;
        src28 <= 16'h1df3;
        src29 <= 16'he62a;
        src30 <= 16'hf429;
        src31 <= 16'h9da1;
        src32 <= 16'h8232;
        src33 <= 16'hbc76;
        src34 <= 16'h7b4a;
        src35 <= 16'h2b5e;
        src36 <= 16'h3f58;
        src37 <= 16'h91d4;
        src38 <= 16'h4498;
        src39 <= 16'hf594;
        src40 <= 16'h1931;
        src41 <= 16'h5a87;
        src42 <= 16'hf55a;
        src43 <= 16'hef3c;
        src44 <= 16'h1c52;
        src45 <= 16'h2475;
        src46 <= 16'h4dad;
        src47 <= 16'h7fea;
        src48 <= 16'h89bb;
        src49 <= 16'hb1d9;
        src50 <= 16'hf675;
        src51 <= 16'hb28c;
        src52 <= 16'hc5a5;
        src53 <= 16'h958c;
        src54 <= 16'h890a;
        src55 <= 16'h92ec;
        src56 <= 16'hfdc9;
        src57 <= 16'hdf12;
        src58 <= 16'hf3ff;
        src59 <= 16'hfafe;
        src60 <= 16'h97d2;
        src61 <= 16'hb42f;
        src62 <= 16'hc598;
        src63 <= 16'h1325;
        src64 <= 16'h7a7d;
        src65 <= 16'h4a97;
        src66 <= 16'h6e8e;
        src67 <= 16'hcbf9;
        src68 <= 16'h2f20;
        src69 <= 16'hc02a;
        src70 <= 16'h3f6c;
        src71 <= 16'h3917;
        src72 <= 16'hbeed;
        src73 <= 16'haa9b;
        src74 <= 16'he6fa;
        src75 <= 16'hca14;
        src76 <= 16'hbbfe;
        src77 <= 16'hf760;
        src78 <= 16'h2c72;
        src79 <= 16'h9383;
        src80 <= 16'hf14f;
        src81 <= 16'hf03c;
        src82 <= 16'he5b0;
        src83 <= 16'hb865;
        src84 <= 16'h7cd1;
        src85 <= 16'h8573;
        src86 <= 16'hbafc;
        src87 <= 16'he4f9;
        src88 <= 16'hf692;
        src89 <= 16'h7a0f;
        src90 <= 16'h4329;
        src91 <= 16'h9f3c;
        src92 <= 16'he53;
        src93 <= 16'h83d0;
        src94 <= 16'hde6a;
        src95 <= 16'h61ac;
        src96 <= 16'h63ce;
        src97 <= 16'h2faf;
        src98 <= 16'h72ff;
        src99 <= 16'h14a3;
        src100 <= 16'h86eb;
        src101 <= 16'h659d;
        src102 <= 16'h15f;
        src103 <= 16'h1bcb;
        src104 <= 16'ha745;
        src105 <= 16'h4808;
        src106 <= 16'h8d08;
        src107 <= 16'hf046;
        src108 <= 16'he231;
        src109 <= 16'hff8;
        src110 <= 16'he56d;
        src111 <= 16'h5e24;
        src112 <= 16'hd387;
        src113 <= 16'he0a5;
        src114 <= 16'h946f;
        src115 <= 16'h770f;
        src116 <= 16'h1dfb;
        src117 <= 16'h8a67;
        src118 <= 16'h651;
        src119 <= 16'h1b4d;
        src120 <= 16'h56f6;
        src121 <= 16'h3bc;
        src122 <= 16'h725c;
        src123 <= 16'h1193;
        src124 <= 16'h9af8;
        src125 <= 16'h839c;
        src126 <= 16'h44aa;
        src127 <= 16'h2c2f;
        exp <= 23'h458151;
        #1
        src0 <= 16'hbe0f;
        src1 <= 16'h94b0;
        src2 <= 16'h84b9;
        src3 <= 16'he65;
        src4 <= 16'h6d7f;
        src5 <= 16'h80d3;
        src6 <= 16'hba76;
        src7 <= 16'hb5bf;
        src8 <= 16'h9741;
        src9 <= 16'h272e;
        src10 <= 16'h54ca;
        src11 <= 16'ha01;
        src12 <= 16'h923;
        src13 <= 16'haf8d;
        src14 <= 16'h606a;
        src15 <= 16'h5d70;
        src16 <= 16'hee4b;
        src17 <= 16'h987e;
        src18 <= 16'ha5d;
        src19 <= 16'h2dcf;
        src20 <= 16'h18c9;
        src21 <= 16'h51a0;
        src22 <= 16'h19a8;
        src23 <= 16'h6fb0;
        src24 <= 16'hcfbc;
        src25 <= 16'h48b5;
        src26 <= 16'h93;
        src27 <= 16'hbc7e;
        src28 <= 16'h690e;
        src29 <= 16'hbb93;
        src30 <= 16'hb50c;
        src31 <= 16'h2f1a;
        src32 <= 16'h4e00;
        src33 <= 16'hedf0;
        src34 <= 16'h4ceb;
        src35 <= 16'hd818;
        src36 <= 16'ha3f1;
        src37 <= 16'h0;
        src38 <= 16'hb0ed;
        src39 <= 16'h3263;
        src40 <= 16'h90dc;
        src41 <= 16'hbd66;
        src42 <= 16'h4b3;
        src43 <= 16'h2e50;
        src44 <= 16'h2e82;
        src45 <= 16'hb1c7;
        src46 <= 16'he7b3;
        src47 <= 16'h9951;
        src48 <= 16'h8717;
        src49 <= 16'h4cfa;
        src50 <= 16'h2345;
        src51 <= 16'hb041;
        src52 <= 16'h6f2;
        src53 <= 16'h54e9;
        src54 <= 16'h6be;
        src55 <= 16'h55e0;
        src56 <= 16'hef8f;
        src57 <= 16'hbee5;
        src58 <= 16'hbc82;
        src59 <= 16'hcb;
        src60 <= 16'h85dd;
        src61 <= 16'hb59f;
        src62 <= 16'h799b;
        src63 <= 16'ha0a6;
        src64 <= 16'ha493;
        src65 <= 16'hc01c;
        src66 <= 16'h682e;
        src67 <= 16'heef0;
        src68 <= 16'hfedf;
        src69 <= 16'h7b9b;
        src70 <= 16'h9425;
        src71 <= 16'h50dc;
        src72 <= 16'h971f;
        src73 <= 16'hcaff;
        src74 <= 16'ha6ed;
        src75 <= 16'h5b01;
        src76 <= 16'he17e;
        src77 <= 16'ha534;
        src78 <= 16'h4ab7;
        src79 <= 16'hd7f9;
        src80 <= 16'hd329;
        src81 <= 16'h9804;
        src82 <= 16'h43be;
        src83 <= 16'h861e;
        src84 <= 16'h6502;
        src85 <= 16'hcdbc;
        src86 <= 16'h7998;
        src87 <= 16'h9326;
        src88 <= 16'hf383;
        src89 <= 16'h71cd;
        src90 <= 16'hac1f;
        src91 <= 16'haad8;
        src92 <= 16'h88c0;
        src93 <= 16'h64ba;
        src94 <= 16'h3ab7;
        src95 <= 16'ha45e;
        src96 <= 16'hd274;
        src97 <= 16'h9f5d;
        src98 <= 16'h6e;
        src99 <= 16'h7f6d;
        src100 <= 16'hdd96;
        src101 <= 16'h59e5;
        src102 <= 16'h91a6;
        src103 <= 16'h965d;
        src104 <= 16'h140a;
        src105 <= 16'h81f7;
        src106 <= 16'hbe4;
        src107 <= 16'hffd4;
        src108 <= 16'h77a1;
        src109 <= 16'ha7ba;
        src110 <= 16'h6b5d;
        src111 <= 16'hdb16;
        src112 <= 16'h1183;
        src113 <= 16'hb95d;
        src114 <= 16'had46;
        src115 <= 16'hde79;
        src116 <= 16'h1cab;
        src117 <= 16'h65c2;
        src118 <= 16'hfac2;
        src119 <= 16'h53a9;
        src120 <= 16'hf3ef;
        src121 <= 16'h856b;
        src122 <= 16'h2036;
        src123 <= 16'h4bba;
        src124 <= 16'h828;
        src125 <= 16'hee9;
        src126 <= 16'h9cd3;
        src127 <= 16'h579a;
        exp <= 23'h3eec7c;
        #1
        src0 <= 16'h5014;
        src1 <= 16'h6aa;
        src2 <= 16'had5;
        src3 <= 16'ha08d;
        src4 <= 16'hf02e;
        src5 <= 16'h3e5d;
        src6 <= 16'hb2b6;
        src7 <= 16'hd428;
        src8 <= 16'hef02;
        src9 <= 16'hd198;
        src10 <= 16'hffc7;
        src11 <= 16'hb62c;
        src12 <= 16'h94a8;
        src13 <= 16'h83a3;
        src14 <= 16'h8116;
        src15 <= 16'h6957;
        src16 <= 16'h74a4;
        src17 <= 16'h903c;
        src18 <= 16'h73ed;
        src19 <= 16'hf670;
        src20 <= 16'h8c40;
        src21 <= 16'h375;
        src22 <= 16'h1389;
        src23 <= 16'he78b;
        src24 <= 16'h2c12;
        src25 <= 16'h25ae;
        src26 <= 16'h4a74;
        src27 <= 16'h1b5e;
        src28 <= 16'h8139;
        src29 <= 16'hf893;
        src30 <= 16'hddfc;
        src31 <= 16'hf94e;
        src32 <= 16'h38fe;
        src33 <= 16'hc180;
        src34 <= 16'hb50e;
        src35 <= 16'h7317;
        src36 <= 16'h8180;
        src37 <= 16'hfc57;
        src38 <= 16'he7fc;
        src39 <= 16'h3b93;
        src40 <= 16'h18b3;
        src41 <= 16'h1cbb;
        src42 <= 16'he383;
        src43 <= 16'h90c5;
        src44 <= 16'h8e4b;
        src45 <= 16'h344;
        src46 <= 16'h7f10;
        src47 <= 16'h974b;
        src48 <= 16'hbf24;
        src49 <= 16'he45b;
        src50 <= 16'h598d;
        src51 <= 16'h7a78;
        src52 <= 16'hc14;
        src53 <= 16'h6dfe;
        src54 <= 16'h3af;
        src55 <= 16'haf0b;
        src56 <= 16'h94ce;
        src57 <= 16'h7c05;
        src58 <= 16'hf174;
        src59 <= 16'h207b;
        src60 <= 16'he80d;
        src61 <= 16'hc91a;
        src62 <= 16'h1c28;
        src63 <= 16'h75dc;
        src64 <= 16'h26b1;
        src65 <= 16'hb1e;
        src66 <= 16'h29e7;
        src67 <= 16'hcec1;
        src68 <= 16'h7d0b;
        src69 <= 16'h3bba;
        src70 <= 16'hc18c;
        src71 <= 16'h77ec;
        src72 <= 16'h8d6f;
        src73 <= 16'hce17;
        src74 <= 16'h94d6;
        src75 <= 16'hf5ce;
        src76 <= 16'hb877;
        src77 <= 16'hc50c;
        src78 <= 16'h9761;
        src79 <= 16'h3b57;
        src80 <= 16'h8cc9;
        src81 <= 16'hc741;
        src82 <= 16'hbf9f;
        src83 <= 16'h1d82;
        src84 <= 16'h6faf;
        src85 <= 16'h8712;
        src86 <= 16'h6740;
        src87 <= 16'ha4e1;
        src88 <= 16'h966d;
        src89 <= 16'hca19;
        src90 <= 16'h2a8;
        src91 <= 16'h8d48;
        src92 <= 16'h497;
        src93 <= 16'h3b29;
        src94 <= 16'h2bcc;
        src95 <= 16'hfc8c;
        src96 <= 16'h9333;
        src97 <= 16'he1bd;
        src98 <= 16'h2278;
        src99 <= 16'hcf99;
        src100 <= 16'hec5d;
        src101 <= 16'hf3d0;
        src102 <= 16'h9a4a;
        src103 <= 16'h1d9;
        src104 <= 16'ha31a;
        src105 <= 16'h508c;
        src106 <= 16'hdf56;
        src107 <= 16'h1c6;
        src108 <= 16'hc2c6;
        src109 <= 16'hddfc;
        src110 <= 16'h5c2c;
        src111 <= 16'hf22b;
        src112 <= 16'h3bae;
        src113 <= 16'h1217;
        src114 <= 16'haf7b;
        src115 <= 16'he7db;
        src116 <= 16'hfa52;
        src117 <= 16'h8f45;
        src118 <= 16'h87b7;
        src119 <= 16'h42f7;
        src120 <= 16'hba0f;
        src121 <= 16'h7b58;
        src122 <= 16'hea31;
        src123 <= 16'h9d80;
        src124 <= 16'h69ee;
        src125 <= 16'h2e44;
        src126 <= 16'hd645;
        src127 <= 16'h93ed;
        exp <= 23'h43d31e;
        #1
        src0 <= 16'h86e2;
        src1 <= 16'hc89;
        src2 <= 16'h9ba8;
        src3 <= 16'hcc8a;
        src4 <= 16'h30d4;
        src5 <= 16'h7b0b;
        src6 <= 16'hee5f;
        src7 <= 16'h2eea;
        src8 <= 16'hce31;
        src9 <= 16'h7f6c;
        src10 <= 16'h49da;
        src11 <= 16'h7437;
        src12 <= 16'h65f8;
        src13 <= 16'h61fc;
        src14 <= 16'h57f5;
        src15 <= 16'h7a1;
        src16 <= 16'hda88;
        src17 <= 16'hc48a;
        src18 <= 16'hd0de;
        src19 <= 16'h902b;
        src20 <= 16'h7579;
        src21 <= 16'hb136;
        src22 <= 16'ha47b;
        src23 <= 16'hdc4f;
        src24 <= 16'h3e47;
        src25 <= 16'hd586;
        src26 <= 16'haf9f;
        src27 <= 16'he43d;
        src28 <= 16'ha1f0;
        src29 <= 16'hc601;
        src30 <= 16'hdcbf;
        src31 <= 16'hbaf7;
        src32 <= 16'h732e;
        src33 <= 16'h6ef7;
        src34 <= 16'had6f;
        src35 <= 16'hafa3;
        src36 <= 16'h5881;
        src37 <= 16'h1c0a;
        src38 <= 16'hdb9;
        src39 <= 16'h2e5d;
        src40 <= 16'hee9;
        src41 <= 16'h2b6f;
        src42 <= 16'hed77;
        src43 <= 16'h8ae8;
        src44 <= 16'h2aa;
        src45 <= 16'h1223;
        src46 <= 16'h2127;
        src47 <= 16'h1125;
        src48 <= 16'h7b0e;
        src49 <= 16'h5deb;
        src50 <= 16'hdc;
        src51 <= 16'hb48b;
        src52 <= 16'h5533;
        src53 <= 16'h5bc6;
        src54 <= 16'h7ddc;
        src55 <= 16'h246f;
        src56 <= 16'h1a0;
        src57 <= 16'h8ad7;
        src58 <= 16'hbd03;
        src59 <= 16'h9c5c;
        src60 <= 16'h9f75;
        src61 <= 16'h7ea7;
        src62 <= 16'h6d;
        src63 <= 16'h9a99;
        src64 <= 16'hd946;
        src65 <= 16'hae58;
        src66 <= 16'h3253;
        src67 <= 16'h43a2;
        src68 <= 16'hddeb;
        src69 <= 16'h7f10;
        src70 <= 16'h3808;
        src71 <= 16'h5975;
        src72 <= 16'hf250;
        src73 <= 16'h5449;
        src74 <= 16'h3e75;
        src75 <= 16'h18e4;
        src76 <= 16'hc1bd;
        src77 <= 16'h2a77;
        src78 <= 16'hbfc7;
        src79 <= 16'h6d8a;
        src80 <= 16'hc041;
        src81 <= 16'hb131;
        src82 <= 16'hdaba;
        src83 <= 16'h2c13;
        src84 <= 16'hd9ce;
        src85 <= 16'h1512;
        src86 <= 16'h5c50;
        src87 <= 16'h9b4a;
        src88 <= 16'hfca;
        src89 <= 16'hde8c;
        src90 <= 16'h54a;
        src91 <= 16'h56b5;
        src92 <= 16'h4bdf;
        src93 <= 16'ha9f6;
        src94 <= 16'hfe08;
        src95 <= 16'hf712;
        src96 <= 16'hffd4;
        src97 <= 16'h42ba;
        src98 <= 16'h3c63;
        src99 <= 16'h13b0;
        src100 <= 16'h44e6;
        src101 <= 16'h9f4e;
        src102 <= 16'hc153;
        src103 <= 16'h660;
        src104 <= 16'hd78f;
        src105 <= 16'he55f;
        src106 <= 16'h5af5;
        src107 <= 16'hb85f;
        src108 <= 16'h59e8;
        src109 <= 16'h1560;
        src110 <= 16'hda5a;
        src111 <= 16'h9f;
        src112 <= 16'hb9ae;
        src113 <= 16'hcbde;
        src114 <= 16'hf9e2;
        src115 <= 16'he987;
        src116 <= 16'h14d1;
        src117 <= 16'h2af1;
        src118 <= 16'hfbe6;
        src119 <= 16'h4208;
        src120 <= 16'he777;
        src121 <= 16'h5e52;
        src122 <= 16'hb8e;
        src123 <= 16'h45ed;
        src124 <= 16'h8945;
        src125 <= 16'h7f6a;
        src126 <= 16'h9120;
        src127 <= 16'h86c3;
        exp <= 23'h3de02a;
        #1
        src0 <= 16'he2ef;
        src1 <= 16'h2a15;
        src2 <= 16'hbbdf;
        src3 <= 16'h6289;
        src4 <= 16'h5bac;
        src5 <= 16'h9fa2;
        src6 <= 16'h33fc;
        src7 <= 16'h409a;
        src8 <= 16'h103e;
        src9 <= 16'hcc68;
        src10 <= 16'hb109;
        src11 <= 16'h8a8e;
        src12 <= 16'h631d;
        src13 <= 16'h2cbc;
        src14 <= 16'hc239;
        src15 <= 16'hebf7;
        src16 <= 16'h4b1d;
        src17 <= 16'h9c63;
        src18 <= 16'h3e5d;
        src19 <= 16'h7cd7;
        src20 <= 16'hb64c;
        src21 <= 16'hbeea;
        src22 <= 16'hc30b;
        src23 <= 16'h927e;
        src24 <= 16'hfe51;
        src25 <= 16'hdcc1;
        src26 <= 16'h5728;
        src27 <= 16'h54da;
        src28 <= 16'hc42a;
        src29 <= 16'h579f;
        src30 <= 16'h3057;
        src31 <= 16'ha306;
        src32 <= 16'h57f3;
        src33 <= 16'h912a;
        src34 <= 16'hb4e1;
        src35 <= 16'heb;
        src36 <= 16'h6dab;
        src37 <= 16'h5667;
        src38 <= 16'h78df;
        src39 <= 16'hc4c0;
        src40 <= 16'h2612;
        src41 <= 16'h6cdb;
        src42 <= 16'hc397;
        src43 <= 16'h7de6;
        src44 <= 16'h76ec;
        src45 <= 16'h8ead;
        src46 <= 16'ha388;
        src47 <= 16'h472a;
        src48 <= 16'h64d5;
        src49 <= 16'h7e3f;
        src50 <= 16'hff24;
        src51 <= 16'h940;
        src52 <= 16'hfe;
        src53 <= 16'h4f9e;
        src54 <= 16'hb80b;
        src55 <= 16'h4a1;
        src56 <= 16'hb745;
        src57 <= 16'h7f0d;
        src58 <= 16'h82e7;
        src59 <= 16'hdf23;
        src60 <= 16'h34b8;
        src61 <= 16'h5424;
        src62 <= 16'h6779;
        src63 <= 16'h4bed;
        src64 <= 16'hdb42;
        src65 <= 16'h25d6;
        src66 <= 16'hd938;
        src67 <= 16'h5a83;
        src68 <= 16'hbd9b;
        src69 <= 16'hd06;
        src70 <= 16'h2dc5;
        src71 <= 16'h2fab;
        src72 <= 16'h6a29;
        src73 <= 16'hd5c7;
        src74 <= 16'hb009;
        src75 <= 16'h49df;
        src76 <= 16'h96a7;
        src77 <= 16'he204;
        src78 <= 16'hdd92;
        src79 <= 16'hc8cf;
        src80 <= 16'hbbf3;
        src81 <= 16'hceec;
        src82 <= 16'h2d3f;
        src83 <= 16'h3403;
        src84 <= 16'hcd42;
        src85 <= 16'he09e;
        src86 <= 16'h84d9;
        src87 <= 16'h6fd9;
        src88 <= 16'hfb20;
        src89 <= 16'h84cf;
        src90 <= 16'hce23;
        src91 <= 16'hd9c6;
        src92 <= 16'h61df;
        src93 <= 16'h6bd8;
        src94 <= 16'h909;
        src95 <= 16'h2912;
        src96 <= 16'hebb3;
        src97 <= 16'h3a7b;
        src98 <= 16'hb7cd;
        src99 <= 16'h1dc5;
        src100 <= 16'h1288;
        src101 <= 16'hd097;
        src102 <= 16'h7578;
        src103 <= 16'h71dc;
        src104 <= 16'hcc1;
        src105 <= 16'hce90;
        src106 <= 16'h1520;
        src107 <= 16'ha24f;
        src108 <= 16'h80cc;
        src109 <= 16'h7cad;
        src110 <= 16'h640b;
        src111 <= 16'h5239;
        src112 <= 16'hf161;
        src113 <= 16'h725;
        src114 <= 16'hb74b;
        src115 <= 16'h3f58;
        src116 <= 16'hf82c;
        src117 <= 16'hc320;
        src118 <= 16'ha079;
        src119 <= 16'h228c;
        src120 <= 16'haa17;
        src121 <= 16'h17be;
        src122 <= 16'hb410;
        src123 <= 16'h4682;
        src124 <= 16'h4909;
        src125 <= 16'hf106;
        src126 <= 16'hf53a;
        src127 <= 16'h670e;
        exp <= 23'h4040fd;
        #1
        src0 <= 16'h1d5f;
        src1 <= 16'h57c8;
        src2 <= 16'h68ab;
        src3 <= 16'h1e77;
        src4 <= 16'h2ac9;
        src5 <= 16'hcacf;
        src6 <= 16'hb37b;
        src7 <= 16'h140f;
        src8 <= 16'h35c3;
        src9 <= 16'h83b0;
        src10 <= 16'h49ed;
        src11 <= 16'he9c7;
        src12 <= 16'he541;
        src13 <= 16'hb610;
        src14 <= 16'h92f8;
        src15 <= 16'h652a;
        src16 <= 16'hb8f8;
        src17 <= 16'h126d;
        src18 <= 16'hb620;
        src19 <= 16'h874e;
        src20 <= 16'h2ed7;
        src21 <= 16'h9f24;
        src22 <= 16'ha0ab;
        src23 <= 16'h1596;
        src24 <= 16'hdb49;
        src25 <= 16'h31ca;
        src26 <= 16'he9d7;
        src27 <= 16'hac94;
        src28 <= 16'he4b6;
        src29 <= 16'ha26c;
        src30 <= 16'hc11f;
        src31 <= 16'hb71c;
        src32 <= 16'h1546;
        src33 <= 16'h39c2;
        src34 <= 16'h3e3f;
        src35 <= 16'hcad4;
        src36 <= 16'hb5b1;
        src37 <= 16'hb29a;
        src38 <= 16'h7690;
        src39 <= 16'haa1a;
        src40 <= 16'h6b4;
        src41 <= 16'h6d1c;
        src42 <= 16'h37f5;
        src43 <= 16'hced8;
        src44 <= 16'h8258;
        src45 <= 16'h4418;
        src46 <= 16'h5f05;
        src47 <= 16'hce47;
        src48 <= 16'h2a68;
        src49 <= 16'h341f;
        src50 <= 16'h39b5;
        src51 <= 16'h8b40;
        src52 <= 16'h760e;
        src53 <= 16'h2eef;
        src54 <= 16'h2545;
        src55 <= 16'hbaf2;
        src56 <= 16'hc362;
        src57 <= 16'hce0b;
        src58 <= 16'hf6b8;
        src59 <= 16'h455c;
        src60 <= 16'h63ce;
        src61 <= 16'hb827;
        src62 <= 16'h6ba9;
        src63 <= 16'ha75e;
        src64 <= 16'h8a7f;
        src65 <= 16'hbc95;
        src66 <= 16'h4df8;
        src67 <= 16'hf8d7;
        src68 <= 16'h4594;
        src69 <= 16'hb0a8;
        src70 <= 16'h6617;
        src71 <= 16'h383a;
        src72 <= 16'h97bb;
        src73 <= 16'hc605;
        src74 <= 16'hf199;
        src75 <= 16'h291a;
        src76 <= 16'hd6fd;
        src77 <= 16'hf367;
        src78 <= 16'h807e;
        src79 <= 16'h19aa;
        src80 <= 16'h8283;
        src81 <= 16'h739b;
        src82 <= 16'hafa3;
        src83 <= 16'hc7c;
        src84 <= 16'hce37;
        src85 <= 16'hff3;
        src86 <= 16'hc04;
        src87 <= 16'h499b;
        src88 <= 16'hdc2a;
        src89 <= 16'h744e;
        src90 <= 16'h80b6;
        src91 <= 16'hffb2;
        src92 <= 16'hb356;
        src93 <= 16'h23af;
        src94 <= 16'h2f47;
        src95 <= 16'hcd90;
        src96 <= 16'h335c;
        src97 <= 16'h7704;
        src98 <= 16'hf4a9;
        src99 <= 16'h22af;
        src100 <= 16'hc57b;
        src101 <= 16'h4819;
        src102 <= 16'h40d;
        src103 <= 16'h5976;
        src104 <= 16'he128;
        src105 <= 16'hefaa;
        src106 <= 16'hcf8;
        src107 <= 16'h55f;
        src108 <= 16'ha5de;
        src109 <= 16'h3636;
        src110 <= 16'hd710;
        src111 <= 16'h2bca;
        src112 <= 16'hb1b3;
        src113 <= 16'h6296;
        src114 <= 16'h260e;
        src115 <= 16'hbd06;
        src116 <= 16'hcbb1;
        src117 <= 16'h3d64;
        src118 <= 16'h34cb;
        src119 <= 16'h3048;
        src120 <= 16'h8086;
        src121 <= 16'hb270;
        src122 <= 16'h7bd8;
        src123 <= 16'h3b85;
        src124 <= 16'he310;
        src125 <= 16'h3d07;
        src126 <= 16'ha3b1;
        src127 <= 16'hc04c;
        exp <= 23'h3eab88;
        #1
        src0 <= 16'h91db;
        src1 <= 16'h73d1;
        src2 <= 16'hdfa2;
        src3 <= 16'h48eb;
        src4 <= 16'hf6e9;
        src5 <= 16'h122f;
        src6 <= 16'hab51;
        src7 <= 16'hca31;
        src8 <= 16'hfa0b;
        src9 <= 16'h8db5;
        src10 <= 16'h357f;
        src11 <= 16'h6f29;
        src12 <= 16'ha31a;
        src13 <= 16'h4b20;
        src14 <= 16'h38f3;
        src15 <= 16'hbcbf;
        src16 <= 16'h4835;
        src17 <= 16'h4355;
        src18 <= 16'h4656;
        src19 <= 16'hb79d;
        src20 <= 16'h2d9c;
        src21 <= 16'h3c71;
        src22 <= 16'hcb1e;
        src23 <= 16'h6b6b;
        src24 <= 16'he61;
        src25 <= 16'hf93d;
        src26 <= 16'h82d6;
        src27 <= 16'h792d;
        src28 <= 16'hd11c;
        src29 <= 16'hc581;
        src30 <= 16'hbd7d;
        src31 <= 16'heda9;
        src32 <= 16'h24fb;
        src33 <= 16'hbb77;
        src34 <= 16'h7dc6;
        src35 <= 16'h182c;
        src36 <= 16'h1198;
        src37 <= 16'h67e0;
        src38 <= 16'hf818;
        src39 <= 16'h670d;
        src40 <= 16'h45f1;
        src41 <= 16'h3cb3;
        src42 <= 16'hf403;
        src43 <= 16'h4655;
        src44 <= 16'hd4ae;
        src45 <= 16'h2980;
        src46 <= 16'h41f8;
        src47 <= 16'hb0ff;
        src48 <= 16'h8cbb;
        src49 <= 16'hae6c;
        src50 <= 16'hd375;
        src51 <= 16'hbe87;
        src52 <= 16'h8941;
        src53 <= 16'h4a1c;
        src54 <= 16'h4a7d;
        src55 <= 16'h3b7c;
        src56 <= 16'h373f;
        src57 <= 16'h7e35;
        src58 <= 16'h30c4;
        src59 <= 16'h16b7;
        src60 <= 16'h315a;
        src61 <= 16'h3cbe;
        src62 <= 16'h3c67;
        src63 <= 16'h43a8;
        src64 <= 16'h59bb;
        src65 <= 16'hae31;
        src66 <= 16'h9dde;
        src67 <= 16'hcb8d;
        src68 <= 16'h1ae9;
        src69 <= 16'h5f8d;
        src70 <= 16'h6d59;
        src71 <= 16'hab06;
        src72 <= 16'he3ed;
        src73 <= 16'h25fa;
        src74 <= 16'hccfc;
        src75 <= 16'h48a9;
        src76 <= 16'h6f7e;
        src77 <= 16'hbb45;
        src78 <= 16'hb57f;
        src79 <= 16'h1eab;
        src80 <= 16'h34d1;
        src81 <= 16'h366f;
        src82 <= 16'hf271;
        src83 <= 16'h9ca6;
        src84 <= 16'hcdcb;
        src85 <= 16'h73d4;
        src86 <= 16'h2dda;
        src87 <= 16'hf503;
        src88 <= 16'h91d5;
        src89 <= 16'h14a9;
        src90 <= 16'ha1af;
        src91 <= 16'h8f06;
        src92 <= 16'h7535;
        src93 <= 16'h9e22;
        src94 <= 16'hd33e;
        src95 <= 16'h7a47;
        src96 <= 16'h7863;
        src97 <= 16'hae40;
        src98 <= 16'h112b;
        src99 <= 16'h9645;
        src100 <= 16'h30b4;
        src101 <= 16'h5c6f;
        src102 <= 16'hf2af;
        src103 <= 16'h5942;
        src104 <= 16'he2cd;
        src105 <= 16'h5dff;
        src106 <= 16'h8ac1;
        src107 <= 16'hccb6;
        src108 <= 16'hc902;
        src109 <= 16'hf4a;
        src110 <= 16'h8be3;
        src111 <= 16'h61d3;
        src112 <= 16'h353;
        src113 <= 16'hebb4;
        src114 <= 16'h8cf9;
        src115 <= 16'h4d7a;
        src116 <= 16'hbc8d;
        src117 <= 16'hb712;
        src118 <= 16'h5733;
        src119 <= 16'h5c52;
        src120 <= 16'h749;
        src121 <= 16'h5e05;
        src122 <= 16'hac48;
        src123 <= 16'ha952;
        src124 <= 16'hb62b;
        src125 <= 16'h9abd;
        src126 <= 16'h3323;
        src127 <= 16'h5cd4;
        exp <= 23'h3e86a7;
        #1
        src0 <= 16'h954c;
        src1 <= 16'hc689;
        src2 <= 16'h91fc;
        src3 <= 16'h4464;
        src4 <= 16'hd8bd;
        src5 <= 16'he7fd;
        src6 <= 16'h5cea;
        src7 <= 16'h3888;
        src8 <= 16'ha6ff;
        src9 <= 16'hb79a;
        src10 <= 16'h1b1d;
        src11 <= 16'hab2e;
        src12 <= 16'hcd6b;
        src13 <= 16'he440;
        src14 <= 16'hd05c;
        src15 <= 16'hcab8;
        src16 <= 16'hc305;
        src17 <= 16'hbf70;
        src18 <= 16'hd43;
        src19 <= 16'h7e63;
        src20 <= 16'h50d0;
        src21 <= 16'h957;
        src22 <= 16'h3cea;
        src23 <= 16'h4bbd;
        src24 <= 16'h8d74;
        src25 <= 16'h6964;
        src26 <= 16'hccad;
        src27 <= 16'h7e3f;
        src28 <= 16'h731c;
        src29 <= 16'h7139;
        src30 <= 16'h96f7;
        src31 <= 16'h5676;
        src32 <= 16'h52d4;
        src33 <= 16'hf928;
        src34 <= 16'h4d30;
        src35 <= 16'hfbd8;
        src36 <= 16'h61c1;
        src37 <= 16'h4f16;
        src38 <= 16'h93c7;
        src39 <= 16'h3be8;
        src40 <= 16'hefd;
        src41 <= 16'h979b;
        src42 <= 16'hcaaa;
        src43 <= 16'he6b;
        src44 <= 16'h3dda;
        src45 <= 16'h7b5d;
        src46 <= 16'h8668;
        src47 <= 16'he992;
        src48 <= 16'h6cf9;
        src49 <= 16'hb45e;
        src50 <= 16'hd600;
        src51 <= 16'h539;
        src52 <= 16'hd3f2;
        src53 <= 16'ha1d5;
        src54 <= 16'h636e;
        src55 <= 16'hf9da;
        src56 <= 16'hc072;
        src57 <= 16'h80b1;
        src58 <= 16'h9161;
        src59 <= 16'h5308;
        src60 <= 16'h32b8;
        src61 <= 16'h7038;
        src62 <= 16'hb3df;
        src63 <= 16'h9808;
        src64 <= 16'h4504;
        src65 <= 16'hd491;
        src66 <= 16'hb361;
        src67 <= 16'hc06f;
        src68 <= 16'hc4a9;
        src69 <= 16'h5dc8;
        src70 <= 16'h11ac;
        src71 <= 16'h4886;
        src72 <= 16'hef8a;
        src73 <= 16'ha925;
        src74 <= 16'h4db4;
        src75 <= 16'h6111;
        src76 <= 16'h8692;
        src77 <= 16'hfaa7;
        src78 <= 16'h5502;
        src79 <= 16'h2541;
        src80 <= 16'hf914;
        src81 <= 16'hab1e;
        src82 <= 16'h6fe7;
        src83 <= 16'h7d95;
        src84 <= 16'h9327;
        src85 <= 16'h679;
        src86 <= 16'h97ab;
        src87 <= 16'h3c27;
        src88 <= 16'hd5b0;
        src89 <= 16'h211f;
        src90 <= 16'hfed7;
        src91 <= 16'hdb13;
        src92 <= 16'hc1bb;
        src93 <= 16'h85d8;
        src94 <= 16'ha36b;
        src95 <= 16'h5321;
        src96 <= 16'h3525;
        src97 <= 16'h894d;
        src98 <= 16'h5b2f;
        src99 <= 16'h17ee;
        src100 <= 16'h3be0;
        src101 <= 16'hca15;
        src102 <= 16'h3d92;
        src103 <= 16'hfc8a;
        src104 <= 16'h6bf6;
        src105 <= 16'he39;
        src106 <= 16'h24e;
        src107 <= 16'h7f8b;
        src108 <= 16'h7789;
        src109 <= 16'h1f29;
        src110 <= 16'heb7;
        src111 <= 16'h5f1f;
        src112 <= 16'ha9cd;
        src113 <= 16'hdf5b;
        src114 <= 16'he2af;
        src115 <= 16'h9406;
        src116 <= 16'hd315;
        src117 <= 16'hc71;
        src118 <= 16'h9c75;
        src119 <= 16'h87fc;
        src120 <= 16'h30de;
        src121 <= 16'hc20c;
        src122 <= 16'h2b45;
        src123 <= 16'h8372;
        src124 <= 16'h3294;
        src125 <= 16'h7092;
        src126 <= 16'h7551;
        src127 <= 16'h701;
        exp <= 23'h4032ea;
        #1
        src0 <= 16'h6d24;
        src1 <= 16'hd3fa;
        src2 <= 16'h6aa1;
        src3 <= 16'h7794;
        src4 <= 16'ha360;
        src5 <= 16'h1316;
        src6 <= 16'h28c3;
        src7 <= 16'ha304;
        src8 <= 16'h5b72;
        src9 <= 16'h1acd;
        src10 <= 16'ha44;
        src11 <= 16'h586e;
        src12 <= 16'h558e;
        src13 <= 16'h52b0;
        src14 <= 16'hdcb5;
        src15 <= 16'hc20d;
        src16 <= 16'h30ff;
        src17 <= 16'h2250;
        src18 <= 16'hd42d;
        src19 <= 16'hb8b6;
        src20 <= 16'ha45d;
        src21 <= 16'h931a;
        src22 <= 16'h7ac1;
        src23 <= 16'h5d18;
        src24 <= 16'hb1bc;
        src25 <= 16'h3f95;
        src26 <= 16'hd735;
        src27 <= 16'h3311;
        src28 <= 16'haa6f;
        src29 <= 16'h95aa;
        src30 <= 16'hb874;
        src31 <= 16'hcc56;
        src32 <= 16'h7ce2;
        src33 <= 16'h39cb;
        src34 <= 16'hff0c;
        src35 <= 16'h82fc;
        src36 <= 16'h32f8;
        src37 <= 16'h8212;
        src38 <= 16'h2bf7;
        src39 <= 16'h6377;
        src40 <= 16'h1986;
        src41 <= 16'h715c;
        src42 <= 16'hcd7;
        src43 <= 16'ha75c;
        src44 <= 16'hb772;
        src45 <= 16'hb0ee;
        src46 <= 16'h7912;
        src47 <= 16'h4729;
        src48 <= 16'haa79;
        src49 <= 16'h85ca;
        src50 <= 16'h96b4;
        src51 <= 16'h6441;
        src52 <= 16'h185d;
        src53 <= 16'h6451;
        src54 <= 16'h54f0;
        src55 <= 16'hbc71;
        src56 <= 16'hd376;
        src57 <= 16'h2464;
        src58 <= 16'h51df;
        src59 <= 16'hfe70;
        src60 <= 16'h37f6;
        src61 <= 16'h93a3;
        src62 <= 16'hade2;
        src63 <= 16'hcc39;
        src64 <= 16'h4393;
        src65 <= 16'h911;
        src66 <= 16'h43f1;
        src67 <= 16'hb706;
        src68 <= 16'h4cc0;
        src69 <= 16'h99dd;
        src70 <= 16'haa68;
        src71 <= 16'h8a6c;
        src72 <= 16'h23c;
        src73 <= 16'h8e40;
        src74 <= 16'h416b;
        src75 <= 16'hbecb;
        src76 <= 16'h2553;
        src77 <= 16'h2d01;
        src78 <= 16'h3ea3;
        src79 <= 16'hc660;
        src80 <= 16'hcc08;
        src81 <= 16'h3777;
        src82 <= 16'h8dbb;
        src83 <= 16'hf6de;
        src84 <= 16'hcd58;
        src85 <= 16'ha258;
        src86 <= 16'hefe9;
        src87 <= 16'h6e2c;
        src88 <= 16'h9b68;
        src89 <= 16'h96d;
        src90 <= 16'h13ac;
        src91 <= 16'h2f15;
        src92 <= 16'h9129;
        src93 <= 16'h4486;
        src94 <= 16'h868d;
        src95 <= 16'hff51;
        src96 <= 16'h522c;
        src97 <= 16'haef4;
        src98 <= 16'h2fde;
        src99 <= 16'hbd6f;
        src100 <= 16'hedc5;
        src101 <= 16'h2761;
        src102 <= 16'h6c92;
        src103 <= 16'hc541;
        src104 <= 16'hda71;
        src105 <= 16'ha47e;
        src106 <= 16'h8f57;
        src107 <= 16'h3704;
        src108 <= 16'h1c88;
        src109 <= 16'h214b;
        src110 <= 16'h80f3;
        src111 <= 16'hc276;
        src112 <= 16'he77b;
        src113 <= 16'h90d0;
        src114 <= 16'hb9d7;
        src115 <= 16'ha24c;
        src116 <= 16'h251a;
        src117 <= 16'h4c43;
        src118 <= 16'hba0f;
        src119 <= 16'hac8d;
        src120 <= 16'h95fd;
        src121 <= 16'hc08e;
        src122 <= 16'h5a3f;
        src123 <= 16'ha611;
        src124 <= 16'h3abf;
        src125 <= 16'h4f12;
        src126 <= 16'hdb01;
        src127 <= 16'hde94;
        exp <= 23'h3ec827;
        #1
        src0 <= 16'hd932;
        src1 <= 16'hd87;
        src2 <= 16'hf8ad;
        src3 <= 16'h9a28;
        src4 <= 16'h6a7e;
        src5 <= 16'h13a6;
        src6 <= 16'h1e2e;
        src7 <= 16'h86ad;
        src8 <= 16'h821b;
        src9 <= 16'hb09;
        src10 <= 16'h7cc;
        src11 <= 16'h6161;
        src12 <= 16'ha569;
        src13 <= 16'h1b4c;
        src14 <= 16'hd7cf;
        src15 <= 16'hf93b;
        src16 <= 16'ha73f;
        src17 <= 16'h41d5;
        src18 <= 16'hb31f;
        src19 <= 16'hd299;
        src20 <= 16'hd5da;
        src21 <= 16'h79db;
        src22 <= 16'h4668;
        src23 <= 16'h4896;
        src24 <= 16'h275e;
        src25 <= 16'hb7b5;
        src26 <= 16'h4a26;
        src27 <= 16'hc13d;
        src28 <= 16'h4607;
        src29 <= 16'hacd6;
        src30 <= 16'h208f;
        src31 <= 16'hec06;
        src32 <= 16'hbf8b;
        src33 <= 16'h2497;
        src34 <= 16'h72e8;
        src35 <= 16'ha4e1;
        src36 <= 16'hdb5d;
        src37 <= 16'h87ab;
        src38 <= 16'hc19f;
        src39 <= 16'hf499;
        src40 <= 16'h1e1e;
        src41 <= 16'hd383;
        src42 <= 16'h5168;
        src43 <= 16'h91f;
        src44 <= 16'hc495;
        src45 <= 16'hc004;
        src46 <= 16'hdaa2;
        src47 <= 16'h9fff;
        src48 <= 16'h6f7c;
        src49 <= 16'h2a36;
        src50 <= 16'hb71f;
        src51 <= 16'hc83f;
        src52 <= 16'h868a;
        src53 <= 16'h39f9;
        src54 <= 16'h68e7;
        src55 <= 16'h9d5d;
        src56 <= 16'h44ad;
        src57 <= 16'h7777;
        src58 <= 16'hfdd0;
        src59 <= 16'h2532;
        src60 <= 16'h4cce;
        src61 <= 16'h76ed;
        src62 <= 16'hc22c;
        src63 <= 16'h6d47;
        src64 <= 16'h4bb0;
        src65 <= 16'hdabf;
        src66 <= 16'hfe83;
        src67 <= 16'h2d85;
        src68 <= 16'h7404;
        src69 <= 16'h88d3;
        src70 <= 16'heacf;
        src71 <= 16'h143e;
        src72 <= 16'hb513;
        src73 <= 16'hce7f;
        src74 <= 16'h359b;
        src75 <= 16'he75b;
        src76 <= 16'he68c;
        src77 <= 16'h8cc;
        src78 <= 16'h8e01;
        src79 <= 16'h700a;
        src80 <= 16'hdd0a;
        src81 <= 16'hc52b;
        src82 <= 16'haa06;
        src83 <= 16'h7190;
        src84 <= 16'h463f;
        src85 <= 16'h1adf;
        src86 <= 16'h2f81;
        src87 <= 16'he895;
        src88 <= 16'hd66b;
        src89 <= 16'hdf64;
        src90 <= 16'he16c;
        src91 <= 16'hda7;
        src92 <= 16'haf7;
        src93 <= 16'hf1b8;
        src94 <= 16'h7fa;
        src95 <= 16'hf1d5;
        src96 <= 16'h71c4;
        src97 <= 16'h9ce8;
        src98 <= 16'h636c;
        src99 <= 16'h749a;
        src100 <= 16'h1a37;
        src101 <= 16'hdb4e;
        src102 <= 16'h7ba3;
        src103 <= 16'h5540;
        src104 <= 16'he049;
        src105 <= 16'h94c8;
        src106 <= 16'h480e;
        src107 <= 16'h427e;
        src108 <= 16'h171c;
        src109 <= 16'h1fa9;
        src110 <= 16'h36ce;
        src111 <= 16'h5a96;
        src112 <= 16'heeca;
        src113 <= 16'h265b;
        src114 <= 16'hf05a;
        src115 <= 16'h9af7;
        src116 <= 16'hdb98;
        src117 <= 16'hbd8;
        src118 <= 16'h1b30;
        src119 <= 16'h97f6;
        src120 <= 16'h2ef0;
        src121 <= 16'h5f1c;
        src122 <= 16'h544b;
        src123 <= 16'hba7b;
        src124 <= 16'hdabd;
        src125 <= 16'hfd87;
        src126 <= 16'hfd23;
        src127 <= 16'h66fd;
        exp <= 23'h41a683;
        #1
        src0 <= 16'h406f;
        src1 <= 16'h183;
        src2 <= 16'h69af;
        src3 <= 16'hdc3a;
        src4 <= 16'h56eb;
        src5 <= 16'h1745;
        src6 <= 16'hdeed;
        src7 <= 16'h43a;
        src8 <= 16'hbad8;
        src9 <= 16'h2595;
        src10 <= 16'hbbd5;
        src11 <= 16'h2713;
        src12 <= 16'ha197;
        src13 <= 16'h24af;
        src14 <= 16'h3101;
        src15 <= 16'hd4d3;
        src16 <= 16'h7e78;
        src17 <= 16'hf3b9;
        src18 <= 16'hfe8e;
        src19 <= 16'he380;
        src20 <= 16'hd323;
        src21 <= 16'h3665;
        src22 <= 16'hb9a8;
        src23 <= 16'hf08;
        src24 <= 16'h77dd;
        src25 <= 16'h3a92;
        src26 <= 16'h5354;
        src27 <= 16'ha87b;
        src28 <= 16'h6446;
        src29 <= 16'h754e;
        src30 <= 16'h7d24;
        src31 <= 16'hfd98;
        src32 <= 16'h1abb;
        src33 <= 16'h31da;
        src34 <= 16'h7ed8;
        src35 <= 16'hca67;
        src36 <= 16'h3e5e;
        src37 <= 16'h4260;
        src38 <= 16'hf531;
        src39 <= 16'habf9;
        src40 <= 16'hd0e0;
        src41 <= 16'h7d73;
        src42 <= 16'h1710;
        src43 <= 16'h38e8;
        src44 <= 16'h3f3e;
        src45 <= 16'h1e2;
        src46 <= 16'h56c5;
        src47 <= 16'h9ade;
        src48 <= 16'h16c4;
        src49 <= 16'hd7a8;
        src50 <= 16'h3f5b;
        src51 <= 16'h5234;
        src52 <= 16'hd9e0;
        src53 <= 16'he6da;
        src54 <= 16'ha1af;
        src55 <= 16'h776e;
        src56 <= 16'h72b0;
        src57 <= 16'h9618;
        src58 <= 16'h8fbc;
        src59 <= 16'hecb1;
        src60 <= 16'h83b8;
        src61 <= 16'hca54;
        src62 <= 16'h9a24;
        src63 <= 16'h3c58;
        src64 <= 16'hef6d;
        src65 <= 16'h64a7;
        src66 <= 16'h65a2;
        src67 <= 16'h166;
        src68 <= 16'h791a;
        src69 <= 16'h2e3a;
        src70 <= 16'h87c1;
        src71 <= 16'hc831;
        src72 <= 16'hfd38;
        src73 <= 16'h3c8;
        src74 <= 16'h239;
        src75 <= 16'h9036;
        src76 <= 16'ha726;
        src77 <= 16'hde44;
        src78 <= 16'h707c;
        src79 <= 16'h9c60;
        src80 <= 16'hdf2e;
        src81 <= 16'he354;
        src82 <= 16'hdeca;
        src83 <= 16'h6ebb;
        src84 <= 16'hd894;
        src85 <= 16'h466;
        src86 <= 16'hdfc2;
        src87 <= 16'ha3c3;
        src88 <= 16'h5bf9;
        src89 <= 16'h7381;
        src90 <= 16'he08a;
        src91 <= 16'h34fb;
        src92 <= 16'h465e;
        src93 <= 16'hdabb;
        src94 <= 16'h88c3;
        src95 <= 16'h80d8;
        src96 <= 16'h5fdd;
        src97 <= 16'h582b;
        src98 <= 16'h46fe;
        src99 <= 16'ha44;
        src100 <= 16'h65c5;
        src101 <= 16'he549;
        src102 <= 16'h7d68;
        src103 <= 16'h1284;
        src104 <= 16'h1fdb;
        src105 <= 16'h7970;
        src106 <= 16'h1472;
        src107 <= 16'h38ac;
        src108 <= 16'hc4c5;
        src109 <= 16'h2c0a;
        src110 <= 16'hf9e2;
        src111 <= 16'h37;
        src112 <= 16'h8c65;
        src113 <= 16'he8a3;
        src114 <= 16'hcffa;
        src115 <= 16'h76e5;
        src116 <= 16'he7c0;
        src117 <= 16'hbe4b;
        src118 <= 16'hac77;
        src119 <= 16'h86e2;
        src120 <= 16'hd8c5;
        src121 <= 16'hc9be;
        src122 <= 16'hb81e;
        src123 <= 16'h8095;
        src124 <= 16'h870c;
        src125 <= 16'h33f4;
        src126 <= 16'hd52e;
        src127 <= 16'h19c3;
        exp <= 23'h404656;
        #1
        src0 <= 16'h8eb3;
        src1 <= 16'had97;
        src2 <= 16'h13b3;
        src3 <= 16'hb5d7;
        src4 <= 16'h286d;
        src5 <= 16'hc3ea;
        src6 <= 16'hd1ab;
        src7 <= 16'he89f;
        src8 <= 16'h1dba;
        src9 <= 16'hd6c6;
        src10 <= 16'hdee9;
        src11 <= 16'h59b4;
        src12 <= 16'hd215;
        src13 <= 16'h3ec1;
        src14 <= 16'hb0a4;
        src15 <= 16'h88aa;
        src16 <= 16'h85bd;
        src17 <= 16'he2de;
        src18 <= 16'hc50b;
        src19 <= 16'ha0c4;
        src20 <= 16'h3435;
        src21 <= 16'h207e;
        src22 <= 16'h3e11;
        src23 <= 16'heb67;
        src24 <= 16'hbf74;
        src25 <= 16'h6df8;
        src26 <= 16'hd979;
        src27 <= 16'hda19;
        src28 <= 16'h2808;
        src29 <= 16'h66ca;
        src30 <= 16'h75b9;
        src31 <= 16'h623e;
        src32 <= 16'h648e;
        src33 <= 16'hbd48;
        src34 <= 16'ha821;
        src35 <= 16'h42e4;
        src36 <= 16'he709;
        src37 <= 16'he873;
        src38 <= 16'h4ed3;
        src39 <= 16'h94dc;
        src40 <= 16'hd506;
        src41 <= 16'hd932;
        src42 <= 16'hc2f2;
        src43 <= 16'h3792;
        src44 <= 16'he29d;
        src45 <= 16'h4f9c;
        src46 <= 16'hf013;
        src47 <= 16'h7755;
        src48 <= 16'h827d;
        src49 <= 16'h50e6;
        src50 <= 16'h2231;
        src51 <= 16'h9f1a;
        src52 <= 16'h58bb;
        src53 <= 16'hc0e7;
        src54 <= 16'h34bd;
        src55 <= 16'h5fce;
        src56 <= 16'h258e;
        src57 <= 16'hdde5;
        src58 <= 16'h812d;
        src59 <= 16'h9cee;
        src60 <= 16'h30c1;
        src61 <= 16'he86;
        src62 <= 16'ha92d;
        src63 <= 16'haa8f;
        src64 <= 16'h454b;
        src65 <= 16'h3343;
        src66 <= 16'h3b0c;
        src67 <= 16'h7efb;
        src68 <= 16'h9958;
        src69 <= 16'h34dc;
        src70 <= 16'h88ee;
        src71 <= 16'h6ad6;
        src72 <= 16'hf50c;
        src73 <= 16'h14d5;
        src74 <= 16'h87e6;
        src75 <= 16'haed8;
        src76 <= 16'h8192;
        src77 <= 16'h3cd3;
        src78 <= 16'h4e7;
        src79 <= 16'h4f02;
        src80 <= 16'h8972;
        src81 <= 16'h69be;
        src82 <= 16'h7001;
        src83 <= 16'h858a;
        src84 <= 16'hc78e;
        src85 <= 16'h6683;
        src86 <= 16'heb18;
        src87 <= 16'he5;
        src88 <= 16'hf37d;
        src89 <= 16'h4fd3;
        src90 <= 16'hea0a;
        src91 <= 16'h2c6;
        src92 <= 16'h1efd;
        src93 <= 16'h50be;
        src94 <= 16'h3ab6;
        src95 <= 16'h3442;
        src96 <= 16'h2e25;
        src97 <= 16'h46fe;
        src98 <= 16'h6fb;
        src99 <= 16'h772b;
        src100 <= 16'h4ce5;
        src101 <= 16'hf80c;
        src102 <= 16'hded;
        src103 <= 16'h3265;
        src104 <= 16'h4d1e;
        src105 <= 16'hca5d;
        src106 <= 16'h877b;
        src107 <= 16'h5dd1;
        src108 <= 16'h3cf3;
        src109 <= 16'he95f;
        src110 <= 16'h19c1;
        src111 <= 16'hb8a7;
        src112 <= 16'h17c;
        src113 <= 16'hdc80;
        src114 <= 16'h1b45;
        src115 <= 16'h6a2f;
        src116 <= 16'h9c89;
        src117 <= 16'hc310;
        src118 <= 16'hc235;
        src119 <= 16'ha6b8;
        src120 <= 16'hea16;
        src121 <= 16'h5d48;
        src122 <= 16'hd432;
        src123 <= 16'hec21;
        src124 <= 16'heed5;
        src125 <= 16'hc1c2;
        src126 <= 16'hbee5;
        src127 <= 16'hb6f0;
        exp <= 23'h40d317;
        #1
        src0 <= 16'hca4b;
        src1 <= 16'h7dad;
        src2 <= 16'h748d;
        src3 <= 16'ha19;
        src4 <= 16'h9faa;
        src5 <= 16'h3102;
        src6 <= 16'h5fd5;
        src7 <= 16'ha3e5;
        src8 <= 16'hd54c;
        src9 <= 16'h73a7;
        src10 <= 16'h6ed9;
        src11 <= 16'h2fe2;
        src12 <= 16'hb4cc;
        src13 <= 16'hf7d2;
        src14 <= 16'h54ba;
        src15 <= 16'haace;
        src16 <= 16'hea61;
        src17 <= 16'hb1a9;
        src18 <= 16'ha267;
        src19 <= 16'hbe08;
        src20 <= 16'h81a5;
        src21 <= 16'hc8eb;
        src22 <= 16'h76da;
        src23 <= 16'h7b8a;
        src24 <= 16'h9283;
        src25 <= 16'h1f37;
        src26 <= 16'hcff4;
        src27 <= 16'h9bf1;
        src28 <= 16'hc618;
        src29 <= 16'h7d6c;
        src30 <= 16'hdba;
        src31 <= 16'h10d0;
        src32 <= 16'h4d2c;
        src33 <= 16'ha5e2;
        src34 <= 16'ha5b1;
        src35 <= 16'hdb2c;
        src36 <= 16'h23ab;
        src37 <= 16'h5897;
        src38 <= 16'hf65a;
        src39 <= 16'h806f;
        src40 <= 16'h474b;
        src41 <= 16'h212c;
        src42 <= 16'ha787;
        src43 <= 16'h4e06;
        src44 <= 16'h6e56;
        src45 <= 16'h4bd4;
        src46 <= 16'hfcde;
        src47 <= 16'h5e76;
        src48 <= 16'hf959;
        src49 <= 16'hec1c;
        src50 <= 16'h4a29;
        src51 <= 16'hb9;
        src52 <= 16'hd68b;
        src53 <= 16'h9ab1;
        src54 <= 16'hb678;
        src55 <= 16'hf6c2;
        src56 <= 16'habbd;
        src57 <= 16'h8fe8;
        src58 <= 16'h36a8;
        src59 <= 16'hff2c;
        src60 <= 16'ha3b;
        src61 <= 16'h1c96;
        src62 <= 16'hcc48;
        src63 <= 16'he463;
        src64 <= 16'h2d03;
        src65 <= 16'hc62;
        src66 <= 16'h7989;
        src67 <= 16'hd105;
        src68 <= 16'h6b02;
        src69 <= 16'hfa02;
        src70 <= 16'h7548;
        src71 <= 16'hf881;
        src72 <= 16'haf21;
        src73 <= 16'h943a;
        src74 <= 16'h151a;
        src75 <= 16'hfe20;
        src76 <= 16'h7685;
        src77 <= 16'h4be1;
        src78 <= 16'h4987;
        src79 <= 16'h3ec8;
        src80 <= 16'h8191;
        src81 <= 16'h1a7a;
        src82 <= 16'he05a;
        src83 <= 16'hf564;
        src84 <= 16'h7f20;
        src85 <= 16'h57da;
        src86 <= 16'h5860;
        src87 <= 16'h1549;
        src88 <= 16'h856;
        src89 <= 16'h51c8;
        src90 <= 16'h983e;
        src91 <= 16'h6165;
        src92 <= 16'h46e;
        src93 <= 16'h9d52;
        src94 <= 16'h67bd;
        src95 <= 16'h43df;
        src96 <= 16'h41aa;
        src97 <= 16'h7ab1;
        src98 <= 16'h1eb6;
        src99 <= 16'hc9c;
        src100 <= 16'h29fc;
        src101 <= 16'h7be2;
        src102 <= 16'h4719;
        src103 <= 16'ha1e2;
        src104 <= 16'h9cbf;
        src105 <= 16'h7fe4;
        src106 <= 16'h5c25;
        src107 <= 16'h6551;
        src108 <= 16'h782a;
        src109 <= 16'hfd65;
        src110 <= 16'h7138;
        src111 <= 16'hdfae;
        src112 <= 16'h7ef3;
        src113 <= 16'hea79;
        src114 <= 16'h64fa;
        src115 <= 16'h16bb;
        src116 <= 16'h2d62;
        src117 <= 16'h2c3d;
        src118 <= 16'h2e7b;
        src119 <= 16'hfc42;
        src120 <= 16'h5992;
        src121 <= 16'h4cd6;
        src122 <= 16'hda94;
        src123 <= 16'h3af;
        src124 <= 16'h2ded;
        src125 <= 16'h9794;
        src126 <= 16'hc645;
        src127 <= 16'haf68;
        exp <= 23'h3eee29;
        #1
        src0 <= 16'h79b7;
        src1 <= 16'h50a8;
        src2 <= 16'h27f5;
        src3 <= 16'hb84d;
        src4 <= 16'hc627;
        src5 <= 16'hf83;
        src6 <= 16'h781;
        src7 <= 16'h2fb1;
        src8 <= 16'h7732;
        src9 <= 16'h3f21;
        src10 <= 16'h21a3;
        src11 <= 16'h18b6;
        src12 <= 16'hcb9;
        src13 <= 16'h43e5;
        src14 <= 16'h397c;
        src15 <= 16'h455a;
        src16 <= 16'h9f31;
        src17 <= 16'hf1a;
        src18 <= 16'hd686;
        src19 <= 16'h458;
        src20 <= 16'h7702;
        src21 <= 16'hdc02;
        src22 <= 16'hb4dc;
        src23 <= 16'h5e44;
        src24 <= 16'h1935;
        src25 <= 16'h8e51;
        src26 <= 16'h3b4c;
        src27 <= 16'h6216;
        src28 <= 16'h54be;
        src29 <= 16'hee6a;
        src30 <= 16'h4234;
        src31 <= 16'h3f5b;
        src32 <= 16'h5750;
        src33 <= 16'hb00f;
        src34 <= 16'h2d9f;
        src35 <= 16'haa7;
        src36 <= 16'h9273;
        src37 <= 16'hfac2;
        src38 <= 16'ha308;
        src39 <= 16'h25a2;
        src40 <= 16'h5bbb;
        src41 <= 16'h5f5d;
        src42 <= 16'h6bdd;
        src43 <= 16'h93ad;
        src44 <= 16'hff63;
        src45 <= 16'he711;
        src46 <= 16'h94e5;
        src47 <= 16'h7e15;
        src48 <= 16'h1dac;
        src49 <= 16'hf7c4;
        src50 <= 16'h1db6;
        src51 <= 16'h2da4;
        src52 <= 16'h56f3;
        src53 <= 16'h988;
        src54 <= 16'h8d98;
        src55 <= 16'h80bb;
        src56 <= 16'ha4dc;
        src57 <= 16'ha0eb;
        src58 <= 16'h5839;
        src59 <= 16'h952e;
        src60 <= 16'h89a7;
        src61 <= 16'hd969;
        src62 <= 16'h27a8;
        src63 <= 16'hdfaf;
        src64 <= 16'hb532;
        src65 <= 16'h832d;
        src66 <= 16'h6261;
        src67 <= 16'hd295;
        src68 <= 16'he684;
        src69 <= 16'h587e;
        src70 <= 16'h244b;
        src71 <= 16'he810;
        src72 <= 16'h3123;
        src73 <= 16'h1a85;
        src74 <= 16'h450f;
        src75 <= 16'h7cec;
        src76 <= 16'hea38;
        src77 <= 16'h4f23;
        src78 <= 16'hcab7;
        src79 <= 16'h2845;
        src80 <= 16'h431;
        src81 <= 16'hc8a9;
        src82 <= 16'h1f8a;
        src83 <= 16'he5d2;
        src84 <= 16'h4771;
        src85 <= 16'hd986;
        src86 <= 16'hfc5;
        src87 <= 16'h9a9c;
        src88 <= 16'h1392;
        src89 <= 16'h987;
        src90 <= 16'hf026;
        src91 <= 16'h4143;
        src92 <= 16'h756c;
        src93 <= 16'h73cd;
        src94 <= 16'hcb5c;
        src95 <= 16'hbc8b;
        src96 <= 16'h97fc;
        src97 <= 16'h231d;
        src98 <= 16'h52be;
        src99 <= 16'h8ed3;
        src100 <= 16'hc165;
        src101 <= 16'h32f1;
        src102 <= 16'h5492;
        src103 <= 16'h5e0e;
        src104 <= 16'haf7f;
        src105 <= 16'h7bda;
        src106 <= 16'hb8b3;
        src107 <= 16'h337;
        src108 <= 16'hff15;
        src109 <= 16'h697b;
        src110 <= 16'h33cf;
        src111 <= 16'hb025;
        src112 <= 16'h2f6c;
        src113 <= 16'h62e5;
        src114 <= 16'he6cb;
        src115 <= 16'h7e0f;
        src116 <= 16'h1f5a;
        src117 <= 16'h88bb;
        src118 <= 16'h38a5;
        src119 <= 16'hdd06;
        src120 <= 16'hdd2d;
        src121 <= 16'h90e6;
        src122 <= 16'h5180;
        src123 <= 16'h1a42;
        src124 <= 16'hc7b4;
        src125 <= 16'h8237;
        src126 <= 16'hae20;
        src127 <= 16'h21ea;
        exp <= 23'h399742;
        #1
        src0 <= 16'h5886;
        src1 <= 16'hc57;
        src2 <= 16'h7a3;
        src3 <= 16'h29d5;
        src4 <= 16'h93a7;
        src5 <= 16'hbf55;
        src6 <= 16'hf83b;
        src7 <= 16'hdbb4;
        src8 <= 16'heda0;
        src9 <= 16'h54ce;
        src10 <= 16'hf17f;
        src11 <= 16'hd0b3;
        src12 <= 16'h5181;
        src13 <= 16'h9529;
        src14 <= 16'h48c8;
        src15 <= 16'h81a6;
        src16 <= 16'h6944;
        src17 <= 16'he93e;
        src18 <= 16'h3bff;
        src19 <= 16'h208d;
        src20 <= 16'h6ee6;
        src21 <= 16'h235a;
        src22 <= 16'h7deb;
        src23 <= 16'hfc08;
        src24 <= 16'h72d8;
        src25 <= 16'h9127;
        src26 <= 16'h3832;
        src27 <= 16'h758c;
        src28 <= 16'hf853;
        src29 <= 16'hb41d;
        src30 <= 16'h4e95;
        src31 <= 16'hf2b4;
        src32 <= 16'hcc90;
        src33 <= 16'hd532;
        src34 <= 16'hc2a1;
        src35 <= 16'hc48;
        src36 <= 16'hc971;
        src37 <= 16'h5b11;
        src38 <= 16'hea91;
        src39 <= 16'h8db5;
        src40 <= 16'h6209;
        src41 <= 16'h64e6;
        src42 <= 16'h4b0b;
        src43 <= 16'h4d18;
        src44 <= 16'h2440;
        src45 <= 16'hb1d7;
        src46 <= 16'h4666;
        src47 <= 16'h6cfa;
        src48 <= 16'h9145;
        src49 <= 16'ha2ea;
        src50 <= 16'h2037;
        src51 <= 16'h6237;
        src52 <= 16'hb703;
        src53 <= 16'hbae9;
        src54 <= 16'he06c;
        src55 <= 16'hee1b;
        src56 <= 16'ha5e7;
        src57 <= 16'h415b;
        src58 <= 16'h5d0c;
        src59 <= 16'h2708;
        src60 <= 16'hfa87;
        src61 <= 16'h3f01;
        src62 <= 16'ha17c;
        src63 <= 16'h4984;
        src64 <= 16'hd0fb;
        src65 <= 16'hd063;
        src66 <= 16'hb4f6;
        src67 <= 16'h10ad;
        src68 <= 16'hc1e1;
        src69 <= 16'hf721;
        src70 <= 16'hf083;
        src71 <= 16'h3dfe;
        src72 <= 16'hdc02;
        src73 <= 16'h9626;
        src74 <= 16'h9892;
        src75 <= 16'hcf25;
        src76 <= 16'h5833;
        src77 <= 16'hc2df;
        src78 <= 16'h77d7;
        src79 <= 16'hb91;
        src80 <= 16'h6a71;
        src81 <= 16'h63a7;
        src82 <= 16'hd112;
        src83 <= 16'hf15;
        src84 <= 16'h287d;
        src85 <= 16'hc897;
        src86 <= 16'habf0;
        src87 <= 16'hd011;
        src88 <= 16'hb99f;
        src89 <= 16'h44af;
        src90 <= 16'hc0fd;
        src91 <= 16'h3208;
        src92 <= 16'heb40;
        src93 <= 16'hfd1d;
        src94 <= 16'h7fa1;
        src95 <= 16'h377;
        src96 <= 16'he764;
        src97 <= 16'hdb9e;
        src98 <= 16'h2cc5;
        src99 <= 16'h7bdf;
        src100 <= 16'hb977;
        src101 <= 16'h6bea;
        src102 <= 16'h4cc7;
        src103 <= 16'hb588;
        src104 <= 16'h8126;
        src105 <= 16'hc2f3;
        src106 <= 16'had69;
        src107 <= 16'h9235;
        src108 <= 16'h3276;
        src109 <= 16'h53f2;
        src110 <= 16'h1bfe;
        src111 <= 16'hafc;
        src112 <= 16'h80b5;
        src113 <= 16'h2710;
        src114 <= 16'hf6ba;
        src115 <= 16'h77da;
        src116 <= 16'h7f5c;
        src117 <= 16'hbaa;
        src118 <= 16'h6dc2;
        src119 <= 16'h626;
        src120 <= 16'ha357;
        src121 <= 16'hc4fa;
        src122 <= 16'h9570;
        src123 <= 16'h8c0;
        src124 <= 16'ha252;
        src125 <= 16'h1b70;
        src126 <= 16'h310e;
        src127 <= 16'hc26e;
        exp <= 23'h421b07;
        #1
        src0 <= 16'h51af;
        src1 <= 16'h847a;
        src2 <= 16'hafe3;
        src3 <= 16'h9dd7;
        src4 <= 16'h3669;
        src5 <= 16'hd56c;
        src6 <= 16'h7571;
        src7 <= 16'h6989;
        src8 <= 16'h42a9;
        src9 <= 16'h3176;
        src10 <= 16'h3d26;
        src11 <= 16'haca4;
        src12 <= 16'hac90;
        src13 <= 16'h6161;
        src14 <= 16'h2cbd;
        src15 <= 16'h72f2;
        src16 <= 16'hf1dc;
        src17 <= 16'h5740;
        src18 <= 16'h67ab;
        src19 <= 16'hab1a;
        src20 <= 16'h68bb;
        src21 <= 16'ha51f;
        src22 <= 16'hd69;
        src23 <= 16'h8214;
        src24 <= 16'h9bff;
        src25 <= 16'hed17;
        src26 <= 16'hce0e;
        src27 <= 16'h4cd3;
        src28 <= 16'h255;
        src29 <= 16'h86a2;
        src30 <= 16'hd2e7;
        src31 <= 16'he92e;
        src32 <= 16'hfda5;
        src33 <= 16'h5c80;
        src34 <= 16'hbe32;
        src35 <= 16'h5f8d;
        src36 <= 16'hec18;
        src37 <= 16'hbcbf;
        src38 <= 16'h9c3c;
        src39 <= 16'h6615;
        src40 <= 16'h5cf0;
        src41 <= 16'h764e;
        src42 <= 16'h9a82;
        src43 <= 16'h40ed;
        src44 <= 16'h2c95;
        src45 <= 16'h4e71;
        src46 <= 16'h43a1;
        src47 <= 16'h4d58;
        src48 <= 16'hda6d;
        src49 <= 16'hb523;
        src50 <= 16'hd670;
        src51 <= 16'h4317;
        src52 <= 16'hc0ac;
        src53 <= 16'h398f;
        src54 <= 16'hafab;
        src55 <= 16'hba06;
        src56 <= 16'he24b;
        src57 <= 16'h6c6a;
        src58 <= 16'hbf72;
        src59 <= 16'heb05;
        src60 <= 16'hb526;
        src61 <= 16'h41b1;
        src62 <= 16'he425;
        src63 <= 16'he825;
        src64 <= 16'h810b;
        src65 <= 16'ha2f0;
        src66 <= 16'h2c47;
        src67 <= 16'haa99;
        src68 <= 16'h69b;
        src69 <= 16'h6f19;
        src70 <= 16'hcb0f;
        src71 <= 16'h5b65;
        src72 <= 16'h9153;
        src73 <= 16'h8b34;
        src74 <= 16'h2dfa;
        src75 <= 16'h84c6;
        src76 <= 16'hfbb3;
        src77 <= 16'h4346;
        src78 <= 16'h1eb7;
        src79 <= 16'ha0a0;
        src80 <= 16'h372f;
        src81 <= 16'h293f;
        src82 <= 16'hd050;
        src83 <= 16'h91fa;
        src84 <= 16'h514e;
        src85 <= 16'h26b3;
        src86 <= 16'h39ec;
        src87 <= 16'hea17;
        src88 <= 16'h4d51;
        src89 <= 16'h4b87;
        src90 <= 16'h9dc7;
        src91 <= 16'h23a5;
        src92 <= 16'he46;
        src93 <= 16'h6167;
        src94 <= 16'hc68f;
        src95 <= 16'h2336;
        src96 <= 16'h32b6;
        src97 <= 16'hfa36;
        src98 <= 16'h50fe;
        src99 <= 16'hd6be;
        src100 <= 16'he49c;
        src101 <= 16'h2de7;
        src102 <= 16'h3d0d;
        src103 <= 16'ha41b;
        src104 <= 16'h848;
        src105 <= 16'h6348;
        src106 <= 16'h3b69;
        src107 <= 16'h5ce1;
        src108 <= 16'h5ae5;
        src109 <= 16'hf4c6;
        src110 <= 16'h77e;
        src111 <= 16'h84e5;
        src112 <= 16'h2b74;
        src113 <= 16'h7247;
        src114 <= 16'hdf0b;
        src115 <= 16'h160b;
        src116 <= 16'hbeb8;
        src117 <= 16'hfe22;
        src118 <= 16'h9bd0;
        src119 <= 16'h2bf;
        src120 <= 16'ha199;
        src121 <= 16'h2de0;
        src122 <= 16'h34ba;
        src123 <= 16'hf620;
        src124 <= 16'h5db7;
        src125 <= 16'h6f6c;
        src126 <= 16'h71df;
        src127 <= 16'h34f9;
        exp <= 23'h3e9f4d;
        #1
        src0 <= 16'h1c7;
        src1 <= 16'h17f5;
        src2 <= 16'ha019;
        src3 <= 16'hc270;
        src4 <= 16'h3fde;
        src5 <= 16'h3cd0;
        src6 <= 16'h5db;
        src7 <= 16'h9607;
        src8 <= 16'h30cc;
        src9 <= 16'h722;
        src10 <= 16'hf159;
        src11 <= 16'h626e;
        src12 <= 16'hef1a;
        src13 <= 16'h6517;
        src14 <= 16'h51a4;
        src15 <= 16'h46da;
        src16 <= 16'h573d;
        src17 <= 16'haa3e;
        src18 <= 16'h161c;
        src19 <= 16'h273e;
        src20 <= 16'h936d;
        src21 <= 16'hc410;
        src22 <= 16'h7869;
        src23 <= 16'h3360;
        src24 <= 16'h2b9d;
        src25 <= 16'h8f2d;
        src26 <= 16'h938f;
        src27 <= 16'hbce5;
        src28 <= 16'h46b5;
        src29 <= 16'h2b21;
        src30 <= 16'hf24c;
        src31 <= 16'h31c5;
        src32 <= 16'hd73d;
        src33 <= 16'h2e6e;
        src34 <= 16'h4e88;
        src35 <= 16'h229e;
        src36 <= 16'h54b5;
        src37 <= 16'h307e;
        src38 <= 16'h70af;
        src39 <= 16'h4042;
        src40 <= 16'h51a5;
        src41 <= 16'hc3ec;
        src42 <= 16'h543;
        src43 <= 16'h44d0;
        src44 <= 16'hc0a5;
        src45 <= 16'hf995;
        src46 <= 16'hff9c;
        src47 <= 16'hfda2;
        src48 <= 16'hcc63;
        src49 <= 16'h778c;
        src50 <= 16'h4dc8;
        src51 <= 16'hb2c7;
        src52 <= 16'he1ea;
        src53 <= 16'hd4bc;
        src54 <= 16'hc133;
        src55 <= 16'h764f;
        src56 <= 16'ha5b1;
        src57 <= 16'hf671;
        src58 <= 16'he8a1;
        src59 <= 16'h4061;
        src60 <= 16'h60f2;
        src61 <= 16'hda9a;
        src62 <= 16'h13ea;
        src63 <= 16'h4313;
        src64 <= 16'hdfcb;
        src65 <= 16'h7f01;
        src66 <= 16'h4f71;
        src67 <= 16'h364a;
        src68 <= 16'h3e6f;
        src69 <= 16'haac9;
        src70 <= 16'hc1f8;
        src71 <= 16'h8add;
        src72 <= 16'hefaa;
        src73 <= 16'h9668;
        src74 <= 16'h122e;
        src75 <= 16'hb196;
        src76 <= 16'h1639;
        src77 <= 16'h6271;
        src78 <= 16'h8cd3;
        src79 <= 16'h5d38;
        src80 <= 16'h5a17;
        src81 <= 16'hd40e;
        src82 <= 16'h3cac;
        src83 <= 16'h8fc0;
        src84 <= 16'h59a9;
        src85 <= 16'h4e97;
        src86 <= 16'hb444;
        src87 <= 16'h3aac;
        src88 <= 16'h6c54;
        src89 <= 16'hce56;
        src90 <= 16'h7fa9;
        src91 <= 16'h109c;
        src92 <= 16'hd84e;
        src93 <= 16'h5f10;
        src94 <= 16'hcbf;
        src95 <= 16'h9972;
        src96 <= 16'hddb6;
        src97 <= 16'h3ed0;
        src98 <= 16'h86d9;
        src99 <= 16'h9dad;
        src100 <= 16'h680e;
        src101 <= 16'h6ec4;
        src102 <= 16'h23f4;
        src103 <= 16'h32bb;
        src104 <= 16'he568;
        src105 <= 16'h198b;
        src106 <= 16'h8133;
        src107 <= 16'hc28c;
        src108 <= 16'h6cf9;
        src109 <= 16'hd5db;
        src110 <= 16'h62cd;
        src111 <= 16'hab87;
        src112 <= 16'h5e74;
        src113 <= 16'hbec6;
        src114 <= 16'h9b53;
        src115 <= 16'h147a;
        src116 <= 16'h1280;
        src117 <= 16'hede0;
        src118 <= 16'h25db;
        src119 <= 16'h3790;
        src120 <= 16'hf3e4;
        src121 <= 16'hf7ec;
        src122 <= 16'h37a0;
        src123 <= 16'h21a4;
        src124 <= 16'h309b;
        src125 <= 16'hc6e;
        src126 <= 16'he7a3;
        src127 <= 16'h2a0a;
        exp <= 23'h3c013e;
        #1
        src0 <= 16'h5582;
        src1 <= 16'h91c6;
        src2 <= 16'hae52;
        src3 <= 16'he2d1;
        src4 <= 16'h8803;
        src5 <= 16'he0c7;
        src6 <= 16'h8eb6;
        src7 <= 16'h70bf;
        src8 <= 16'h16d;
        src9 <= 16'ha115;
        src10 <= 16'hbf4d;
        src11 <= 16'h4b09;
        src12 <= 16'h393a;
        src13 <= 16'h3aa;
        src14 <= 16'hf73;
        src15 <= 16'h5ff8;
        src16 <= 16'h3bdf;
        src17 <= 16'hac7b;
        src18 <= 16'hd93c;
        src19 <= 16'h7944;
        src20 <= 16'hc3b4;
        src21 <= 16'h454c;
        src22 <= 16'hcc74;
        src23 <= 16'h5c4e;
        src24 <= 16'h3c8d;
        src25 <= 16'hf575;
        src26 <= 16'h63dd;
        src27 <= 16'h4ece;
        src28 <= 16'h5aa2;
        src29 <= 16'hd518;
        src30 <= 16'hed0;
        src31 <= 16'h38e4;
        src32 <= 16'hea19;
        src33 <= 16'hc2bc;
        src34 <= 16'haf53;
        src35 <= 16'hb69;
        src36 <= 16'he5d4;
        src37 <= 16'h814d;
        src38 <= 16'h3fc;
        src39 <= 16'ha497;
        src40 <= 16'hf5a2;
        src41 <= 16'h1035;
        src42 <= 16'h27a9;
        src43 <= 16'hb32b;
        src44 <= 16'hb862;
        src45 <= 16'h586;
        src46 <= 16'h561;
        src47 <= 16'h8189;
        src48 <= 16'h92f7;
        src49 <= 16'h12ca;
        src50 <= 16'h4f59;
        src51 <= 16'h2417;
        src52 <= 16'hafcb;
        src53 <= 16'h60cd;
        src54 <= 16'h216e;
        src55 <= 16'h58d3;
        src56 <= 16'hc52b;
        src57 <= 16'h8b4b;
        src58 <= 16'h5ddb;
        src59 <= 16'he8af;
        src60 <= 16'hb6d3;
        src61 <= 16'hc8fb;
        src62 <= 16'h9aee;
        src63 <= 16'hc433;
        src64 <= 16'hc9f0;
        src65 <= 16'hac0;
        src66 <= 16'ha105;
        src67 <= 16'h72b8;
        src68 <= 16'h1cd7;
        src69 <= 16'h1244;
        src70 <= 16'h5744;
        src71 <= 16'hd149;
        src72 <= 16'hfa8e;
        src73 <= 16'h38ba;
        src74 <= 16'h5748;
        src75 <= 16'ha81e;
        src76 <= 16'h13bf;
        src77 <= 16'hcd50;
        src78 <= 16'h8f38;
        src79 <= 16'haca3;
        src80 <= 16'h5824;
        src81 <= 16'hd627;
        src82 <= 16'h5cbd;
        src83 <= 16'h26e8;
        src84 <= 16'hcd7d;
        src85 <= 16'h1d80;
        src86 <= 16'hf8d4;
        src87 <= 16'he1c7;
        src88 <= 16'hf9cf;
        src89 <= 16'h2e7c;
        src90 <= 16'h3b93;
        src91 <= 16'hefd5;
        src92 <= 16'h523c;
        src93 <= 16'h1aca;
        src94 <= 16'he08a;
        src95 <= 16'h9b3;
        src96 <= 16'hb497;
        src97 <= 16'h275b;
        src98 <= 16'h514a;
        src99 <= 16'h1a1b;
        src100 <= 16'hdd4e;
        src101 <= 16'h49f9;
        src102 <= 16'hfc4e;
        src103 <= 16'hb74d;
        src104 <= 16'h1e12;
        src105 <= 16'h48d1;
        src106 <= 16'hc15;
        src107 <= 16'hc493;
        src108 <= 16'h7ff2;
        src109 <= 16'hb68a;
        src110 <= 16'h8283;
        src111 <= 16'h6dd7;
        src112 <= 16'hbd08;
        src113 <= 16'h73ab;
        src114 <= 16'hb48;
        src115 <= 16'he82a;
        src116 <= 16'ha269;
        src117 <= 16'hfa00;
        src118 <= 16'hbf7c;
        src119 <= 16'h6700;
        src120 <= 16'hb2de;
        src121 <= 16'h7225;
        src122 <= 16'h6e0e;
        src123 <= 16'h5c0e;
        src124 <= 16'h32d3;
        src125 <= 16'hf0fc;
        src126 <= 16'h3259;
        src127 <= 16'hf688;
        exp <= 23'h3f0ee1;
        #1
        src0 <= 16'he314;
        src1 <= 16'hf7f0;
        src2 <= 16'hc64e;
        src3 <= 16'hf202;
        src4 <= 16'hceba;
        src5 <= 16'hc522;
        src6 <= 16'hfd13;
        src7 <= 16'hfee3;
        src8 <= 16'h11d4;
        src9 <= 16'h9d7a;
        src10 <= 16'h1a8b;
        src11 <= 16'hde82;
        src12 <= 16'h97f4;
        src13 <= 16'hb440;
        src14 <= 16'h6bcc;
        src15 <= 16'hf292;
        src16 <= 16'hd33c;
        src17 <= 16'h25c0;
        src18 <= 16'h667;
        src19 <= 16'hf5d2;
        src20 <= 16'hf45b;
        src21 <= 16'hc123;
        src22 <= 16'h6654;
        src23 <= 16'hf85d;
        src24 <= 16'h49c6;
        src25 <= 16'h10b7;
        src26 <= 16'h97c6;
        src27 <= 16'h5599;
        src28 <= 16'h53b2;
        src29 <= 16'h26a;
        src30 <= 16'h8e5c;
        src31 <= 16'h534c;
        src32 <= 16'hb0b0;
        src33 <= 16'hbc06;
        src34 <= 16'h9dbd;
        src35 <= 16'hc0c1;
        src36 <= 16'h7073;
        src37 <= 16'ha22d;
        src38 <= 16'hfdd4;
        src39 <= 16'ha40e;
        src40 <= 16'hbe18;
        src41 <= 16'hca01;
        src42 <= 16'h4769;
        src43 <= 16'he94a;
        src44 <= 16'hd848;
        src45 <= 16'h5c76;
        src46 <= 16'h252;
        src47 <= 16'hdfb2;
        src48 <= 16'h6053;
        src49 <= 16'h815a;
        src50 <= 16'h1c2e;
        src51 <= 16'h6b40;
        src52 <= 16'h8e29;
        src53 <= 16'h6d4e;
        src54 <= 16'h9961;
        src55 <= 16'hfd80;
        src56 <= 16'h4742;
        src57 <= 16'h58f5;
        src58 <= 16'hd3a5;
        src59 <= 16'hc06b;
        src60 <= 16'he0e7;
        src61 <= 16'h8592;
        src62 <= 16'hf44c;
        src63 <= 16'hc29e;
        src64 <= 16'h4f10;
        src65 <= 16'haf8c;
        src66 <= 16'ha0b4;
        src67 <= 16'hede4;
        src68 <= 16'he685;
        src69 <= 16'h7c10;
        src70 <= 16'h194d;
        src71 <= 16'h184a;
        src72 <= 16'h7e1b;
        src73 <= 16'hdaec;
        src74 <= 16'hdb4;
        src75 <= 16'h9bd;
        src76 <= 16'h8bc7;
        src77 <= 16'hc129;
        src78 <= 16'h994d;
        src79 <= 16'h9a57;
        src80 <= 16'hd616;
        src81 <= 16'h8c1b;
        src82 <= 16'h7e8c;
        src83 <= 16'haeb1;
        src84 <= 16'h7c87;
        src85 <= 16'h9982;
        src86 <= 16'h41dc;
        src87 <= 16'haf89;
        src88 <= 16'hbb;
        src89 <= 16'ha084;
        src90 <= 16'h9552;
        src91 <= 16'h3df6;
        src92 <= 16'hedee;
        src93 <= 16'hfb77;
        src94 <= 16'hb33c;
        src95 <= 16'h94a4;
        src96 <= 16'h5c19;
        src97 <= 16'h449d;
        src98 <= 16'ha76;
        src99 <= 16'hb6b4;
        src100 <= 16'hd6ca;
        src101 <= 16'h66b4;
        src102 <= 16'h792f;
        src103 <= 16'hd5f9;
        src104 <= 16'h9bad;
        src105 <= 16'he42c;
        src106 <= 16'h8d4e;
        src107 <= 16'h3581;
        src108 <= 16'h44b0;
        src109 <= 16'h6dbd;
        src110 <= 16'h231a;
        src111 <= 16'hff4;
        src112 <= 16'h8036;
        src113 <= 16'h78d2;
        src114 <= 16'h2164;
        src115 <= 16'h6458;
        src116 <= 16'h5e1;
        src117 <= 16'h5d8c;
        src118 <= 16'h56e2;
        src119 <= 16'hdcb7;
        src120 <= 16'hb876;
        src121 <= 16'had84;
        src122 <= 16'h88aa;
        src123 <= 16'h57e1;
        src124 <= 16'h82c6;
        src125 <= 16'h8cc5;
        src126 <= 16'h38b4;
        src127 <= 16'hdf4f;
        exp <= 23'h468512;
        #1
        src0 <= 16'h605d;
        src1 <= 16'ha76c;
        src2 <= 16'h9887;
        src3 <= 16'hbcc6;
        src4 <= 16'h85e;
        src5 <= 16'hd7ea;
        src6 <= 16'hcb26;
        src7 <= 16'h8f53;
        src8 <= 16'hb18a;
        src9 <= 16'h2ac1;
        src10 <= 16'hfdfa;
        src11 <= 16'h7c2e;
        src12 <= 16'haf05;
        src13 <= 16'hfa1d;
        src14 <= 16'h66bb;
        src15 <= 16'h8b07;
        src16 <= 16'hbe1a;
        src17 <= 16'h23ea;
        src18 <= 16'h1c97;
        src19 <= 16'h8f9e;
        src20 <= 16'h9f6;
        src21 <= 16'h6e46;
        src22 <= 16'hebb9;
        src23 <= 16'hcd96;
        src24 <= 16'h4184;
        src25 <= 16'hac57;
        src26 <= 16'h112d;
        src27 <= 16'h3e03;
        src28 <= 16'hc381;
        src29 <= 16'hb65d;
        src30 <= 16'h2d22;
        src31 <= 16'heab5;
        src32 <= 16'h7474;
        src33 <= 16'h8a26;
        src34 <= 16'h5e1f;
        src35 <= 16'h47e6;
        src36 <= 16'h48c8;
        src37 <= 16'h84c0;
        src38 <= 16'hff71;
        src39 <= 16'h3e08;
        src40 <= 16'h5e47;
        src41 <= 16'h6c32;
        src42 <= 16'hace9;
        src43 <= 16'h4745;
        src44 <= 16'h649d;
        src45 <= 16'h5eee;
        src46 <= 16'h91fe;
        src47 <= 16'hfdff;
        src48 <= 16'hb5c0;
        src49 <= 16'h26d8;
        src50 <= 16'h766;
        src51 <= 16'h6abd;
        src52 <= 16'h3615;
        src53 <= 16'h56dc;
        src54 <= 16'h2640;
        src55 <= 16'hcb3c;
        src56 <= 16'h8bfc;
        src57 <= 16'h3f65;
        src58 <= 16'hdba3;
        src59 <= 16'he3b0;
        src60 <= 16'h8756;
        src61 <= 16'h4a25;
        src62 <= 16'ha5dc;
        src63 <= 16'hb8c2;
        src64 <= 16'h35c8;
        src65 <= 16'h2742;
        src66 <= 16'h1ff6;
        src67 <= 16'h996f;
        src68 <= 16'h2214;
        src69 <= 16'h1396;
        src70 <= 16'hb846;
        src71 <= 16'h80e3;
        src72 <= 16'hd3c1;
        src73 <= 16'h24e;
        src74 <= 16'h110;
        src75 <= 16'hce55;
        src76 <= 16'h6b19;
        src77 <= 16'h470c;
        src78 <= 16'h3726;
        src79 <= 16'h4e67;
        src80 <= 16'h884c;
        src81 <= 16'h19f9;
        src82 <= 16'hba4d;
        src83 <= 16'hbe68;
        src84 <= 16'hcec0;
        src85 <= 16'hb759;
        src86 <= 16'h5b99;
        src87 <= 16'hfdb6;
        src88 <= 16'he636;
        src89 <= 16'he658;
        src90 <= 16'hd673;
        src91 <= 16'h7b5f;
        src92 <= 16'h1759;
        src93 <= 16'h1a5c;
        src94 <= 16'hcb6b;
        src95 <= 16'h2e4c;
        src96 <= 16'h5fd5;
        src97 <= 16'h2a10;
        src98 <= 16'h3a02;
        src99 <= 16'h2461;
        src100 <= 16'h1575;
        src101 <= 16'hbda8;
        src102 <= 16'h4a69;
        src103 <= 16'h3f51;
        src104 <= 16'h3d99;
        src105 <= 16'h7daa;
        src106 <= 16'h3016;
        src107 <= 16'h3b9c;
        src108 <= 16'h60eb;
        src109 <= 16'hfee9;
        src110 <= 16'h1016;
        src111 <= 16'h917b;
        src112 <= 16'h9209;
        src113 <= 16'hfff4;
        src114 <= 16'hac50;
        src115 <= 16'h5dcc;
        src116 <= 16'hfbf5;
        src117 <= 16'hb866;
        src118 <= 16'ha8db;
        src119 <= 16'h4d0;
        src120 <= 16'h505b;
        src121 <= 16'h711d;
        src122 <= 16'hf623;
        src123 <= 16'h4b85;
        src124 <= 16'hb7d8;
        src125 <= 16'hd485;
        src126 <= 16'he8ee;
        src127 <= 16'hd126;
        exp <= 23'h3ebd35;
        #1
        src0 <= 16'haefc;
        src1 <= 16'had3e;
        src2 <= 16'hcd36;
        src3 <= 16'h212f;
        src4 <= 16'h6606;
        src5 <= 16'h81d2;
        src6 <= 16'h292e;
        src7 <= 16'h5a5d;
        src8 <= 16'h19b6;
        src9 <= 16'h8c97;
        src10 <= 16'h9bc6;
        src11 <= 16'hca06;
        src12 <= 16'h28eb;
        src13 <= 16'h6bf2;
        src14 <= 16'hf2f3;
        src15 <= 16'he6de;
        src16 <= 16'h920b;
        src17 <= 16'h1ec5;
        src18 <= 16'h2d6;
        src19 <= 16'h853d;
        src20 <= 16'h828c;
        src21 <= 16'hff66;
        src22 <= 16'h1eb1;
        src23 <= 16'h9ab1;
        src24 <= 16'h89c;
        src25 <= 16'ha011;
        src26 <= 16'h6300;
        src27 <= 16'h1e37;
        src28 <= 16'h79a6;
        src29 <= 16'h4b0c;
        src30 <= 16'h58b6;
        src31 <= 16'hd781;
        src32 <= 16'h915d;
        src33 <= 16'hf62b;
        src34 <= 16'h5282;
        src35 <= 16'h214e;
        src36 <= 16'he112;
        src37 <= 16'h6d3d;
        src38 <= 16'hdce1;
        src39 <= 16'he803;
        src40 <= 16'h43f2;
        src41 <= 16'h111b;
        src42 <= 16'h5f52;
        src43 <= 16'hf03b;
        src44 <= 16'hccdd;
        src45 <= 16'h7075;
        src46 <= 16'hd916;
        src47 <= 16'hbab3;
        src48 <= 16'hbaa2;
        src49 <= 16'hb212;
        src50 <= 16'h26ce;
        src51 <= 16'h996d;
        src52 <= 16'hee8e;
        src53 <= 16'h8791;
        src54 <= 16'h1904;
        src55 <= 16'h7e94;
        src56 <= 16'hd8c2;
        src57 <= 16'h4142;
        src58 <= 16'hf200;
        src59 <= 16'h8466;
        src60 <= 16'hec39;
        src61 <= 16'hd68e;
        src62 <= 16'h315f;
        src63 <= 16'h1e83;
        src64 <= 16'h6be8;
        src65 <= 16'hfdec;
        src66 <= 16'hae42;
        src67 <= 16'h7beb;
        src68 <= 16'hc287;
        src69 <= 16'h9a80;
        src70 <= 16'hf14a;
        src71 <= 16'h813b;
        src72 <= 16'h628e;
        src73 <= 16'he169;
        src74 <= 16'h568c;
        src75 <= 16'h3d98;
        src76 <= 16'h7606;
        src77 <= 16'hc139;
        src78 <= 16'hb49c;
        src79 <= 16'h2842;
        src80 <= 16'hd7a6;
        src81 <= 16'h17ec;
        src82 <= 16'h612;
        src83 <= 16'heccb;
        src84 <= 16'hfca6;
        src85 <= 16'h82fc;
        src86 <= 16'h8d48;
        src87 <= 16'he741;
        src88 <= 16'hba3;
        src89 <= 16'hd950;
        src90 <= 16'h51b9;
        src91 <= 16'h9bab;
        src92 <= 16'h35d;
        src93 <= 16'he78f;
        src94 <= 16'h5f3c;
        src95 <= 16'hb614;
        src96 <= 16'hfe0c;
        src97 <= 16'h4cb2;
        src98 <= 16'h3eb3;
        src99 <= 16'hfeb0;
        src100 <= 16'h9dbd;
        src101 <= 16'h6191;
        src102 <= 16'h8403;
        src103 <= 16'h4cde;
        src104 <= 16'h8756;
        src105 <= 16'h4672;
        src106 <= 16'hfd0a;
        src107 <= 16'he8ef;
        src108 <= 16'hfd8e;
        src109 <= 16'h701a;
        src110 <= 16'h7890;
        src111 <= 16'h8290;
        src112 <= 16'h4998;
        src113 <= 16'ha139;
        src114 <= 16'hec55;
        src115 <= 16'hfd46;
        src116 <= 16'h27a;
        src117 <= 16'hff99;
        src118 <= 16'hc31f;
        src119 <= 16'hef94;
        src120 <= 16'he672;
        src121 <= 16'hdb95;
        src122 <= 16'h224a;
        src123 <= 16'h19d4;
        src124 <= 16'h8a16;
        src125 <= 16'hf61d;
        src126 <= 16'hfd3f;
        src127 <= 16'h843a;
        exp <= 23'h471c94;
        #1
        src0 <= 16'h471;
        src1 <= 16'h833b;
        src2 <= 16'hf698;
        src3 <= 16'h57c4;
        src4 <= 16'ha7ad;
        src5 <= 16'h42e4;
        src6 <= 16'h4aae;
        src7 <= 16'h944f;
        src8 <= 16'hd136;
        src9 <= 16'heac0;
        src10 <= 16'he360;
        src11 <= 16'h4203;
        src12 <= 16'hb578;
        src13 <= 16'h794e;
        src14 <= 16'hbfcd;
        src15 <= 16'hfd2e;
        src16 <= 16'h1225;
        src17 <= 16'h91a2;
        src18 <= 16'hf77c;
        src19 <= 16'h552b;
        src20 <= 16'h5070;
        src21 <= 16'he87a;
        src22 <= 16'h9d1d;
        src23 <= 16'h8480;
        src24 <= 16'ha4ad;
        src25 <= 16'h70ce;
        src26 <= 16'h8dc7;
        src27 <= 16'h7d3d;
        src28 <= 16'h4e02;
        src29 <= 16'haba8;
        src30 <= 16'he325;
        src31 <= 16'he89c;
        src32 <= 16'hcbb6;
        src33 <= 16'h4af2;
        src34 <= 16'h57dd;
        src35 <= 16'hbd7a;
        src36 <= 16'h3a6f;
        src37 <= 16'h7352;
        src38 <= 16'hde0f;
        src39 <= 16'hd795;
        src40 <= 16'hf64f;
        src41 <= 16'hfbe1;
        src42 <= 16'h5478;
        src43 <= 16'h81f6;
        src44 <= 16'h46e;
        src45 <= 16'h41e2;
        src46 <= 16'h4688;
        src47 <= 16'h1abb;
        src48 <= 16'h7941;
        src49 <= 16'h3505;
        src50 <= 16'h86c6;
        src51 <= 16'h9708;
        src52 <= 16'h5e3b;
        src53 <= 16'h1887;
        src54 <= 16'h5f50;
        src55 <= 16'hfa27;
        src56 <= 16'h1348;
        src57 <= 16'h1b4f;
        src58 <= 16'haa12;
        src59 <= 16'h5ae9;
        src60 <= 16'h7f5e;
        src61 <= 16'hf8a;
        src62 <= 16'h5744;
        src63 <= 16'h8ecd;
        src64 <= 16'h3eef;
        src65 <= 16'h79fb;
        src66 <= 16'h78f6;
        src67 <= 16'h838e;
        src68 <= 16'hd145;
        src69 <= 16'hecfc;
        src70 <= 16'h21da;
        src71 <= 16'h7f70;
        src72 <= 16'h3037;
        src73 <= 16'he99a;
        src74 <= 16'h4008;
        src75 <= 16'ha618;
        src76 <= 16'h2935;
        src77 <= 16'had3e;
        src78 <= 16'h84de;
        src79 <= 16'h25ee;
        src80 <= 16'hd770;
        src81 <= 16'h7cdc;
        src82 <= 16'h4a11;
        src83 <= 16'hfeb5;
        src84 <= 16'h9f66;
        src85 <= 16'hc73a;
        src86 <= 16'ha8ef;
        src87 <= 16'haf78;
        src88 <= 16'h50f6;
        src89 <= 16'h7913;
        src90 <= 16'hc7a3;
        src91 <= 16'hba34;
        src92 <= 16'ha8b7;
        src93 <= 16'h3da2;
        src94 <= 16'hc925;
        src95 <= 16'hed41;
        src96 <= 16'h70a1;
        src97 <= 16'h77fa;
        src98 <= 16'h2f87;
        src99 <= 16'h1dfb;
        src100 <= 16'h8b69;
        src101 <= 16'hb16b;
        src102 <= 16'h5526;
        src103 <= 16'h47f3;
        src104 <= 16'h68c2;
        src105 <= 16'h44a9;
        src106 <= 16'hc878;
        src107 <= 16'h5792;
        src108 <= 16'heb2c;
        src109 <= 16'h3c18;
        src110 <= 16'h752b;
        src111 <= 16'h3fb1;
        src112 <= 16'hec60;
        src113 <= 16'hf597;
        src114 <= 16'h3d90;
        src115 <= 16'hb1f5;
        src116 <= 16'h8bdf;
        src117 <= 16'h9089;
        src118 <= 16'h2f85;
        src119 <= 16'hf8cd;
        src120 <= 16'hf812;
        src121 <= 16'h4a89;
        src122 <= 16'h93bb;
        src123 <= 16'h2daa;
        src124 <= 16'hc9d2;
        src125 <= 16'h703c;
        src126 <= 16'h42ae;
        src127 <= 16'ha3cc;
        exp <= 23'h42b13a;
        #1
        src0 <= 16'ha593;
        src1 <= 16'hc998;
        src2 <= 16'hf82e;
        src3 <= 16'h209;
        src4 <= 16'hc607;
        src5 <= 16'h8009;
        src6 <= 16'ha4b7;
        src7 <= 16'h3889;
        src8 <= 16'h9bb0;
        src9 <= 16'hd832;
        src10 <= 16'h8d06;
        src11 <= 16'hf798;
        src12 <= 16'hbb81;
        src13 <= 16'hec77;
        src14 <= 16'hc2e0;
        src15 <= 16'hc9ac;
        src16 <= 16'h63bf;
        src17 <= 16'hf20;
        src18 <= 16'h3c58;
        src19 <= 16'hd497;
        src20 <= 16'hae3a;
        src21 <= 16'h4d82;
        src22 <= 16'hf913;
        src23 <= 16'h6add;
        src24 <= 16'hf5b6;
        src25 <= 16'hca97;
        src26 <= 16'hf73a;
        src27 <= 16'ha9ed;
        src28 <= 16'h30c3;
        src29 <= 16'h7afd;
        src30 <= 16'h9ccd;
        src31 <= 16'hea11;
        src32 <= 16'h1a22;
        src33 <= 16'hfb32;
        src34 <= 16'h2c9e;
        src35 <= 16'h19a8;
        src36 <= 16'he347;
        src37 <= 16'h2af5;
        src38 <= 16'hb6b2;
        src39 <= 16'h61b8;
        src40 <= 16'hc78c;
        src41 <= 16'ha1ce;
        src42 <= 16'h18f8;
        src43 <= 16'hb595;
        src44 <= 16'h388;
        src45 <= 16'hfe40;
        src46 <= 16'h47b6;
        src47 <= 16'h8a52;
        src48 <= 16'h5b82;
        src49 <= 16'he691;
        src50 <= 16'h8130;
        src51 <= 16'hff2c;
        src52 <= 16'h6761;
        src53 <= 16'h7166;
        src54 <= 16'hd864;
        src55 <= 16'hda9d;
        src56 <= 16'h6a4d;
        src57 <= 16'h2ac2;
        src58 <= 16'h5fef;
        src59 <= 16'h7bab;
        src60 <= 16'hd0c6;
        src61 <= 16'h6309;
        src62 <= 16'h8eb1;
        src63 <= 16'hb841;
        src64 <= 16'h6969;
        src65 <= 16'hca8;
        src66 <= 16'hc954;
        src67 <= 16'h6be3;
        src68 <= 16'hc373;
        src69 <= 16'h654f;
        src70 <= 16'h8af1;
        src71 <= 16'h4a50;
        src72 <= 16'h4c95;
        src73 <= 16'h48bd;
        src74 <= 16'h2bed;
        src75 <= 16'h6642;
        src76 <= 16'hb046;
        src77 <= 16'h6f42;
        src78 <= 16'he521;
        src79 <= 16'hbbf0;
        src80 <= 16'h36e1;
        src81 <= 16'hff09;
        src82 <= 16'h7c63;
        src83 <= 16'h7514;
        src84 <= 16'he435;
        src85 <= 16'h8d4a;
        src86 <= 16'h906b;
        src87 <= 16'h70a0;
        src88 <= 16'h9cd8;
        src89 <= 16'h811b;
        src90 <= 16'hc87f;
        src91 <= 16'h1e35;
        src92 <= 16'hc986;
        src93 <= 16'h1315;
        src94 <= 16'h4886;
        src95 <= 16'h7aa2;
        src96 <= 16'h45d2;
        src97 <= 16'h94c;
        src98 <= 16'h2976;
        src99 <= 16'ha28d;
        src100 <= 16'h57f0;
        src101 <= 16'h50b1;
        src102 <= 16'h1d4d;
        src103 <= 16'h3987;
        src104 <= 16'h1b4f;
        src105 <= 16'h6a8d;
        src106 <= 16'hb083;
        src107 <= 16'hd54c;
        src108 <= 16'h4b99;
        src109 <= 16'hb871;
        src110 <= 16'hf8be;
        src111 <= 16'h5f9e;
        src112 <= 16'ha730;
        src113 <= 16'h435f;
        src114 <= 16'h1be3;
        src115 <= 16'h9c3e;
        src116 <= 16'h6a9;
        src117 <= 16'h659f;
        src118 <= 16'h30c9;
        src119 <= 16'hd8c5;
        src120 <= 16'h37a3;
        src121 <= 16'h315f;
        src122 <= 16'h4c64;
        src123 <= 16'hf1ff;
        src124 <= 16'h8b3d;
        src125 <= 16'hed9c;
        src126 <= 16'h5d1f;
        src127 <= 16'h74cd;
        exp <= 23'h4255eb;
        #1
        src0 <= 16'h8149;
        src1 <= 16'he503;
        src2 <= 16'hbae1;
        src3 <= 16'ha275;
        src4 <= 16'he400;
        src5 <= 16'h66cd;
        src6 <= 16'h625c;
        src7 <= 16'hd8d2;
        src8 <= 16'hb912;
        src9 <= 16'he95c;
        src10 <= 16'h5976;
        src11 <= 16'hbbdd;
        src12 <= 16'hebe6;
        src13 <= 16'h19cd;
        src14 <= 16'hb483;
        src15 <= 16'h8376;
        src16 <= 16'h705d;
        src17 <= 16'heb1b;
        src18 <= 16'h9bc2;
        src19 <= 16'h9d6a;
        src20 <= 16'h229c;
        src21 <= 16'h299e;
        src22 <= 16'h7c64;
        src23 <= 16'h4711;
        src24 <= 16'h30c8;
        src25 <= 16'he025;
        src26 <= 16'h8dbc;
        src27 <= 16'h8303;
        src28 <= 16'hc258;
        src29 <= 16'h9ba6;
        src30 <= 16'h611e;
        src31 <= 16'h91d8;
        src32 <= 16'hf7eb;
        src33 <= 16'hce92;
        src34 <= 16'h91dd;
        src35 <= 16'h29c8;
        src36 <= 16'hf599;
        src37 <= 16'h62d2;
        src38 <= 16'h8c01;
        src39 <= 16'he3b7;
        src40 <= 16'hc343;
        src41 <= 16'h66ab;
        src42 <= 16'h2e15;
        src43 <= 16'h2bee;
        src44 <= 16'h17f0;
        src45 <= 16'haf55;
        src46 <= 16'h8a97;
        src47 <= 16'h4038;
        src48 <= 16'hc312;
        src49 <= 16'h1674;
        src50 <= 16'h104d;
        src51 <= 16'h9b1f;
        src52 <= 16'h46ea;
        src53 <= 16'h4ab3;
        src54 <= 16'h2caf;
        src55 <= 16'h10e1;
        src56 <= 16'hc660;
        src57 <= 16'ha26e;
        src58 <= 16'h10e9;
        src59 <= 16'he143;
        src60 <= 16'hb7f5;
        src61 <= 16'ha2c;
        src62 <= 16'h1d19;
        src63 <= 16'h249d;
        src64 <= 16'hf618;
        src65 <= 16'h5571;
        src66 <= 16'h19ee;
        src67 <= 16'hb985;
        src68 <= 16'h57d7;
        src69 <= 16'h5760;
        src70 <= 16'ha7d3;
        src71 <= 16'hc559;
        src72 <= 16'hda4f;
        src73 <= 16'haaa6;
        src74 <= 16'hc814;
        src75 <= 16'h97a4;
        src76 <= 16'h744b;
        src77 <= 16'h69c8;
        src78 <= 16'hc38;
        src79 <= 16'h8419;
        src80 <= 16'h495;
        src81 <= 16'h78ea;
        src82 <= 16'h1124;
        src83 <= 16'ha150;
        src84 <= 16'h6ab4;
        src85 <= 16'hbfa1;
        src86 <= 16'h80ea;
        src87 <= 16'h192e;
        src88 <= 16'h3244;
        src89 <= 16'h3c3;
        src90 <= 16'h7506;
        src91 <= 16'h20c0;
        src92 <= 16'hbb45;
        src93 <= 16'hc16a;
        src94 <= 16'ha88f;
        src95 <= 16'hd88;
        src96 <= 16'hbd38;
        src97 <= 16'hef24;
        src98 <= 16'hb7;
        src99 <= 16'he46;
        src100 <= 16'he82b;
        src101 <= 16'h7815;
        src102 <= 16'hf585;
        src103 <= 16'h8551;
        src104 <= 16'hffd3;
        src105 <= 16'h57bd;
        src106 <= 16'hc847;
        src107 <= 16'h6df6;
        src108 <= 16'hc5db;
        src109 <= 16'h9123;
        src110 <= 16'hd21b;
        src111 <= 16'h8251;
        src112 <= 16'h9bd3;
        src113 <= 16'h5ea7;
        src114 <= 16'hfa62;
        src115 <= 16'h3d7d;
        src116 <= 16'hf451;
        src117 <= 16'hbb6d;
        src118 <= 16'he801;
        src119 <= 16'h22b5;
        src120 <= 16'hcb2f;
        src121 <= 16'hc3b8;
        src122 <= 16'h34e0;
        src123 <= 16'h9907;
        src124 <= 16'haada;
        src125 <= 16'hd0d9;
        src126 <= 16'h9b8a;
        src127 <= 16'h2bb5;
        exp <= 23'h4246cd;
        #1
        src0 <= 16'h5e23;
        src1 <= 16'hf811;
        src2 <= 16'h4da7;
        src3 <= 16'h9e63;
        src4 <= 16'ha3ab;
        src5 <= 16'hfe;
        src6 <= 16'hd4d1;
        src7 <= 16'he26b;
        src8 <= 16'hc97e;
        src9 <= 16'hbba6;
        src10 <= 16'h689c;
        src11 <= 16'hbb5b;
        src12 <= 16'h88d;
        src13 <= 16'hdb6a;
        src14 <= 16'hd7b2;
        src15 <= 16'hfcee;
        src16 <= 16'ha4f8;
        src17 <= 16'h8879;
        src18 <= 16'h7be9;
        src19 <= 16'h3e69;
        src20 <= 16'h21e8;
        src21 <= 16'h4296;
        src22 <= 16'h8ab3;
        src23 <= 16'hc31f;
        src24 <= 16'hddc8;
        src25 <= 16'hf8fb;
        src26 <= 16'h2025;
        src27 <= 16'h29c0;
        src28 <= 16'heeb6;
        src29 <= 16'hb102;
        src30 <= 16'h9318;
        src31 <= 16'h16c3;
        src32 <= 16'ha5a;
        src33 <= 16'hfc22;
        src34 <= 16'h81cb;
        src35 <= 16'h6a3;
        src36 <= 16'h95c7;
        src37 <= 16'h97dc;
        src38 <= 16'hdd01;
        src39 <= 16'hec8c;
        src40 <= 16'hd9f9;
        src41 <= 16'hc568;
        src42 <= 16'h289e;
        src43 <= 16'h2fd1;
        src44 <= 16'hb008;
        src45 <= 16'hb5ee;
        src46 <= 16'he3e2;
        src47 <= 16'hfacf;
        src48 <= 16'h6d8e;
        src49 <= 16'h69e;
        src50 <= 16'hd852;
        src51 <= 16'h7f4;
        src52 <= 16'h686f;
        src53 <= 16'he389;
        src54 <= 16'h7078;
        src55 <= 16'hb44f;
        src56 <= 16'h29e3;
        src57 <= 16'h63f0;
        src58 <= 16'hebce;
        src59 <= 16'hd34b;
        src60 <= 16'h2273;
        src61 <= 16'h5bb0;
        src62 <= 16'hd7f4;
        src63 <= 16'hc059;
        src64 <= 16'hc282;
        src65 <= 16'h4b66;
        src66 <= 16'hd531;
        src67 <= 16'ha994;
        src68 <= 16'hfc73;
        src69 <= 16'h3899;
        src70 <= 16'h410c;
        src71 <= 16'h9956;
        src72 <= 16'hce1a;
        src73 <= 16'hd6c1;
        src74 <= 16'h3c5a;
        src75 <= 16'h9eb8;
        src76 <= 16'h6f46;
        src77 <= 16'h7fbc;
        src78 <= 16'h5282;
        src79 <= 16'h230;
        src80 <= 16'h6300;
        src81 <= 16'h83cc;
        src82 <= 16'h4b51;
        src83 <= 16'hd6e7;
        src84 <= 16'h27;
        src85 <= 16'h178d;
        src86 <= 16'h1fd0;
        src87 <= 16'h5af5;
        src88 <= 16'h251a;
        src89 <= 16'h29cd;
        src90 <= 16'h47cd;
        src91 <= 16'hf061;
        src92 <= 16'hdf18;
        src93 <= 16'h8a83;
        src94 <= 16'h270c;
        src95 <= 16'h6018;
        src96 <= 16'h7289;
        src97 <= 16'h1cc4;
        src98 <= 16'hee0d;
        src99 <= 16'hf084;
        src100 <= 16'he574;
        src101 <= 16'he432;
        src102 <= 16'h40c4;
        src103 <= 16'hc50f;
        src104 <= 16'hfe83;
        src105 <= 16'h80d9;
        src106 <= 16'hb8b4;
        src107 <= 16'hb6fc;
        src108 <= 16'h92e6;
        src109 <= 16'hd56b;
        src110 <= 16'h20cc;
        src111 <= 16'h6f17;
        src112 <= 16'h6c50;
        src113 <= 16'h4e03;
        src114 <= 16'h5bfb;
        src115 <= 16'h9cfb;
        src116 <= 16'hd798;
        src117 <= 16'h32c6;
        src118 <= 16'h7177;
        src119 <= 16'h75dd;
        src120 <= 16'ha860;
        src121 <= 16'h3747;
        src122 <= 16'h178a;
        src123 <= 16'h244;
        src124 <= 16'hc0d;
        src125 <= 16'hd285;
        src126 <= 16'h3d7f;
        src127 <= 16'hfff2;
        exp <= 23'h434158;
        #1
        src0 <= 16'he67a;
        src1 <= 16'h4b6e;
        src2 <= 16'h6c67;
        src3 <= 16'h1aeb;
        src4 <= 16'h128a;
        src5 <= 16'h371c;
        src6 <= 16'h4e44;
        src7 <= 16'ha7f6;
        src8 <= 16'h92ba;
        src9 <= 16'h7b31;
        src10 <= 16'hc6e4;
        src11 <= 16'h1d59;
        src12 <= 16'h14b0;
        src13 <= 16'h44a3;
        src14 <= 16'h3ea7;
        src15 <= 16'h73f1;
        src16 <= 16'hc743;
        src17 <= 16'h5a38;
        src18 <= 16'hc20d;
        src19 <= 16'hee14;
        src20 <= 16'h25f4;
        src21 <= 16'h2433;
        src22 <= 16'he0c7;
        src23 <= 16'h191e;
        src24 <= 16'hb4aa;
        src25 <= 16'h9b4b;
        src26 <= 16'h867d;
        src27 <= 16'hc345;
        src28 <= 16'hbe23;
        src29 <= 16'h94a8;
        src30 <= 16'h52;
        src31 <= 16'h9110;
        src32 <= 16'h3cb4;
        src33 <= 16'h835b;
        src34 <= 16'haab6;
        src35 <= 16'hfebb;
        src36 <= 16'hf3c6;
        src37 <= 16'h977c;
        src38 <= 16'had56;
        src39 <= 16'h5a62;
        src40 <= 16'hb34d;
        src41 <= 16'h8749;
        src42 <= 16'h3da5;
        src43 <= 16'h1ca9;
        src44 <= 16'hdd14;
        src45 <= 16'h5aa5;
        src46 <= 16'h9bf1;
        src47 <= 16'h1a8c;
        src48 <= 16'hb837;
        src49 <= 16'h8875;
        src50 <= 16'hb017;
        src51 <= 16'h5b5f;
        src52 <= 16'hb68d;
        src53 <= 16'h25c0;
        src54 <= 16'he9a2;
        src55 <= 16'hb5d0;
        src56 <= 16'h818b;
        src57 <= 16'hb7f5;
        src58 <= 16'hb978;
        src59 <= 16'h4e40;
        src60 <= 16'he469;
        src61 <= 16'h46a4;
        src62 <= 16'hb45b;
        src63 <= 16'h110e;
        src64 <= 16'hc48a;
        src65 <= 16'hcabe;
        src66 <= 16'hcafb;
        src67 <= 16'h25cf;
        src68 <= 16'h6e3a;
        src69 <= 16'ha273;
        src70 <= 16'h6848;
        src71 <= 16'ha95e;
        src72 <= 16'h5952;
        src73 <= 16'haf19;
        src74 <= 16'h3041;
        src75 <= 16'h48c4;
        src76 <= 16'hea0a;
        src77 <= 16'h69e7;
        src78 <= 16'h1c7a;
        src79 <= 16'haa88;
        src80 <= 16'h7abf;
        src81 <= 16'hb009;
        src82 <= 16'h4f28;
        src83 <= 16'h28bb;
        src84 <= 16'hccd7;
        src85 <= 16'hc995;
        src86 <= 16'h38bd;
        src87 <= 16'h2830;
        src88 <= 16'h7270;
        src89 <= 16'h82be;
        src90 <= 16'ha635;
        src91 <= 16'haa01;
        src92 <= 16'h7a24;
        src93 <= 16'hb92c;
        src94 <= 16'hb944;
        src95 <= 16'h5414;
        src96 <= 16'h7cf9;
        src97 <= 16'h2f52;
        src98 <= 16'h2d29;
        src99 <= 16'h4af;
        src100 <= 16'h7ef9;
        src101 <= 16'h1419;
        src102 <= 16'hfb45;
        src103 <= 16'h2e98;
        src104 <= 16'hd5e3;
        src105 <= 16'h8afa;
        src106 <= 16'hc6fd;
        src107 <= 16'h567;
        src108 <= 16'hd0c1;
        src109 <= 16'he29c;
        src110 <= 16'hb9e6;
        src111 <= 16'h7a58;
        src112 <= 16'hda9d;
        src113 <= 16'h7f66;
        src114 <= 16'h964b;
        src115 <= 16'h533e;
        src116 <= 16'hb031;
        src117 <= 16'h4101;
        src118 <= 16'h3671;
        src119 <= 16'h14ef;
        src120 <= 16'hc161;
        src121 <= 16'hb487;
        src122 <= 16'hd8f7;
        src123 <= 16'h3f82;
        src124 <= 16'h43d7;
        src125 <= 16'h18f2;
        src126 <= 16'h7170;
        src127 <= 16'h6d4f;
        exp <= 23'h3f5ca9;
        #1
        src0 <= 16'h84d5;
        src1 <= 16'h26c8;
        src2 <= 16'h44ea;
        src3 <= 16'hfee9;
        src4 <= 16'h1933;
        src5 <= 16'hc07a;
        src6 <= 16'hf24e;
        src7 <= 16'hceeb;
        src8 <= 16'h622a;
        src9 <= 16'h588a;
        src10 <= 16'h3b1e;
        src11 <= 16'hb7cd;
        src12 <= 16'hd149;
        src13 <= 16'hf25d;
        src14 <= 16'h3816;
        src15 <= 16'h8b88;
        src16 <= 16'h91bb;
        src17 <= 16'hc912;
        src18 <= 16'h73bf;
        src19 <= 16'h4148;
        src20 <= 16'h665f;
        src21 <= 16'h6d7a;
        src22 <= 16'hb291;
        src23 <= 16'hfc39;
        src24 <= 16'h693a;
        src25 <= 16'h6b2f;
        src26 <= 16'hc5a;
        src27 <= 16'h22b5;
        src28 <= 16'h2ee2;
        src29 <= 16'h4cf8;
        src30 <= 16'ha963;
        src31 <= 16'hf3cb;
        src32 <= 16'hf578;
        src33 <= 16'h88ae;
        src34 <= 16'he7df;
        src35 <= 16'h6327;
        src36 <= 16'h4edc;
        src37 <= 16'h884b;
        src38 <= 16'h406b;
        src39 <= 16'h724f;
        src40 <= 16'h8ae0;
        src41 <= 16'h3668;
        src42 <= 16'hbe5e;
        src43 <= 16'hdf10;
        src44 <= 16'haf6a;
        src45 <= 16'h50d;
        src46 <= 16'hef94;
        src47 <= 16'h27d6;
        src48 <= 16'h4d7;
        src49 <= 16'hafe0;
        src50 <= 16'h1e77;
        src51 <= 16'hd77a;
        src52 <= 16'h7fb5;
        src53 <= 16'he715;
        src54 <= 16'h7911;
        src55 <= 16'heeda;
        src56 <= 16'hb646;
        src57 <= 16'h6eb5;
        src58 <= 16'h3f67;
        src59 <= 16'hac49;
        src60 <= 16'hac64;
        src61 <= 16'hfdcc;
        src62 <= 16'hc7c2;
        src63 <= 16'hc81a;
        src64 <= 16'h9698;
        src65 <= 16'hb32d;
        src66 <= 16'hde5a;
        src67 <= 16'hadc8;
        src68 <= 16'hc5e4;
        src69 <= 16'h7259;
        src70 <= 16'h5e13;
        src71 <= 16'h998d;
        src72 <= 16'h8f3a;
        src73 <= 16'h4f58;
        src74 <= 16'hc674;
        src75 <= 16'h68b1;
        src76 <= 16'h299d;
        src77 <= 16'hcd8b;
        src78 <= 16'hbd44;
        src79 <= 16'h1625;
        src80 <= 16'hc50a;
        src81 <= 16'h8d23;
        src82 <= 16'h9a17;
        src83 <= 16'h18f0;
        src84 <= 16'h78f8;
        src85 <= 16'hfbf2;
        src86 <= 16'h75d9;
        src87 <= 16'h46c4;
        src88 <= 16'hf2d7;
        src89 <= 16'h3491;
        src90 <= 16'h763c;
        src91 <= 16'hfc34;
        src92 <= 16'hca43;
        src93 <= 16'hbcab;
        src94 <= 16'he544;
        src95 <= 16'h8a8b;
        src96 <= 16'h8a1d;
        src97 <= 16'h286f;
        src98 <= 16'hb938;
        src99 <= 16'hf4a7;
        src100 <= 16'h7879;
        src101 <= 16'h5c8c;
        src102 <= 16'hcf5b;
        src103 <= 16'h97ac;
        src104 <= 16'h3031;
        src105 <= 16'h1b66;
        src106 <= 16'hce21;
        src107 <= 16'he2c1;
        src108 <= 16'hccaa;
        src109 <= 16'hb769;
        src110 <= 16'h8c0c;
        src111 <= 16'h8bc1;
        src112 <= 16'hde07;
        src113 <= 16'hc0f2;
        src114 <= 16'h668d;
        src115 <= 16'hdded;
        src116 <= 16'h7d61;
        src117 <= 16'hb2d5;
        src118 <= 16'h7797;
        src119 <= 16'hba40;
        src120 <= 16'h29ae;
        src121 <= 16'h8f34;
        src122 <= 16'h47cd;
        src123 <= 16'h8c16;
        src124 <= 16'h60d0;
        src125 <= 16'hb8a1;
        src126 <= 16'hb73a;
        src127 <= 16'h2e77;
        exp <= 23'h475b7b;
        #1
        src0 <= 16'h2d55;
        src1 <= 16'h27ff;
        src2 <= 16'h5ce7;
        src3 <= 16'h9459;
        src4 <= 16'hea9e;
        src5 <= 16'h2a90;
        src6 <= 16'h8d8;
        src7 <= 16'h7886;
        src8 <= 16'h5aad;
        src9 <= 16'h5b55;
        src10 <= 16'hd11b;
        src11 <= 16'h28cb;
        src12 <= 16'he90c;
        src13 <= 16'h340a;
        src14 <= 16'h380a;
        src15 <= 16'h1feb;
        src16 <= 16'h5338;
        src17 <= 16'h9461;
        src18 <= 16'h2234;
        src19 <= 16'hd127;
        src20 <= 16'hfa6;
        src21 <= 16'h7d48;
        src22 <= 16'h569b;
        src23 <= 16'hcec4;
        src24 <= 16'he0a6;
        src25 <= 16'h2a69;
        src26 <= 16'ha617;
        src27 <= 16'h3aad;
        src28 <= 16'h9eee;
        src29 <= 16'h4dde;
        src30 <= 16'hefd2;
        src31 <= 16'h5910;
        src32 <= 16'hd212;
        src33 <= 16'h62d0;
        src34 <= 16'h211c;
        src35 <= 16'h81cb;
        src36 <= 16'h76fa;
        src37 <= 16'hf937;
        src38 <= 16'hc5aa;
        src39 <= 16'h225b;
        src40 <= 16'he860;
        src41 <= 16'hefed;
        src42 <= 16'h5af0;
        src43 <= 16'h8868;
        src44 <= 16'h6739;
        src45 <= 16'hd394;
        src46 <= 16'hee34;
        src47 <= 16'h5627;
        src48 <= 16'h2a99;
        src49 <= 16'h95cc;
        src50 <= 16'he5af;
        src51 <= 16'h12da;
        src52 <= 16'hc3b0;
        src53 <= 16'h714d;
        src54 <= 16'hc0b7;
        src55 <= 16'he8b0;
        src56 <= 16'h569;
        src57 <= 16'h531b;
        src58 <= 16'he2f6;
        src59 <= 16'hc499;
        src60 <= 16'h95e3;
        src61 <= 16'h8e77;
        src62 <= 16'h67d3;
        src63 <= 16'h91a2;
        src64 <= 16'h4ee1;
        src65 <= 16'hac0b;
        src66 <= 16'ha5e0;
        src67 <= 16'he504;
        src68 <= 16'ha2f0;
        src69 <= 16'h7afe;
        src70 <= 16'h2e88;
        src71 <= 16'h302e;
        src72 <= 16'hffd6;
        src73 <= 16'h3369;
        src74 <= 16'hc9f8;
        src75 <= 16'hf7e9;
        src76 <= 16'hc510;
        src77 <= 16'heece;
        src78 <= 16'h3839;
        src79 <= 16'heda1;
        src80 <= 16'h905c;
        src81 <= 16'hb6cc;
        src82 <= 16'h4240;
        src83 <= 16'h4d78;
        src84 <= 16'hae9;
        src85 <= 16'h1a73;
        src86 <= 16'h755;
        src87 <= 16'h7050;
        src88 <= 16'hc188;
        src89 <= 16'hc467;
        src90 <= 16'hf698;
        src91 <= 16'heca4;
        src92 <= 16'hbc0b;
        src93 <= 16'hc374;
        src94 <= 16'h1bf4;
        src95 <= 16'h82d9;
        src96 <= 16'h394f;
        src97 <= 16'hc856;
        src98 <= 16'h1e8f;
        src99 <= 16'h469e;
        src100 <= 16'hdc3e;
        src101 <= 16'h3a57;
        src102 <= 16'h8eed;
        src103 <= 16'hb3b7;
        src104 <= 16'hf4e3;
        src105 <= 16'habf6;
        src106 <= 16'h4db9;
        src107 <= 16'h9ae0;
        src108 <= 16'h23e2;
        src109 <= 16'h90a9;
        src110 <= 16'h3c5e;
        src111 <= 16'hcdf8;
        src112 <= 16'heeea;
        src113 <= 16'h54ee;
        src114 <= 16'hbc39;
        src115 <= 16'h3841;
        src116 <= 16'h4fd7;
        src117 <= 16'he2e;
        src118 <= 16'hbb40;
        src119 <= 16'hd309;
        src120 <= 16'h48df;
        src121 <= 16'h3ddd;
        src122 <= 16'h26fe;
        src123 <= 16'ha3d;
        src124 <= 16'h9553;
        src125 <= 16'h8181;
        src126 <= 16'he74b;
        src127 <= 16'h101f;
        exp <= 23'h4090ac;
        #1
        src0 <= 16'hde1e;
        src1 <= 16'h8864;
        src2 <= 16'he4dd;
        src3 <= 16'h72ff;
        src4 <= 16'h9b0c;
        src5 <= 16'h3cbf;
        src6 <= 16'hb032;
        src7 <= 16'h1b23;
        src8 <= 16'hc3da;
        src9 <= 16'h9282;
        src10 <= 16'h4153;
        src11 <= 16'h4fa3;
        src12 <= 16'hc928;
        src13 <= 16'h7ec9;
        src14 <= 16'hb71e;
        src15 <= 16'h989c;
        src16 <= 16'h996;
        src17 <= 16'h41e9;
        src18 <= 16'h87ea;
        src19 <= 16'hef21;
        src20 <= 16'h2e4c;
        src21 <= 16'h979f;
        src22 <= 16'h8f34;
        src23 <= 16'hf37;
        src24 <= 16'h489c;
        src25 <= 16'h4b70;
        src26 <= 16'hdc94;
        src27 <= 16'hb1a5;
        src28 <= 16'h4d3;
        src29 <= 16'he5f3;
        src30 <= 16'h369f;
        src31 <= 16'h5152;
        src32 <= 16'hca95;
        src33 <= 16'hf9af;
        src34 <= 16'h8875;
        src35 <= 16'h81ed;
        src36 <= 16'h7ab7;
        src37 <= 16'h9d7c;
        src38 <= 16'hdda1;
        src39 <= 16'he4d3;
        src40 <= 16'h2cd6;
        src41 <= 16'hc0fa;
        src42 <= 16'h10ee;
        src43 <= 16'hb0df;
        src44 <= 16'h8d9f;
        src45 <= 16'h9fde;
        src46 <= 16'hc3f7;
        src47 <= 16'ha7a0;
        src48 <= 16'hdda7;
        src49 <= 16'hbaad;
        src50 <= 16'h29af;
        src51 <= 16'hb6e5;
        src52 <= 16'h14d;
        src53 <= 16'h8dbf;
        src54 <= 16'h178f;
        src55 <= 16'h76f7;
        src56 <= 16'h737;
        src57 <= 16'h774e;
        src58 <= 16'h8c8a;
        src59 <= 16'h7ef5;
        src60 <= 16'hc00f;
        src61 <= 16'h6411;
        src62 <= 16'h88c8;
        src63 <= 16'h3ade;
        src64 <= 16'h583d;
        src65 <= 16'h6a9c;
        src66 <= 16'he59d;
        src67 <= 16'h5d7b;
        src68 <= 16'h32a5;
        src69 <= 16'hbeca;
        src70 <= 16'hb5a4;
        src71 <= 16'hfcf5;
        src72 <= 16'hcee7;
        src73 <= 16'h2a7a;
        src74 <= 16'ha4f9;
        src75 <= 16'h1a21;
        src76 <= 16'h82a7;
        src77 <= 16'h7427;
        src78 <= 16'hc49d;
        src79 <= 16'h4db;
        src80 <= 16'hff6c;
        src81 <= 16'hfa9;
        src82 <= 16'h7a93;
        src83 <= 16'h3876;
        src84 <= 16'hcfc1;
        src85 <= 16'h384;
        src86 <= 16'hff5b;
        src87 <= 16'h78ab;
        src88 <= 16'h9289;
        src89 <= 16'h7a29;
        src90 <= 16'h38b1;
        src91 <= 16'h5584;
        src92 <= 16'hd540;
        src93 <= 16'hff2f;
        src94 <= 16'hd331;
        src95 <= 16'hacad;
        src96 <= 16'h70f;
        src97 <= 16'h344d;
        src98 <= 16'h4792;
        src99 <= 16'haa7a;
        src100 <= 16'hb1ae;
        src101 <= 16'ha1f3;
        src102 <= 16'h7cfd;
        src103 <= 16'hd8dc;
        src104 <= 16'hf03d;
        src105 <= 16'h381a;
        src106 <= 16'h96ce;
        src107 <= 16'h82b7;
        src108 <= 16'ha086;
        src109 <= 16'h8f7c;
        src110 <= 16'h9a5e;
        src111 <= 16'h67f0;
        src112 <= 16'h758f;
        src113 <= 16'hd958;
        src114 <= 16'h61e3;
        src115 <= 16'h86e7;
        src116 <= 16'he5e1;
        src117 <= 16'hef73;
        src118 <= 16'hfebe;
        src119 <= 16'hda0;
        src120 <= 16'hb747;
        src121 <= 16'hc3fa;
        src122 <= 16'h7419;
        src123 <= 16'h54c1;
        src124 <= 16'ha358;
        src125 <= 16'hb7f3;
        src126 <= 16'h511e;
        src127 <= 16'h9279;
        exp <= 23'h439d5e;
        #1
        src0 <= 16'hcd7;
        src1 <= 16'h107c;
        src2 <= 16'h8e6f;
        src3 <= 16'hf9fe;
        src4 <= 16'ha4db;
        src5 <= 16'h3f69;
        src6 <= 16'h6727;
        src7 <= 16'hd090;
        src8 <= 16'hfbb3;
        src9 <= 16'hb695;
        src10 <= 16'hc7ee;
        src11 <= 16'h84ef;
        src12 <= 16'h4ab8;
        src13 <= 16'hb52d;
        src14 <= 16'h54cc;
        src15 <= 16'hcfc6;
        src16 <= 16'h9774;
        src17 <= 16'hd7e1;
        src18 <= 16'h1374;
        src19 <= 16'he18b;
        src20 <= 16'h75ad;
        src21 <= 16'hfe3f;
        src22 <= 16'h3571;
        src23 <= 16'h993b;
        src24 <= 16'he2d7;
        src25 <= 16'h6ea0;
        src26 <= 16'hf126;
        src27 <= 16'h38ad;
        src28 <= 16'h1d36;
        src29 <= 16'h54b2;
        src30 <= 16'h9995;
        src31 <= 16'he49d;
        src32 <= 16'h481c;
        src33 <= 16'h2737;
        src34 <= 16'h6514;
        src35 <= 16'hffcd;
        src36 <= 16'hd86c;
        src37 <= 16'hc624;
        src38 <= 16'ha470;
        src39 <= 16'hbcf6;
        src40 <= 16'ha0d;
        src41 <= 16'haaee;
        src42 <= 16'h699c;
        src43 <= 16'h8a4f;
        src44 <= 16'hd8fa;
        src45 <= 16'he1ae;
        src46 <= 16'hdd95;
        src47 <= 16'hbcaa;
        src48 <= 16'hef50;
        src49 <= 16'h21e8;
        src50 <= 16'hd32f;
        src51 <= 16'h6d01;
        src52 <= 16'hc582;
        src53 <= 16'h35cd;
        src54 <= 16'hc5f;
        src55 <= 16'h461;
        src56 <= 16'h5c73;
        src57 <= 16'h4a60;
        src58 <= 16'h1f79;
        src59 <= 16'h79d;
        src60 <= 16'h594a;
        src61 <= 16'he171;
        src62 <= 16'hfa58;
        src63 <= 16'he70d;
        src64 <= 16'hbd30;
        src65 <= 16'h4c15;
        src66 <= 16'hab5b;
        src67 <= 16'h5c7a;
        src68 <= 16'h87a2;
        src69 <= 16'heb9e;
        src70 <= 16'h187c;
        src71 <= 16'hc2d4;
        src72 <= 16'ha1d2;
        src73 <= 16'h83a0;
        src74 <= 16'h50d7;
        src75 <= 16'h9010;
        src76 <= 16'h766e;
        src77 <= 16'hfddf;
        src78 <= 16'h78f0;
        src79 <= 16'h9506;
        src80 <= 16'h2127;
        src81 <= 16'h17d4;
        src82 <= 16'h193;
        src83 <= 16'he38e;
        src84 <= 16'h761f;
        src85 <= 16'hddb0;
        src86 <= 16'h5e73;
        src87 <= 16'h994f;
        src88 <= 16'h8ca7;
        src89 <= 16'h121d;
        src90 <= 16'haf37;
        src91 <= 16'heb20;
        src92 <= 16'hfde3;
        src93 <= 16'hf3b5;
        src94 <= 16'h91ab;
        src95 <= 16'hd5a6;
        src96 <= 16'hb292;
        src97 <= 16'hfdda;
        src98 <= 16'h67b3;
        src99 <= 16'h2644;
        src100 <= 16'h5a47;
        src101 <= 16'h6e6d;
        src102 <= 16'hf4ad;
        src103 <= 16'hcb3c;
        src104 <= 16'h5024;
        src105 <= 16'h57c7;
        src106 <= 16'h6935;
        src107 <= 16'hf857;
        src108 <= 16'h260a;
        src109 <= 16'h15d9;
        src110 <= 16'h16e9;
        src111 <= 16'hcd23;
        src112 <= 16'h706f;
        src113 <= 16'h4974;
        src114 <= 16'h5754;
        src115 <= 16'hcf34;
        src116 <= 16'h6fb5;
        src117 <= 16'h5c80;
        src118 <= 16'he932;
        src119 <= 16'hd7e5;
        src120 <= 16'hc3b2;
        src121 <= 16'hc368;
        src122 <= 16'h1202;
        src123 <= 16'h2fe4;
        src124 <= 16'h5c3d;
        src125 <= 16'hc54a;
        src126 <= 16'h6018;
        src127 <= 16'h4950;
        exp <= 23'h44e721;
        #1
        src0 <= 16'h363a;
        src1 <= 16'h23f0;
        src2 <= 16'hd1ff;
        src3 <= 16'hc4fa;
        src4 <= 16'h3b42;
        src5 <= 16'h1f62;
        src6 <= 16'h1bd9;
        src7 <= 16'hacdf;
        src8 <= 16'hee57;
        src9 <= 16'h1d3a;
        src10 <= 16'hb427;
        src11 <= 16'h8a71;
        src12 <= 16'ha5bf;
        src13 <= 16'h40b3;
        src14 <= 16'h793f;
        src15 <= 16'hca72;
        src16 <= 16'h1a1c;
        src17 <= 16'h6770;
        src18 <= 16'h96c5;
        src19 <= 16'hf06e;
        src20 <= 16'h9b2b;
        src21 <= 16'h37e5;
        src22 <= 16'hfa99;
        src23 <= 16'h1c36;
        src24 <= 16'he1a5;
        src25 <= 16'hb10b;
        src26 <= 16'hc42;
        src27 <= 16'h6d25;
        src28 <= 16'hd206;
        src29 <= 16'h9a16;
        src30 <= 16'hd6d1;
        src31 <= 16'hc788;
        src32 <= 16'h9d31;
        src33 <= 16'h405f;
        src34 <= 16'ha33e;
        src35 <= 16'h9185;
        src36 <= 16'h5b5c;
        src37 <= 16'hac8;
        src38 <= 16'hdb90;
        src39 <= 16'h16df;
        src40 <= 16'h2599;
        src41 <= 16'h64a7;
        src42 <= 16'hec11;
        src43 <= 16'h8fc2;
        src44 <= 16'h7076;
        src45 <= 16'h967c;
        src46 <= 16'hc3e9;
        src47 <= 16'hbe44;
        src48 <= 16'hf43b;
        src49 <= 16'he1e2;
        src50 <= 16'hb6c7;
        src51 <= 16'h79bd;
        src52 <= 16'h9ac4;
        src53 <= 16'hc84b;
        src54 <= 16'hba54;
        src55 <= 16'ha434;
        src56 <= 16'h67b9;
        src57 <= 16'h64db;
        src58 <= 16'h134f;
        src59 <= 16'h8ed0;
        src60 <= 16'h5c00;
        src61 <= 16'h75c2;
        src62 <= 16'hf51a;
        src63 <= 16'h9da1;
        src64 <= 16'h3b34;
        src65 <= 16'hb95b;
        src66 <= 16'h2edd;
        src67 <= 16'h743f;
        src68 <= 16'h44d4;
        src69 <= 16'h715a;
        src70 <= 16'h2983;
        src71 <= 16'h6fb2;
        src72 <= 16'hf4a5;
        src73 <= 16'h9dbd;
        src74 <= 16'h3979;
        src75 <= 16'ha8d9;
        src76 <= 16'h857d;
        src77 <= 16'h9078;
        src78 <= 16'hd0aa;
        src79 <= 16'h9d28;
        src80 <= 16'hd63d;
        src81 <= 16'hf176;
        src82 <= 16'h26eb;
        src83 <= 16'h5a33;
        src84 <= 16'h1a63;
        src85 <= 16'hdc03;
        src86 <= 16'hc13b;
        src87 <= 16'hb41;
        src88 <= 16'h7174;
        src89 <= 16'hdd6b;
        src90 <= 16'he121;
        src91 <= 16'h8298;
        src92 <= 16'h3900;
        src93 <= 16'h6efb;
        src94 <= 16'h4dcd;
        src95 <= 16'h8c66;
        src96 <= 16'h482e;
        src97 <= 16'h5375;
        src98 <= 16'hc223;
        src99 <= 16'he8d4;
        src100 <= 16'h704b;
        src101 <= 16'hc62f;
        src102 <= 16'h9f48;
        src103 <= 16'he909;
        src104 <= 16'h54;
        src105 <= 16'h345a;
        src106 <= 16'h467e;
        src107 <= 16'hee71;
        src108 <= 16'h5a7a;
        src109 <= 16'h907e;
        src110 <= 16'h8c1f;
        src111 <= 16'h8276;
        src112 <= 16'h597e;
        src113 <= 16'h8f;
        src114 <= 16'h6a29;
        src115 <= 16'h4533;
        src116 <= 16'h1e00;
        src117 <= 16'h8561;
        src118 <= 16'h6605;
        src119 <= 16'haf8a;
        src120 <= 16'h4ad9;
        src121 <= 16'h7880;
        src122 <= 16'h14c;
        src123 <= 16'hee75;
        src124 <= 16'h1c94;
        src125 <= 16'h3e38;
        src126 <= 16'h6703;
        src127 <= 16'h59bd;
        exp <= 23'h404105;
        #1
        src0 <= 16'hba74;
        src1 <= 16'ha701;
        src2 <= 16'h9554;
        src3 <= 16'h150;
        src4 <= 16'h5679;
        src5 <= 16'h67c1;
        src6 <= 16'hba2;
        src7 <= 16'hc18e;
        src8 <= 16'h3974;
        src9 <= 16'hd2e7;
        src10 <= 16'he228;
        src11 <= 16'h82ff;
        src12 <= 16'hf296;
        src13 <= 16'hac28;
        src14 <= 16'h334;
        src15 <= 16'h794a;
        src16 <= 16'h3ae8;
        src17 <= 16'h1c75;
        src18 <= 16'h8ba1;
        src19 <= 16'hd8a5;
        src20 <= 16'h7d59;
        src21 <= 16'h941;
        src22 <= 16'h6ae9;
        src23 <= 16'h7675;
        src24 <= 16'hab49;
        src25 <= 16'h5eaf;
        src26 <= 16'hbdfc;
        src27 <= 16'hf143;
        src28 <= 16'h64e6;
        src29 <= 16'hd0fe;
        src30 <= 16'he37e;
        src31 <= 16'hd4d5;
        src32 <= 16'h3ca;
        src33 <= 16'h1436;
        src34 <= 16'h8c86;
        src35 <= 16'hd649;
        src36 <= 16'h1aae;
        src37 <= 16'h208c;
        src38 <= 16'h3264;
        src39 <= 16'h82ff;
        src40 <= 16'hd8d5;
        src41 <= 16'h59ad;
        src42 <= 16'hbcab;
        src43 <= 16'hf102;
        src44 <= 16'h33a6;
        src45 <= 16'h7c2d;
        src46 <= 16'hc4db;
        src47 <= 16'h163f;
        src48 <= 16'h8307;
        src49 <= 16'h3641;
        src50 <= 16'h2452;
        src51 <= 16'h1287;
        src52 <= 16'hb0df;
        src53 <= 16'h4a70;
        src54 <= 16'he54e;
        src55 <= 16'h10b1;
        src56 <= 16'ha781;
        src57 <= 16'h2a83;
        src58 <= 16'hc659;
        src59 <= 16'had18;
        src60 <= 16'he117;
        src61 <= 16'h5c8a;
        src62 <= 16'hdaa9;
        src63 <= 16'hcdb7;
        src64 <= 16'h1d2b;
        src65 <= 16'h3a34;
        src66 <= 16'h53fe;
        src67 <= 16'h8bbe;
        src68 <= 16'h6dec;
        src69 <= 16'h5b9a;
        src70 <= 16'h2539;
        src71 <= 16'h7240;
        src72 <= 16'h9305;
        src73 <= 16'he73c;
        src74 <= 16'h379b;
        src75 <= 16'he3af;
        src76 <= 16'ha59f;
        src77 <= 16'hec1;
        src78 <= 16'h8f95;
        src79 <= 16'h4c21;
        src80 <= 16'ha348;
        src81 <= 16'hea0d;
        src82 <= 16'hfe92;
        src83 <= 16'hb83e;
        src84 <= 16'ha5c2;
        src85 <= 16'he4f;
        src86 <= 16'h321f;
        src87 <= 16'h2278;
        src88 <= 16'h8162;
        src89 <= 16'h57d4;
        src90 <= 16'h8bb;
        src91 <= 16'hf38e;
        src92 <= 16'h1784;
        src93 <= 16'h9189;
        src94 <= 16'h6c91;
        src95 <= 16'h114b;
        src96 <= 16'hfca2;
        src97 <= 16'h7a6f;
        src98 <= 16'h48af;
        src99 <= 16'h4ba;
        src100 <= 16'h264c;
        src101 <= 16'h91fb;
        src102 <= 16'h5c35;
        src103 <= 16'h5a8a;
        src104 <= 16'h6992;
        src105 <= 16'h2b5;
        src106 <= 16'h9dd9;
        src107 <= 16'h1862;
        src108 <= 16'hcd39;
        src109 <= 16'hc78a;
        src110 <= 16'hdc49;
        src111 <= 16'h25a1;
        src112 <= 16'h5e8d;
        src113 <= 16'h79ed;
        src114 <= 16'h8caf;
        src115 <= 16'h7dcc;
        src116 <= 16'h91ba;
        src117 <= 16'he8b6;
        src118 <= 16'h715;
        src119 <= 16'h4da1;
        src120 <= 16'h21f;
        src121 <= 16'h5e0a;
        src122 <= 16'h2c57;
        src123 <= 16'hfce4;
        src124 <= 16'h8966;
        src125 <= 16'h4152;
        src126 <= 16'hc90c;
        src127 <= 16'h4797;
        exp <= 23'h3bc930;
        #1
        src0 <= 16'h48a7;
        src1 <= 16'had5c;
        src2 <= 16'ha8c7;
        src3 <= 16'h8736;
        src4 <= 16'h7fed;
        src5 <= 16'h16f8;
        src6 <= 16'h12db;
        src7 <= 16'hbff1;
        src8 <= 16'hc3d3;
        src9 <= 16'h11f7;
        src10 <= 16'h718b;
        src11 <= 16'h86b0;
        src12 <= 16'h8d2;
        src13 <= 16'hb046;
        src14 <= 16'h79ef;
        src15 <= 16'he4bd;
        src16 <= 16'hd449;
        src17 <= 16'hfb93;
        src18 <= 16'hb848;
        src19 <= 16'hf802;
        src20 <= 16'h9948;
        src21 <= 16'h1038;
        src22 <= 16'h62df;
        src23 <= 16'h90;
        src24 <= 16'h7fbb;
        src25 <= 16'ha602;
        src26 <= 16'hb54f;
        src27 <= 16'h49cf;
        src28 <= 16'h6c8;
        src29 <= 16'hc639;
        src30 <= 16'hdf18;
        src31 <= 16'h9efc;
        src32 <= 16'h5b0c;
        src33 <= 16'h5189;
        src34 <= 16'h922c;
        src35 <= 16'h14b5;
        src36 <= 16'h87e6;
        src37 <= 16'h1043;
        src38 <= 16'h158f;
        src39 <= 16'hfdb2;
        src40 <= 16'h8d77;
        src41 <= 16'h562b;
        src42 <= 16'h7dae;
        src43 <= 16'h5a87;
        src44 <= 16'h385f;
        src45 <= 16'hfcef;
        src46 <= 16'h7bbf;
        src47 <= 16'hd0c4;
        src48 <= 16'ha5d5;
        src49 <= 16'h32e3;
        src50 <= 16'h769e;
        src51 <= 16'h1c1a;
        src52 <= 16'h8702;
        src53 <= 16'h7b9;
        src54 <= 16'h183b;
        src55 <= 16'h2490;
        src56 <= 16'h7d16;
        src57 <= 16'h12b5;
        src58 <= 16'h149;
        src59 <= 16'h4239;
        src60 <= 16'h8fa4;
        src61 <= 16'hb00;
        src62 <= 16'hcba4;
        src63 <= 16'h92cc;
        src64 <= 16'h2125;
        src65 <= 16'h9891;
        src66 <= 16'hae2c;
        src67 <= 16'he74c;
        src68 <= 16'hf340;
        src69 <= 16'hd875;
        src70 <= 16'h8552;
        src71 <= 16'h1885;
        src72 <= 16'h2cb;
        src73 <= 16'h5c22;
        src74 <= 16'hdddf;
        src75 <= 16'h8807;
        src76 <= 16'hcf32;
        src77 <= 16'h8d65;
        src78 <= 16'h27ef;
        src79 <= 16'h9a4d;
        src80 <= 16'h1815;
        src81 <= 16'hbe50;
        src82 <= 16'h30ad;
        src83 <= 16'h563e;
        src84 <= 16'h63fe;
        src85 <= 16'hc254;
        src86 <= 16'h40ca;
        src87 <= 16'h624a;
        src88 <= 16'hc1e6;
        src89 <= 16'h3a78;
        src90 <= 16'h2c12;
        src91 <= 16'h2ad2;
        src92 <= 16'hb04;
        src93 <= 16'h6564;
        src94 <= 16'h8d25;
        src95 <= 16'he913;
        src96 <= 16'h5adb;
        src97 <= 16'h9638;
        src98 <= 16'hc024;
        src99 <= 16'haa87;
        src100 <= 16'hbcfb;
        src101 <= 16'h93e9;
        src102 <= 16'h7184;
        src103 <= 16'hfb46;
        src104 <= 16'he25b;
        src105 <= 16'h6f7d;
        src106 <= 16'h69eb;
        src107 <= 16'he3c;
        src108 <= 16'hcae9;
        src109 <= 16'h61bd;
        src110 <= 16'h2fe3;
        src111 <= 16'hbef7;
        src112 <= 16'hc588;
        src113 <= 16'h5e63;
        src114 <= 16'h5fd6;
        src115 <= 16'hd554;
        src116 <= 16'h434e;
        src117 <= 16'h3e38;
        src118 <= 16'h503b;
        src119 <= 16'hb046;
        src120 <= 16'hf57f;
        src121 <= 16'haa32;
        src122 <= 16'he971;
        src123 <= 16'h3708;
        src124 <= 16'h1cc9;
        src125 <= 16'hfbf8;
        src126 <= 16'hc7cd;
        src127 <= 16'hc3a0;
        exp <= 23'h3dedb5;
        #1
        src0 <= 16'hf77d;
        src1 <= 16'hd052;
        src2 <= 16'h9d17;
        src3 <= 16'h51bb;
        src4 <= 16'h5ad6;
        src5 <= 16'h8f12;
        src6 <= 16'hd00;
        src7 <= 16'h1da7;
        src8 <= 16'he405;
        src9 <= 16'haed9;
        src10 <= 16'hed1b;
        src11 <= 16'hc744;
        src12 <= 16'h3e60;
        src13 <= 16'h87cb;
        src14 <= 16'hbd2b;
        src15 <= 16'h938d;
        src16 <= 16'h13d2;
        src17 <= 16'h1533;
        src18 <= 16'h2fd;
        src19 <= 16'h4bc0;
        src20 <= 16'h670e;
        src21 <= 16'h89b8;
        src22 <= 16'he9fb;
        src23 <= 16'h487d;
        src24 <= 16'he985;
        src25 <= 16'hd603;
        src26 <= 16'hc06e;
        src27 <= 16'h1de8;
        src28 <= 16'h7bed;
        src29 <= 16'h1f5c;
        src30 <= 16'h8f81;
        src31 <= 16'h8536;
        src32 <= 16'h714c;
        src33 <= 16'h93d6;
        src34 <= 16'hf613;
        src35 <= 16'hc4d4;
        src36 <= 16'he283;
        src37 <= 16'h2e3;
        src38 <= 16'h79fd;
        src39 <= 16'h817e;
        src40 <= 16'hc40;
        src41 <= 16'h84fe;
        src42 <= 16'he831;
        src43 <= 16'hca1;
        src44 <= 16'hd190;
        src45 <= 16'hac98;
        src46 <= 16'h16cb;
        src47 <= 16'h835a;
        src48 <= 16'hcad2;
        src49 <= 16'hb899;
        src50 <= 16'h80ce;
        src51 <= 16'h8009;
        src52 <= 16'h1961;
        src53 <= 16'h4954;
        src54 <= 16'h4a7a;
        src55 <= 16'hded6;
        src56 <= 16'h34e3;
        src57 <= 16'ha572;
        src58 <= 16'h7354;
        src59 <= 16'h674e;
        src60 <= 16'h45b7;
        src61 <= 16'h76d2;
        src62 <= 16'hf530;
        src63 <= 16'ha3e6;
        src64 <= 16'h1d35;
        src65 <= 16'h80e2;
        src66 <= 16'h4832;
        src67 <= 16'hfe6e;
        src68 <= 16'h4003;
        src69 <= 16'h7e89;
        src70 <= 16'h5ccf;
        src71 <= 16'hb4a2;
        src72 <= 16'hd4be;
        src73 <= 16'hde71;
        src74 <= 16'hb5ae;
        src75 <= 16'h2c25;
        src76 <= 16'he5d8;
        src77 <= 16'he5b8;
        src78 <= 16'ha3ea;
        src79 <= 16'h8675;
        src80 <= 16'he29d;
        src81 <= 16'hcb60;
        src82 <= 16'hf3a7;
        src83 <= 16'h4213;
        src84 <= 16'h1a;
        src85 <= 16'h2e96;
        src86 <= 16'h1d25;
        src87 <= 16'hc441;
        src88 <= 16'hfa0d;
        src89 <= 16'h3702;
        src90 <= 16'hd70d;
        src91 <= 16'h8e43;
        src92 <= 16'he8ff;
        src93 <= 16'hfb56;
        src94 <= 16'h7882;
        src95 <= 16'ha24c;
        src96 <= 16'hbfc7;
        src97 <= 16'h24ff;
        src98 <= 16'h250e;
        src99 <= 16'h16;
        src100 <= 16'heed7;
        src101 <= 16'hde9b;
        src102 <= 16'h3ef9;
        src103 <= 16'hedd3;
        src104 <= 16'h497a;
        src105 <= 16'h909a;
        src106 <= 16'hf41;
        src107 <= 16'h33be;
        src108 <= 16'h3cc;
        src109 <= 16'h64f8;
        src110 <= 16'h2b9b;
        src111 <= 16'ha3bf;
        src112 <= 16'h2437;
        src113 <= 16'h7cbb;
        src114 <= 16'h19d1;
        src115 <= 16'hb63e;
        src116 <= 16'hf332;
        src117 <= 16'hf82f;
        src118 <= 16'hb3c1;
        src119 <= 16'h6e16;
        src120 <= 16'h7bff;
        src121 <= 16'h829;
        src122 <= 16'h5af1;
        src123 <= 16'hc139;
        src124 <= 16'h6c67;
        src125 <= 16'h1dd3;
        src126 <= 16'hb936;
        src127 <= 16'hf3c5;
        exp <= 23'h41e45f;
        #1
        src0 <= 16'ha072;
        src1 <= 16'h7035;
        src2 <= 16'h61e0;
        src3 <= 16'h2b0a;
        src4 <= 16'haef9;
        src5 <= 16'h773;
        src6 <= 16'he8aa;
        src7 <= 16'hacbf;
        src8 <= 16'h4687;
        src9 <= 16'h501c;
        src10 <= 16'h7e7f;
        src11 <= 16'h79bd;
        src12 <= 16'hc387;
        src13 <= 16'h5b7e;
        src14 <= 16'h8064;
        src15 <= 16'h368f;
        src16 <= 16'h2916;
        src17 <= 16'h10d0;
        src18 <= 16'h9940;
        src19 <= 16'h332;
        src20 <= 16'h7acf;
        src21 <= 16'h4af4;
        src22 <= 16'h6bb9;
        src23 <= 16'h9162;
        src24 <= 16'h978b;
        src25 <= 16'hf237;
        src26 <= 16'h2a88;
        src27 <= 16'h689c;
        src28 <= 16'h43e8;
        src29 <= 16'h90bd;
        src30 <= 16'h8f65;
        src31 <= 16'hbf25;
        src32 <= 16'hcf4c;
        src33 <= 16'h4831;
        src34 <= 16'he5b;
        src35 <= 16'h7367;
        src36 <= 16'h4f42;
        src37 <= 16'ha06a;
        src38 <= 16'h8d40;
        src39 <= 16'h4187;
        src40 <= 16'h8993;
        src41 <= 16'hef65;
        src42 <= 16'hba7a;
        src43 <= 16'h54bf;
        src44 <= 16'h5eb4;
        src45 <= 16'hd657;
        src46 <= 16'he393;
        src47 <= 16'hd814;
        src48 <= 16'h1d0d;
        src49 <= 16'h1e61;
        src50 <= 16'hb5e7;
        src51 <= 16'hd081;
        src52 <= 16'h26a5;
        src53 <= 16'h29f2;
        src54 <= 16'h91a8;
        src55 <= 16'hf1d3;
        src56 <= 16'h3add;
        src57 <= 16'h1384;
        src58 <= 16'h2b30;
        src59 <= 16'hc653;
        src60 <= 16'h6290;
        src61 <= 16'h9239;
        src62 <= 16'haa37;
        src63 <= 16'h883a;
        src64 <= 16'h1bc8;
        src65 <= 16'h674d;
        src66 <= 16'h10e3;
        src67 <= 16'h32c2;
        src68 <= 16'h3587;
        src69 <= 16'h4ad5;
        src70 <= 16'h7daa;
        src71 <= 16'h32a5;
        src72 <= 16'h3b58;
        src73 <= 16'h5c3c;
        src74 <= 16'hbe9b;
        src75 <= 16'h78b8;
        src76 <= 16'h5e18;
        src77 <= 16'h12b1;
        src78 <= 16'h54d7;
        src79 <= 16'haa4d;
        src80 <= 16'hc00a;
        src81 <= 16'hb66e;
        src82 <= 16'hed18;
        src83 <= 16'h420e;
        src84 <= 16'hf06d;
        src85 <= 16'h93ab;
        src86 <= 16'hbd2a;
        src87 <= 16'h4f2f;
        src88 <= 16'h125a;
        src89 <= 16'hcf36;
        src90 <= 16'h2a25;
        src91 <= 16'h1210;
        src92 <= 16'h4e47;
        src93 <= 16'ha0c0;
        src94 <= 16'h1e96;
        src95 <= 16'ha3cb;
        src96 <= 16'h965a;
        src97 <= 16'hbeaf;
        src98 <= 16'hbfa3;
        src99 <= 16'hc71e;
        src100 <= 16'hede0;
        src101 <= 16'hb50;
        src102 <= 16'h1661;
        src103 <= 16'h901d;
        src104 <= 16'h7590;
        src105 <= 16'h6aa6;
        src106 <= 16'h9cbf;
        src107 <= 16'had3f;
        src108 <= 16'h60a0;
        src109 <= 16'h7701;
        src110 <= 16'hf014;
        src111 <= 16'h3094;
        src112 <= 16'h9214;
        src113 <= 16'ha87a;
        src114 <= 16'hb5e;
        src115 <= 16'h4806;
        src116 <= 16'habaa;
        src117 <= 16'ha987;
        src118 <= 16'h693d;
        src119 <= 16'h124;
        src120 <= 16'h2fb9;
        src121 <= 16'h8757;
        src122 <= 16'hcd1f;
        src123 <= 16'h8a43;
        src124 <= 16'h517c;
        src125 <= 16'h77aa;
        src126 <= 16'he3c1;
        src127 <= 16'h2033;
        exp <= 23'h3af79d;
        #1
        src0 <= 16'h2883;
        src1 <= 16'hbd5;
        src2 <= 16'hf295;
        src3 <= 16'h1f64;
        src4 <= 16'hc7ca;
        src5 <= 16'hbad6;
        src6 <= 16'h6a69;
        src7 <= 16'hf4c0;
        src8 <= 16'hd365;
        src9 <= 16'hd7b5;
        src10 <= 16'h8c83;
        src11 <= 16'h2ee4;
        src12 <= 16'ha1ae;
        src13 <= 16'hd5cc;
        src14 <= 16'hf541;
        src15 <= 16'h5c61;
        src16 <= 16'hc182;
        src17 <= 16'hb7dd;
        src18 <= 16'hf00e;
        src19 <= 16'hbb4d;
        src20 <= 16'hdb59;
        src21 <= 16'h9f62;
        src22 <= 16'h3aae;
        src23 <= 16'hc064;
        src24 <= 16'hadac;
        src25 <= 16'he0b1;
        src26 <= 16'h744;
        src27 <= 16'h3878;
        src28 <= 16'hb924;
        src29 <= 16'hf2c9;
        src30 <= 16'hc535;
        src31 <= 16'h41c0;
        src32 <= 16'h8e4c;
        src33 <= 16'h9fe2;
        src34 <= 16'hd988;
        src35 <= 16'hecac;
        src36 <= 16'hac01;
        src37 <= 16'hc26f;
        src38 <= 16'h4707;
        src39 <= 16'h151b;
        src40 <= 16'hfc98;
        src41 <= 16'h6e98;
        src42 <= 16'h2f50;
        src43 <= 16'hb45a;
        src44 <= 16'h82a0;
        src45 <= 16'h3ef6;
        src46 <= 16'h7809;
        src47 <= 16'h18d8;
        src48 <= 16'hb72;
        src49 <= 16'hce92;
        src50 <= 16'hbc30;
        src51 <= 16'h616f;
        src52 <= 16'h33a9;
        src53 <= 16'h92ed;
        src54 <= 16'h1a6c;
        src55 <= 16'hce2;
        src56 <= 16'hfad1;
        src57 <= 16'hc2f9;
        src58 <= 16'h97e8;
        src59 <= 16'h6e53;
        src60 <= 16'hba42;
        src61 <= 16'h559e;
        src62 <= 16'h22a4;
        src63 <= 16'h4fc6;
        src64 <= 16'h689d;
        src65 <= 16'h66f2;
        src66 <= 16'h777b;
        src67 <= 16'h336e;
        src68 <= 16'hfd;
        src69 <= 16'h75f9;
        src70 <= 16'he03f;
        src71 <= 16'h7717;
        src72 <= 16'h137d;
        src73 <= 16'heee6;
        src74 <= 16'h6ec8;
        src75 <= 16'hb6ca;
        src76 <= 16'h87f8;
        src77 <= 16'hcf99;
        src78 <= 16'h327f;
        src79 <= 16'hd90d;
        src80 <= 16'h5c7b;
        src81 <= 16'hd89d;
        src82 <= 16'hb0b9;
        src83 <= 16'h46c9;
        src84 <= 16'h1260;
        src85 <= 16'hd09b;
        src86 <= 16'h6f45;
        src87 <= 16'h8c5e;
        src88 <= 16'h9a60;
        src89 <= 16'ha392;
        src90 <= 16'h97d0;
        src91 <= 16'h50f7;
        src92 <= 16'hbb0;
        src93 <= 16'h8ec0;
        src94 <= 16'h41e6;
        src95 <= 16'h59a9;
        src96 <= 16'hcc4d;
        src97 <= 16'h329e;
        src98 <= 16'hc4c9;
        src99 <= 16'hc700;
        src100 <= 16'hbc99;
        src101 <= 16'h9f05;
        src102 <= 16'h9057;
        src103 <= 16'hf6a1;
        src104 <= 16'hdbb1;
        src105 <= 16'h55c3;
        src106 <= 16'h2fd0;
        src107 <= 16'h6005;
        src108 <= 16'hd6e0;
        src109 <= 16'h37b4;
        src110 <= 16'haaff;
        src111 <= 16'h568;
        src112 <= 16'h1515;
        src113 <= 16'h8b5a;
        src114 <= 16'h7c6e;
        src115 <= 16'h4828;
        src116 <= 16'h618e;
        src117 <= 16'h7812;
        src118 <= 16'he0ca;
        src119 <= 16'habb2;
        src120 <= 16'ha7db;
        src121 <= 16'h12ca;
        src122 <= 16'h6618;
        src123 <= 16'he6c2;
        src124 <= 16'hc8dd;
        src125 <= 16'h1f56;
        src126 <= 16'hd258;
        src127 <= 16'h4783;
        exp <= 23'h42fd56;
        #1
        src0 <= 16'h4313;
        src1 <= 16'h44d4;
        src2 <= 16'h1da3;
        src3 <= 16'hf1f8;
        src4 <= 16'h5bb3;
        src5 <= 16'h7b3e;
        src6 <= 16'h84;
        src7 <= 16'h41ce;
        src8 <= 16'h868d;
        src9 <= 16'h41f4;
        src10 <= 16'h342d;
        src11 <= 16'h7b6c;
        src12 <= 16'h4903;
        src13 <= 16'ha816;
        src14 <= 16'h695f;
        src15 <= 16'h7edc;
        src16 <= 16'h8a72;
        src17 <= 16'heffa;
        src18 <= 16'h60c6;
        src19 <= 16'hdb14;
        src20 <= 16'h2dcb;
        src21 <= 16'hf168;
        src22 <= 16'h1c4a;
        src23 <= 16'hfe63;
        src24 <= 16'hd057;
        src25 <= 16'h1d5b;
        src26 <= 16'hb639;
        src27 <= 16'h3f8;
        src28 <= 16'hf121;
        src29 <= 16'hd0b5;
        src30 <= 16'h891;
        src31 <= 16'he2ed;
        src32 <= 16'ha3ab;
        src33 <= 16'h3a85;
        src34 <= 16'h9e7d;
        src35 <= 16'hb14d;
        src36 <= 16'he856;
        src37 <= 16'hacb0;
        src38 <= 16'h26b;
        src39 <= 16'hb07b;
        src40 <= 16'h2dcf;
        src41 <= 16'h70cc;
        src42 <= 16'ha14e;
        src43 <= 16'hfb01;
        src44 <= 16'h2a5f;
        src45 <= 16'he7dd;
        src46 <= 16'h36b5;
        src47 <= 16'h5ca6;
        src48 <= 16'h3e3d;
        src49 <= 16'h6c71;
        src50 <= 16'hc31e;
        src51 <= 16'hf256;
        src52 <= 16'hf26c;
        src53 <= 16'hd698;
        src54 <= 16'h2074;
        src55 <= 16'hd7d4;
        src56 <= 16'h9786;
        src57 <= 16'he158;
        src58 <= 16'h2e0e;
        src59 <= 16'h39f5;
        src60 <= 16'hb25;
        src61 <= 16'hc176;
        src62 <= 16'h5b4c;
        src63 <= 16'hf64a;
        src64 <= 16'h9c93;
        src65 <= 16'h6a00;
        src66 <= 16'hd76c;
        src67 <= 16'h9f9;
        src68 <= 16'h60e1;
        src69 <= 16'hc27c;
        src70 <= 16'h8dbb;
        src71 <= 16'h31a;
        src72 <= 16'h85cd;
        src73 <= 16'hc7bc;
        src74 <= 16'hd228;
        src75 <= 16'hfdde;
        src76 <= 16'hac2d;
        src77 <= 16'h41c5;
        src78 <= 16'h8e89;
        src79 <= 16'hb20d;
        src80 <= 16'h1a1a;
        src81 <= 16'hbf1a;
        src82 <= 16'h216e;
        src83 <= 16'h2ed3;
        src84 <= 16'haeb9;
        src85 <= 16'h37ec;
        src86 <= 16'h713c;
        src87 <= 16'hada1;
        src88 <= 16'hbda5;
        src89 <= 16'h371e;
        src90 <= 16'ha1e7;
        src91 <= 16'h1387;
        src92 <= 16'h6224;
        src93 <= 16'haa1e;
        src94 <= 16'h4921;
        src95 <= 16'h6eb7;
        src96 <= 16'h3af3;
        src97 <= 16'hbec3;
        src98 <= 16'h8fa8;
        src99 <= 16'h5ef2;
        src100 <= 16'h9666;
        src101 <= 16'h65ac;
        src102 <= 16'h4310;
        src103 <= 16'h60e4;
        src104 <= 16'h4b1e;
        src105 <= 16'h4a99;
        src106 <= 16'h3c4b;
        src107 <= 16'hf477;
        src108 <= 16'hb770;
        src109 <= 16'he72a;
        src110 <= 16'hfc19;
        src111 <= 16'hd4af;
        src112 <= 16'hf04;
        src113 <= 16'hf243;
        src114 <= 16'h6250;
        src115 <= 16'h6509;
        src116 <= 16'hf01e;
        src117 <= 16'h9132;
        src118 <= 16'h816d;
        src119 <= 16'h809e;
        src120 <= 16'hb3d5;
        src121 <= 16'h17d9;
        src122 <= 16'haaa6;
        src123 <= 16'h1d6f;
        src124 <= 16'he1c9;
        src125 <= 16'h989f;
        src126 <= 16'ha041;
        src127 <= 16'h9744;
        exp <= 23'h4193d6;
        #1
        src0 <= 16'hda4a;
        src1 <= 16'h457a;
        src2 <= 16'h8bd3;
        src3 <= 16'haa4d;
        src4 <= 16'h3ea9;
        src5 <= 16'heb09;
        src6 <= 16'hfcdc;
        src7 <= 16'hc6fc;
        src8 <= 16'he6d8;
        src9 <= 16'haa57;
        src10 <= 16'he060;
        src11 <= 16'h8da3;
        src12 <= 16'hbd5c;
        src13 <= 16'hb89a;
        src14 <= 16'h7cb2;
        src15 <= 16'h7b06;
        src16 <= 16'h1860;
        src17 <= 16'hae10;
        src18 <= 16'hf71;
        src19 <= 16'h550d;
        src20 <= 16'h1d36;
        src21 <= 16'h6ebc;
        src22 <= 16'h8e73;
        src23 <= 16'h8e7e;
        src24 <= 16'hf320;
        src25 <= 16'ha2f2;
        src26 <= 16'h2519;
        src27 <= 16'h789c;
        src28 <= 16'haae;
        src29 <= 16'h1a72;
        src30 <= 16'h15d4;
        src31 <= 16'hf3ec;
        src32 <= 16'hdfed;
        src33 <= 16'hc660;
        src34 <= 16'hb255;
        src35 <= 16'h47ba;
        src36 <= 16'hce29;
        src37 <= 16'ha4e;
        src38 <= 16'hb6a6;
        src39 <= 16'hc692;
        src40 <= 16'hd714;
        src41 <= 16'h38f4;
        src42 <= 16'h8a10;
        src43 <= 16'h6c5c;
        src44 <= 16'ha012;
        src45 <= 16'h253c;
        src46 <= 16'hedd1;
        src47 <= 16'h607c;
        src48 <= 16'h5786;
        src49 <= 16'he1c6;
        src50 <= 16'hc826;
        src51 <= 16'hda26;
        src52 <= 16'h2e5b;
        src53 <= 16'he105;
        src54 <= 16'h9cfb;
        src55 <= 16'h4903;
        src56 <= 16'h67da;
        src57 <= 16'hca90;
        src58 <= 16'h9ddd;
        src59 <= 16'h4222;
        src60 <= 16'h420b;
        src61 <= 16'hf686;
        src62 <= 16'h9260;
        src63 <= 16'hbda0;
        src64 <= 16'h8e66;
        src65 <= 16'h9ed0;
        src66 <= 16'h66e4;
        src67 <= 16'hd40b;
        src68 <= 16'h84c8;
        src69 <= 16'h574c;
        src70 <= 16'h3b6c;
        src71 <= 16'hb5e8;
        src72 <= 16'he25;
        src73 <= 16'h2bf9;
        src74 <= 16'hbde1;
        src75 <= 16'hc67d;
        src76 <= 16'he688;
        src77 <= 16'h91b0;
        src78 <= 16'h2a9a;
        src79 <= 16'hcf0b;
        src80 <= 16'hf2aa;
        src81 <= 16'he30b;
        src82 <= 16'ha44a;
        src83 <= 16'hf217;
        src84 <= 16'hdf09;
        src85 <= 16'hd7d7;
        src86 <= 16'h9efd;
        src87 <= 16'h2810;
        src88 <= 16'h13ce;
        src89 <= 16'h2870;
        src90 <= 16'hed93;
        src91 <= 16'h8f0c;
        src92 <= 16'h1440;
        src93 <= 16'hbcb9;
        src94 <= 16'h1604;
        src95 <= 16'hccca;
        src96 <= 16'h476;
        src97 <= 16'hb8ff;
        src98 <= 16'h5155;
        src99 <= 16'h613a;
        src100 <= 16'hb840;
        src101 <= 16'h4fce;
        src102 <= 16'h1f5f;
        src103 <= 16'hb8d9;
        src104 <= 16'hbf26;
        src105 <= 16'hcd5;
        src106 <= 16'h4bee;
        src107 <= 16'had10;
        src108 <= 16'hab3c;
        src109 <= 16'h5614;
        src110 <= 16'h25ca;
        src111 <= 16'hdd43;
        src112 <= 16'h2d2c;
        src113 <= 16'h1618;
        src114 <= 16'h59a9;
        src115 <= 16'h17ba;
        src116 <= 16'h6921;
        src117 <= 16'h9d38;
        src118 <= 16'h7f8c;
        src119 <= 16'hfb42;
        src120 <= 16'h208e;
        src121 <= 16'h5384;
        src122 <= 16'h94c9;
        src123 <= 16'hecf9;
        src124 <= 16'hcfe8;
        src125 <= 16'h90f2;
        src126 <= 16'h82a5;
        src127 <= 16'h4347;
        exp <= 23'h438b65;
        #1
        src0 <= 16'h2a7f;
        src1 <= 16'hedf4;
        src2 <= 16'h7e1e;
        src3 <= 16'h7075;
        src4 <= 16'hec2e;
        src5 <= 16'h693e;
        src6 <= 16'hda62;
        src7 <= 16'hf7d5;
        src8 <= 16'hfada;
        src9 <= 16'h723e;
        src10 <= 16'h2c4c;
        src11 <= 16'h477c;
        src12 <= 16'h23ef;
        src13 <= 16'h2fe1;
        src14 <= 16'h2b43;
        src15 <= 16'hafaa;
        src16 <= 16'h7e31;
        src17 <= 16'ha2b2;
        src18 <= 16'haba3;
        src19 <= 16'hcf97;
        src20 <= 16'h36b1;
        src21 <= 16'hff1f;
        src22 <= 16'h6f5c;
        src23 <= 16'h482e;
        src24 <= 16'ha7ba;
        src25 <= 16'hc303;
        src26 <= 16'h865f;
        src27 <= 16'h5671;
        src28 <= 16'h4c92;
        src29 <= 16'hea3a;
        src30 <= 16'he278;
        src31 <= 16'hce28;
        src32 <= 16'h2159;
        src33 <= 16'hdc5c;
        src34 <= 16'h391b;
        src35 <= 16'hb151;
        src36 <= 16'h1d6b;
        src37 <= 16'h9512;
        src38 <= 16'hcc1b;
        src39 <= 16'h7321;
        src40 <= 16'h1685;
        src41 <= 16'h30b9;
        src42 <= 16'h99a3;
        src43 <= 16'h692f;
        src44 <= 16'hbf95;
        src45 <= 16'h19cd;
        src46 <= 16'h717a;
        src47 <= 16'h8751;
        src48 <= 16'hb304;
        src49 <= 16'h2fd2;
        src50 <= 16'h4277;
        src51 <= 16'hc1b0;
        src52 <= 16'hab5c;
        src53 <= 16'h1cbb;
        src54 <= 16'hc2a9;
        src55 <= 16'hfb9b;
        src56 <= 16'h5db6;
        src57 <= 16'h1fbb;
        src58 <= 16'hc4f2;
        src59 <= 16'hed86;
        src60 <= 16'hce7d;
        src61 <= 16'h762e;
        src62 <= 16'h54c;
        src63 <= 16'h918f;
        src64 <= 16'hb70a;
        src65 <= 16'h781d;
        src66 <= 16'hfdd1;
        src67 <= 16'h2212;
        src68 <= 16'h2452;
        src69 <= 16'h31ab;
        src70 <= 16'h6412;
        src71 <= 16'h1f16;
        src72 <= 16'h28f8;
        src73 <= 16'ha02d;
        src74 <= 16'h80cf;
        src75 <= 16'hc224;
        src76 <= 16'h8c4a;
        src77 <= 16'he40a;
        src78 <= 16'h3e90;
        src79 <= 16'hfe29;
        src80 <= 16'hae6b;
        src81 <= 16'h3dcf;
        src82 <= 16'haf08;
        src83 <= 16'hd137;
        src84 <= 16'h34b5;
        src85 <= 16'h7e71;
        src86 <= 16'hba5f;
        src87 <= 16'hdb90;
        src88 <= 16'h3587;
        src89 <= 16'hb5b2;
        src90 <= 16'hfe65;
        src91 <= 16'h4bdb;
        src92 <= 16'hdf0a;
        src93 <= 16'h1fd2;
        src94 <= 16'hc094;
        src95 <= 16'h2ed6;
        src96 <= 16'haaa1;
        src97 <= 16'h39e6;
        src98 <= 16'h79c8;
        src99 <= 16'h9b84;
        src100 <= 16'h30a4;
        src101 <= 16'he537;
        src102 <= 16'hf14a;
        src103 <= 16'h4563;
        src104 <= 16'he80b;
        src105 <= 16'h6d06;
        src106 <= 16'he99e;
        src107 <= 16'hd650;
        src108 <= 16'h632a;
        src109 <= 16'h5a28;
        src110 <= 16'he12c;
        src111 <= 16'h6285;
        src112 <= 16'h4f25;
        src113 <= 16'hb35b;
        src114 <= 16'hfa38;
        src115 <= 16'hbe1f;
        src116 <= 16'h3270;
        src117 <= 16'h41b2;
        src118 <= 16'h7821;
        src119 <= 16'h629d;
        src120 <= 16'h30de;
        src121 <= 16'h9390;
        src122 <= 16'h7a4;
        src123 <= 16'hf80;
        src124 <= 16'hb93e;
        src125 <= 16'hf503;
        src126 <= 16'h8022;
        src127 <= 16'ha64e;
        exp <= 23'h43368c;
        #1
        src0 <= 16'h4b77;
        src1 <= 16'hb09a;
        src2 <= 16'he88e;
        src3 <= 16'hb47;
        src4 <= 16'hf449;
        src5 <= 16'h3f82;
        src6 <= 16'h4124;
        src7 <= 16'hdc0c;
        src8 <= 16'h74c;
        src9 <= 16'h17f;
        src10 <= 16'hf3d2;
        src11 <= 16'h96dc;
        src12 <= 16'h769b;
        src13 <= 16'h8fa0;
        src14 <= 16'he46b;
        src15 <= 16'h40b8;
        src16 <= 16'h4f9;
        src17 <= 16'hcdff;
        src18 <= 16'hb10e;
        src19 <= 16'ha004;
        src20 <= 16'hf897;
        src21 <= 16'h6494;
        src22 <= 16'h41b1;
        src23 <= 16'h4c42;
        src24 <= 16'h28c4;
        src25 <= 16'h11bb;
        src26 <= 16'hc6fa;
        src27 <= 16'hfb29;
        src28 <= 16'h770b;
        src29 <= 16'h78;
        src30 <= 16'hc586;
        src31 <= 16'h9f60;
        src32 <= 16'h3a9b;
        src33 <= 16'h58e;
        src34 <= 16'h676c;
        src35 <= 16'h94f7;
        src36 <= 16'h4fc;
        src37 <= 16'hab1a;
        src38 <= 16'haff9;
        src39 <= 16'h1f62;
        src40 <= 16'h1343;
        src41 <= 16'hb621;
        src42 <= 16'ha091;
        src43 <= 16'h1eea;
        src44 <= 16'hd21;
        src45 <= 16'h15d6;
        src46 <= 16'h93be;
        src47 <= 16'h3e8b;
        src48 <= 16'h5739;
        src49 <= 16'hcc2f;
        src50 <= 16'h4ff6;
        src51 <= 16'h8eeb;
        src52 <= 16'hbc6f;
        src53 <= 16'h830a;
        src54 <= 16'he628;
        src55 <= 16'h22f9;
        src56 <= 16'hfc47;
        src57 <= 16'h6ae6;
        src58 <= 16'hbe97;
        src59 <= 16'he59d;
        src60 <= 16'h7f1c;
        src61 <= 16'h1587;
        src62 <= 16'h6c7d;
        src63 <= 16'h8f34;
        src64 <= 16'h4a31;
        src65 <= 16'hf71f;
        src66 <= 16'h314f;
        src67 <= 16'h9035;
        src68 <= 16'hbb4a;
        src69 <= 16'hb35e;
        src70 <= 16'h504d;
        src71 <= 16'h1be6;
        src72 <= 16'h4eb2;
        src73 <= 16'h6235;
        src74 <= 16'h217c;
        src75 <= 16'heed7;
        src76 <= 16'hfe2d;
        src77 <= 16'h58b1;
        src78 <= 16'hff6;
        src79 <= 16'h4671;
        src80 <= 16'h54a1;
        src81 <= 16'h3946;
        src82 <= 16'h649e;
        src83 <= 16'h6587;
        src84 <= 16'hdf4a;
        src85 <= 16'h518a;
        src86 <= 16'hb237;
        src87 <= 16'he724;
        src88 <= 16'hd1a4;
        src89 <= 16'ha60e;
        src90 <= 16'h8c8f;
        src91 <= 16'h706b;
        src92 <= 16'hd44a;
        src93 <= 16'hdfc8;
        src94 <= 16'h680b;
        src95 <= 16'h3528;
        src96 <= 16'hb74;
        src97 <= 16'h9f6c;
        src98 <= 16'h8ad0;
        src99 <= 16'h842;
        src100 <= 16'h4316;
        src101 <= 16'h49c6;
        src102 <= 16'h4504;
        src103 <= 16'h2ba3;
        src104 <= 16'h3797;
        src105 <= 16'h9f95;
        src106 <= 16'h3be7;
        src107 <= 16'h80a2;
        src108 <= 16'h30bc;
        src109 <= 16'h4a47;
        src110 <= 16'h6112;
        src111 <= 16'hd429;
        src112 <= 16'hd4eb;
        src113 <= 16'he31e;
        src114 <= 16'h28b7;
        src115 <= 16'ha56a;
        src116 <= 16'h4e63;
        src117 <= 16'hec8e;
        src118 <= 16'h83db;
        src119 <= 16'hda05;
        src120 <= 16'h26b0;
        src121 <= 16'hde49;
        src122 <= 16'h3b7e;
        src123 <= 16'hca7b;
        src124 <= 16'h4c6;
        src125 <= 16'h779f;
        src126 <= 16'hdd94;
        src127 <= 16'h852f;
        exp <= 23'h3cc576;
        #1
        src0 <= 16'hdbe2;
        src1 <= 16'hc23a;
        src2 <= 16'h95be;
        src3 <= 16'h859f;
        src4 <= 16'hf417;
        src5 <= 16'h74a3;
        src6 <= 16'hf10a;
        src7 <= 16'h8e37;
        src8 <= 16'h25d1;
        src9 <= 16'hfba2;
        src10 <= 16'hb30;
        src11 <= 16'hca43;
        src12 <= 16'h4144;
        src13 <= 16'h2b59;
        src14 <= 16'h96ac;
        src15 <= 16'ha86d;
        src16 <= 16'h85ae;
        src17 <= 16'h9d74;
        src18 <= 16'hc752;
        src19 <= 16'h245;
        src20 <= 16'hf109;
        src21 <= 16'h65c8;
        src22 <= 16'hca55;
        src23 <= 16'h363d;
        src24 <= 16'h96f9;
        src25 <= 16'hadc8;
        src26 <= 16'h6248;
        src27 <= 16'h2074;
        src28 <= 16'h3ec4;
        src29 <= 16'h12a2;
        src30 <= 16'h50b7;
        src31 <= 16'hd10;
        src32 <= 16'h6c19;
        src33 <= 16'hc446;
        src34 <= 16'ha4fd;
        src35 <= 16'h392e;
        src36 <= 16'hde4;
        src37 <= 16'he67f;
        src38 <= 16'h202f;
        src39 <= 16'hcb26;
        src40 <= 16'haf21;
        src41 <= 16'hfc14;
        src42 <= 16'h7a5d;
        src43 <= 16'he12e;
        src44 <= 16'h231;
        src45 <= 16'h707d;
        src46 <= 16'h4b6f;
        src47 <= 16'hcd7a;
        src48 <= 16'hb8e1;
        src49 <= 16'h3bf9;
        src50 <= 16'hb182;
        src51 <= 16'h1e73;
        src52 <= 16'hba2b;
        src53 <= 16'h3390;
        src54 <= 16'h3912;
        src55 <= 16'hefed;
        src56 <= 16'h8aba;
        src57 <= 16'hd5d4;
        src58 <= 16'h8feb;
        src59 <= 16'hb9a3;
        src60 <= 16'he52a;
        src61 <= 16'hb2d4;
        src62 <= 16'hf3fd;
        src63 <= 16'h4a06;
        src64 <= 16'he98a;
        src65 <= 16'hb0ba;
        src66 <= 16'h5be2;
        src67 <= 16'h5848;
        src68 <= 16'h480d;
        src69 <= 16'h9ce1;
        src70 <= 16'h8955;
        src71 <= 16'h2d26;
        src72 <= 16'h6ae0;
        src73 <= 16'had04;
        src74 <= 16'h9cca;
        src75 <= 16'h686a;
        src76 <= 16'h4184;
        src77 <= 16'ha446;
        src78 <= 16'hdd3d;
        src79 <= 16'hbbfb;
        src80 <= 16'h1bb6;
        src81 <= 16'h38f8;
        src82 <= 16'hdf12;
        src83 <= 16'h495e;
        src84 <= 16'he378;
        src85 <= 16'ha08f;
        src86 <= 16'hcb97;
        src87 <= 16'h6ecb;
        src88 <= 16'h2ed6;
        src89 <= 16'h9e83;
        src90 <= 16'hb3a4;
        src91 <= 16'h9ee2;
        src92 <= 16'hca11;
        src93 <= 16'h304d;
        src94 <= 16'h706e;
        src95 <= 16'hbb65;
        src96 <= 16'h7dc9;
        src97 <= 16'hf447;
        src98 <= 16'h1b97;
        src99 <= 16'h2fcc;
        src100 <= 16'h9cb8;
        src101 <= 16'h8e48;
        src102 <= 16'h7274;
        src103 <= 16'h4a4e;
        src104 <= 16'h8e27;
        src105 <= 16'h6586;
        src106 <= 16'h1d94;
        src107 <= 16'h83d6;
        src108 <= 16'hcbcc;
        src109 <= 16'hdcea;
        src110 <= 16'hf6de;
        src111 <= 16'h481e;
        src112 <= 16'hd3ea;
        src113 <= 16'hd2cd;
        src114 <= 16'h8dc4;
        src115 <= 16'h5696;
        src116 <= 16'h43b7;
        src117 <= 16'h8a2b;
        src118 <= 16'h60f;
        src119 <= 16'hcb2f;
        src120 <= 16'h5f82;
        src121 <= 16'h4fc1;
        src122 <= 16'h9705;
        src123 <= 16'h57a3;
        src124 <= 16'h5ac7;
        src125 <= 16'h8d;
        src126 <= 16'hee47;
        src127 <= 16'h15fe;
        exp <= 23'h422c50;
        #1
        src0 <= 16'h3cb1;
        src1 <= 16'hd9dd;
        src2 <= 16'hbeec;
        src3 <= 16'h2362;
        src4 <= 16'h7efb;
        src5 <= 16'h47fe;
        src6 <= 16'h89bc;
        src7 <= 16'h5aad;
        src8 <= 16'hc9d7;
        src9 <= 16'h9713;
        src10 <= 16'h2459;
        src11 <= 16'haa57;
        src12 <= 16'h377d;
        src13 <= 16'h88df;
        src14 <= 16'hc49c;
        src15 <= 16'h94dd;
        src16 <= 16'hc39b;
        src17 <= 16'h2ef5;
        src18 <= 16'h984a;
        src19 <= 16'h1d27;
        src20 <= 16'hce2c;
        src21 <= 16'h9bd7;
        src22 <= 16'hcd00;
        src23 <= 16'hdb9f;
        src24 <= 16'h5726;
        src25 <= 16'h8822;
        src26 <= 16'h2341;
        src27 <= 16'h2223;
        src28 <= 16'h7b9c;
        src29 <= 16'h2380;
        src30 <= 16'hbf10;
        src31 <= 16'h800b;
        src32 <= 16'h37b0;
        src33 <= 16'hc1bb;
        src34 <= 16'hddb;
        src35 <= 16'h30fe;
        src36 <= 16'h8f56;
        src37 <= 16'h7fe7;
        src38 <= 16'hde3e;
        src39 <= 16'h633a;
        src40 <= 16'he8f5;
        src41 <= 16'hd5d5;
        src42 <= 16'h4558;
        src43 <= 16'h4c26;
        src44 <= 16'hbed3;
        src45 <= 16'h326c;
        src46 <= 16'hdebf;
        src47 <= 16'he6f;
        src48 <= 16'h77f0;
        src49 <= 16'hb551;
        src50 <= 16'h63cd;
        src51 <= 16'h5ca9;
        src52 <= 16'hf202;
        src53 <= 16'hc48f;
        src54 <= 16'h4b18;
        src55 <= 16'h28be;
        src56 <= 16'h1b05;
        src57 <= 16'h23c2;
        src58 <= 16'h1565;
        src59 <= 16'h7794;
        src60 <= 16'h5a95;
        src61 <= 16'h95fa;
        src62 <= 16'hb615;
        src63 <= 16'h87f5;
        src64 <= 16'h1f26;
        src65 <= 16'h29b1;
        src66 <= 16'hefa7;
        src67 <= 16'h4d4;
        src68 <= 16'h9134;
        src69 <= 16'hcff4;
        src70 <= 16'ha4cc;
        src71 <= 16'h42f;
        src72 <= 16'h97cc;
        src73 <= 16'he229;
        src74 <= 16'h771d;
        src75 <= 16'hc2c2;
        src76 <= 16'h35c0;
        src77 <= 16'h5332;
        src78 <= 16'h8f81;
        src79 <= 16'hdd7;
        src80 <= 16'ha241;
        src81 <= 16'h6a1f;
        src82 <= 16'h6163;
        src83 <= 16'h137a;
        src84 <= 16'h1867;
        src85 <= 16'h326d;
        src86 <= 16'hb49;
        src87 <= 16'ha189;
        src88 <= 16'h532a;
        src89 <= 16'hcf27;
        src90 <= 16'he0b;
        src91 <= 16'h677f;
        src92 <= 16'hbddb;
        src93 <= 16'h1f05;
        src94 <= 16'he20e;
        src95 <= 16'h494a;
        src96 <= 16'hd74;
        src97 <= 16'h886c;
        src98 <= 16'h6b85;
        src99 <= 16'h4c1d;
        src100 <= 16'h3df8;
        src101 <= 16'h3670;
        src102 <= 16'h7a18;
        src103 <= 16'h38a3;
        src104 <= 16'hd18;
        src105 <= 16'h1ea3;
        src106 <= 16'h63be;
        src107 <= 16'hcc68;
        src108 <= 16'h74c6;
        src109 <= 16'h19d8;
        src110 <= 16'h9237;
        src111 <= 16'h1f4a;
        src112 <= 16'h8c8;
        src113 <= 16'hb17b;
        src114 <= 16'h26c5;
        src115 <= 16'h8297;
        src116 <= 16'h481e;
        src117 <= 16'h3265;
        src118 <= 16'h17f1;
        src119 <= 16'h7b2a;
        src120 <= 16'h4eaa;
        src121 <= 16'h9d;
        src122 <= 16'h583d;
        src123 <= 16'hbb7a;
        src124 <= 16'h75ff;
        src125 <= 16'h266f;
        src126 <= 16'hdbf6;
        src127 <= 16'h1619;
        exp <= 23'h36233e;
        #1
        src0 <= 16'h8a81;
        src1 <= 16'ha1f;
        src2 <= 16'h645a;
        src3 <= 16'hd76d;
        src4 <= 16'h6d3c;
        src5 <= 16'he274;
        src6 <= 16'he13b;
        src7 <= 16'h33c1;
        src8 <= 16'h2e4f;
        src9 <= 16'h5767;
        src10 <= 16'ha112;
        src11 <= 16'hf7f0;
        src12 <= 16'hcb40;
        src13 <= 16'h3f9d;
        src14 <= 16'h1afe;
        src15 <= 16'hd5f0;
        src16 <= 16'ha456;
        src17 <= 16'hf027;
        src18 <= 16'hc1f5;
        src19 <= 16'h310b;
        src20 <= 16'hfe70;
        src21 <= 16'hca06;
        src22 <= 16'hb089;
        src23 <= 16'h9c31;
        src24 <= 16'h650f;
        src25 <= 16'h395b;
        src26 <= 16'h7a67;
        src27 <= 16'hb1ea;
        src28 <= 16'h65a1;
        src29 <= 16'h94c3;
        src30 <= 16'h835b;
        src31 <= 16'hb8d7;
        src32 <= 16'h43e6;
        src33 <= 16'h1007;
        src34 <= 16'hd5c2;
        src35 <= 16'hf940;
        src36 <= 16'hc896;
        src37 <= 16'h284b;
        src38 <= 16'h682e;
        src39 <= 16'h749a;
        src40 <= 16'h9d13;
        src41 <= 16'he726;
        src42 <= 16'h51;
        src43 <= 16'h531d;
        src44 <= 16'hbcd3;
        src45 <= 16'he63d;
        src46 <= 16'h15bb;
        src47 <= 16'h3b8f;
        src48 <= 16'hc260;
        src49 <= 16'h1645;
        src50 <= 16'h4bd4;
        src51 <= 16'haccd;
        src52 <= 16'h2bec;
        src53 <= 16'h579f;
        src54 <= 16'heec3;
        src55 <= 16'h513f;
        src56 <= 16'h680f;
        src57 <= 16'hd674;
        src58 <= 16'h19bb;
        src59 <= 16'h4243;
        src60 <= 16'ha056;
        src61 <= 16'hb107;
        src62 <= 16'hbd3e;
        src63 <= 16'h277b;
        src64 <= 16'hd467;
        src65 <= 16'h27f5;
        src66 <= 16'h2efd;
        src67 <= 16'h3168;
        src68 <= 16'ha2f1;
        src69 <= 16'hf414;
        src70 <= 16'hbbe0;
        src71 <= 16'he1dc;
        src72 <= 16'hbcef;
        src73 <= 16'h8c3;
        src74 <= 16'ha5f0;
        src75 <= 16'h3cf0;
        src76 <= 16'he9e9;
        src77 <= 16'h8133;
        src78 <= 16'hafa2;
        src79 <= 16'hdf51;
        src80 <= 16'hd587;
        src81 <= 16'h3f01;
        src82 <= 16'hfe4a;
        src83 <= 16'ha0f2;
        src84 <= 16'h994f;
        src85 <= 16'h5a62;
        src86 <= 16'hd8f8;
        src87 <= 16'h7457;
        src88 <= 16'hf2e6;
        src89 <= 16'h63b5;
        src90 <= 16'h7012;
        src91 <= 16'hb0c5;
        src92 <= 16'h9e6a;
        src93 <= 16'h4192;
        src94 <= 16'h3fa3;
        src95 <= 16'h2ce4;
        src96 <= 16'h30a;
        src97 <= 16'hf3ea;
        src98 <= 16'h80c1;
        src99 <= 16'hcff8;
        src100 <= 16'hf923;
        src101 <= 16'h2ddc;
        src102 <= 16'he001;
        src103 <= 16'h3e95;
        src104 <= 16'h2a90;
        src105 <= 16'hfdb3;
        src106 <= 16'hfb3d;
        src107 <= 16'h7d33;
        src108 <= 16'h2117;
        src109 <= 16'h7463;
        src110 <= 16'h79e0;
        src111 <= 16'h8226;
        src112 <= 16'h631c;
        src113 <= 16'h5c7f;
        src114 <= 16'h39ff;
        src115 <= 16'hfbeb;
        src116 <= 16'h77bd;
        src117 <= 16'h1a25;
        src118 <= 16'h9fe8;
        src119 <= 16'hf8cc;
        src120 <= 16'hb4c;
        src121 <= 16'h5666;
        src122 <= 16'h842e;
        src123 <= 16'ha1be;
        src124 <= 16'h5a7a;
        src125 <= 16'h5b26;
        src126 <= 16'hd704;
        src127 <= 16'hf41b;
        exp <= 23'h43e460;
        #1
        src0 <= 16'h36d0;
        src1 <= 16'hc45b;
        src2 <= 16'hf484;
        src3 <= 16'hc337;
        src4 <= 16'h9262;
        src5 <= 16'h7024;
        src6 <= 16'ha1e7;
        src7 <= 16'h6d60;
        src8 <= 16'h6b8;
        src9 <= 16'hc28a;
        src10 <= 16'h59a0;
        src11 <= 16'hce50;
        src12 <= 16'h3411;
        src13 <= 16'ha443;
        src14 <= 16'h37d3;
        src15 <= 16'hf23d;
        src16 <= 16'hba4d;
        src17 <= 16'h9990;
        src18 <= 16'hc9f9;
        src19 <= 16'hb15;
        src20 <= 16'h76b0;
        src21 <= 16'h2b45;
        src22 <= 16'h1e03;
        src23 <= 16'h9724;
        src24 <= 16'h1a84;
        src25 <= 16'h7e53;
        src26 <= 16'hae2b;
        src27 <= 16'hec4b;
        src28 <= 16'hfd15;
        src29 <= 16'hbb76;
        src30 <= 16'hc6d6;
        src31 <= 16'hd7ec;
        src32 <= 16'h3628;
        src33 <= 16'hb70d;
        src34 <= 16'hbc3c;
        src35 <= 16'hf79c;
        src36 <= 16'hb1f1;
        src37 <= 16'h9dd4;
        src38 <= 16'h8408;
        src39 <= 16'he89;
        src40 <= 16'hb441;
        src41 <= 16'h72ca;
        src42 <= 16'hd4b4;
        src43 <= 16'hbe1d;
        src44 <= 16'hbbd0;
        src45 <= 16'ha10;
        src46 <= 16'h1161;
        src47 <= 16'h12e0;
        src48 <= 16'h2fff;
        src49 <= 16'hb061;
        src50 <= 16'hffa8;
        src51 <= 16'h30a7;
        src52 <= 16'h462f;
        src53 <= 16'h5a0e;
        src54 <= 16'h5d1e;
        src55 <= 16'h461;
        src56 <= 16'h3dc5;
        src57 <= 16'hbed7;
        src58 <= 16'hbaab;
        src59 <= 16'h9972;
        src60 <= 16'h272;
        src61 <= 16'hb88e;
        src62 <= 16'h3eea;
        src63 <= 16'ha397;
        src64 <= 16'hcd33;
        src65 <= 16'h5fe6;
        src66 <= 16'hbd7e;
        src67 <= 16'h178f;
        src68 <= 16'ha59b;
        src69 <= 16'h8785;
        src70 <= 16'hc9e0;
        src71 <= 16'haa1;
        src72 <= 16'h1765;
        src73 <= 16'h1e3b;
        src74 <= 16'h5c5a;
        src75 <= 16'he09c;
        src76 <= 16'hefdd;
        src77 <= 16'hac4d;
        src78 <= 16'h370e;
        src79 <= 16'hc24b;
        src80 <= 16'h392e;
        src81 <= 16'h63f2;
        src82 <= 16'h90e3;
        src83 <= 16'h1bd1;
        src84 <= 16'h67a4;
        src85 <= 16'hcd54;
        src86 <= 16'he098;
        src87 <= 16'hb9b0;
        src88 <= 16'he5c0;
        src89 <= 16'h3427;
        src90 <= 16'h91ff;
        src91 <= 16'hb7aa;
        src92 <= 16'h5b0c;
        src93 <= 16'hb398;
        src94 <= 16'h68f2;
        src95 <= 16'h1a0e;
        src96 <= 16'h4033;
        src97 <= 16'hbfed;
        src98 <= 16'h1c3c;
        src99 <= 16'hbefa;
        src100 <= 16'h594;
        src101 <= 16'hf645;
        src102 <= 16'h441;
        src103 <= 16'h8196;
        src104 <= 16'h9ef9;
        src105 <= 16'h8e2d;
        src106 <= 16'h100d;
        src107 <= 16'h7538;
        src108 <= 16'h128d;
        src109 <= 16'hacdf;
        src110 <= 16'hffe8;
        src111 <= 16'h635e;
        src112 <= 16'hca5a;
        src113 <= 16'h9a43;
        src114 <= 16'hbe29;
        src115 <= 16'hd366;
        src116 <= 16'hdaef;
        src117 <= 16'hb9ab;
        src118 <= 16'hec7b;
        src119 <= 16'he3db;
        src120 <= 16'h73b8;
        src121 <= 16'h1062;
        src122 <= 16'h301;
        src123 <= 16'hcd53;
        src124 <= 16'h43e;
        src125 <= 16'h2258;
        src126 <= 16'h444f;
        src127 <= 16'h5d9f;
        exp <= 23'h40af48;
        #1
        src0 <= 16'h2d23;
        src1 <= 16'h8db7;
        src2 <= 16'h21a2;
        src3 <= 16'hd9db;
        src4 <= 16'h4f13;
        src5 <= 16'h6303;
        src6 <= 16'hd51a;
        src7 <= 16'hbfa0;
        src8 <= 16'h551c;
        src9 <= 16'h263a;
        src10 <= 16'he1f0;
        src11 <= 16'h187c;
        src12 <= 16'h4470;
        src13 <= 16'h40;
        src14 <= 16'h531e;
        src15 <= 16'h2777;
        src16 <= 16'h83ce;
        src17 <= 16'h11c6;
        src18 <= 16'h2862;
        src19 <= 16'h6799;
        src20 <= 16'h4d99;
        src21 <= 16'hfc0c;
        src22 <= 16'h3fbf;
        src23 <= 16'hbeb9;
        src24 <= 16'h88a1;
        src25 <= 16'h23ad;
        src26 <= 16'hf4c9;
        src27 <= 16'h135;
        src28 <= 16'hc6d4;
        src29 <= 16'hdd08;
        src30 <= 16'h8526;
        src31 <= 16'h4cd;
        src32 <= 16'h98e7;
        src33 <= 16'h8779;
        src34 <= 16'h7086;
        src35 <= 16'h91f9;
        src36 <= 16'h23cf;
        src37 <= 16'h18c0;
        src38 <= 16'h2e56;
        src39 <= 16'h5556;
        src40 <= 16'he90e;
        src41 <= 16'hd8a8;
        src42 <= 16'hd11a;
        src43 <= 16'h5464;
        src44 <= 16'h7db0;
        src45 <= 16'ha579;
        src46 <= 16'h24f2;
        src47 <= 16'hd138;
        src48 <= 16'hc1c6;
        src49 <= 16'hcf87;
        src50 <= 16'h57f;
        src51 <= 16'hbcfe;
        src52 <= 16'heb3b;
        src53 <= 16'hd362;
        src54 <= 16'h6705;
        src55 <= 16'hfbd;
        src56 <= 16'hf37b;
        src57 <= 16'hc4e8;
        src58 <= 16'h703f;
        src59 <= 16'hf489;
        src60 <= 16'hdb1e;
        src61 <= 16'h79c6;
        src62 <= 16'hdc26;
        src63 <= 16'hc431;
        src64 <= 16'h362d;
        src65 <= 16'h4893;
        src66 <= 16'h7983;
        src67 <= 16'hfe79;
        src68 <= 16'hd0e7;
        src69 <= 16'h72bc;
        src70 <= 16'h832e;
        src71 <= 16'hfcb3;
        src72 <= 16'hdb9a;
        src73 <= 16'h7f59;
        src74 <= 16'hc93e;
        src75 <= 16'h2353;
        src76 <= 16'hb903;
        src77 <= 16'hd340;
        src78 <= 16'hf481;
        src79 <= 16'h45d7;
        src80 <= 16'he791;
        src81 <= 16'ha4c7;
        src82 <= 16'hebe3;
        src83 <= 16'h8b9f;
        src84 <= 16'hd04c;
        src85 <= 16'h97f7;
        src86 <= 16'h8e54;
        src87 <= 16'h7c85;
        src88 <= 16'h21e0;
        src89 <= 16'h7dea;
        src90 <= 16'hb930;
        src91 <= 16'h89af;
        src92 <= 16'hd640;
        src93 <= 16'hc0b6;
        src94 <= 16'h2d68;
        src95 <= 16'hf797;
        src96 <= 16'h21f0;
        src97 <= 16'he430;
        src98 <= 16'h5e1d;
        src99 <= 16'hb1c5;
        src100 <= 16'h6bd9;
        src101 <= 16'h913f;
        src102 <= 16'hb5b2;
        src103 <= 16'h80ff;
        src104 <= 16'hd13d;
        src105 <= 16'hd4e2;
        src106 <= 16'he625;
        src107 <= 16'hf501;
        src108 <= 16'hceaa;
        src109 <= 16'h56ee;
        src110 <= 16'h2ceb;
        src111 <= 16'hbfe2;
        src112 <= 16'h53c7;
        src113 <= 16'h34e3;
        src114 <= 16'he75f;
        src115 <= 16'h5774;
        src116 <= 16'hb834;
        src117 <= 16'h16df;
        src118 <= 16'hbc8a;
        src119 <= 16'hb3b4;
        src120 <= 16'hd545;
        src121 <= 16'h6607;
        src122 <= 16'h76dc;
        src123 <= 16'h79a1;
        src124 <= 16'ha4f3;
        src125 <= 16'h5d14;
        src126 <= 16'h7a18;
        src127 <= 16'hf9bc;
        exp <= 23'h4652ff;
        #1
        src0 <= 16'h46f2;
        src1 <= 16'h69d5;
        src2 <= 16'heae;
        src3 <= 16'hbda8;
        src4 <= 16'h1e72;
        src5 <= 16'hc942;
        src6 <= 16'h546e;
        src7 <= 16'h672;
        src8 <= 16'ha23f;
        src9 <= 16'ha3b;
        src10 <= 16'ha167;
        src11 <= 16'hfe6e;
        src12 <= 16'h48d2;
        src13 <= 16'hb5e9;
        src14 <= 16'hd8b0;
        src15 <= 16'he927;
        src16 <= 16'h6209;
        src17 <= 16'hd2bc;
        src18 <= 16'h4b4c;
        src19 <= 16'hff97;
        src20 <= 16'haed4;
        src21 <= 16'h885f;
        src22 <= 16'h492a;
        src23 <= 16'hc1e8;
        src24 <= 16'hd898;
        src25 <= 16'hd32f;
        src26 <= 16'h2630;
        src27 <= 16'heda4;
        src28 <= 16'hbb9c;
        src29 <= 16'h4e69;
        src30 <= 16'haea2;
        src31 <= 16'h25e6;
        src32 <= 16'h34f1;
        src33 <= 16'he7dc;
        src34 <= 16'hd19e;
        src35 <= 16'ha264;
        src36 <= 16'h52ec;
        src37 <= 16'ha887;
        src38 <= 16'hced1;
        src39 <= 16'hce91;
        src40 <= 16'hf3f0;
        src41 <= 16'h8244;
        src42 <= 16'hc9e8;
        src43 <= 16'hd930;
        src44 <= 16'hd5b0;
        src45 <= 16'hb4e9;
        src46 <= 16'h97bb;
        src47 <= 16'h8208;
        src48 <= 16'h7b53;
        src49 <= 16'h60e5;
        src50 <= 16'h1c02;
        src51 <= 16'hfe42;
        src52 <= 16'h407e;
        src53 <= 16'h1c17;
        src54 <= 16'h3e59;
        src55 <= 16'h85f9;
        src56 <= 16'hdbd8;
        src57 <= 16'h40b3;
        src58 <= 16'h723d;
        src59 <= 16'h3dee;
        src60 <= 16'h31e8;
        src61 <= 16'he58;
        src62 <= 16'h9086;
        src63 <= 16'h9ee;
        src64 <= 16'hcc74;
        src65 <= 16'h6d45;
        src66 <= 16'hd572;
        src67 <= 16'h37;
        src68 <= 16'h506a;
        src69 <= 16'hb35b;
        src70 <= 16'h6773;
        src71 <= 16'h7868;
        src72 <= 16'hfac7;
        src73 <= 16'hca8f;
        src74 <= 16'h84d9;
        src75 <= 16'h64cc;
        src76 <= 16'h45c8;
        src77 <= 16'h64c3;
        src78 <= 16'ha82b;
        src79 <= 16'h7b72;
        src80 <= 16'h6e08;
        src81 <= 16'h1087;
        src82 <= 16'hf37e;
        src83 <= 16'h9675;
        src84 <= 16'h7fef;
        src85 <= 16'h4100;
        src86 <= 16'hc22d;
        src87 <= 16'h605;
        src88 <= 16'hd762;
        src89 <= 16'h8f8f;
        src90 <= 16'h7d65;
        src91 <= 16'hb69b;
        src92 <= 16'h6d27;
        src93 <= 16'h640c;
        src94 <= 16'h56c0;
        src95 <= 16'h3b9d;
        src96 <= 16'h5be;
        src97 <= 16'h987a;
        src98 <= 16'hb252;
        src99 <= 16'hce7b;
        src100 <= 16'h1142;
        src101 <= 16'hed60;
        src102 <= 16'h7097;
        src103 <= 16'h95a;
        src104 <= 16'h86f1;
        src105 <= 16'h1306;
        src106 <= 16'h4543;
        src107 <= 16'hbef4;
        src108 <= 16'h3925;
        src109 <= 16'hf386;
        src110 <= 16'hb77d;
        src111 <= 16'hb92b;
        src112 <= 16'h174f;
        src113 <= 16'he926;
        src114 <= 16'h81ac;
        src115 <= 16'h7b8d;
        src116 <= 16'hb669;
        src117 <= 16'heceb;
        src118 <= 16'h6c24;
        src119 <= 16'hb448;
        src120 <= 16'h9e6e;
        src121 <= 16'hb585;
        src122 <= 16'hc432;
        src123 <= 16'h27d7;
        src124 <= 16'h3e49;
        src125 <= 16'hfc65;
        src126 <= 16'hb4bb;
        src127 <= 16'h5edb;
        exp <= 23'h42f5d0;
        #1
        src0 <= 16'hb364;
        src1 <= 16'hb141;
        src2 <= 16'hecf4;
        src3 <= 16'h3679;
        src4 <= 16'h8aeb;
        src5 <= 16'hd3da;
        src6 <= 16'h6cfb;
        src7 <= 16'h7844;
        src8 <= 16'h4a6c;
        src9 <= 16'haade;
        src10 <= 16'hdec3;
        src11 <= 16'h92ee;
        src12 <= 16'h3c43;
        src13 <= 16'ha1c5;
        src14 <= 16'hb164;
        src15 <= 16'h48af;
        src16 <= 16'h38db;
        src17 <= 16'h8472;
        src18 <= 16'h7742;
        src19 <= 16'ha927;
        src20 <= 16'habd8;
        src21 <= 16'h88ee;
        src22 <= 16'h7c76;
        src23 <= 16'h7ca2;
        src24 <= 16'h4d29;
        src25 <= 16'had75;
        src26 <= 16'hf15a;
        src27 <= 16'hc351;
        src28 <= 16'he254;
        src29 <= 16'h7472;
        src30 <= 16'h5bcd;
        src31 <= 16'hbc14;
        src32 <= 16'h5a14;
        src33 <= 16'hbccb;
        src34 <= 16'h4c16;
        src35 <= 16'hc04d;
        src36 <= 16'h4d5a;
        src37 <= 16'h93b6;
        src38 <= 16'hc33f;
        src39 <= 16'h7c66;
        src40 <= 16'hc7e5;
        src41 <= 16'h8bae;
        src42 <= 16'h218a;
        src43 <= 16'hb;
        src44 <= 16'h2c12;
        src45 <= 16'h7d2a;
        src46 <= 16'h4094;
        src47 <= 16'h397b;
        src48 <= 16'h724f;
        src49 <= 16'h34dc;
        src50 <= 16'h3585;
        src51 <= 16'h3cb3;
        src52 <= 16'h4dc3;
        src53 <= 16'hc29b;
        src54 <= 16'h2b9c;
        src55 <= 16'hbfe8;
        src56 <= 16'h4498;
        src57 <= 16'h1462;
        src58 <= 16'h4534;
        src59 <= 16'h9dad;
        src60 <= 16'h2a12;
        src61 <= 16'he44e;
        src62 <= 16'h425c;
        src63 <= 16'h68be;
        src64 <= 16'h8802;
        src65 <= 16'h2a97;
        src66 <= 16'hdca2;
        src67 <= 16'hab2a;
        src68 <= 16'h9611;
        src69 <= 16'h62ac;
        src70 <= 16'h37da;
        src71 <= 16'h72a0;
        src72 <= 16'hf73e;
        src73 <= 16'hfdce;
        src74 <= 16'h14c9;
        src75 <= 16'h3c3e;
        src76 <= 16'hdc13;
        src77 <= 16'hd5a6;
        src78 <= 16'h8dea;
        src79 <= 16'ha991;
        src80 <= 16'h3811;
        src81 <= 16'h4a6;
        src82 <= 16'hff68;
        src83 <= 16'h8149;
        src84 <= 16'h5693;
        src85 <= 16'h7b56;
        src86 <= 16'hf272;
        src87 <= 16'h370d;
        src88 <= 16'hf27a;
        src89 <= 16'ha12e;
        src90 <= 16'hd240;
        src91 <= 16'h3b9a;
        src92 <= 16'h5da6;
        src93 <= 16'h9e00;
        src94 <= 16'h9016;
        src95 <= 16'hcdd0;
        src96 <= 16'hf1ae;
        src97 <= 16'h4aa;
        src98 <= 16'h9771;
        src99 <= 16'h33f6;
        src100 <= 16'h6fc0;
        src101 <= 16'h1d85;
        src102 <= 16'hf215;
        src103 <= 16'h3401;
        src104 <= 16'hd046;
        src105 <= 16'hce6c;
        src106 <= 16'h5e66;
        src107 <= 16'he89d;
        src108 <= 16'h28bc;
        src109 <= 16'h268b;
        src110 <= 16'ha0e0;
        src111 <= 16'hde18;
        src112 <= 16'h1837;
        src113 <= 16'hdd5;
        src114 <= 16'ha801;
        src115 <= 16'hfa6;
        src116 <= 16'h43bb;
        src117 <= 16'h10bc;
        src118 <= 16'he850;
        src119 <= 16'hdeac;
        src120 <= 16'ha135;
        src121 <= 16'h59c;
        src122 <= 16'h2290;
        src123 <= 16'h4cb8;
        src124 <= 16'h5dab;
        src125 <= 16'h67c9;
        src126 <= 16'hf31d;
        src127 <= 16'h9977;
        exp <= 23'h3f66ca;
        #1
        src0 <= 16'h63d1;
        src1 <= 16'h6e63;
        src2 <= 16'h6101;
        src3 <= 16'h1218;
        src4 <= 16'h9e97;
        src5 <= 16'h4657;
        src6 <= 16'h5ae3;
        src7 <= 16'h889b;
        src8 <= 16'h7c37;
        src9 <= 16'hb131;
        src10 <= 16'h78ca;
        src11 <= 16'h62dc;
        src12 <= 16'h5e92;
        src13 <= 16'h2288;
        src14 <= 16'h7deb;
        src15 <= 16'he20a;
        src16 <= 16'hdfd7;
        src17 <= 16'h1c95;
        src18 <= 16'h3cdb;
        src19 <= 16'he96;
        src20 <= 16'h5f4e;
        src21 <= 16'h2a78;
        src22 <= 16'h3a95;
        src23 <= 16'ha78b;
        src24 <= 16'hb335;
        src25 <= 16'h3b1;
        src26 <= 16'h81f5;
        src27 <= 16'h288a;
        src28 <= 16'h3265;
        src29 <= 16'ha469;
        src30 <= 16'hf70b;
        src31 <= 16'hbafc;
        src32 <= 16'h78b8;
        src33 <= 16'h1806;
        src34 <= 16'he8d7;
        src35 <= 16'h37ec;
        src36 <= 16'hc5b;
        src37 <= 16'h35ef;
        src38 <= 16'h2b38;
        src39 <= 16'h8af5;
        src40 <= 16'h5805;
        src41 <= 16'h2944;
        src42 <= 16'h757c;
        src43 <= 16'h31e7;
        src44 <= 16'h7354;
        src45 <= 16'hedb5;
        src46 <= 16'hffd7;
        src47 <= 16'hd49a;
        src48 <= 16'h6ac2;
        src49 <= 16'he61d;
        src50 <= 16'h750b;
        src51 <= 16'hfcab;
        src52 <= 16'h582f;
        src53 <= 16'h7112;
        src54 <= 16'h5505;
        src55 <= 16'hbcf;
        src56 <= 16'he91f;
        src57 <= 16'h4bfa;
        src58 <= 16'h38c7;
        src59 <= 16'hc9d5;
        src60 <= 16'ha6fa;
        src61 <= 16'ha74c;
        src62 <= 16'h9c24;
        src63 <= 16'hce3d;
        src64 <= 16'h9bb2;
        src65 <= 16'h3f28;
        src66 <= 16'h9e1b;
        src67 <= 16'h3b7b;
        src68 <= 16'hce87;
        src69 <= 16'ha19;
        src70 <= 16'hf8d5;
        src71 <= 16'hfbde;
        src72 <= 16'hfbf4;
        src73 <= 16'hd986;
        src74 <= 16'h52de;
        src75 <= 16'hd79d;
        src76 <= 16'he841;
        src77 <= 16'h3625;
        src78 <= 16'h5596;
        src79 <= 16'ha429;
        src80 <= 16'h2be;
        src81 <= 16'h31ef;
        src82 <= 16'h7b4e;
        src83 <= 16'h3358;
        src84 <= 16'h72d6;
        src85 <= 16'h49de;
        src86 <= 16'heccb;
        src87 <= 16'h4219;
        src88 <= 16'hcf61;
        src89 <= 16'he21b;
        src90 <= 16'h64db;
        src91 <= 16'h18d4;
        src92 <= 16'h1f3e;
        src93 <= 16'h4335;
        src94 <= 16'h15b7;
        src95 <= 16'h41b;
        src96 <= 16'h10e6;
        src97 <= 16'hf327;
        src98 <= 16'h1e3f;
        src99 <= 16'h5b2a;
        src100 <= 16'h5d14;
        src101 <= 16'hbc7e;
        src102 <= 16'h27;
        src103 <= 16'hd678;
        src104 <= 16'hf470;
        src105 <= 16'h50c2;
        src106 <= 16'h498a;
        src107 <= 16'h1788;
        src108 <= 16'ha2c4;
        src109 <= 16'hb6bd;
        src110 <= 16'h2159;
        src111 <= 16'h43d6;
        src112 <= 16'hfdc;
        src113 <= 16'h3770;
        src114 <= 16'h71b6;
        src115 <= 16'he441;
        src116 <= 16'hf9d1;
        src117 <= 16'h3509;
        src118 <= 16'h6cdc;
        src119 <= 16'he686;
        src120 <= 16'h768c;
        src121 <= 16'hdc5b;
        src122 <= 16'hf67c;
        src123 <= 16'h19d6;
        src124 <= 16'hbfda;
        src125 <= 16'h226c;
        src126 <= 16'h56f1;
        src127 <= 16'h565c;
        exp <= 23'h3b7415;
        #1
        src0 <= 16'hc63a;
        src1 <= 16'h3381;
        src2 <= 16'hdf22;
        src3 <= 16'ha542;
        src4 <= 16'h85e2;
        src5 <= 16'h7a8f;
        src6 <= 16'hb87f;
        src7 <= 16'hf911;
        src8 <= 16'h6bb8;
        src9 <= 16'h46d1;
        src10 <= 16'h3d1b;
        src11 <= 16'h7fbc;
        src12 <= 16'h856c;
        src13 <= 16'h77f9;
        src14 <= 16'h3bca;
        src15 <= 16'hb4ce;
        src16 <= 16'h4b76;
        src17 <= 16'h65f3;
        src18 <= 16'h4c65;
        src19 <= 16'h94c5;
        src20 <= 16'hb2a8;
        src21 <= 16'hede4;
        src22 <= 16'h6d93;
        src23 <= 16'hb62b;
        src24 <= 16'h9add;
        src25 <= 16'h5673;
        src26 <= 16'haec6;
        src27 <= 16'he4d9;
        src28 <= 16'h4bd4;
        src29 <= 16'hcf9c;
        src30 <= 16'h2f2b;
        src31 <= 16'h70fd;
        src32 <= 16'h6a4;
        src33 <= 16'haf8;
        src34 <= 16'hc038;
        src35 <= 16'hc8e7;
        src36 <= 16'h3af7;
        src37 <= 16'hf476;
        src38 <= 16'h77a4;
        src39 <= 16'hd3d4;
        src40 <= 16'h979;
        src41 <= 16'h820;
        src42 <= 16'ha8eb;
        src43 <= 16'hbb86;
        src44 <= 16'hcb54;
        src45 <= 16'hea2d;
        src46 <= 16'h849c;
        src47 <= 16'hebd;
        src48 <= 16'hed5e;
        src49 <= 16'he176;
        src50 <= 16'h5474;
        src51 <= 16'he955;
        src52 <= 16'h1387;
        src53 <= 16'h47bc;
        src54 <= 16'h8c34;
        src55 <= 16'h32d8;
        src56 <= 16'hd0dc;
        src57 <= 16'hba36;
        src58 <= 16'h20fe;
        src59 <= 16'hc273;
        src60 <= 16'h8605;
        src61 <= 16'h71de;
        src62 <= 16'hfc52;
        src63 <= 16'h48cc;
        src64 <= 16'hd22e;
        src65 <= 16'hc307;
        src66 <= 16'hb685;
        src67 <= 16'h66f5;
        src68 <= 16'h2228;
        src69 <= 16'h657d;
        src70 <= 16'hfc56;
        src71 <= 16'h6601;
        src72 <= 16'h2e56;
        src73 <= 16'hf75e;
        src74 <= 16'h7f64;
        src75 <= 16'h9bae;
        src76 <= 16'h2843;
        src77 <= 16'h2ae9;
        src78 <= 16'hf676;
        src79 <= 16'ha363;
        src80 <= 16'ha9fe;
        src81 <= 16'h575;
        src82 <= 16'hd652;
        src83 <= 16'h50e8;
        src84 <= 16'hc347;
        src85 <= 16'hfa20;
        src86 <= 16'h9ef8;
        src87 <= 16'h4068;
        src88 <= 16'haa56;
        src89 <= 16'hef4d;
        src90 <= 16'h7396;
        src91 <= 16'hd6f6;
        src92 <= 16'h8d54;
        src93 <= 16'h6670;
        src94 <= 16'h83f6;
        src95 <= 16'hdfd6;
        src96 <= 16'h37f7;
        src97 <= 16'he529;
        src98 <= 16'h4708;
        src99 <= 16'h81f0;
        src100 <= 16'h99aa;
        src101 <= 16'hd926;
        src102 <= 16'h5228;
        src103 <= 16'h6f03;
        src104 <= 16'h286e;
        src105 <= 16'h7467;
        src106 <= 16'hc64e;
        src107 <= 16'hdf57;
        src108 <= 16'h3b01;
        src109 <= 16'h15f2;
        src110 <= 16'h2c3f;
        src111 <= 16'h1188;
        src112 <= 16'h203c;
        src113 <= 16'h64cf;
        src114 <= 16'h1a8c;
        src115 <= 16'hd974;
        src116 <= 16'h5180;
        src117 <= 16'hd025;
        src118 <= 16'h69b3;
        src119 <= 16'hf2dd;
        src120 <= 16'h1edc;
        src121 <= 16'hde9f;
        src122 <= 16'hb1f;
        src123 <= 16'hf5b9;
        src124 <= 16'he286;
        src125 <= 16'he27c;
        src126 <= 16'hac9;
        src127 <= 16'h3e35;
        exp <= 23'h433458;
        #1
        src0 <= 16'h965c;
        src1 <= 16'h4540;
        src2 <= 16'h7cfd;
        src3 <= 16'hd035;
        src4 <= 16'he30f;
        src5 <= 16'h79a5;
        src6 <= 16'h10b;
        src7 <= 16'heba0;
        src8 <= 16'hbfb;
        src9 <= 16'h79c2;
        src10 <= 16'h7201;
        src11 <= 16'hb4a6;
        src12 <= 16'hfa05;
        src13 <= 16'h78ae;
        src14 <= 16'h3e0b;
        src15 <= 16'h98;
        src16 <= 16'hb233;
        src17 <= 16'hf44a;
        src18 <= 16'h7dd9;
        src19 <= 16'h4026;
        src20 <= 16'h19b3;
        src21 <= 16'h84b3;
        src22 <= 16'h2655;
        src23 <= 16'h97a8;
        src24 <= 16'h3f4a;
        src25 <= 16'h6fcc;
        src26 <= 16'h5e8e;
        src27 <= 16'he50;
        src28 <= 16'hd6c3;
        src29 <= 16'hc61a;
        src30 <= 16'h26e6;
        src31 <= 16'h966e;
        src32 <= 16'h3bbb;
        src33 <= 16'h2f3;
        src34 <= 16'h59fd;
        src35 <= 16'h327b;
        src36 <= 16'h11c8;
        src37 <= 16'hae4b;
        src38 <= 16'hd70d;
        src39 <= 16'h6cff;
        src40 <= 16'h9aae;
        src41 <= 16'hcf4e;
        src42 <= 16'h576b;
        src43 <= 16'hd88e;
        src44 <= 16'hcb90;
        src45 <= 16'h509b;
        src46 <= 16'h4fa1;
        src47 <= 16'h5ab2;
        src48 <= 16'hc019;
        src49 <= 16'h1be6;
        src50 <= 16'h821a;
        src51 <= 16'h8628;
        src52 <= 16'h2732;
        src53 <= 16'h718c;
        src54 <= 16'he343;
        src55 <= 16'heaca;
        src56 <= 16'he206;
        src57 <= 16'hbfeb;
        src58 <= 16'hf776;
        src59 <= 16'h69fc;
        src60 <= 16'h1675;
        src61 <= 16'h7e5;
        src62 <= 16'ha096;
        src63 <= 16'hc223;
        src64 <= 16'h9ba0;
        src65 <= 16'h717;
        src66 <= 16'hec8d;
        src67 <= 16'hc01c;
        src68 <= 16'h90cd;
        src69 <= 16'hca1f;
        src70 <= 16'hf150;
        src71 <= 16'h320;
        src72 <= 16'hbc2d;
        src73 <= 16'haf37;
        src74 <= 16'h226;
        src75 <= 16'h2361;
        src76 <= 16'h2d92;
        src77 <= 16'ha040;
        src78 <= 16'ha97f;
        src79 <= 16'hc265;
        src80 <= 16'hcb1c;
        src81 <= 16'h72d3;
        src82 <= 16'h90ed;
        src83 <= 16'h8d2f;
        src84 <= 16'hff89;
        src85 <= 16'hbbbc;
        src86 <= 16'hd94;
        src87 <= 16'hb9a5;
        src88 <= 16'h768f;
        src89 <= 16'hdff4;
        src90 <= 16'hcbd5;
        src91 <= 16'h9ac5;
        src92 <= 16'hedae;
        src93 <= 16'ha2a9;
        src94 <= 16'h6cd0;
        src95 <= 16'h7cab;
        src96 <= 16'h1ee0;
        src97 <= 16'hccda;
        src98 <= 16'h5d54;
        src99 <= 16'h602b;
        src100 <= 16'hfc54;
        src101 <= 16'h67ea;
        src102 <= 16'hf6c5;
        src103 <= 16'ha7c0;
        src104 <= 16'hec60;
        src105 <= 16'h1f7e;
        src106 <= 16'h4f66;
        src107 <= 16'ha3cc;
        src108 <= 16'h841c;
        src109 <= 16'h9c39;
        src110 <= 16'h61cb;
        src111 <= 16'h4462;
        src112 <= 16'h5e6c;
        src113 <= 16'he217;
        src114 <= 16'h6a95;
        src115 <= 16'hb1c2;
        src116 <= 16'hd187;
        src117 <= 16'hf6e9;
        src118 <= 16'h27ab;
        src119 <= 16'h9749;
        src120 <= 16'hd00e;
        src121 <= 16'h497b;
        src122 <= 16'hb461;
        src123 <= 16'h2ba2;
        src124 <= 16'h9b78;
        src125 <= 16'he073;
        src126 <= 16'hfa6e;
        src127 <= 16'h6f1a;
        exp <= 23'h43b9c5;
        #1
        src0 <= 16'h840f;
        src1 <= 16'h12ff;
        src2 <= 16'h8513;
        src3 <= 16'h313d;
        src4 <= 16'h3096;
        src5 <= 16'h8a17;
        src6 <= 16'hdc43;
        src7 <= 16'hd47e;
        src8 <= 16'h2de;
        src9 <= 16'h43c1;
        src10 <= 16'hb526;
        src11 <= 16'hc26d;
        src12 <= 16'hba74;
        src13 <= 16'h6aa5;
        src14 <= 16'hf8a1;
        src15 <= 16'h4ed9;
        src16 <= 16'h606c;
        src17 <= 16'h30d2;
        src18 <= 16'h1e12;
        src19 <= 16'hff60;
        src20 <= 16'h107a;
        src21 <= 16'hb24d;
        src22 <= 16'h112e;
        src23 <= 16'h26d5;
        src24 <= 16'ha36f;
        src25 <= 16'h8ccb;
        src26 <= 16'h5565;
        src27 <= 16'heba;
        src28 <= 16'h36b4;
        src29 <= 16'ha993;
        src30 <= 16'h3b54;
        src31 <= 16'hdaa;
        src32 <= 16'h7e8a;
        src33 <= 16'h8406;
        src34 <= 16'h43d6;
        src35 <= 16'hd3c9;
        src36 <= 16'h67e6;
        src37 <= 16'h4176;
        src38 <= 16'ha7dc;
        src39 <= 16'hd92;
        src40 <= 16'hd310;
        src41 <= 16'h1a31;
        src42 <= 16'h66d5;
        src43 <= 16'hb2f5;
        src44 <= 16'ha12e;
        src45 <= 16'h5506;
        src46 <= 16'hd44e;
        src47 <= 16'h9995;
        src48 <= 16'h38ca;
        src49 <= 16'h9ece;
        src50 <= 16'h89f8;
        src51 <= 16'hb9d5;
        src52 <= 16'h1f01;
        src53 <= 16'h9bc8;
        src54 <= 16'hea91;
        src55 <= 16'h882c;
        src56 <= 16'h379e;
        src57 <= 16'h24c3;
        src58 <= 16'h9ad7;
        src59 <= 16'h9cfd;
        src60 <= 16'h48a9;
        src61 <= 16'hadcd;
        src62 <= 16'he94d;
        src63 <= 16'h5bec;
        src64 <= 16'h7916;
        src65 <= 16'h96ab;
        src66 <= 16'hac62;
        src67 <= 16'h8446;
        src68 <= 16'hbedc;
        src69 <= 16'h8f1b;
        src70 <= 16'h52e5;
        src71 <= 16'h3e29;
        src72 <= 16'hb4ac;
        src73 <= 16'hb6b0;
        src74 <= 16'hc0eb;
        src75 <= 16'h8a63;
        src76 <= 16'h5c1a;
        src77 <= 16'h6464;
        src78 <= 16'h93eb;
        src79 <= 16'hf5fc;
        src80 <= 16'hfa7d;
        src81 <= 16'ha94e;
        src82 <= 16'hb409;
        src83 <= 16'h5a38;
        src84 <= 16'h8a6f;
        src85 <= 16'h979b;
        src86 <= 16'hf6e0;
        src87 <= 16'h637;
        src88 <= 16'hfeb8;
        src89 <= 16'h8087;
        src90 <= 16'habaf;
        src91 <= 16'h3832;
        src92 <= 16'hec67;
        src93 <= 16'h396c;
        src94 <= 16'h401a;
        src95 <= 16'h7c01;
        src96 <= 16'hb55d;
        src97 <= 16'h2a1d;
        src98 <= 16'haddd;
        src99 <= 16'habf1;
        src100 <= 16'h69d;
        src101 <= 16'hf558;
        src102 <= 16'hd5f0;
        src103 <= 16'hdeb8;
        src104 <= 16'hbb55;
        src105 <= 16'h8844;
        src106 <= 16'h29d8;
        src107 <= 16'h5c2a;
        src108 <= 16'h9ac8;
        src109 <= 16'hc4cd;
        src110 <= 16'hd12e;
        src111 <= 16'h740d;
        src112 <= 16'h287e;
        src113 <= 16'h71c8;
        src114 <= 16'hcd18;
        src115 <= 16'h362e;
        src116 <= 16'he011;
        src117 <= 16'hd03e;
        src118 <= 16'h9efe;
        src119 <= 16'h3f1;
        src120 <= 16'h2819;
        src121 <= 16'h1723;
        src122 <= 16'h42fc;
        src123 <= 16'hf639;
        src124 <= 16'h71a0;
        src125 <= 16'h2918;
        src126 <= 16'hd530;
        src127 <= 16'h721f;
        exp <= 23'h4021dd;
        #1
        src0 <= 16'h8452;
        src1 <= 16'hc671;
        src2 <= 16'h1391;
        src3 <= 16'h3bb;
        src4 <= 16'h6fde;
        src5 <= 16'h7f04;
        src6 <= 16'h8fcf;
        src7 <= 16'h2b00;
        src8 <= 16'h920c;
        src9 <= 16'h6292;
        src10 <= 16'h10da;
        src11 <= 16'ha86f;
        src12 <= 16'he52e;
        src13 <= 16'h468f;
        src14 <= 16'h5770;
        src15 <= 16'hb6a9;
        src16 <= 16'ha4a5;
        src17 <= 16'h6ff9;
        src18 <= 16'h908b;
        src19 <= 16'h2067;
        src20 <= 16'h2776;
        src21 <= 16'haa4f;
        src22 <= 16'hba28;
        src23 <= 16'hf082;
        src24 <= 16'hc032;
        src25 <= 16'he2a6;
        src26 <= 16'h1a78;
        src27 <= 16'he511;
        src28 <= 16'ha3a3;
        src29 <= 16'h5601;
        src30 <= 16'hd1da;
        src31 <= 16'h9065;
        src32 <= 16'h7592;
        src33 <= 16'h9a00;
        src34 <= 16'h535;
        src35 <= 16'hffb;
        src36 <= 16'h343d;
        src37 <= 16'h2e12;
        src38 <= 16'ha43c;
        src39 <= 16'h1070;
        src40 <= 16'h47b4;
        src41 <= 16'h16be;
        src42 <= 16'h74c2;
        src43 <= 16'hff4b;
        src44 <= 16'hf3fb;
        src45 <= 16'hf871;
        src46 <= 16'h6086;
        src47 <= 16'hdb70;
        src48 <= 16'h434e;
        src49 <= 16'h350a;
        src50 <= 16'hba3;
        src51 <= 16'hdfe6;
        src52 <= 16'h17b4;
        src53 <= 16'hddd7;
        src54 <= 16'hc421;
        src55 <= 16'h897f;
        src56 <= 16'hb4a9;
        src57 <= 16'hfc88;
        src58 <= 16'h23c0;
        src59 <= 16'hef34;
        src60 <= 16'hcb60;
        src61 <= 16'h6874;
        src62 <= 16'h196e;
        src63 <= 16'h96d4;
        src64 <= 16'h5a50;
        src65 <= 16'h6645;
        src66 <= 16'hb3a1;
        src67 <= 16'h8059;
        src68 <= 16'h85ff;
        src69 <= 16'h80ea;
        src70 <= 16'h7bcf;
        src71 <= 16'h582b;
        src72 <= 16'he79a;
        src73 <= 16'heb81;
        src74 <= 16'h5574;
        src75 <= 16'h1ac3;
        src76 <= 16'hf7fc;
        src77 <= 16'ha114;
        src78 <= 16'hafa5;
        src79 <= 16'h1ed4;
        src80 <= 16'h2f9b;
        src81 <= 16'h4f44;
        src82 <= 16'h976;
        src83 <= 16'hf292;
        src84 <= 16'h239a;
        src85 <= 16'hee2;
        src86 <= 16'h86f5;
        src87 <= 16'h25aa;
        src88 <= 16'h5cb9;
        src89 <= 16'hda9a;
        src90 <= 16'h10f8;
        src91 <= 16'h5078;
        src92 <= 16'h74c0;
        src93 <= 16'h1eca;
        src94 <= 16'hade0;
        src95 <= 16'h9182;
        src96 <= 16'hca92;
        src97 <= 16'h1903;
        src98 <= 16'h7d61;
        src99 <= 16'h9026;
        src100 <= 16'h9e6d;
        src101 <= 16'hcc22;
        src102 <= 16'h959a;
        src103 <= 16'h69e7;
        src104 <= 16'h2484;
        src105 <= 16'he9bf;
        src106 <= 16'h2c3f;
        src107 <= 16'hdb60;
        src108 <= 16'h7812;
        src109 <= 16'ha42c;
        src110 <= 16'h9576;
        src111 <= 16'h13d0;
        src112 <= 16'h1e8b;
        src113 <= 16'h9dc2;
        src114 <= 16'hcfbc;
        src115 <= 16'h32a;
        src116 <= 16'h82b2;
        src117 <= 16'hda48;
        src118 <= 16'hf0b3;
        src119 <= 16'h321;
        src120 <= 16'hefb0;
        src121 <= 16'hc20f;
        src122 <= 16'h2d1c;
        src123 <= 16'h3af1;
        src124 <= 16'h85ee;
        src125 <= 16'h26a5;
        src126 <= 16'he19e;
        src127 <= 16'hfc5a;
        exp <= 23'h3eb48d;
        #1
        src0 <= 16'he380;
        src1 <= 16'hd15a;
        src2 <= 16'h91d1;
        src3 <= 16'ha79d;
        src4 <= 16'h7423;
        src5 <= 16'he3d1;
        src6 <= 16'hec86;
        src7 <= 16'h7917;
        src8 <= 16'h7cce;
        src9 <= 16'h61e;
        src10 <= 16'hbf2f;
        src11 <= 16'h1861;
        src12 <= 16'h11ac;
        src13 <= 16'hd4e5;
        src14 <= 16'h2484;
        src15 <= 16'hc1f1;
        src16 <= 16'hd7fa;
        src17 <= 16'h871c;
        src18 <= 16'h5962;
        src19 <= 16'hff3b;
        src20 <= 16'h8d57;
        src21 <= 16'h2182;
        src22 <= 16'he8f1;
        src23 <= 16'hbe00;
        src24 <= 16'h83d3;
        src25 <= 16'h7a0e;
        src26 <= 16'h295c;
        src27 <= 16'h94ab;
        src28 <= 16'he365;
        src29 <= 16'hb8ec;
        src30 <= 16'hc80d;
        src31 <= 16'hf149;
        src32 <= 16'hcc79;
        src33 <= 16'h6ae0;
        src34 <= 16'h8c86;
        src35 <= 16'h8cd8;
        src36 <= 16'h9771;
        src37 <= 16'h6f84;
        src38 <= 16'hdfc0;
        src39 <= 16'h7f78;
        src40 <= 16'hd49f;
        src41 <= 16'h7ce;
        src42 <= 16'he254;
        src43 <= 16'hcc9;
        src44 <= 16'h1166;
        src45 <= 16'h46c7;
        src46 <= 16'hc0f0;
        src47 <= 16'h4d8f;
        src48 <= 16'h7a89;
        src49 <= 16'h131c;
        src50 <= 16'hd1c;
        src51 <= 16'hf4a2;
        src52 <= 16'h3723;
        src53 <= 16'h78a7;
        src54 <= 16'h642;
        src55 <= 16'hcb80;
        src56 <= 16'h6cc1;
        src57 <= 16'hd232;
        src58 <= 16'h15b3;
        src59 <= 16'h64a7;
        src60 <= 16'h767b;
        src61 <= 16'h5724;
        src62 <= 16'h3d95;
        src63 <= 16'h7045;
        src64 <= 16'h135a;
        src65 <= 16'h48fc;
        src66 <= 16'hdb57;
        src67 <= 16'h5971;
        src68 <= 16'h680d;
        src69 <= 16'h1be4;
        src70 <= 16'hfc3f;
        src71 <= 16'h773d;
        src72 <= 16'h23d3;
        src73 <= 16'h5e69;
        src74 <= 16'h111;
        src75 <= 16'h8bec;
        src76 <= 16'hff7e;
        src77 <= 16'h3e8;
        src78 <= 16'h9acb;
        src79 <= 16'hce82;
        src80 <= 16'h62eb;
        src81 <= 16'h68c8;
        src82 <= 16'h7c43;
        src83 <= 16'h56a0;
        src84 <= 16'h1219;
        src85 <= 16'h5149;
        src86 <= 16'h144;
        src87 <= 16'h648c;
        src88 <= 16'h5787;
        src89 <= 16'h484b;
        src90 <= 16'hb228;
        src91 <= 16'he561;
        src92 <= 16'h773c;
        src93 <= 16'he78b;
        src94 <= 16'h4c26;
        src95 <= 16'h20e0;
        src96 <= 16'h595d;
        src97 <= 16'h9ab0;
        src98 <= 16'ha075;
        src99 <= 16'heca5;
        src100 <= 16'h895f;
        src101 <= 16'h3f56;
        src102 <= 16'h3de4;
        src103 <= 16'hf25c;
        src104 <= 16'h31f0;
        src105 <= 16'hf462;
        src106 <= 16'he7d0;
        src107 <= 16'h1e00;
        src108 <= 16'hfddf;
        src109 <= 16'h1753;
        src110 <= 16'h18fc;
        src111 <= 16'h7c5a;
        src112 <= 16'h2d35;
        src113 <= 16'hf195;
        src114 <= 16'h2199;
        src115 <= 16'h8211;
        src116 <= 16'hd126;
        src117 <= 16'hebb3;
        src118 <= 16'h23c;
        src119 <= 16'he8db;
        src120 <= 16'h2c9f;
        src121 <= 16'h6d17;
        src122 <= 16'hc371;
        src123 <= 16'he1dc;
        src124 <= 16'h3e8b;
        src125 <= 16'h1552;
        src126 <= 16'h52ec;
        src127 <= 16'h1382;
        exp <= 23'h3e4515;
        #1
        src0 <= 16'hec59;
        src1 <= 16'h8be4;
        src2 <= 16'hd99e;
        src3 <= 16'h211c;
        src4 <= 16'h4a8;
        src5 <= 16'h3ee6;
        src6 <= 16'h585f;
        src7 <= 16'h4659;
        src8 <= 16'h445f;
        src9 <= 16'h33e2;
        src10 <= 16'hb47b;
        src11 <= 16'h3ccf;
        src12 <= 16'h532c;
        src13 <= 16'hb21e;
        src14 <= 16'ha4a9;
        src15 <= 16'hb82c;
        src16 <= 16'h3be6;
        src17 <= 16'ha08e;
        src18 <= 16'h7651;
        src19 <= 16'hf5fb;
        src20 <= 16'h62fd;
        src21 <= 16'h68b0;
        src22 <= 16'hc908;
        src23 <= 16'h1af6;
        src24 <= 16'h124c;
        src25 <= 16'hf9e1;
        src26 <= 16'h9e31;
        src27 <= 16'h922a;
        src28 <= 16'ha73;
        src29 <= 16'h293c;
        src30 <= 16'hb605;
        src31 <= 16'hde6;
        src32 <= 16'hfedb;
        src33 <= 16'h2560;
        src34 <= 16'h25dd;
        src35 <= 16'h68b9;
        src36 <= 16'he85c;
        src37 <= 16'ha46;
        src38 <= 16'ha876;
        src39 <= 16'hc0a2;
        src40 <= 16'ha2ba;
        src41 <= 16'h5ce8;
        src42 <= 16'he091;
        src43 <= 16'h83f5;
        src44 <= 16'hf08f;
        src45 <= 16'he957;
        src46 <= 16'h4f31;
        src47 <= 16'he4cc;
        src48 <= 16'h7464;
        src49 <= 16'h80bc;
        src50 <= 16'h9d98;
        src51 <= 16'h1859;
        src52 <= 16'h86db;
        src53 <= 16'h4ae5;
        src54 <= 16'hbd1c;
        src55 <= 16'hfa24;
        src56 <= 16'hc4cd;
        src57 <= 16'h7107;
        src58 <= 16'h4669;
        src59 <= 16'h5459;
        src60 <= 16'h70d0;
        src61 <= 16'h59fa;
        src62 <= 16'h98f9;
        src63 <= 16'h3987;
        src64 <= 16'hebd9;
        src65 <= 16'h83e3;
        src66 <= 16'hf9c6;
        src67 <= 16'h9702;
        src68 <= 16'hd110;
        src69 <= 16'h7fe7;
        src70 <= 16'hf774;
        src71 <= 16'hab06;
        src72 <= 16'h22e3;
        src73 <= 16'h18eb;
        src74 <= 16'h7c6b;
        src75 <= 16'h466d;
        src76 <= 16'h8670;
        src77 <= 16'h438b;
        src78 <= 16'h5206;
        src79 <= 16'habaf;
        src80 <= 16'hfd7f;
        src81 <= 16'h6c11;
        src82 <= 16'he2de;
        src83 <= 16'h5644;
        src84 <= 16'hc2b;
        src85 <= 16'h5c0d;
        src86 <= 16'h2b6f;
        src87 <= 16'h1cb9;
        src88 <= 16'hc825;
        src89 <= 16'h5f4;
        src90 <= 16'h62e3;
        src91 <= 16'h8bc9;
        src92 <= 16'h4e43;
        src93 <= 16'h8c1c;
        src94 <= 16'hf134;
        src95 <= 16'h7d99;
        src96 <= 16'h9dd8;
        src97 <= 16'h844a;
        src98 <= 16'hda06;
        src99 <= 16'hb114;
        src100 <= 16'h3180;
        src101 <= 16'hcdf2;
        src102 <= 16'h955;
        src103 <= 16'hacd3;
        src104 <= 16'hef7d;
        src105 <= 16'hfc7a;
        src106 <= 16'hfd48;
        src107 <= 16'h25f0;
        src108 <= 16'hdbdf;
        src109 <= 16'h5393;
        src110 <= 16'hef0;
        src111 <= 16'h16bc;
        src112 <= 16'hc1f1;
        src113 <= 16'h78f8;
        src114 <= 16'h6b11;
        src115 <= 16'he8ae;
        src116 <= 16'hdb1;
        src117 <= 16'hd12b;
        src118 <= 16'hf151;
        src119 <= 16'h6fe3;
        src120 <= 16'h1722;
        src121 <= 16'h8362;
        src122 <= 16'h3f9a;
        src123 <= 16'had14;
        src124 <= 16'h42fd;
        src125 <= 16'h1820;
        src126 <= 16'h7258;
        src127 <= 16'hed44;
        exp <= 23'h405b0f;
        #1
        src0 <= 16'h6574;
        src1 <= 16'hf734;
        src2 <= 16'h91fe;
        src3 <= 16'h17db;
        src4 <= 16'h80ea;
        src5 <= 16'h658e;
        src6 <= 16'h2899;
        src7 <= 16'h2921;
        src8 <= 16'h46ad;
        src9 <= 16'ha086;
        src10 <= 16'hc50e;
        src11 <= 16'h210f;
        src12 <= 16'hdaab;
        src13 <= 16'h818d;
        src14 <= 16'h962e;
        src15 <= 16'h4888;
        src16 <= 16'h4597;
        src17 <= 16'h2952;
        src18 <= 16'hb884;
        src19 <= 16'h50cb;
        src20 <= 16'h2eec;
        src21 <= 16'h6578;
        src22 <= 16'h94a1;
        src23 <= 16'hfae8;
        src24 <= 16'h16c8;
        src25 <= 16'h4317;
        src26 <= 16'h6ebf;
        src27 <= 16'hcfea;
        src28 <= 16'h4688;
        src29 <= 16'h6772;
        src30 <= 16'h6754;
        src31 <= 16'hd12f;
        src32 <= 16'h488c;
        src33 <= 16'he4e1;
        src34 <= 16'h886b;
        src35 <= 16'h8147;
        src36 <= 16'ha8cf;
        src37 <= 16'hbcff;
        src38 <= 16'hd505;
        src39 <= 16'he8b9;
        src40 <= 16'hbe15;
        src41 <= 16'h109b;
        src42 <= 16'h98ec;
        src43 <= 16'hb25e;
        src44 <= 16'h5abe;
        src45 <= 16'hcc15;
        src46 <= 16'h798f;
        src47 <= 16'hf992;
        src48 <= 16'hb180;
        src49 <= 16'hee59;
        src50 <= 16'he898;
        src51 <= 16'h4326;
        src52 <= 16'h8edb;
        src53 <= 16'hdfb8;
        src54 <= 16'hd3a2;
        src55 <= 16'hbce;
        src56 <= 16'hf530;
        src57 <= 16'h6dfb;
        src58 <= 16'h19ee;
        src59 <= 16'h373b;
        src60 <= 16'h1220;
        src61 <= 16'hba54;
        src62 <= 16'h18fb;
        src63 <= 16'he63a;
        src64 <= 16'h4151;
        src65 <= 16'hd599;
        src66 <= 16'hb8e4;
        src67 <= 16'he844;
        src68 <= 16'h6621;
        src69 <= 16'h143f;
        src70 <= 16'h58e;
        src71 <= 16'hc373;
        src72 <= 16'hdedf;
        src73 <= 16'h84f4;
        src74 <= 16'hb276;
        src75 <= 16'he8e8;
        src76 <= 16'heb22;
        src77 <= 16'hd86e;
        src78 <= 16'h81b1;
        src79 <= 16'hd247;
        src80 <= 16'h73ff;
        src81 <= 16'ha2e5;
        src82 <= 16'hd8c5;
        src83 <= 16'h42b9;
        src84 <= 16'h2d15;
        src85 <= 16'hd481;
        src86 <= 16'h3712;
        src87 <= 16'h9856;
        src88 <= 16'h7570;
        src89 <= 16'h7ee4;
        src90 <= 16'h8244;
        src91 <= 16'h9a5d;
        src92 <= 16'h4c6c;
        src93 <= 16'ha227;
        src94 <= 16'h9591;
        src95 <= 16'h4499;
        src96 <= 16'h815c;
        src97 <= 16'h8be0;
        src98 <= 16'h209b;
        src99 <= 16'h1692;
        src100 <= 16'h2c79;
        src101 <= 16'h305a;
        src102 <= 16'h3336;
        src103 <= 16'hdcdf;
        src104 <= 16'h5a23;
        src105 <= 16'ha94b;
        src106 <= 16'h9307;
        src107 <= 16'h5297;
        src108 <= 16'hc185;
        src109 <= 16'hdc1a;
        src110 <= 16'hd2a;
        src111 <= 16'hd317;
        src112 <= 16'h5de4;
        src113 <= 16'h8f53;
        src114 <= 16'hb622;
        src115 <= 16'h630;
        src116 <= 16'hf46f;
        src117 <= 16'ha25c;
        src118 <= 16'h299c;
        src119 <= 16'h96f2;
        src120 <= 16'h2cec;
        src121 <= 16'h2231;
        src122 <= 16'hcc49;
        src123 <= 16'h5a5f;
        src124 <= 16'hadc0;
        src125 <= 16'h1a41;
        src126 <= 16'hb2d1;
        src127 <= 16'h6aea;
        exp <= 23'h416e29;
        #1
        src0 <= 16'h6193;
        src1 <= 16'h2063;
        src2 <= 16'hbe30;
        src3 <= 16'h7861;
        src4 <= 16'h166c;
        src5 <= 16'h6b65;
        src6 <= 16'h68f5;
        src7 <= 16'hf9d7;
        src8 <= 16'h89df;
        src9 <= 16'h6b;
        src10 <= 16'h572b;
        src11 <= 16'h9477;
        src12 <= 16'hbb02;
        src13 <= 16'h722c;
        src14 <= 16'h24cc;
        src15 <= 16'h7959;
        src16 <= 16'hac5b;
        src17 <= 16'h30b7;
        src18 <= 16'h4dac;
        src19 <= 16'he9c7;
        src20 <= 16'hfb09;
        src21 <= 16'hbfb9;
        src22 <= 16'h2624;
        src23 <= 16'h48b;
        src24 <= 16'h5510;
        src25 <= 16'hfc54;
        src26 <= 16'h8f33;
        src27 <= 16'hb7c7;
        src28 <= 16'hb4d8;
        src29 <= 16'hd0a6;
        src30 <= 16'hdd3a;
        src31 <= 16'h5852;
        src32 <= 16'h3416;
        src33 <= 16'h7203;
        src34 <= 16'h1e80;
        src35 <= 16'hc9f4;
        src36 <= 16'hdf58;
        src37 <= 16'h9cdb;
        src38 <= 16'hd044;
        src39 <= 16'h8a8c;
        src40 <= 16'h4719;
        src41 <= 16'hb0dd;
        src42 <= 16'h1b87;
        src43 <= 16'hf50c;
        src44 <= 16'h54f9;
        src45 <= 16'hff4a;
        src46 <= 16'h3de1;
        src47 <= 16'haecd;
        src48 <= 16'hac33;
        src49 <= 16'h60a0;
        src50 <= 16'h2f8b;
        src51 <= 16'hb6ae;
        src52 <= 16'h3a59;
        src53 <= 16'h380d;
        src54 <= 16'h909e;
        src55 <= 16'hc557;
        src56 <= 16'hc16b;
        src57 <= 16'h7450;
        src58 <= 16'hb5f0;
        src59 <= 16'he079;
        src60 <= 16'hef65;
        src61 <= 16'he3c;
        src62 <= 16'hee5;
        src63 <= 16'h98c0;
        src64 <= 16'hd589;
        src65 <= 16'h4de7;
        src66 <= 16'h9f0c;
        src67 <= 16'h10bf;
        src68 <= 16'h23e6;
        src69 <= 16'hbd2e;
        src70 <= 16'h776d;
        src71 <= 16'h775a;
        src72 <= 16'h5026;
        src73 <= 16'hf254;
        src74 <= 16'hf7a6;
        src75 <= 16'h7562;
        src76 <= 16'h6f64;
        src77 <= 16'h7d4e;
        src78 <= 16'hd3ac;
        src79 <= 16'h2298;
        src80 <= 16'h7b03;
        src81 <= 16'h58b0;
        src82 <= 16'haf;
        src83 <= 16'h8e46;
        src84 <= 16'ha7fe;
        src85 <= 16'h285b;
        src86 <= 16'h7013;
        src87 <= 16'he02f;
        src88 <= 16'h3171;
        src89 <= 16'ha338;
        src90 <= 16'h90b8;
        src91 <= 16'hb384;
        src92 <= 16'h57de;
        src93 <= 16'h84ba;
        src94 <= 16'h67c6;
        src95 <= 16'h45ca;
        src96 <= 16'h1ce1;
        src97 <= 16'h2a3f;
        src98 <= 16'h59ef;
        src99 <= 16'h36c0;
        src100 <= 16'h7da;
        src101 <= 16'h4a65;
        src102 <= 16'h6783;
        src103 <= 16'h77e0;
        src104 <= 16'hbaaf;
        src105 <= 16'hf2f8;
        src106 <= 16'hb8c;
        src107 <= 16'h2db6;
        src108 <= 16'hf0eb;
        src109 <= 16'he9a9;
        src110 <= 16'h3108;
        src111 <= 16'h8ade;
        src112 <= 16'h2849;
        src113 <= 16'h6633;
        src114 <= 16'h4c6;
        src115 <= 16'hfdef;
        src116 <= 16'h8388;
        src117 <= 16'hfeca;
        src118 <= 16'ha9e7;
        src119 <= 16'h3f55;
        src120 <= 16'hcfc;
        src121 <= 16'h4e07;
        src122 <= 16'h532d;
        src123 <= 16'h1654;
        src124 <= 16'h52fc;
        src125 <= 16'h2ba0;
        src126 <= 16'h5486;
        src127 <= 16'hb27b;
        exp <= 23'h3d312e;
        #1
        src0 <= 16'hf118;
        src1 <= 16'h8035;
        src2 <= 16'he1ec;
        src3 <= 16'h30b1;
        src4 <= 16'h7648;
        src5 <= 16'h34e7;
        src6 <= 16'h3af0;
        src7 <= 16'h774;
        src8 <= 16'h3231;
        src9 <= 16'h9445;
        src10 <= 16'h78a5;
        src11 <= 16'h4175;
        src12 <= 16'h6e60;
        src13 <= 16'h277c;
        src14 <= 16'h76d4;
        src15 <= 16'hdf7c;
        src16 <= 16'he114;
        src17 <= 16'h1ac3;
        src18 <= 16'h1795;
        src19 <= 16'h6e29;
        src20 <= 16'h9415;
        src21 <= 16'ha70;
        src22 <= 16'h21ba;
        src23 <= 16'h9875;
        src24 <= 16'hbd42;
        src25 <= 16'h946;
        src26 <= 16'h871c;
        src27 <= 16'hfa95;
        src28 <= 16'h5c6f;
        src29 <= 16'h634f;
        src30 <= 16'hc66f;
        src31 <= 16'hffc0;
        src32 <= 16'hfdd;
        src33 <= 16'h97e4;
        src34 <= 16'h1891;
        src35 <= 16'hc075;
        src36 <= 16'h7634;
        src37 <= 16'h8fd0;
        src38 <= 16'h30f7;
        src39 <= 16'h42f2;
        src40 <= 16'h307a;
        src41 <= 16'h4970;
        src42 <= 16'hadff;
        src43 <= 16'h3fd;
        src44 <= 16'h4859;
        src45 <= 16'he357;
        src46 <= 16'hcaac;
        src47 <= 16'hda22;
        src48 <= 16'h7663;
        src49 <= 16'h525f;
        src50 <= 16'h1ff0;
        src51 <= 16'h433c;
        src52 <= 16'hd757;
        src53 <= 16'haa90;
        src54 <= 16'hea0d;
        src55 <= 16'h2c75;
        src56 <= 16'h95ba;
        src57 <= 16'h80e9;
        src58 <= 16'h55a;
        src59 <= 16'h722f;
        src60 <= 16'hf044;
        src61 <= 16'h2196;
        src62 <= 16'h3a5a;
        src63 <= 16'ha875;
        src64 <= 16'h3951;
        src65 <= 16'he2c5;
        src66 <= 16'hce25;
        src67 <= 16'hc68;
        src68 <= 16'h45df;
        src69 <= 16'h7fa8;
        src70 <= 16'hb0ca;
        src71 <= 16'h32fe;
        src72 <= 16'hd5f9;
        src73 <= 16'hc32b;
        src74 <= 16'hf71c;
        src75 <= 16'h8f36;
        src76 <= 16'h4d5;
        src77 <= 16'hfaf2;
        src78 <= 16'h205d;
        src79 <= 16'h9695;
        src80 <= 16'hbe92;
        src81 <= 16'h78f9;
        src82 <= 16'hf209;
        src83 <= 16'h2320;
        src84 <= 16'h2911;
        src85 <= 16'h76ce;
        src86 <= 16'hc4b;
        src87 <= 16'h43dd;
        src88 <= 16'h98ef;
        src89 <= 16'h1329;
        src90 <= 16'hc00a;
        src91 <= 16'hb80a;
        src92 <= 16'h49d2;
        src93 <= 16'h7ce3;
        src94 <= 16'h8824;
        src95 <= 16'h147e;
        src96 <= 16'h58dc;
        src97 <= 16'h786d;
        src98 <= 16'h8c92;
        src99 <= 16'hd3d6;
        src100 <= 16'h894f;
        src101 <= 16'h70c3;
        src102 <= 16'hfdbc;
        src103 <= 16'h8f0f;
        src104 <= 16'h43a4;
        src105 <= 16'hee36;
        src106 <= 16'h131e;
        src107 <= 16'h8f63;
        src108 <= 16'h66be;
        src109 <= 16'habf4;
        src110 <= 16'h3236;
        src111 <= 16'h6edd;
        src112 <= 16'haa98;
        src113 <= 16'h44c;
        src114 <= 16'hbe79;
        src115 <= 16'h228e;
        src116 <= 16'h708c;
        src117 <= 16'h9eb9;
        src118 <= 16'hb4cc;
        src119 <= 16'h21c7;
        src120 <= 16'h75f9;
        src121 <= 16'h5ecf;
        src122 <= 16'h6a3b;
        src123 <= 16'h3466;
        src124 <= 16'h8a36;
        src125 <= 16'h8bf9;
        src126 <= 16'h3e9d;
        src127 <= 16'he383;
        exp <= 23'h3b6174;
        #1
        src0 <= 16'hae43;
        src1 <= 16'h1644;
        src2 <= 16'hc0ad;
        src3 <= 16'hf8ba;
        src4 <= 16'h21ad;
        src5 <= 16'h25f2;
        src6 <= 16'hade6;
        src7 <= 16'hd4ae;
        src8 <= 16'hdc67;
        src9 <= 16'h4d15;
        src10 <= 16'h7229;
        src11 <= 16'h5ad5;
        src12 <= 16'h202d;
        src13 <= 16'h8479;
        src14 <= 16'hf9fe;
        src15 <= 16'hdb8f;
        src16 <= 16'h379a;
        src17 <= 16'h9015;
        src18 <= 16'h5038;
        src19 <= 16'h191c;
        src20 <= 16'h4acb;
        src21 <= 16'haeab;
        src22 <= 16'h4bd;
        src23 <= 16'hea21;
        src24 <= 16'h6e80;
        src25 <= 16'h2632;
        src26 <= 16'h693;
        src27 <= 16'h1587;
        src28 <= 16'h5b88;
        src29 <= 16'he58f;
        src30 <= 16'h943d;
        src31 <= 16'h73e3;
        src32 <= 16'hfb42;
        src33 <= 16'h1228;
        src34 <= 16'hdd8;
        src35 <= 16'h6852;
        src36 <= 16'hf0b9;
        src37 <= 16'h6b95;
        src38 <= 16'hbbe;
        src39 <= 16'hb5e1;
        src40 <= 16'h28da;
        src41 <= 16'h84d3;
        src42 <= 16'h4cb8;
        src43 <= 16'hd603;
        src44 <= 16'h56a8;
        src45 <= 16'h9b1;
        src46 <= 16'hd8ca;
        src47 <= 16'hcd72;
        src48 <= 16'h549e;
        src49 <= 16'hb24a;
        src50 <= 16'hac4b;
        src51 <= 16'hb1fd;
        src52 <= 16'ha8fb;
        src53 <= 16'hc1f7;
        src54 <= 16'hfbf5;
        src55 <= 16'hd48e;
        src56 <= 16'hd74b;
        src57 <= 16'ha6b0;
        src58 <= 16'he712;
        src59 <= 16'h1cf2;
        src60 <= 16'h44f1;
        src61 <= 16'h18d4;
        src62 <= 16'h6f6d;
        src63 <= 16'h7d4d;
        src64 <= 16'h7035;
        src65 <= 16'h1471;
        src66 <= 16'h867e;
        src67 <= 16'h5601;
        src68 <= 16'hddb5;
        src69 <= 16'h829b;
        src70 <= 16'h4124;
        src71 <= 16'hd032;
        src72 <= 16'hf23d;
        src73 <= 16'h68ea;
        src74 <= 16'h4bb5;
        src75 <= 16'h3330;
        src76 <= 16'h6fe5;
        src77 <= 16'h72f8;
        src78 <= 16'hdf51;
        src79 <= 16'h9b51;
        src80 <= 16'h95e9;
        src81 <= 16'hfc2d;
        src82 <= 16'h14;
        src83 <= 16'ha495;
        src84 <= 16'h52b3;
        src85 <= 16'h5825;
        src86 <= 16'h9dfd;
        src87 <= 16'hee61;
        src88 <= 16'h330b;
        src89 <= 16'h7715;
        src90 <= 16'h62dc;
        src91 <= 16'h2ec5;
        src92 <= 16'hf88;
        src93 <= 16'h9f93;
        src94 <= 16'h2a3e;
        src95 <= 16'hee01;
        src96 <= 16'hf23d;
        src97 <= 16'hef77;
        src98 <= 16'h1a96;
        src99 <= 16'hc543;
        src100 <= 16'h1f62;
        src101 <= 16'h9944;
        src102 <= 16'h95d7;
        src103 <= 16'h53a1;
        src104 <= 16'h6305;
        src105 <= 16'h9bde;
        src106 <= 16'hb45;
        src107 <= 16'h2bfa;
        src108 <= 16'h5cc2;
        src109 <= 16'h437f;
        src110 <= 16'hdc72;
        src111 <= 16'hb638;
        src112 <= 16'he7d0;
        src113 <= 16'hc31c;
        src114 <= 16'h210c;
        src115 <= 16'hc9ad;
        src116 <= 16'h3a59;
        src117 <= 16'hfd55;
        src118 <= 16'he5;
        src119 <= 16'haf45;
        src120 <= 16'hfde6;
        src121 <= 16'h6eea;
        src122 <= 16'he737;
        src123 <= 16'hd335;
        src124 <= 16'h7975;
        src125 <= 16'hcbd2;
        src126 <= 16'h7a1f;
        src127 <= 16'h1477;
        exp <= 23'h40727d;
        #1
        src0 <= 16'he1d9;
        src1 <= 16'h8736;
        src2 <= 16'h45aa;
        src3 <= 16'h20f1;
        src4 <= 16'hda01;
        src5 <= 16'h4fac;
        src6 <= 16'hd264;
        src7 <= 16'h922b;
        src8 <= 16'h5bb9;
        src9 <= 16'hae5e;
        src10 <= 16'hf2aa;
        src11 <= 16'h372b;
        src12 <= 16'hbf64;
        src13 <= 16'h860a;
        src14 <= 16'h6ec8;
        src15 <= 16'h3957;
        src16 <= 16'h1254;
        src17 <= 16'ha0e7;
        src18 <= 16'hf4d;
        src19 <= 16'h854f;
        src20 <= 16'hbeea;
        src21 <= 16'ha64d;
        src22 <= 16'h5b0f;
        src23 <= 16'h454d;
        src24 <= 16'h1c02;
        src25 <= 16'h87aa;
        src26 <= 16'hc37a;
        src27 <= 16'hbef8;
        src28 <= 16'h1caa;
        src29 <= 16'h2185;
        src30 <= 16'hd8cf;
        src31 <= 16'h1a4e;
        src32 <= 16'h70c6;
        src33 <= 16'h5d97;
        src34 <= 16'h53ad;
        src35 <= 16'hbb73;
        src36 <= 16'hc3e2;
        src37 <= 16'hd409;
        src38 <= 16'hffd9;
        src39 <= 16'h39d;
        src40 <= 16'hcb5e;
        src41 <= 16'h6b57;
        src42 <= 16'h43fc;
        src43 <= 16'h727a;
        src44 <= 16'he23d;
        src45 <= 16'h245e;
        src46 <= 16'hae8;
        src47 <= 16'h7cce;
        src48 <= 16'hbc04;
        src49 <= 16'h30ee;
        src50 <= 16'h4494;
        src51 <= 16'h62d2;
        src52 <= 16'hd558;
        src53 <= 16'h81c;
        src54 <= 16'h6c13;
        src55 <= 16'hbb29;
        src56 <= 16'hd12a;
        src57 <= 16'h21dc;
        src58 <= 16'h3029;
        src59 <= 16'he268;
        src60 <= 16'h2054;
        src61 <= 16'ha977;
        src62 <= 16'he84;
        src63 <= 16'hf29d;
        src64 <= 16'h3cda;
        src65 <= 16'hd80e;
        src66 <= 16'hf917;
        src67 <= 16'ha2de;
        src68 <= 16'h38b6;
        src69 <= 16'h8e;
        src70 <= 16'h82a9;
        src71 <= 16'h1615;
        src72 <= 16'hbdf9;
        src73 <= 16'h3cd9;
        src74 <= 16'hb391;
        src75 <= 16'h661c;
        src76 <= 16'h91c6;
        src77 <= 16'h4e7f;
        src78 <= 16'haa66;
        src79 <= 16'hd124;
        src80 <= 16'hb773;
        src81 <= 16'h6f50;
        src82 <= 16'h9c39;
        src83 <= 16'h85dc;
        src84 <= 16'hfcb;
        src85 <= 16'hf525;
        src86 <= 16'h4104;
        src87 <= 16'hafb;
        src88 <= 16'h8a32;
        src89 <= 16'h7cb7;
        src90 <= 16'h79be;
        src91 <= 16'h5383;
        src92 <= 16'h74c7;
        src93 <= 16'h119;
        src94 <= 16'he24c;
        src95 <= 16'hb48e;
        src96 <= 16'h298b;
        src97 <= 16'he7fd;
        src98 <= 16'h32b6;
        src99 <= 16'h6afa;
        src100 <= 16'h3c34;
        src101 <= 16'h2f3;
        src102 <= 16'hd46a;
        src103 <= 16'h5b01;
        src104 <= 16'h5a56;
        src105 <= 16'h7afd;
        src106 <= 16'he674;
        src107 <= 16'h3707;
        src108 <= 16'h7a6a;
        src109 <= 16'he3b0;
        src110 <= 16'hac82;
        src111 <= 16'hbadf;
        src112 <= 16'ha10f;
        src113 <= 16'h14ab;
        src114 <= 16'h80ac;
        src115 <= 16'h5f79;
        src116 <= 16'h4774;
        src117 <= 16'h6b32;
        src118 <= 16'h3d19;
        src119 <= 16'h7ae;
        src120 <= 16'hfdd1;
        src121 <= 16'h186c;
        src122 <= 16'h581f;
        src123 <= 16'hdb76;
        src124 <= 16'h629c;
        src125 <= 16'h8f04;
        src126 <= 16'hc889;
        src127 <= 16'hc70c;
        exp <= 23'h3d1e56;
        #1
        src0 <= 16'h9bc1;
        src1 <= 16'ha0bb;
        src2 <= 16'h65da;
        src3 <= 16'hb299;
        src4 <= 16'h9c05;
        src5 <= 16'h1a0;
        src6 <= 16'hbe1f;
        src7 <= 16'h7b07;
        src8 <= 16'h3929;
        src9 <= 16'h860a;
        src10 <= 16'h6873;
        src11 <= 16'h6d8a;
        src12 <= 16'h8532;
        src13 <= 16'hf7c3;
        src14 <= 16'h8bff;
        src15 <= 16'h60b2;
        src16 <= 16'ha127;
        src17 <= 16'hbdb2;
        src18 <= 16'ha2da;
        src19 <= 16'h8978;
        src20 <= 16'ha6ae;
        src21 <= 16'hc4ed;
        src22 <= 16'h4376;
        src23 <= 16'h82c1;
        src24 <= 16'hd666;
        src25 <= 16'h5274;
        src26 <= 16'h6f8d;
        src27 <= 16'h54e1;
        src28 <= 16'h1b5e;
        src29 <= 16'hba3b;
        src30 <= 16'h16ae;
        src31 <= 16'h8dfa;
        src32 <= 16'h6fc8;
        src33 <= 16'h9144;
        src34 <= 16'h6322;
        src35 <= 16'hb5da;
        src36 <= 16'ha907;
        src37 <= 16'h4bc8;
        src38 <= 16'h2d4f;
        src39 <= 16'hf542;
        src40 <= 16'h1293;
        src41 <= 16'h9ac9;
        src42 <= 16'h33d4;
        src43 <= 16'h8436;
        src44 <= 16'hde9c;
        src45 <= 16'hf2dd;
        src46 <= 16'h95;
        src47 <= 16'hd877;
        src48 <= 16'hae1f;
        src49 <= 16'h9d67;
        src50 <= 16'h99a3;
        src51 <= 16'ha76a;
        src52 <= 16'hf293;
        src53 <= 16'h5fe3;
        src54 <= 16'hdd38;
        src55 <= 16'h2f9d;
        src56 <= 16'h527b;
        src57 <= 16'hd5fc;
        src58 <= 16'hde1d;
        src59 <= 16'he8c4;
        src60 <= 16'h964c;
        src61 <= 16'he21e;
        src62 <= 16'hf6c7;
        src63 <= 16'hee0e;
        src64 <= 16'h42e2;
        src65 <= 16'h3880;
        src66 <= 16'h4623;
        src67 <= 16'hc92e;
        src68 <= 16'h7de3;
        src69 <= 16'h6bff;
        src70 <= 16'h707e;
        src71 <= 16'h74d5;
        src72 <= 16'hac2f;
        src73 <= 16'h238e;
        src74 <= 16'h119e;
        src75 <= 16'h74bb;
        src76 <= 16'ha113;
        src77 <= 16'ha7a3;
        src78 <= 16'hcc67;
        src79 <= 16'hb759;
        src80 <= 16'hfd4d;
        src81 <= 16'hfb64;
        src82 <= 16'h91b;
        src83 <= 16'h3bd2;
        src84 <= 16'h88d7;
        src85 <= 16'h34a9;
        src86 <= 16'hcbe6;
        src87 <= 16'hc98d;
        src88 <= 16'hbeed;
        src89 <= 16'h1626;
        src90 <= 16'h999b;
        src91 <= 16'h4644;
        src92 <= 16'h616f;
        src93 <= 16'h52fc;
        src94 <= 16'h4c63;
        src95 <= 16'h850a;
        src96 <= 16'h9b22;
        src97 <= 16'h15cc;
        src98 <= 16'h3e7d;
        src99 <= 16'h29df;
        src100 <= 16'h2e80;
        src101 <= 16'hec49;
        src102 <= 16'hd2de;
        src103 <= 16'h4376;
        src104 <= 16'h1541;
        src105 <= 16'h171a;
        src106 <= 16'h652;
        src107 <= 16'hd771;
        src108 <= 16'hbaf6;
        src109 <= 16'h99ba;
        src110 <= 16'h4d80;
        src111 <= 16'h3bad;
        src112 <= 16'hc2bf;
        src113 <= 16'hb0d9;
        src114 <= 16'h74a9;
        src115 <= 16'h62b2;
        src116 <= 16'h1e7b;
        src117 <= 16'h7e75;
        src118 <= 16'h5e8b;
        src119 <= 16'hc39d;
        src120 <= 16'heee0;
        src121 <= 16'h1bdf;
        src122 <= 16'heebe;
        src123 <= 16'ha742;
        src124 <= 16'h5ee5;
        src125 <= 16'hbf51;
        src126 <= 16'ha814;
        src127 <= 16'h754a;
        exp <= 23'h42296d;
        #1
        src0 <= 16'hc98a;
        src1 <= 16'h3052;
        src2 <= 16'hb275;
        src3 <= 16'h6769;
        src4 <= 16'h508c;
        src5 <= 16'h676;
        src6 <= 16'h58b;
        src7 <= 16'h9ed5;
        src8 <= 16'h1b1f;
        src9 <= 16'h5b98;
        src10 <= 16'h271a;
        src11 <= 16'hb0;
        src12 <= 16'h2c35;
        src13 <= 16'he891;
        src14 <= 16'h29c8;
        src15 <= 16'h42eb;
        src16 <= 16'hae7f;
        src17 <= 16'ha77f;
        src18 <= 16'h6baf;
        src19 <= 16'hbaab;
        src20 <= 16'h66cd;
        src21 <= 16'he5c0;
        src22 <= 16'h2f1c;
        src23 <= 16'h1b90;
        src24 <= 16'h751a;
        src25 <= 16'hf030;
        src26 <= 16'h2ea2;
        src27 <= 16'hda4a;
        src28 <= 16'h9fb4;
        src29 <= 16'hb5dd;
        src30 <= 16'h1a9c;
        src31 <= 16'h301;
        src32 <= 16'h8099;
        src33 <= 16'h10cc;
        src34 <= 16'he661;
        src35 <= 16'ha8c5;
        src36 <= 16'h9d5d;
        src37 <= 16'h3d51;
        src38 <= 16'hf4f4;
        src39 <= 16'h4adf;
        src40 <= 16'h4827;
        src41 <= 16'hed9a;
        src42 <= 16'hb0ae;
        src43 <= 16'hd959;
        src44 <= 16'hbb60;
        src45 <= 16'h2d82;
        src46 <= 16'h661b;
        src47 <= 16'h4f4a;
        src48 <= 16'hbf5c;
        src49 <= 16'h1d73;
        src50 <= 16'h239b;
        src51 <= 16'hd753;
        src52 <= 16'h12c1;
        src53 <= 16'h4c1a;
        src54 <= 16'had89;
        src55 <= 16'h4e97;
        src56 <= 16'hbe37;
        src57 <= 16'h9826;
        src58 <= 16'h4e59;
        src59 <= 16'h6d65;
        src60 <= 16'hf1ea;
        src61 <= 16'hf08a;
        src62 <= 16'h6fcd;
        src63 <= 16'h7088;
        src64 <= 16'hfbf2;
        src65 <= 16'hf8c4;
        src66 <= 16'h2440;
        src67 <= 16'hf9b6;
        src68 <= 16'ha6e4;
        src69 <= 16'h8170;
        src70 <= 16'h3469;
        src71 <= 16'h2ffa;
        src72 <= 16'hfa12;
        src73 <= 16'h39fd;
        src74 <= 16'hb1aa;
        src75 <= 16'h3158;
        src76 <= 16'hb3d1;
        src77 <= 16'hf78c;
        src78 <= 16'hc3e7;
        src79 <= 16'ha390;
        src80 <= 16'h70f;
        src81 <= 16'h245d;
        src82 <= 16'h36c0;
        src83 <= 16'h3c01;
        src84 <= 16'hc950;
        src85 <= 16'hc2c2;
        src86 <= 16'h93b6;
        src87 <= 16'he;
        src88 <= 16'h89f5;
        src89 <= 16'h7637;
        src90 <= 16'hfed0;
        src91 <= 16'h1e0e;
        src92 <= 16'h28be;
        src93 <= 16'hda6e;
        src94 <= 16'h1e33;
        src95 <= 16'hcca6;
        src96 <= 16'h22bf;
        src97 <= 16'hf737;
        src98 <= 16'hd5c9;
        src99 <= 16'h3f24;
        src100 <= 16'h6ce7;
        src101 <= 16'h23e9;
        src102 <= 16'hf879;
        src103 <= 16'h351f;
        src104 <= 16'hb980;
        src105 <= 16'hf6fe;
        src106 <= 16'h3735;
        src107 <= 16'ha121;
        src108 <= 16'h3c18;
        src109 <= 16'hb5d1;
        src110 <= 16'h931b;
        src111 <= 16'h1353;
        src112 <= 16'h1639;
        src113 <= 16'h70c8;
        src114 <= 16'hde27;
        src115 <= 16'h856d;
        src116 <= 16'ha074;
        src117 <= 16'had40;
        src118 <= 16'h1a75;
        src119 <= 16'h6cb5;
        src120 <= 16'h856b;
        src121 <= 16'h3eed;
        src122 <= 16'h6339;
        src123 <= 16'h1f4f;
        src124 <= 16'h92a9;
        src125 <= 16'h574c;
        src126 <= 16'h8b60;
        src127 <= 16'h169d;
        exp <= 23'h3cf7d7;
        #1
        src0 <= 16'h1440;
        src1 <= 16'hebf9;
        src2 <= 16'h9d3c;
        src3 <= 16'h4b0d;
        src4 <= 16'hb7f5;
        src5 <= 16'h822c;
        src6 <= 16'h2212;
        src7 <= 16'h427f;
        src8 <= 16'h7de0;
        src9 <= 16'h6930;
        src10 <= 16'h6f07;
        src11 <= 16'h9f1a;
        src12 <= 16'h56b0;
        src13 <= 16'he520;
        src14 <= 16'h4e2b;
        src15 <= 16'hc7ef;
        src16 <= 16'hc113;
        src17 <= 16'hc3c6;
        src18 <= 16'h69d1;
        src19 <= 16'ha7f7;
        src20 <= 16'hd3f0;
        src21 <= 16'hb393;
        src22 <= 16'hea42;
        src23 <= 16'h712f;
        src24 <= 16'hd1b7;
        src25 <= 16'h8cf6;
        src26 <= 16'h5f2f;
        src27 <= 16'hb071;
        src28 <= 16'hd691;
        src29 <= 16'h2ff1;
        src30 <= 16'h8c9e;
        src31 <= 16'h72fc;
        src32 <= 16'hc008;
        src33 <= 16'h934d;
        src34 <= 16'h530f;
        src35 <= 16'hc580;
        src36 <= 16'h7de8;
        src37 <= 16'h9804;
        src38 <= 16'hd77b;
        src39 <= 16'hff75;
        src40 <= 16'h2df3;
        src41 <= 16'hd262;
        src42 <= 16'hdbeb;
        src43 <= 16'h95dd;
        src44 <= 16'he87a;
        src45 <= 16'h9189;
        src46 <= 16'h92e7;
        src47 <= 16'h741;
        src48 <= 16'h2ea2;
        src49 <= 16'hbd7f;
        src50 <= 16'hf11c;
        src51 <= 16'h7bc8;
        src52 <= 16'h71a4;
        src53 <= 16'h2c60;
        src54 <= 16'hfee0;
        src55 <= 16'hffc;
        src56 <= 16'h6c29;
        src57 <= 16'hf9ce;
        src58 <= 16'haa5d;
        src59 <= 16'h6ce8;
        src60 <= 16'h6adc;
        src61 <= 16'h7ef3;
        src62 <= 16'h1482;
        src63 <= 16'hef69;
        src64 <= 16'hcc18;
        src65 <= 16'h7ccf;
        src66 <= 16'hf6f2;
        src67 <= 16'ha756;
        src68 <= 16'h652f;
        src69 <= 16'hd94c;
        src70 <= 16'hbffd;
        src71 <= 16'h7dad;
        src72 <= 16'h7c22;
        src73 <= 16'hbb4a;
        src74 <= 16'hff95;
        src75 <= 16'h3d9b;
        src76 <= 16'h5c67;
        src77 <= 16'h2723;
        src78 <= 16'h5b75;
        src79 <= 16'h4f6e;
        src80 <= 16'hb5b7;
        src81 <= 16'hd833;
        src82 <= 16'h3302;
        src83 <= 16'h192c;
        src84 <= 16'h693e;
        src85 <= 16'h648f;
        src86 <= 16'h6643;
        src87 <= 16'h6d8;
        src88 <= 16'h3473;
        src89 <= 16'h561c;
        src90 <= 16'h236a;
        src91 <= 16'ha643;
        src92 <= 16'h3e8f;
        src93 <= 16'h5e5c;
        src94 <= 16'h58ea;
        src95 <= 16'h73f0;
        src96 <= 16'h98f5;
        src97 <= 16'ha6c5;
        src98 <= 16'h8ce1;
        src99 <= 16'hbbb4;
        src100 <= 16'hcbdd;
        src101 <= 16'hd8b7;
        src102 <= 16'h9a91;
        src103 <= 16'h729b;
        src104 <= 16'hd5a1;
        src105 <= 16'hb502;
        src106 <= 16'h44e9;
        src107 <= 16'hfb4f;
        src108 <= 16'h9612;
        src109 <= 16'he51c;
        src110 <= 16'h7399;
        src111 <= 16'h7fad;
        src112 <= 16'h689b;
        src113 <= 16'h825d;
        src114 <= 16'h86a6;
        src115 <= 16'hdfe8;
        src116 <= 16'h41c9;
        src117 <= 16'h57c0;
        src118 <= 16'h3956;
        src119 <= 16'had8b;
        src120 <= 16'h85b0;
        src121 <= 16'hdb72;
        src122 <= 16'h3541;
        src123 <= 16'hcbb9;
        src124 <= 16'h7b57;
        src125 <= 16'hed4d;
        src126 <= 16'ha325;
        src127 <= 16'heac3;
        exp <= 23'h468384;
        #1
        src0 <= 16'hebd9;
        src1 <= 16'hbb24;
        src2 <= 16'h5072;
        src3 <= 16'h1b23;
        src4 <= 16'h9bb;
        src5 <= 16'h9419;
        src6 <= 16'h4536;
        src7 <= 16'h8c3a;
        src8 <= 16'hdaaa;
        src9 <= 16'h6d96;
        src10 <= 16'h9414;
        src11 <= 16'h92f0;
        src12 <= 16'h8115;
        src13 <= 16'h2bca;
        src14 <= 16'h8073;
        src15 <= 16'h77ab;
        src16 <= 16'h7952;
        src17 <= 16'h6a1b;
        src18 <= 16'h63dc;
        src19 <= 16'h6af5;
        src20 <= 16'h4927;
        src21 <= 16'ha1d1;
        src22 <= 16'h47d0;
        src23 <= 16'h9d29;
        src24 <= 16'h51cc;
        src25 <= 16'he926;
        src26 <= 16'hb426;
        src27 <= 16'h558d;
        src28 <= 16'h96bd;
        src29 <= 16'h5668;
        src30 <= 16'he1a3;
        src31 <= 16'h677c;
        src32 <= 16'h975b;
        src33 <= 16'h25e3;
        src34 <= 16'h6b25;
        src35 <= 16'h6535;
        src36 <= 16'h761;
        src37 <= 16'hc808;
        src38 <= 16'h449d;
        src39 <= 16'h9374;
        src40 <= 16'h2b27;
        src41 <= 16'h1ced;
        src42 <= 16'h6723;
        src43 <= 16'hf6d7;
        src44 <= 16'hf6c8;
        src45 <= 16'habe3;
        src46 <= 16'h2a8b;
        src47 <= 16'h77c1;
        src48 <= 16'h9e72;
        src49 <= 16'hb303;
        src50 <= 16'hd2c5;
        src51 <= 16'h662e;
        src52 <= 16'hc2ff;
        src53 <= 16'hb714;
        src54 <= 16'h3c6f;
        src55 <= 16'h228c;
        src56 <= 16'h43d1;
        src57 <= 16'hac99;
        src58 <= 16'h2904;
        src59 <= 16'h430f;
        src60 <= 16'ha93e;
        src61 <= 16'h5eab;
        src62 <= 16'hdf9;
        src63 <= 16'hacd3;
        src64 <= 16'hbe9f;
        src65 <= 16'hc269;
        src66 <= 16'h269a;
        src67 <= 16'hb2f3;
        src68 <= 16'h12d6;
        src69 <= 16'h9c7;
        src70 <= 16'h3faa;
        src71 <= 16'hbe64;
        src72 <= 16'he6b3;
        src73 <= 16'hb36b;
        src74 <= 16'hddb8;
        src75 <= 16'hd502;
        src76 <= 16'h5ee2;
        src77 <= 16'hb213;
        src78 <= 16'hafae;
        src79 <= 16'hc9a1;
        src80 <= 16'h782c;
        src81 <= 16'h27ca;
        src82 <= 16'h7d1b;
        src83 <= 16'hc0b9;
        src84 <= 16'h2294;
        src85 <= 16'hbdd1;
        src86 <= 16'had9f;
        src87 <= 16'h4b66;
        src88 <= 16'h9e02;
        src89 <= 16'h3d28;
        src90 <= 16'hdb56;
        src91 <= 16'h6e89;
        src92 <= 16'h8d28;
        src93 <= 16'he230;
        src94 <= 16'h101b;
        src95 <= 16'h39af;
        src96 <= 16'h6836;
        src97 <= 16'haa89;
        src98 <= 16'hdd87;
        src99 <= 16'h6dea;
        src100 <= 16'h5ba7;
        src101 <= 16'ha930;
        src102 <= 16'hfc11;
        src103 <= 16'h2461;
        src104 <= 16'h16d4;
        src105 <= 16'h59fe;
        src106 <= 16'hd692;
        src107 <= 16'h8600;
        src108 <= 16'hd55d;
        src109 <= 16'h3583;
        src110 <= 16'he838;
        src111 <= 16'h5456;
        src112 <= 16'h775c;
        src113 <= 16'h4621;
        src114 <= 16'h411b;
        src115 <= 16'hb28;
        src116 <= 16'h76f3;
        src117 <= 16'h2b9b;
        src118 <= 16'h6321;
        src119 <= 16'haa23;
        src120 <= 16'ha6d3;
        src121 <= 16'h69e9;
        src122 <= 16'hf51d;
        src123 <= 16'ha78c;
        src124 <= 16'h5619;
        src125 <= 16'hb9;
        src126 <= 16'hc788;
        src127 <= 16'hd97d;
        exp <= 23'h3f0ec2;
        #1
        src0 <= 16'hbc46;
        src1 <= 16'h3865;
        src2 <= 16'h97bf;
        src3 <= 16'hc40a;
        src4 <= 16'hcd4;
        src5 <= 16'h6e53;
        src6 <= 16'hd96d;
        src7 <= 16'h7a42;
        src8 <= 16'h6b3f;
        src9 <= 16'h23a0;
        src10 <= 16'h9d2d;
        src11 <= 16'h6852;
        src12 <= 16'h2a19;
        src13 <= 16'hce08;
        src14 <= 16'hf04a;
        src15 <= 16'hdb44;
        src16 <= 16'h7f96;
        src17 <= 16'h9e5c;
        src18 <= 16'hefd;
        src19 <= 16'heffa;
        src20 <= 16'hed;
        src21 <= 16'h50cb;
        src22 <= 16'hd9e9;
        src23 <= 16'hcca1;
        src24 <= 16'hd25f;
        src25 <= 16'h9084;
        src26 <= 16'he8a7;
        src27 <= 16'h4f74;
        src28 <= 16'hec51;
        src29 <= 16'h327b;
        src30 <= 16'h8bcc;
        src31 <= 16'he556;
        src32 <= 16'hf6ec;
        src33 <= 16'hdf62;
        src34 <= 16'he30e;
        src35 <= 16'hf47d;
        src36 <= 16'h8f28;
        src37 <= 16'h1965;
        src38 <= 16'hed1;
        src39 <= 16'hdf93;
        src40 <= 16'ha3dd;
        src41 <= 16'h98cd;
        src42 <= 16'h188d;
        src43 <= 16'h19a0;
        src44 <= 16'h31fe;
        src45 <= 16'haa91;
        src46 <= 16'h4a2e;
        src47 <= 16'h8f5;
        src48 <= 16'h9874;
        src49 <= 16'h53e2;
        src50 <= 16'h8515;
        src51 <= 16'h9db6;
        src52 <= 16'hd3fd;
        src53 <= 16'h8796;
        src54 <= 16'h6394;
        src55 <= 16'h97b;
        src56 <= 16'h25d9;
        src57 <= 16'h716d;
        src58 <= 16'hbdf8;
        src59 <= 16'hbec7;
        src60 <= 16'ha101;
        src61 <= 16'h4916;
        src62 <= 16'he9f2;
        src63 <= 16'hce74;
        src64 <= 16'h3608;
        src65 <= 16'h2a58;
        src66 <= 16'h374f;
        src67 <= 16'h2fac;
        src68 <= 16'h4bdd;
        src69 <= 16'h7b24;
        src70 <= 16'h2c33;
        src71 <= 16'hc887;
        src72 <= 16'h43e;
        src73 <= 16'h1482;
        src74 <= 16'h63ca;
        src75 <= 16'h1dd2;
        src76 <= 16'h2594;
        src77 <= 16'hc93b;
        src78 <= 16'h5233;
        src79 <= 16'h4446;
        src80 <= 16'h2df3;
        src81 <= 16'h4d53;
        src82 <= 16'hbd4e;
        src83 <= 16'hc041;
        src84 <= 16'h391;
        src85 <= 16'hd59b;
        src86 <= 16'hf582;
        src87 <= 16'h12c7;
        src88 <= 16'h5872;
        src89 <= 16'h222a;
        src90 <= 16'hc076;
        src91 <= 16'hedf4;
        src92 <= 16'h55e8;
        src93 <= 16'ha661;
        src94 <= 16'h233f;
        src95 <= 16'hcebb;
        src96 <= 16'hf38c;
        src97 <= 16'h5a0f;
        src98 <= 16'h487;
        src99 <= 16'h5b8b;
        src100 <= 16'h18c4;
        src101 <= 16'h62fc;
        src102 <= 16'h8c7d;
        src103 <= 16'h4b11;
        src104 <= 16'h2ad6;
        src105 <= 16'h8b66;
        src106 <= 16'h4f2e;
        src107 <= 16'h8636;
        src108 <= 16'h1b5b;
        src109 <= 16'h6e21;
        src110 <= 16'h49e0;
        src111 <= 16'h4256;
        src112 <= 16'h2f6f;
        src113 <= 16'h8361;
        src114 <= 16'h635f;
        src115 <= 16'hb706;
        src116 <= 16'ha592;
        src117 <= 16'h7ae6;
        src118 <= 16'h4508;
        src119 <= 16'hdc46;
        src120 <= 16'he861;
        src121 <= 16'h4830;
        src122 <= 16'h5ca5;
        src123 <= 16'hd78a;
        src124 <= 16'h7150;
        src125 <= 16'ha8a3;
        src126 <= 16'hf50;
        src127 <= 16'h755e;
        exp <= 23'h3c71fc;
        #1
        src0 <= 16'h6f5c;
        src1 <= 16'h3c19;
        src2 <= 16'h2fee;
        src3 <= 16'ha00d;
        src4 <= 16'h7424;
        src5 <= 16'ha69c;
        src6 <= 16'hb96e;
        src7 <= 16'hb9b1;
        src8 <= 16'h7e;
        src9 <= 16'h63a3;
        src10 <= 16'hdf12;
        src11 <= 16'hd478;
        src12 <= 16'h810c;
        src13 <= 16'h2723;
        src14 <= 16'h4143;
        src15 <= 16'h32c7;
        src16 <= 16'h8659;
        src17 <= 16'heaf2;
        src18 <= 16'hba98;
        src19 <= 16'h10ef;
        src20 <= 16'h938b;
        src21 <= 16'h1c38;
        src22 <= 16'hc314;
        src23 <= 16'h751a;
        src24 <= 16'h1a15;
        src25 <= 16'h722;
        src26 <= 16'h2527;
        src27 <= 16'heb15;
        src28 <= 16'h6604;
        src29 <= 16'h76cf;
        src30 <= 16'hc7c2;
        src31 <= 16'ha459;
        src32 <= 16'hd280;
        src33 <= 16'h7ddc;
        src34 <= 16'h4cad;
        src35 <= 16'h3039;
        src36 <= 16'hbe43;
        src37 <= 16'hf7af;
        src38 <= 16'hf2ca;
        src39 <= 16'h12ba;
        src40 <= 16'h6756;
        src41 <= 16'h2b8f;
        src42 <= 16'h16d8;
        src43 <= 16'h837e;
        src44 <= 16'h1f7b;
        src45 <= 16'h2e7d;
        src46 <= 16'h3e3c;
        src47 <= 16'h9676;
        src48 <= 16'h8026;
        src49 <= 16'h264e;
        src50 <= 16'h91c0;
        src51 <= 16'h88bf;
        src52 <= 16'hd71d;
        src53 <= 16'h5d56;
        src54 <= 16'h3422;
        src55 <= 16'h2615;
        src56 <= 16'hb154;
        src57 <= 16'h70a6;
        src58 <= 16'hafc2;
        src59 <= 16'h10d;
        src60 <= 16'hbc1b;
        src61 <= 16'hd8bc;
        src62 <= 16'h99ea;
        src63 <= 16'hd0fd;
        src64 <= 16'h6251;
        src65 <= 16'h2ecb;
        src66 <= 16'hef10;
        src67 <= 16'h4ab1;
        src68 <= 16'h8580;
        src69 <= 16'hcc0e;
        src70 <= 16'h4d28;
        src71 <= 16'h35ae;
        src72 <= 16'h801c;
        src73 <= 16'h8126;
        src74 <= 16'h9c48;
        src75 <= 16'hf67c;
        src76 <= 16'h10b8;
        src77 <= 16'h517;
        src78 <= 16'hc0cb;
        src79 <= 16'h5978;
        src80 <= 16'h2de8;
        src81 <= 16'hd4f2;
        src82 <= 16'h8d3c;
        src83 <= 16'hbaaa;
        src84 <= 16'h343c;
        src85 <= 16'ha89d;
        src86 <= 16'h905;
        src87 <= 16'h7d06;
        src88 <= 16'hebed;
        src89 <= 16'h4f66;
        src90 <= 16'h1dc5;
        src91 <= 16'h23be;
        src92 <= 16'he1a5;
        src93 <= 16'h9a9c;
        src94 <= 16'hc961;
        src95 <= 16'h184b;
        src96 <= 16'h53e7;
        src97 <= 16'hc330;
        src98 <= 16'h2126;
        src99 <= 16'hf607;
        src100 <= 16'h52fe;
        src101 <= 16'hfbc1;
        src102 <= 16'h889a;
        src103 <= 16'h59dd;
        src104 <= 16'h178b;
        src105 <= 16'h14b;
        src106 <= 16'h9f45;
        src107 <= 16'h3c42;
        src108 <= 16'h10ac;
        src109 <= 16'h101f;
        src110 <= 16'ha78b;
        src111 <= 16'h6e6e;
        src112 <= 16'h562c;
        src113 <= 16'h4dde;
        src114 <= 16'h434b;
        src115 <= 16'hfb4a;
        src116 <= 16'h7007;
        src117 <= 16'he685;
        src118 <= 16'h74cb;
        src119 <= 16'h9659;
        src120 <= 16'h5a7a;
        src121 <= 16'heeac;
        src122 <= 16'he3f1;
        src123 <= 16'hf45c;
        src124 <= 16'hc77;
        src125 <= 16'h626d;
        src126 <= 16'hdac9;
        src127 <= 16'hc5f1;
        exp <= 23'h3cc2d3;
        #1
        src0 <= 16'hbcf0;
        src1 <= 16'h82e4;
        src2 <= 16'h4607;
        src3 <= 16'hdb45;
        src4 <= 16'h186f;
        src5 <= 16'h569;
        src6 <= 16'h8c58;
        src7 <= 16'h6590;
        src8 <= 16'hc46d;
        src9 <= 16'h6a36;
        src10 <= 16'hd6e7;
        src11 <= 16'h98b;
        src12 <= 16'h6ed8;
        src13 <= 16'haf6;
        src14 <= 16'h5c4f;
        src15 <= 16'he701;
        src16 <= 16'h67e1;
        src17 <= 16'h55a4;
        src18 <= 16'h2e4e;
        src19 <= 16'h47db;
        src20 <= 16'hef0d;
        src21 <= 16'hb163;
        src22 <= 16'ha297;
        src23 <= 16'h5311;
        src24 <= 16'h9a9f;
        src25 <= 16'hbc06;
        src26 <= 16'hef9c;
        src27 <= 16'h1c7a;
        src28 <= 16'hd924;
        src29 <= 16'hf979;
        src30 <= 16'hb7b;
        src31 <= 16'haa21;
        src32 <= 16'h32c4;
        src33 <= 16'h229a;
        src34 <= 16'h3354;
        src35 <= 16'haf32;
        src36 <= 16'h65ec;
        src37 <= 16'he3d3;
        src38 <= 16'h5335;
        src39 <= 16'h1ded;
        src40 <= 16'hb065;
        src41 <= 16'hd770;
        src42 <= 16'hf0f1;
        src43 <= 16'h75e5;
        src44 <= 16'h43f7;
        src45 <= 16'h9e38;
        src46 <= 16'h41fb;
        src47 <= 16'h8cdf;
        src48 <= 16'ha3eb;
        src49 <= 16'h8691;
        src50 <= 16'h659c;
        src51 <= 16'h790f;
        src52 <= 16'h5fcb;
        src53 <= 16'hb8e7;
        src54 <= 16'h7da1;
        src55 <= 16'h8998;
        src56 <= 16'hb1e6;
        src57 <= 16'h52a8;
        src58 <= 16'hf199;
        src59 <= 16'h1254;
        src60 <= 16'hce70;
        src61 <= 16'hdf73;
        src62 <= 16'h6f76;
        src63 <= 16'hc5bf;
        src64 <= 16'ha498;
        src65 <= 16'h865b;
        src66 <= 16'h37e6;
        src67 <= 16'hc142;
        src68 <= 16'h8024;
        src69 <= 16'hb744;
        src70 <= 16'hcab7;
        src71 <= 16'hf581;
        src72 <= 16'h7138;
        src73 <= 16'he882;
        src74 <= 16'haaa1;
        src75 <= 16'hacc2;
        src76 <= 16'h49d1;
        src77 <= 16'hd407;
        src78 <= 16'h45d;
        src79 <= 16'hfc57;
        src80 <= 16'h9f99;
        src81 <= 16'hc295;
        src82 <= 16'hca47;
        src83 <= 16'h68ae;
        src84 <= 16'hbb08;
        src85 <= 16'h995d;
        src86 <= 16'hf70d;
        src87 <= 16'he1f7;
        src88 <= 16'h5240;
        src89 <= 16'hcc4f;
        src90 <= 16'heb66;
        src91 <= 16'h37f2;
        src92 <= 16'hb840;
        src93 <= 16'h19fa;
        src94 <= 16'h8365;
        src95 <= 16'hd0a2;
        src96 <= 16'h1539;
        src97 <= 16'hb72d;
        src98 <= 16'h2fff;
        src99 <= 16'h3815;
        src100 <= 16'h49b0;
        src101 <= 16'h8ff3;
        src102 <= 16'hc30e;
        src103 <= 16'hd3c4;
        src104 <= 16'hf703;
        src105 <= 16'h61d9;
        src106 <= 16'hf49c;
        src107 <= 16'hf8d;
        src108 <= 16'hd148;
        src109 <= 16'hfcb;
        src110 <= 16'h947;
        src111 <= 16'h835e;
        src112 <= 16'h3a42;
        src113 <= 16'h4ef4;
        src114 <= 16'h80d0;
        src115 <= 16'h43b5;
        src116 <= 16'ha2d7;
        src117 <= 16'h2f6;
        src118 <= 16'hd2ea;
        src119 <= 16'hbcc1;
        src120 <= 16'h7a99;
        src121 <= 16'h7455;
        src122 <= 16'h2403;
        src123 <= 16'h9188;
        src124 <= 16'h9d1f;
        src125 <= 16'h6a01;
        src126 <= 16'h42a7;
        src127 <= 16'h7700;
        exp <= 23'h430722;
        #1
        src0 <= 16'h127;
        src1 <= 16'he022;
        src2 <= 16'h26cf;
        src3 <= 16'hcbcf;
        src4 <= 16'h656b;
        src5 <= 16'hbcc6;
        src6 <= 16'ha137;
        src7 <= 16'h10bc;
        src8 <= 16'ha59b;
        src9 <= 16'hb99c;
        src10 <= 16'h9af2;
        src11 <= 16'h5724;
        src12 <= 16'hb844;
        src13 <= 16'hddce;
        src14 <= 16'hcb4d;
        src15 <= 16'h9dfa;
        src16 <= 16'h6c69;
        src17 <= 16'h7440;
        src18 <= 16'he3b5;
        src19 <= 16'h69ec;
        src20 <= 16'hed6c;
        src21 <= 16'he93e;
        src22 <= 16'h193c;
        src23 <= 16'hc21c;
        src24 <= 16'he98;
        src25 <= 16'hcf7a;
        src26 <= 16'he69d;
        src27 <= 16'haf3f;
        src28 <= 16'h2b38;
        src29 <= 16'hac11;
        src30 <= 16'ha3d4;
        src31 <= 16'h2bc5;
        src32 <= 16'h18d1;
        src33 <= 16'h8294;
        src34 <= 16'h5b76;
        src35 <= 16'hcf59;
        src36 <= 16'h35e8;
        src37 <= 16'hda19;
        src38 <= 16'h2d5;
        src39 <= 16'hd9b;
        src40 <= 16'hb1ac;
        src41 <= 16'ha94c;
        src42 <= 16'h30e9;
        src43 <= 16'h33a1;
        src44 <= 16'h2fdd;
        src45 <= 16'h98d;
        src46 <= 16'h7fd3;
        src47 <= 16'hbcc2;
        src48 <= 16'hec4f;
        src49 <= 16'h2180;
        src50 <= 16'h5eda;
        src51 <= 16'hebf4;
        src52 <= 16'h3827;
        src53 <= 16'he97c;
        src54 <= 16'hbee1;
        src55 <= 16'h6143;
        src56 <= 16'he3bc;
        src57 <= 16'h355a;
        src58 <= 16'h25ce;
        src59 <= 16'ha2c1;
        src60 <= 16'haa1a;
        src61 <= 16'h165d;
        src62 <= 16'h2e4d;
        src63 <= 16'hceac;
        src64 <= 16'h7d6a;
        src65 <= 16'hb111;
        src66 <= 16'h985;
        src67 <= 16'ha11e;
        src68 <= 16'hcdd0;
        src69 <= 16'hb280;
        src70 <= 16'h5575;
        src71 <= 16'h4448;
        src72 <= 16'h6f23;
        src73 <= 16'hcce3;
        src74 <= 16'hc2e;
        src75 <= 16'hf0e6;
        src76 <= 16'hbecd;
        src77 <= 16'h87ea;
        src78 <= 16'h5165;
        src79 <= 16'hbd11;
        src80 <= 16'h5968;
        src81 <= 16'h395e;
        src82 <= 16'hf157;
        src83 <= 16'hceaa;
        src84 <= 16'hd9d2;
        src85 <= 16'h39d6;
        src86 <= 16'hf4cb;
        src87 <= 16'h2a5f;
        src88 <= 16'h5e38;
        src89 <= 16'haf4f;
        src90 <= 16'haf42;
        src91 <= 16'he5f9;
        src92 <= 16'h227f;
        src93 <= 16'h913c;
        src94 <= 16'hd395;
        src95 <= 16'h8348;
        src96 <= 16'he31e;
        src97 <= 16'h3752;
        src98 <= 16'hc194;
        src99 <= 16'h3ac5;
        src100 <= 16'hb8d4;
        src101 <= 16'h1b8d;
        src102 <= 16'h37c8;
        src103 <= 16'h437f;
        src104 <= 16'h1dcf;
        src105 <= 16'h2228;
        src106 <= 16'hcf93;
        src107 <= 16'hca7;
        src108 <= 16'h3ea4;
        src109 <= 16'h1971;
        src110 <= 16'h6853;
        src111 <= 16'h5574;
        src112 <= 16'hd949;
        src113 <= 16'h4d50;
        src114 <= 16'hee1d;
        src115 <= 16'hf68e;
        src116 <= 16'hb865;
        src117 <= 16'hf7e3;
        src118 <= 16'hdaab;
        src119 <= 16'he37;
        src120 <= 16'h751b;
        src121 <= 16'hdd60;
        src122 <= 16'hd21c;
        src123 <= 16'hbd7e;
        src124 <= 16'ha2c6;
        src125 <= 16'hb4ff;
        src126 <= 16'h140f;
        src127 <= 16'h3fc2;
        exp <= 23'h41c868;
        #1
        $finish;
    end
endmodule

