module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [16:0] src18;
    reg [15:0] src19;
    reg [14:0] src20;
    reg [13:0] src21;
    reg [12:0] src22;
    reg [11:0] src23;
    reg [10:0] src24;
    reg [9:0] src25;
    reg [8:0] src26;
    reg [7:0] src27;
    reg [6:0] src28;
    reg [5:0] src29;
    reg [4:0] src30;
    reg [3:0] src31;
    reg [2:0] src32;
    reg [1:0] src33;
    reg [0:0] src34;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [35:0] srcsum;
    wire [35:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3])<<31) + ((src32[0] + src32[1] + src32[2])<<32) + ((src33[0] + src33[1])<<33) + ((src34[0])<<34);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6602093003adf0bc19fbbff911d53bfba78dacfe9c8ecb53f4e5b19355e349feabfd2c2f43dbb6d0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2702fcb2db6ffcde1b3154b26921900505577f097a8888276dc61b0fd8af91d8d3669bf96370c87e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6861b7d044de2303dbf5fbc6a6b4fa04a168d4a51d7f1977ec4a3f7387570eab535d6e4f9efdd4e3a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f3eb88446eb101fa0fcaf1cb3c7226c1a753622750833efb2899fab0dc7c5f16cdcf90d59b15e7f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd626dd512b03ba553e00b2fdbaf964a78b1ac0527608215aa39f041014ff501ac2e3c1806105f6e88;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d2d6ec44c8c48a28ff7ce9edf49f45d950f1273b203a1a87ead9b03493c8f00db2611dcbbe94522d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52c97e2c19fa4d44cd5650aeb4cd95d066c63fb0ca1db7491593808d6635a5747644dc505b660465e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h769851591a8fe2b13375d7ca03e56edb897b29de37ad2a065d5322294990ea734dc9b986bd7d79890;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71101550c76125770fef2313e257263ce264ade42f3963071ac805f39edd94d02b65bbf76bc90eb68;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8c5da82103cb84b740f2c81ed65439f5edd9921be5cb559cbde7272ac2bbd5c3e7b386e908c93ed3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d7238954c7cfc10d9c0af5a17ba79ad5247a1c6529950d5c974d691a054ae469234f5162d178fd25;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6dd4a94223af3d09e8417c8a61adcd487695eb1488ee0a4101498dc28cef3d1d5cfaa23519606d399;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0eaae82619509941e831fd4455d989ef7c35554beb13d0b8fbf6e37b26657777c7e432f07142874e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf478e53d652b21f21667d0b2cd53791690344db4bf1b2e2fcc337f48cabfb92fd31ceb2de08118838;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80f402d26d26b1433bcd685df0d9f83b4ba843f607c961bc2160b79468932ab002f0fd24b9ac4fb80;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha9ba176b17f361a71c58436a8f88ac574e219798420ceb36c99a2abf86733a01c0309021f0bb795de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he462b61a24f0e613828c73599a1e6fb0efc5241a665e1a675fbe4ecbc798b35e4f0822f773a75286f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b6c31ef81cbe6d6acc70d5f451b6edd1f980092e52582569839e040a87becb89f8d3f9e59d00759c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3379cc6052326b91493a2d2d797767d34d62c9e5614288dd73a8157eb790eb132067a21064feb03d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc6b07715ca08e9e6a3a13b2bcbab8346f34f1dbb15d1a0243383944c02359546e89e9d6244fde3d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5dd15ba108b82ae6c32a7da2ba9c2e36488d316b438df04ca1529b9152e573b4d7d46952c5622ebb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ccb9a8a7c4932932c8ae4432a64324a579a7ad87a29870db916761c07506df03227c4f63f32a6993;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10145b26670ade00a75fc0ed1f6b627a6d3005025ab0593028ca07207fc552d50a9ff669bfa8b3e98;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8011a666d69ed17abf7a50686066a72de18ad9ec0339cdc1502cfbf4de979a861da14ca1fe79f33d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd176bc1546fc841214aa2f9c7d2eb3bf95cdc269025f043ac577d9772c445a83a9a9ba24ffba43ff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34124d28920280e8a55d82864704a678a5a27c06fef2f8353e982d5d1be96bf8a0caf962f317817aa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48ee1cdde68885a018d7f738caa5ebbe9dd09b67be72a53934df1b1d73ce0f741f1363078838f209f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habdefd297b6c902d18cf2c8d514f472205fb11fba2d49696bbcd61c79fd02cac3d97d086723264ff8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcea9c7b4c37eeaffd1bc3babfc6b9fc359530467fb22d89308ca954fb219e659d9ee238a4c436ddb7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82af10a1f99854e019b69180dbd4d843b04a8141e9f200b0a7ce4e717c92a54fd51a17f7329545ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77522dd57cbeb75fff905b673049852bdbc8a614eec3864bd0b47aebb9c24c5ab04c842516fd48f9c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b9731fd9114fd5ac3c8afcc7ab5a9c8d14f1015bbccbbc2dd5f0dbac974063dc9b232b2552e6a4ab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42bbbf830ac907d2ab5b9a6307cde8864fd93b56618862d57224564260bee8ed6d5272b0a9a049ce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19860c3d0883aca1404ee2489acd3f1bd95d5a7d10d7d22ea73be7ef06690c8925cfac0c8938d212c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h205847415be69c870658786b34e0ca1846650ad9196c3489b787f7137f2a2eb8a44e865bbb62cef04;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h277b71c3805913f496b744e2c00c6f79f3336279a1e75451d0d1caebb5b4ca872183e306866934f0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce1ec447e357ae1f7568348fbc2e2ccf6dd8c15f7a6efa160b55c64b5e4787a81eaab0c0f392b9d5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0f07fc0d77b0354c58499a324afd3b683f1727ed1ae38068a3120f9f7e1302e603f9ab4d73e3cfae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf04b8bbf336e67a6fbbf69f880533f902e65c3d6966689ff4e6464ecdc4597606a3a20543159d186;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6ba8e31e867e8d8a52cb81047b530a4c413e6598421ed5592f92efb69cc13462b91a1beff0b364dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bd58695b052ea357950ee79267989d4aaf65903289c1d893627b1b8fab2f09b2530f5d897e29584a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f0352dd46aff418d065ed3c9157cbe5b0667b69b30423f05a5afadec230bd8d7091acaf1395808d1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he92697823a411361117aed002c11f3b0ca42833705230b1cb23c895fc33d802d637bfd7ebe8df0031;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b1940f04aaebf719aa6247ee81d9a7a1b5617799ca316e5d7944541270e87db2f5d44314ff72520f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53af1d88e7e23e9841f5ae5def7b77f183d01ca20dd12f513a2c995fd311aaa3abd085dd7209f0e83;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f1f94b8b8877d85b4504cdfe9c2c13d2a804018ab4b165ad6f393d606a4bdf9e46bd9693108cf349;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb33fc253ca6c0fc3b8aa06ebe1702bea09b0526a915dc425930104708be974dd0c625e0709c8ccfa6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e43068ba5df4905b54bfbf7b0ceafbfe2aa23a0a57217ecafddf13c7177a8e945403f3d685b4f973;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b2e2331083f55e020cddcded1d7aae8f7f3ed7e76b90b9f2b33d9c4eda4fd263a5034a5f24bf4bea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d76074e1cf177dd0bd853bb2ff00b5ff6b911b4ae945e695a7823c2ae5d65391eac9625f46a86ea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87fa4b7edf069374a62b8f52c03796722eab1a67862f04bf5af64142d5c315e7345e91f676f464154;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8cf2d9f43b2826ea6ad7a95dd30f0b85e82c20d3c01bfeebcd47f884725d5b58e566a932cb5fe87e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf9dd3c9f957d580640848542f784c30f7c16fc59be33550ef99379a131d4f2faf99528de6f48b96c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8aacdff1eda9448097c88844d11cdb6acaf5cb9d6f6156fabe308ba29d811e26a8c602e1f9f5e074;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d7d306bd450c488cafddb06dc01ba7e0360a5765c7be9393491f23a543d81943a7d02e57943bc710;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc88537a7309afd8ebe76d17fd45c6b7e89cbe483507603b6b0fb6a6b9bb9bb40f880660f48a0d5c7d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6b317f768fbaf4b8dabe5a27fb185675da6c7d47470046b3b6f13b0cd46499cce4f611d1ace40b68;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc618a700acb2708a70b6d326af7a4bb06e5cf477df99d723bc2352028d2724d219c525b1546727611;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd47b44b5f318915ae6330aeac930ca8bb3c110eb5ca1eabfb8e4eb91340f8cc1a363b8e970edf2dbd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa15dfb51e5313079f44c0bf9b591fdc18a317419465654f33729003874bd866447506b04cffd5a78;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7400d54c0d99e7ad6dc29cc47ea1f47e97498bbe3db0249d86c6f4a05b0a67039a6f06cbfadb8bb70;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h659c21fd7bb4097e63a58db83ec69b245c6949b45d6159b114b3b8115838aaa1a674a6d5471fc47e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc881d4a49f2983d2734281a7df7bab7a4edafe08b96a506103438fb5351cb68bc69d09a7f9c394fe5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde416e41f44733af9da1f131f2eae193c7416b1bac6c7511d804b8045d29e5e7384b6a5a7e6f1a77a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe63537944f507f8d890790ac710ebd76b2bc0f5c12da80b90c53ef080a2d480d04ac6816f250d7f9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h688bea3d4209c2dcb919a8e3fbcebe953abf9cb83c87f599cd6ce4f4ab35ea9aa04f2cf45f2283e67;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f14a16ff81d353a08f7d670cf003360e5e12666f17e72d89f7029e2bf5de62dd146c74c7635dc42b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a84ab37d2df48d6b7ddfc05315771c432cb7067f053ad1b2e2917bbbeca0fa0f49f0278265fc6fec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h642d56f14e5b50728dd0117528e28ecd69f3f03d722a1ef53ed2725e2003b382a6517c9e89280ce14;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7eceefbf8b5b7213ddbb738020f0d7e5dc513435e6d610e367e2331ea55d0cdfcd221e2dd43b9cdc1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6af7a6b73c31531c4b1d9438653474e33fa9b955c9bb71f77f11399d8faf86a76829ed0ea678b7258;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81f7e738dd77869f1cc2600f61296a8d2460233e5cf1579242e3b7c04e21d6bbf3ea244da5ed00f74;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f0f9f082605a69d5b192a95a7acba86f7fe7ad63f5f8f1aa43eec5b90a5aa582ac8bc1ac1e87d59c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85ab20e62fdf49814cbf942956741fcc08ac136f7161191b927e71d96a984af97c17f819322924d5b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7d3a7beb0e3a67e1061b97312dce06e3a2d72244a7f0f9905b055dbf319ec406e3fcc7d0a86ab882;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34c8b46880b1eaeb326274100bee1a6655da051edd3a42c565f3a99abb255efe486600268ceb0a905;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd19072f794c854f6389e2e8da9d75e127f5b36a569ddc6db500d1a50371182ff4e0c7da62002425eb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb9c82473ecab35bf260f425db468474152d0622b7ee517f54abcd9afba673f402bb69da49a041490;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha77fd58baeaf69bb9bfe5cc778941dafc2c716654968e40c8d009ea3b151526dbaa3cc0e382109096;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0571fb0069abfcb3c48193d02f1b8a8b6a39798c64ec7e1cc0aebe9f7e77d73385316d6ed02d3ccc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc12030bdfde2b03723c12c9b5380c74a1229c9bb7aa1a8b530bf18714d6f906c8e761cb009fa7304e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30c5c86e87d2c81982663ed35571426aab1e0135ff791b775c60ce98ba443727bc059b0e5a9fd250;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a20d2efc73fc7aba8a1f8878401423ed69a7f80ab78799d539f4c51079b589ee46661b701aaff016;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4ae068e0b8616994e4399ac914df5c08bb8893cf63ca6c8ad93c00593840892a771ef1f9944b8227;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d805486a20ff95b6ff9fc1d87a292c14579c8732acda0b48afd33f717364c99248914c7a6927677e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7885f1041bc64f6987a2669f2e91399202f2762a2f46bedaf77eb3d8b586612c8bc852e6990f8490;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7750d8bf9c7fd46fe58350f1ef966ea80fd1cf0f5c4d9671b4d38cebeae4d759fb32c571566f05b00;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9302068580a1399b1a4a46b9a3efe5cdfffba0372019e520f6af53a9c66cbaac9158491079603413e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h533db76de6bd866fd57ccc49e2ec3661c2bcbb9a8b210a16994dc6792a7f95d99cd802c4b98bd9bc2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h727f9c81a365419cd2acde7edd44d5479fc6e2bdc9421a98dfae0ca12cc899679220f621cd18a4ce4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29be843e80b2ddd01de932f1611d7ebcea38d0d2ecc8f9b9e637526659d03698cc88a2bba6c5d5ec3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7edd54204137f3b6ed53005c7cfe39be4dbac1967423a5bb9c89746172b072dcd29c0bd8560ad0b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7457753b5585d2fc67fb8af864b789fefe71ac88e508bccd06274ac292776654084b7c788c3b7d5fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97bec5023486f427f3a73c40158aebf2e48cbe410c0e4553f0a1f85679d9f0772d9a01bff755cdae5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8a1a5afd0426af7605faebc460e174d2896a5046d481d0b9bee1934641986c370fdc80d82f037f62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93ff409e1778c31cce01739ff473a9f6b7fd3ba835b23f5a9895b036319418e67f4ae7a24f7bc4c6d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7172b26aa583a472dfed050b25e4e37593ce97924e7c3626a0983ed354fa0d31eb5c03e086e48c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7cf2b80dbf9981d8c90bf6b3bd3e2a8bee5e9572b47452e62c6895204957b0f48fbde37ba9f71b37f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a08cd88730d94ac37d217b1a74a29de7cd4aa8460b895565cf8052d6be44707aa6e99bf0fc54f42b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea6c7e7967d1b8e133f6710aaefca00b2d080c57a1cc63335839870d14c24dc5c4cb538094c082cc1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c7b91fc5e08ee64a124599fb253c3e94938306cd452a8a390edaf829560c672655d4e961e78cc3dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb55f36df9832a00226c84b95a3799306785a5e671f651e4c99f9de63942cf368aa9665e44270687;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e664b09858a75cfcdd723b6270c2d8302ad17d6f34638c8c8416131bd2c48e4f9759ae6884fa3d97;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71e88e4748126d919522dc22e161577c0738ba5ea0f3de8806f46ef8602c4e67bb81d227403acb060;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c5f5115c2bd64ac4bcaa36c428b5b2a409bcaca08c182e98d966c425aaa4845a98809a65a5a980de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb589ae09f34c19fc7458f5b83807f41a43c364c64e8654ad8523238ada827f16290afcf0f30d74dd3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf551989197ba0bb191dee29e06a842f25cf694a502abe6b5120ce6e61706d5c768f77c926acad4720;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h780d4671f70fc8fb268f81c895b9463d99aaf1d00e3104818310b02ba6452839a5f9d2edaeb98e6ea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8fe4f9bf65b413fee72e7be62cc522669606e13d271035b878db3ba0e3f6bab8b72de5eddb5300e85;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2c7ddba454ade0f29b7e7eb434cbf0e94adb5fea59d7ea4b3b2080453987e7f6f1fd03bfb1f1186e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h744773927ddc2385ac7be75b856d1cca3152ffe0f4cd4a60ac285cda0574c6a4714db5bf1b5640221;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88fa55013b9167d524860f7a59556b5ace3c85cd1f0db4be27405197bceeb28790340e5f2b00a1fbb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a6548d649ba70fe3a945e2afda3c946ff059a125c018796cbb86f1ad2279874c9dfb49904d2137b3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b4a870df0a2e151268f3fadf4bc40bd675616dc3b282953ce9a9e4aa2dda3f0b4f373bcd52b14175;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h535bb816ba93edf180b2e416446db35492c2c10ef15b8e214eb363bbbc71f8ed504a1a7b7a4087b61;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd25eff9d66c64c22f71d1d2369f432db33bb16c79536b6144a9bae8a69183ed7a0e6a854bbc05713d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e71bb0b14c6a384c608099beb0e8c742e31fd2ec2b6695d2c9abba8feb2f3d7156e2a90e3b617738;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha39f004415579c3bfbd8eef80aa8976f9165adc27864451f507fcda3fd33c5432433d3f6381365e00;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h444635f8acfca496230a432de7961ca6655915237a00906e2cece8e57b81e69af300c89b964d83106;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbeacb06938ae078bade7dd58a6c961578498912f02e01bd614eb0f626e5e39788111b1ed6ce99778c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ae971ee2379df3ac653cab6d5bbcc52a59a6f54fa50754b75d788a52823ade8fea10d15c3fde2b00;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d1d2aa3068f75839f56eb623790aea14a292a24986cd30a9ba24b64381e8d567d1aba57ec3a076b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf15791c5d19ec078f6edfe3f0a94792a82a4fb1be439118be9cdd2aa8b3cfedb644c81c6aaae5becd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf19668a1714b63f5a58d7129ca0d79f2811e357a482247647393ff7217c924a303d6bad71e50a9342;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1fe861e3ad66de21b415b77dea65bbc35665f8bb1e642b2f3792da18962bff31260841e31fd4d72f0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6021d58cdf08c2535ac6b8f78d122b36c9046dfd4456db13261f5cd6252fb594ea1ddfdc1f9435eb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf3b49a1d874e3ddae612507352a8e52ed57d622def1ded7515bca4360a408bc50831fae63c9aa20e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38478f1782f0370704fa99c649cb210ffc8d7c83f8358eb5196c3815f8567c821c39937ddfc7244bd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f228a307267b3dd8df1eb77c0fd9db4bb671db4371b99a491c11959bb53297478c7299a72c0e5f5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b5bcd4672cbff6f4d6a43b4aa61664dd9aa4b13603919d1014dc60a804bc687031183b8f3acd2782;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b4be87d558b02066f4b0f277d2548b080e614ce003818ea2019958113fb14aa247761e579c0863e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94396c5aed45967acc1e14821b0b561afbf69447c0d8b6f3bc15286c2aaf17f468c6a0c1caf4885fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b19c878e2afaf5f7146a3f1f72d0dcfc5a2ebcc6354e7e260eb711c10b5418c253702de930bfd801;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7e637475ded0c9c26a63e518bb6bbb35d8fba1ee28ed87f7668dd17ffc1f8ea778096f8cb1ed10d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he03f058cf12a5e04c67f91b4f02757a70a668cb70ed863190a652a61b873fb726ced0df5e17c7370f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f2ffd0253fba5c1bfe622fd7d43d2c2d3582ef8c50301b4029c6e1bb99ab30180f0eb1e20eb493c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h575343c67c7d41e15257a8b376bb6c35841cb2260725efb2f9459fa6d3300cc43d9c165f0481e9cee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10360a268f9eb5621e7db1983149bfa4b7b8d56183720396d8b246fe56c2270d90c6c80fa9f47db09;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d02e3e8f7df3791229581a339cbb61163c026c40e686530baf4e7040add5195a603d5a9505b17648;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3ad01858ba0fd5254806e2583bfc2fcd03ef0df279d58795a52bf048483af999fea9ad7c5d979b3c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd956a716e6f2efa0d3155f34ec87cc557b6fb8b2d902fefc28f9e16baa840f6da16c852195527c602;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h25fa566d9f9e794c217ff334310f7939f59cc814df9755572a6b3d38330529d7d5d959035c2b0986c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7a7832f6119d1b9cae117d993da0be2e46703e3f1c464023724be31052d95b6fd06a9153d886ff7c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ac963e09ca1440d8db481047113c64a9152573cdc9dfa7c43ac6a2e42b8e5cb110689340cba2b93b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6816deb97ad717e5c865b073cf83a577506614dd58ecb058ae972833a4b363b24e84bc50acad418c7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2d6c835b075a11a6acda0827baab459e96a19da0458dfb156b485f9aadaf0a0910112a8f018ff6f5c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6034c9ce2aa36107ee9ee8738ac78856f5bf7395155b01366f824629549da675c97dbd95bb841f26;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5060e000fcfdaa0e4364712ce5e344c0eeb089646bb13d4fcc3913f800c4db7f53548a853a7f53b3c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde0141f3c3f8e6a595a23c8d98771aa163116f5db8be04690fa39b11aa490afb7121bed8df365dfc9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc23e3fca1f4d9226a631ba332bbdcd8701e233326335fa55c50a655dd9c7c59856b20419b16e2ac69;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39d48329f151d29141300653946c701f8d926baa317282b1891fcba2918c6afa72b298da32688c3e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f15110d69c079bace51743dc1fd3c54558524834e068c393f94c513344670b2b830b9b0768dd4ae5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b8b71153d874a76c9638e1948fc3554e0eb6f55fb877ba2e6a776a826127421b1e61d278dfa53845;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7e0ba724dbbc203838ea3c43e2dd3d81e829ac533d3febb98670cbf3c6624c557f0d1210d41360a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h745ab8e6ddb3e1cdec0c921c3cdbccd052988ce489ab67f5bf6f075fa17a9b566b4a86acd87e69229;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbac3baa5b144cc01f4d5f4cb505acbe8a2f81d764766023eb1f675e6b0565fbd90229a2e695c46652;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3fdb089127dcefaf320131d21d445466bd47175fa1b53ca62539106298c52b3308a842dfab849d7b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c504e5c869dc03f745b9d2e7e9a878c1663d904cab89d208d6369a16d41fbfcdae43fd0a15be7eb0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h827cafbe255c38bfd3354bb46b7bf903920622d7d39a13a7f35c78d7c1cc06f6c97373ff9971287ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8935b503f13029309c356752d588e5f2b6a84609cdeb078857fd2493d69a7716845659e5613645f49;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda77432de40da476b05373f8a16b65310e6318c1ebc7bb6c50e1d475a3535bf86f4e9a846ed942d3e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec41b309bf024d43ee52d60ccd5899c52ae6133771cce7ad41337f5b03337bc3458ca9d74b2ade78f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h540da05d957f4137d29c6d48b057c4a9ea3cf0b77180d212198544b43cbf96a04958b7ba6cbba5b64;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41b40a61d14586603ce4dec88c59f9003222f903342e1fe8d2ea082c16913bee6a6b5d1bafb62a032;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea5532f8a17c1bae264a1835e7e78290f185165f99c7c2f11ace0db0dc6a54719f3ccccf03261134b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6465c266abcbc8d92ad3ef2c008199840ae99c4d2474bf9f0eb539e22d2f678be8b14c1c9671bad8a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6966e098b3e2add8687596331209d8dfc6fedbe3c5dbb95ae748fabc8240e9589613758499c90f879;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ad6105167384945567dd1ed408da302f52b0d2431002cf54f3fd51106580783c51d7ae57bc45a213;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf42491166c2b5f797ca7bcf258021b3c849db44938987d5641ab86302229c7fed1234a2326b6afb7b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbedb7a9de385973279c8e3a3d574f069c34e0f69981dd5db7da2d5427fa850667c0c4827cebc815e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19e5eb9fd1f2720a141ea9d40fd6ea37dec453bb4a9aad12619531ae6b1fbc356ff903d2616ef9271;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he993d67c9b2bcb6a3e0a1d199ed37fbbe834cc0e14575b947a06254b4e0bda7aa6dad2cc0ca860d31;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6e8378d9eb750f226e55f541c699fc2c1375049e7f0a5565380ff794cd2e70700d4424f424b35dd6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22e6063961065cd757ff0121689ec5376913becd59e981dd07e35a26d4f4dacf082028aad0809bbfe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1ce57493c2db19dec39340c8dadbfdfbc86d3af118f6bf5b5c3bd67f86c91e00100b38fe0d14b11b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h832a53c44b43b59efc72343ffe2e0fbefb496594e73246753f62027447b79582211b5a412f8f7854f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9921aeca56724805c06ef2e63632499f0b62b3be576b9bc444188dee28b72dc76678944f0bcb0ab01;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6aa509df05ac664531b04e195e462397c394d26fc9feb2936eee9c0407cab2c61304097ef42ce712;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8288ce2820fcd0dc0c3f32790c5ff5d86470a39c6a7e952d9e468f0db9a35460ee86f4e7a7e79d247;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd60b1c0201e4aa47ce69f66f68d5ba31d6e086184036e98254b856f3d03d8f4d26f2da834f710e919;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdffe5b0f338c8a5a5f747a407888e0ea28b40e8a9d46159435d3df460b5eb84a218ef549063f07d6d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h731a9feccd5f2cdff6d928f53c8691425ab34c3c052d432104117eef88c0ea57d597438c9285783ac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h178d4fcfde0a11f0b8c9e7a18f0b71faeceaa5b623b8c8ea5eaf914e7443eda68abb16fe0555777e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f1d1a8c788031b4c044ac20fd9cb29ce8fdc74b0cb78f61a74297f89c32d3becee144842ed060285;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd84f8984cee066ecd526bb0c0d89d5e2af58ba3cc913a61e731fc7fb9edd34adf752203b6d4901fc5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a6841c8b468e39175fe4dbefc4037ca4b07fe5924f3e9ae204ea508a9bc3a030b0d6c243528e3282;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9335a347dade84b522fb965c770de317bfdda5214872ad73aba1c710dc371feb27de3806b601cfe7e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h753442bd6b7cb6bc99632beb4e9b9cbfff52e0f1bce69186ac03600b58ac3e7d2b343a738fc03044f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc128aa988f503e6f1cdc6052b2d7673becb5e985b313aa536bdbd6caea5360167e21228b1c8d59c2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88baff7e15ca6f185b779a0960cde7b13cc16b1a0a5869edbc23f8667b45b687a30c1655c3467b2cf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9701b69191b568ca6ba01e566aa14fbd4c77f4192f22051606ce68e28e05313348ca832dead7cd923;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9314c0119d91aa43946a6f2795ba19c33e09a0f24f320c9b199a0e45481682ac57a9bbfdf2492fd52;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb356d5303fb39b620c820b3eda8340c2d11df3a6fbb0208d2f51fc319939deff63e1263c2c5c98545;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd54c922b206438c204c2f8ec99a80da6c36e4d88738e6c557b90717f11890089c7e60fe0e2bcd141;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9869c68a64ea6e09c37045d93c49f14a1acfd6f76e77c5a552e329a4943eefc85aabafe5ccfa910c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf623ff0bcbc650f33aa30a63693548b85af65db192e0544a46dd42fb058bda381e08a0680755eb938;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7a0cea0b4b5ea511233595eb94d989889ca7516c58234e3dfe4b193327ad7b077f00444da9e8f414;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h287799be458856a718c816d2d5ad9949fd1b8e2dd84a973ecfbd470e27aa5b70baeb45d3b1cc6b8a2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce8fdf457fa4ea6452bdabb89c9666929c3ab00736b678fc437b3459d55e1578f8f0df3e3195742d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4abf3dfc0513c8b72917f8a8bfd9dd150663a352f4f0aeaa58c6020e08b91f3118d97e7d7baf608c0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha84e550de50d77b701ee2ae812208e399e18bfc3e043970e0de3cd8e96f43ce00e90028099a53f3cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e47a23f9c4dee6e2b5139edce3e2481cc8495fb8721e8482a5bbf5abeb1a6dd21795c549f2c9a880;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88d22c777c27748a7ec77387c9eca3bdb53a2dcd42baa55e1b424865c0f7ad59f487665437e5d9ca3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc65f3189657c7e701028e73533c89f2ce2e0e605c58302354673d331600c37fd6630b131e0f96f005;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89363eeb636007a0c094e6dded835edb49b2ab062df1864690fd0fb3a554dc806022c3bcce9dcf9b6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf5b22071bc3ee492dde43d0f3f661b2b14a903630d61e73b920f331fd3beec1efcb848af2b0c2629c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30f9f55c3ce898e21fd9e87128f28e002c1c34ab5ebdaf4553a0ea29261894b963f6de2bc38c576fe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1d412c6e10b14dfabf302e40b8b30de7bdfa908c30e003308fe2f48ee0ab9897e317e3dbaff0c639;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h938d070985e798978aeb8062b4b6b11a19b96d00ee18f98f0d0df4c9f71e867c63bebbff7b03203f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6ce25a2be4b0fc60a62588ceb15647736147b5bb5ba9729b30204a51378ebb58a681a2f59d6260ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcfeea1e8baedbfc441a092cb35d4e62c149d8612715fb94090a274434aa37a4a6e7820408708aa9c9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2df995b0d066f45fc1d1c6a92d32d306e75ac54e20b5bbe68cc46c5a4987ce93e225bf70ed690f40b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdebe34f9bb0e1e17a586254cbaaa45a1557d1ca26befdb1972718f78a32389f2cc9b11413519d2439;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2317e837a88fe65de3b7596a04026bf0d2c301ae6ca7430ed9c05d386052c1b24e28efae0bb330266;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f5eb8ac40b1ef21914c1106b96f826c015bed0c9c25821ad3d90f63411a3bb9b6685e262db1aaae4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefe697a024d6b32fcbdc79510ac5e6074ab0af70256da22247c0fe27b54a72edc6ce606ff8583053c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbeb36af5be55fbcfc687bf49632781dfac64fb1cfb35e64254bd67a198a8b86d7d21bc708d6259f7f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f82d5520e277137bb57edb9e12b436cce8323c65e675a76b06c498f91b04fbff3ccdd72cd05ea24d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6142e37d3d7ce51b4609b66e25e378f4a11b54f780f726a20906e192fa3ef8a7cc271141004932ba1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha18afc985863da7a25224b29d269aa4e2c9ec4b7d554a5f8e465944344b08e0a8d6a453221d0f7cac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27a0acf567a81859434b64067b26169d2cacc5e7af5022875a5b77e813549bce2f0e79bd07d97880d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b3de78a8d7575d408d6ce88a42e81d42d0eb9b63406af26a2719e014085e3d780007a7763b3dd637;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fe839a2487feda23e156b61ad95ac1f72666dbc579f737b8f5db79d9ab47c7a107ee14719f57f656;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he23886206fa2cf607794fab0a8e258aeaa90c6ee770034bc84a0e70dbd8f882b3767e6793815cc946;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h325c61d6e5fcae4881bdcff6955fd77ea29ca0c70d838a3c1aac08a31ec1cead9c603875b8654c4c7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'head74238b95237261c8c9eab682ea8371d7ca0d09a47aae64fa38afd2524c98140a4cd72763b08f4d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b2ed5d33bf4f4ffbd0fd5fabbecedc6a29aa361d85edc301cdadef56a456add9de8d2897028021f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b39e4917009eb6ba5db666fe771f2643e03d4e1cfbeec595de57c32bc118b9251a26f27b25a4a891;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbdb8293fdede1ca936506a3f1faddf1ab6f7eea27fd25948d4ac71a287fe2d7fbba395ef7371cf739;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3de3a691ff3994f2af3ca1e6e70c60148f3fd4d1d3f143dc8309f5bd345344b6346723b72093021e0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe77cd361ca656a57f41d4b6e4f9ca714a30b016306ee5ff7eecae6498e26e13586abf8053c1e549e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1159a78562ab61436a362fe7dc68c48aed5a9a19574bdaf495f4204c8a6a6f0d3b25a949ec453027;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h220c46c4c85a13282377e1d9b5082a8fb39c15743c94046031a42fe5968c9994642f474fc710a5590;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e091c67c871da90a36d0051e1cc722c0bdbc72c293170dd20c5e3d582f35faa05285920ef44bf946;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf83c42c31bce0e4a524bfcbdf3c2e3fa477ded5015ab595690737d5eed82e5bc5da56de1394341d54;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81d44ce807eb8b6acd1d0630e407c987617a8ce238fd357679a297cc5d88b68945ed94cf8097951ad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha88f59be0b020f91523df73f535b59fad65df7280b87b1e823170cc77b105b28e7db8ca5f3cc013a4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16d6109c2ab05143d7f0dcc2a49f78822b27735b5eb371b299facef2062547d58e6dd024c8de66d6c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0955d4a719cfb9145f4d1f13dc2bf0fa96069ceb5522772c0959c72cd4e600590802a199f86e816f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf018f70047ea6b4a978da9d7147530f776197831984e000ca72c2ca30467860ea861243e0fffe6cc4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac9aaf88142539d88b24ef43f8c101224706202e2b6df6df10ee15b79edf125f4fe6e50aa8e539c98;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87329bc6f9109ceae16a0cf92a42fea460ebd84ecfd5a52d7ecd70a7069ae458840af7fffc98da22;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc76a191cbcd3b26e9bd4032b40663333c22a13cfdb426a4268351f05470c5b76501ba7e1d69eb506;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h959031e86355e2e715989d649fe9e6e78f3c60e83593e2fac16a108b3b60a2219d55f7b0b5743b00d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe31a29a93d9b859377401a76614404c08e645c17476d207f62e4b1aecad233ab04211cdb5bab0624;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe0820a0d2e5dda28123b335ff8ba853feed950d22374d66bea5e69e569090b9fda8f534c5fc9f053;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4ec3ac99a2df3d550a401a77567592d889a946e29d7fcb789267e1f207606721a4c9acf8bb8139ce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7af3bf9b55322974a5ad26350d6ab84c84f5bdf092bd254cdd32b2afc38e78573ad26a9f63aafc29;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a25ea92fa86ed77fee0d1743a5084d8c16d86f7c2e10e09f752491c88bdfe7e32b79ad916dcf57c3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf85348373e59752c3e2f3d2d23960a2244a1743fd3fd5fb865b8a3a16d4e529a452b65a37a1dd1f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43c0f5ae7c6fd92afdbc5e0b778ab6c3a7c8f2bc0c9e08ae0452a1d3c2843e2df347c246034532a32;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h140c70da8462a81d435362b6c1cb9c56c44ece9457fe50645da975610138d7487639ba38cf52a91e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91c38715083340a9afc1d71ea82624244c73b35c4fcaa3c1d7c0ad28c3a0364170196104d3a90af63;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99828b092f5d4fc5b9f9587caa83ac1e421b3b8dfcb5a586aedda44d41b04173db6f3140c09e39695;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcfffc0c15e117e5a9cf1a6fae7d4711bea5f63c908184b99bc57ae9aa9e7c8e8497bc0c66b545a084;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha56920276ae514d416240693f8ed7f559f7850aab9457cd9aa69a8b7daab277a6035172c73a2c1a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha27d370477d454e0cd00c8c82f9ae14db96353a355293bab672d9b108a03d0064c51d80a0bf95bf16;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16bd5637ebf43c0c03087601364589a571120f435b3cd1bd4ba8b22835320d0e385463a04f5b64fbc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3189da71b140e2e1ca5305e03ad9f857be3dc3b267e2ba0cff36b9d5ba12526c7a2511eb057dd1bac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28dc56110db8280d053028484188fb35a5a2e3577e030a83d56bbca13cde9eac9c3967a44dcb1dfdb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ed743baa43d7ddf5e6ea6b869b36db5d26c41f977439639f276316857fbf2268655c5d3e872e46a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ddafc34b231c685a5f8a36c1af346403610a10f23a70dfd33d442b70f97dd699e84ae0477288c8ea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h927624109e0c71b50d7e2b2971f9bded13d92323ef413d39cd0f4d5b8fc15cab5754e4ab093296559;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14b78a0d2fb47f33af27a250f944eb1066462225a8e87999a6288040a748e9c2722c015a0f427d92b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79e1c8893a9daaafe074b78e27815e7a126b3e0a64e8d4ca5f0dc000f05663c03c58d8d00d8a76b00;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h222931a66c6eaf70ce98e140ce5f1fa9990813922d9b00f90a17fc48ebf0e553120208417ee0d5005;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf357926bf833db13e3d5cf02aa3aef34f242869f40db448e5fd8d56e12e58ea1a4571ae85f2f9f9a4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h600ac11cc3ddb6b7e62bb01d97cb090f7eb12f11d203cc71aeebcb106bc2dd9ddebb3a3699449108c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5c1b7e42666a559b4aee5d81ff7a071549789182840acaee2d9e4c20ddf145de98cb194d50192eb1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a80154820b726aa7c433b7a385dd2e7af920918491711ab4568baa79a760507ab119bb9faf9667b8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24e707244ae557c5eb84b0d77a85a584da8dd6bf4faedd37c9cb11b933e863d40b1b2f42c1a9a4691;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h312f12e7c858e92194a60de4b83208bfc794577b6a5ec318fb4c853abae317697e6acf5b1a10bee3a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3768d2ee9896051aeeaf4fe60a37e6635e0eac9b87e4ffba756ec95b266c9d88e70e3fe44442527a0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h661e1cc32ce0230b7e1a229f17eef0772d30793406946837a65d48e1651927426746d63b091745322;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5d9e2b68990fe07b684cc780a73f1dfd12d9de4cd1ff30e5f4f41099ad462194f1c787cd8fcc43c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h215feeea799d6d117742ecc574d5b50226356c09b2a12919d0612c1f2f5d50f317788615f7bea1391;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15bc7a344848dbc75eff11bfbfe1414cbf0ec6c31ecbe26f47c109d4ebce3060bcc156f6588a2e8e0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7425953a81e15c6bcc8802a7a223f460e0b2ab3f1db78eb9c794868409a5e08b83398be520862dee8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43c1602b260cccd3029ff167b75c9eb7a2cab620f49b7f87e730e8e577af2b2cdc401a55e90f3ebd7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1bbc0892466dd3494200b001078ce848f3409f41899e16e405a7631a09bfde866ffdbca4e2caa4530;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d7ac11d8bdf1c5562b3565f4c6afcfa251280ec985dbf9bfb44cb3f78e01b567dd85e8720733e83a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed0cd571e0a501b6344c049aa2bd121bc20f24af80defe605352234abce49c9f19d5d7bb88eede937;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h576cbabf7b98893f483880f1e04fd14ba2dbd1fa6b55bbaa09ac3632f3d545011de0f738d725009e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38fb078e31c168e3dec92254a7bfc9de96967aa96a4ef8427f856acd26e38435d8caeaf76fa62ecaf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37ee87e3bd451265b0bee5aaa0e770cbd863a63fd24bab75ef516333a6b6ac83a3f558d524d79acdd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f064b111441b42c6854a8b41c8b2722cb1055c1735080d95850fea3540685a3ad01444637933dd1b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haff14710a619db90933837c6bbae458111a6ad157f804bff75a63ad85b35878ed0d36396cd661a4d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb88bf977a45bc0d0d9b95c092178ae78493e1fe887ea1d2b0889eb81bb9c1b657cb714d522fe84b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a8e460b7fccca024890972ad5404ebd970e0cfe364ac374957be4f65ac78f0992e487a795fcfc87e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8953f17c48ee84cc7aaa8be9d2eb762cbee6309f6085c45a7eb0db7235f7d3de80876ec6e4fc86a40;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1fc9c525399fd23cd1d0abf001361c0767c1f5bb3196d6f045632c2a71b69c95d184cf497f34f4437;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1046110ad57c1e7cc2e1e9ae29efc12695ace604e8e9992cb95692a96b39531ba95d63cc5a5eeaef4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d1abc62588c92c6264595b710b97d6bf6e557ba9b19be64725b4ad6657358a777ac1a6fced6a6955;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4d6e81c510193f9ff553105f4e5b8e7702e66f39beba8e140748e1f69da82d8a74df9e1a1ede421e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae211f72143c5764437d6c8af0d8b0887b965057fba3da28ad2f4587aeddc75b2e3be6513c0b17903;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d9fc9035442c3fdf93877be6d980112a64b09b1820e701488c0dbe3d52a90d13355c97af37fc201e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40a041959421efb52d6c446f65c387cea15a4bf4177abeff78063042af2abda62f8126cd4510a5e62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd4c85f30709859f53f3e7ae28c3c99ad92f09c3580a00ca1e3ad67009bf22e3261c5259922003662;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9bc4fbef24f20d45826d3cd90b96f63a88c60733a9e93d8cc6bbb2f14cb7ed77e1ffcd9e589d359a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0da7505b5b7154eeae66ad3936eb666efa30979b15bd6b9d4d09e4c379d5b797657e1271e0afdfe0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74aa3d81299748f309741822794ae1997f1184e05f52d0307b2c4b35539ff6f6a3595c856892f2bcd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6676c4dc9d2a017fa76bcd6c01dd6cfe9d5521f9818d642f12248c22ec52179788600832ee994e4f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6416530d215ac6288dfc9dac820bcf2327d6bedfaca58032c2cea1c2a77d89d89f4f3b18e537a3766;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h934d9122b32b305ae97a2f40fe39cc162e8acb9cc4c71dada72ec1835207a32b2824b1359af7e1ae8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c140d9bcb6be385ee6ca8adf80cc92980e32c0f6f9b5c4fcdc6268ddc66f3427fda38c9afba962a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7760f93dac04a634e997735fd6e7ac88b69b99d2a5b239ed9e0f5f48c93c1ab9dc0b35c6b65c2431;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc89e8e970ebf82b4f95a281f268dcfaecb4930c42dc5272113e0e998801e93bdef35a4ab078517db5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd87f14eb19c6e0e63760ea0d7d3159198a63e1966c59a1f85e5db954f9da90361974ac1769369226;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f8a4a3d55b384aa7260cbe16758ffb2384a0b42831746f48e91fe010b47d380db39f0fc2b6d1f696;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h183c2fa145d919108b2af92b1246ddc865929c18cd00d720aec713065ffe276450b80cac7c1e7c96f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1b395acf8026edaa77fbf1c2a9e1ea46c19be0d46a47fc0a430ea3184816a23a76d5eea1bcfe5aaa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3702569757f5591fd2cfd0a1abb568e30bf4eaf0b1985967beb020495ad9ac951bc27d8e251013db0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86d0dd247c88b98fa30e7d8880ebcf4e18a9358b7eca6e4f52f08433c29d94ec434be62cbd3f1c2bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e741117c04f8937f474a0cb3fda8f7cf48476ccd771ff6189ad1003528483117d57b5a76cbba8ed4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe02544ccf512913fb840370c9e7d70570850ed7c868c38fb8306372c34059faac7ed5f2a7b54f1ef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14c7f6108dcaff801867176156292c2d72698ccc58ed6dd44300162dcc7fac4bd85e523f39af94096;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8b11267d0d70115b310070aef83365c77519d7012ef919671de3d737084f5ebeb971ecf6bc70501d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72d4d4bc3a225fb327153547129e879b6b2f5946b00d9817bc85c57db729ae8173bf28462b22a7181;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b6f13b80a7f282aaa96d0ff5fd779a8f9f158541ae5d1ac1de70adf4b9cc5efb2608729060e81f0f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e5db934b2d49bb1d6fca4f3177cacf427c223544412af0205d1559f5944dce793f2c52604a59ca62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf941380625c91da58b534b8c840ee116e0a0f18459887d0081e5785af91a4651905d269b8c56c545;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc06981e8993b2bb72cb9747581ca5ced9b621608b242cf758bd7ae0d86d5eb8d05bd753f3a9ad96f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcfa6523e4adf696cdf3935387144c4e85554f1403f3aecff21042407fd5ab0227f8c62d4f65cfb170;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3554cb0115d8867fda8ed367d7912949ecbd1c1119aaaf36e9a11ed8b1f39755a09372216e0a77d5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2839a24c09edb2fa266e6a8d139aa82ca0ca00275d2e6024f2be40fd53a946cb211c809408742256c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a7910e2dd69d6848b19381a6e3c81e4843c9b3461466b8bc03ebfda4f5cafb31ee44d2a6bf263c01;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd857543144489a4716a1bb9198dd99db8463c7442b180235da46d3f8b36a769ed8a22a316d5abe1b8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8bf902751e6ca69348e8ffa8b57b05c615845c24a5c3d0db13c05ffe89c251c52f15517f262ce23e6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21deb0eca21743f58766fb98ba45b3246ac8f27986ddfe719c9d431f275e3d059f8197fb5342ff909;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14262cebbd397e5540f4d142d4a4faaa903fef3daf089efa43dc6418fe93a8a3fcd7aa09122edb214;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ab8ed7082556496b1a2d3ccbed7066ad5309a6d222eea3b8b12b5b3559f72d693fa431b3aaae523e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1048ed1e043df2be42de7eae61e32713eac774ddbdce24fc32ae6baef2e8d41d156d01a1f44fbdc14;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82d7972095f0137693958affb4dde3a1227a745435335ac1ffb6a9fa8400601e0b64b046abebcbe73;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe50cb24d052249ba6774b0d5ac8d0cd9c4d706eda94d3433ceed9c5914dd6ab7ecd030e965597b6a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b7f5f96a96a23e9708e71aaffc2a9f32d9ebda739cdf693c1f595f57a2cbaeaa18aa7277e0e815c3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3da73428c55996f1c8af703e9b40200178e9fc0e004d3c30e3d060fd2b6d79c263c16d06cd34293a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91b853f02b7b11d167f534d8327816076f78348768cdbe858300cef3a37461d17447d79a96e8be660;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d20cf3994a711161e7ab60227bfb8a6095a4a849d18d9531ab5d23c65a5761430f8e283abd3a9ea3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefe51983957843887ea59a40f258cc1078112757e6ff927755c656c8c46081a90e55c4df86e7f8588;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h923d9f08b376a4f5745aebea55d4ff9d155af663f01a33a6c02a4b61127ee8d0cb8ce521527697029;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5e9bb7898baea2461f47880b2e57cffc714db97e5407b45c1759662ea8ab32a190359e5ee316bec4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24251d19d38a00fcfb4d1706bab45643fe7a8c1ae8cd05ffa2f49d06927098eb2fa6cef02e6514ba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha88864f6bfb313c3f03297db7e0217192f13733f636dcfc996ef8e904ff62ce8ef11ae276dee580cf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h351a7e089513518f8545cf18f533a36af6087cc1c8606d3e68008f40f7cb2f80820ff8abe7f9dba2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d95167f296b166616998cd356533b4bca62cffd1993deb7d810a48ea8820e0b50821a8431d2858be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8276b9fefba36e7101ce9d743faaccdeb9196491df07b63ffde434d090e70e2481cd426c5a5eedf44;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6bb5449ea0add10e2585f910f6bd45417b346ff6f16518d3c0964a3f0c64caba774d757049b4e39c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0c2f69d9edd6eec57634b59bac99bc40027a1f2b8307a475151f2bb11a4a80c4970cc25adb0bb1ba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cd2f1b2af47d6e9f48cfc1da39a606a2e5d541d66747f494eb90985d727d8a4deebad44ca34cac88;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55264ffb0b217e8ce1871247f335f576368c95aa377613860f5ac2e50ad3d85c7a72360393eb23e77;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h253b761d46fae9f8bf934a865dd21d575028b7c4367b9d559ba03531423d7e2a08304d73d9f839546;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h202c7102c958e2b4ea6a511b2e61b9aaf2071a53f31c986f117e9179abe092ac49af00ee772ab1407;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff14022a8a4a1baf7d3e64a25081046c6f65f0a78c616ce384c168609726604890b17178210662ef2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h698ba397b63fd2de0f4eb29b92e9742be1828d40956c7d71bb0d9b8ca7a456f113a5fecd4c2e357a2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19f8cf7ad384f1608d93e4c35f6723af4dc07af9b18088e6987913e96648bd2133e8a7a4274c046e3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed887cd3e14ce01089e9e78587dc86be0e95d7bd963c0f41faa6992a9fff229d7df8074e80ad01e16;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb20f2050f71d2c93b42e6260bb86e0d0142b0406c51db6bf6da76853202cccae8260ff3c3dfc8fa0a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a75a50e64e969a3a231a927c4a687e20804660db60184d70c891fa9cb9337a96f89c59c718bf6e71;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e02d8eb2cf529863ffa1ed93ac7635ddbe555a2c2c5714d4296839ce94f77d7dde66e3f8c7ad53e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h976027e255505ba2f58cfaeb8a864c133df1ef4e8a11653f69474e38736037dc899de55bb8ca8a78b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heff9ba5df7e8d64ae160cbbaf86983c1198bd239caff7d0a6b01f0291dc4d349a5638d1def9e8f271;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he124014cfd93236a2b5fe56150e71d005227ad7573dba56cf06288bf942f2bf63a4b3393259d3afa0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3305d1665f07cedf76b8a610fffdc426f2a16b5e0124dbc465f125abf33baa62773d0cced5c63668d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7085dfd95296cc65cd0d477c7a18f758f4cd7595d6c94c9a33829dc5b47e38d2ba57b8ec5a170b37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8bb976511e68533d79aef034dc7fafedc594ce440585b9a236754a18667487d45fc89bf9743e46a81;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbfdcdda91cb7ca7dbc4f9f3a15479010b13019082b4e3a55e0b4be3518185f336257e34301004a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62fe4446abac00a250c75bd42bc5584b3e9a15dd9c15fdf17a1e7f6be43ec80e22aa74f5a0c0418c6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha645a91d99d3cf82d6e5bfc02355a32f5529dce4f119d96c0362b207f86cbfc6265bda9ba5e877903;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc78ec8dac6a630931d56c4eaaa652d6e3aeaec5be912b71f230c700183062e5e0ad3692bfd46ff294;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8779b065f8d8a771f748b67fe1e790f38d92f9be084a4785804469725edf015462ffa9da7f226db;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8fc1def71fd15b226c7ab014f9bdb61fd89f17be0f2f0c1fc52d919597c0f4fc07064b13538e7587;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe1817230613fe4b6b07f8e3e1a4b136eacedaa55d6a42233578ae77b8be4f31c64e00db97e5781e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h374f7a477c85ab233dfb2fc752351d4d3a8a4ccb3b800a6571cec24cf45b0675b993560a2ea4bd46e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3290aecb3ae57bb6c3f3e6e79dc1d41604ad6d89471f35a429223bf6dcb3644f7b255215e1b39c7d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85433177d509cfc3840d6a6e056bec58ae9e6490addb5671b6a18735342681060f0640ff0bb5ca6e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3e1db07b5b239ff71fae6f968803a4117d046d8dd0a46a24102e4fcb9d71e43b6f895a2c6835e316;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0c36ef401f373f6c8a7d08227113a4a840634b1251170040cb04e0c1f5cdd7973061934c83af8b8f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9fb0c69aa5a6e03ab023843bcca20349ffa04d9e8349ef4b4c1af482c159f54aba5b7655c2b31edc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h674bfaa4c48ce676677b00798188f56fa7e8a2f65b7e2ad8e96074e1a784287e6dba8c193374154f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee1afba28eab4bdc6d9157cfc66027a0b3be89b1170ae671aa331fc336a8702b037de7990b3ec6ad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67b0322abadb7d6e925f070ecb6ae4c17ac09f9738c68f61c285943b609b68684c84208e41f9238fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f08271901725da925d71c974ed79e4289cd95ec14aae5015cd008e190a82cc964821af8fb5dcd6bf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5d1b07da3d337c830e04a41363ae3b8bf6b4ca35fe397e567f40d1cfef86f3133c10862ea2025efd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5866da1542b9ab073b105c2549a8d51624ec3c68da84863e64b905a25d69d57e9a3ddd191e3dc71a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdbc5a392f3a2bf01b9999e408f70d044ad2fadab21901f0d1d56d8a42971bf3caaecb81eb6e823be8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30ad996b9332fcbbe10d0aab54b9323ab8d6752fdb6f45dc4fdb3b05ecb8aaa6014a4a3f53223e295;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb545b47c2d5bc926f35749f6a659f22d8e4df3e513b667213be995d20b4b451f3d8f79b017ce706f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee2a61050032c9cc5e977a9477a66645a0964489b626269b08a2614031bddef9aab79590763c8ff59;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a1181e3557214c48ea1becc5b04f66ed4b19456c4282fa019d54530fad656c2782ea14742f9977a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31aaeb715fef95f96436a20fe5c786b0ce8124f19caf35094f28511d25ec82d41a16c797ccc24df59;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9293cfba9257aae47ac1be32a739f87cdcc9014b147f027dd220433caee7d9a5fad07c68d965a7033;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6fb5e06ed84994a5413075a921aab6983ae1d14559f92ce6a15d63fa7055357eaac752db16e8e944;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he97404adc481f88687af88d0d7d2f644f09083a04e5cf966ce27cd2514e6a745811c7551fa24a879c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6be5efdde2803a3aa5b1fa9722bb5b2e7a893feec63875749f70baae75f209d24a5a32bf1934b9938;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0cfbb2f51d9dc121559d04e78be657ac3d94380ecedce571196b9b7057ca5b0e1dd011b7657e070d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36b531a25f6969f577b5f68870264aea0bf2a53a74cb8e46235b481c394611fd2d893f01ff7670611;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9547e29c0169f524553a4d6a2d742af6ae4c00fc1be4141ba8c8084dfb7b92ea08f5b8f5d89ad5c54;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e9f7f4f399f924f3b6ffa355a0ab19fae9196a04585c50cfb9bf895631e811b04ee4e28bf6b0ec51;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8d13d37c900c59eec5911ca17370caff134a20db67f911072fbe2ebec09b0eb7e5f1aa60fb94ac0f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb01f584353626099ec86c22b5466292d658422a0382958b9304b4744303b6662238070c4a4fac94d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd262f437d7e18d74a05398481aa0f268cb722e1e875da2a2c60500d244dc311a88c76abc3b1d1bf3c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b7815b2296e3d92e741ff3e9d1c258ce7807be8d96ce28f53af75ee58fcf3bfb79ac370737e74c3f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9f85fcb8b5a56f93c17f16025c56d93a00059257a249f8ec8944d9bbc7b3ba9ed9d8a8747c377575;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28f7b3ccfabdf4fccd6b0da97613b9b81c020f04c6500d30f37eca37725d8139536ad5b4a50992c39;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9232fcbdb60172fad24a066de03a4ff1abc3ed03de7fbe339bddf2044d15da3c92381a46b75f73e3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6740d25fe88f7cd15c2fc70fbff9a4aa1b3cfedb253f0d6b2edc2c6b7df4fb76fbfde6e7db1807a7d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb600f357779380b65eb8f388d033820352d4b15203b83fee5d846c58f51a80bc899c37e8b08ce8d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc6f9e2c924a921750c12858576d8eb6a0598da4b2427d8649541decf702603e898a507fcfe87080f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70e278fb1101e900af8d28aa54671fb9a158adb342875bfd2fd3f1c69228bae191fc4777a2dfe4366;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h233cdecd09d4a5e8016f2e920cd570afe63240c5d3a69889992c399fa5cbaa7a7ed89c2572dbff8b5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60f363158e57d982718e9357e0ddb1790d4fc8fdfa2f8ce3e6f1bd11768bb7e36a859ef243ed4deda;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h146cd7f8f7843b611d83f8d65538d078eed21a11997163c99221f69a8ed0dd404d6e28550387d584;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8eae65213c47b101fa2de8682b45d60cc6835ce65e101c6c4c5ecc23fc6029a247ec1f1949996beab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb23c9f20e3d1b0d8a23623658d71af9af4b2f0b59c6782389c540a903e5d7a8c621315fb10124f39a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c99edcf18b0bb3a3c615307f80cca5c38f3d46a443fc87754aa5fbfc3beb2a02f185ae5317c436f2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96e81f34ad0f3ee214637332d232f22b3e125cdd4af6d2b2ce75b7887a9e2b6a85a4ea0386c8c81a4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e61d7bfae9cbadc6e109536fde5211c60686692d8ac6ee6afa091d1bf268879adf9e334f8392398;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda4c3251055f3d9d0814f6ef41f1f60a88fd7f2ba12b6929d38281597b89346b783d6ab1564dab497;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h603c0f473afe8d2d1f40e3f25b88064a49499f7fe04c459749b1c57d4ff1810970b70be30329795bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8248de8f5f7815baf33b65456048e2c2ecef52ff2dd7236775f9dcf161806461a65d0bcd0ec934688;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6fe78603fa46da4ccc4be1a7654f137b828bb9de3f4fa6a1aa3d5cf84ceda68fd6cedff7fb140c71;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4685b9b3a78235d78e90754f45c7ea59f33cb9a1caef3c8ee2da230ed313bae1c4ae5d13f7f598c0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1f617e90ee37fe4dd37b1ff01c54c965e4538a99e913803867ce5d1231896e1e42310e68d11d0cf6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h209ea94a78aaae3217e54e0093d283ea08bfb19d3306fc7277394b6ffbfd613e4cfee6231bc32e2a5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf05b2d150953de7c233e6f8738ee65b16dd03c599043d154ddbe129b583a0a7bb8710bb1e65a677d3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97c7426af3aeebfb278eaa8ddd2f905ab3bda222e189321a1018af63a6cf20f9ce46bec3948211f58;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e3fb0f022cd75cce3cc9a00b686735f103c08071db07a1b6568e0ec3487f41ce2fd6b664ea9b6509;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbefe22dc4bd07a331223ce4ff51666d193126f72de5b1b63e2a05029d7f510c0dcdf97e425b670142;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6df357f66f5b3c9567d5fd2ab37bee204fb2265188519f5b1538c5095c8bdef826b6e6603ebc043a1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he27deae28a79e82dd4ed23f21d13f4fd9ad0dd9bba0abb6221cfff08948fb85f494b4a71195a0cfad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf757dacf2c68ca6c8f63340c5fe84fda0d74c95f54cb3244a73030b7f7d4e75668b0b9d6ee27372b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h307e7dfc80d27c42b08e77ebadd8922aee90f76b6a5a8cae6a9e3243a7a6513763f0e920426265487;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58000e7b7f748884050e515a560ae19585078f92d3c3c6b20c5f25952f03dbc1110bcb3743936f08e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc315fefdba0eb943c91d43cd98941ec9d5321cd0b9252bd9ec17c4f44a5213e210eecf7884fe720c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b67a61572ae223ae36865cfbf194b9e9babf594c8c2fac086ef4704721901de0cd71312cc715c6e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d407b7756e97d1c0cb39f5612c085e05737df3f26b03d01bd3a81dd4a326d3345df06dfed04b40a4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbbf72d09c79bab6cd95ea7080851926ed709f707a5b058882e424714c71edc54ed3df2a7c19e8ab4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c5d4f885445dd818c22736da516cb3f776f8a5d55bead9a7333c5b636e8f67ca16e72ccf07844ff7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h267ef66166824b1d0eb66859b98eda6643cb293cb8817735d2681d47d3fc6883b6e4d53d2a9de087b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe7fca180bd03e7765b2b7ae2279c2e33b92b9c310faf8eab296cdfffaba370df72618715672ecbf7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6e5c53614b55428937ee6efef960a64eacc7edecdfd3ede32636439efdd3101723c336ee50e6d5ec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce4404bcdc806db5996cd2867c1c97b29afefa701988584fa6d064ef632fb278a60464bd8a406e1c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62f00c6a56e1df5829b51528b8f4837c969abf6e0f6544fba36b24e6a30f031ded35450736450b8a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23ebda5e78ed974aa99acc1eae63c8b3578e951af0c1ecf0a54085e88a155de24f7c9990265d6765a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4bf33d04f8d05e5eb7e053e1203cf3ae2ca97f00c158f8e65a8bcbb6152209d3405ff5641fd3e1d5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d18adbfb242cee622ff7a979d5ed54dfba49ab57e6d00fe07043b508008677f3073b8ba866cc9715;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45f3658c122b7f0c04bf0096c736f1c170c5c2c898be256e2d24cd33a6b9f2ef011606309e1111114;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfb6a91941c45d8cab92d9f66302cb1523d42b867067ee7b9b9081d9c1d6ee820aa94bbe0658d8380;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h134c5ed9443a1786315afcc6b8ba2a5a4d667f9a9504bfec6c81f07e1da3d24b7a3078b9d969d95e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he76029edd9fe8af96ded9b332421634b33692849432801a622c9e8a798186ebafaa4148f43510e4bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fc5ed3e369bd5237bc37ac666c8c652bc7fe95ad6f510c21a69096b63b7cedf10ff888ec5362dbb8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0b19c6f37b59157a26123a90c32b78081ad72e2b2ba4430cdd2ab997e426d338f74ea6248ef39105;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba5c3f6b2088a1f695f65adb3f9429f0295a7dcd3ee83f2fdaa77e8ce12bafac9aa1e87e2e7053384;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd39ce0c6e31c1e66505f7cd9dd7a0c387a6cb6e0a29a26a55c62398255c034fcc6b6300b7d0af7cc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90f1d09b8528f93e69fa4a3e39a8335fe94662a41eb16551d9d87571ab15563251b2dbe7bbcf631b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e4336cef481cab24edb00df539b75649078dc822dfc424027f691646531156a083506ce979a7ccda;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he510e7a6f1b36572cfc10e7107689a660b10af90249ba9b7e20eb1115433b711fe3b5c2540628ef7f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcbf58af3417d4de385289c0b013724457c241b1f591cc665a066d23e40b009f401f01cfeddf3cfc5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5afa198da63cfe261c12979c1443eea18aa01612739b7e5995f6dc79f328f5573f6eeeffff48bdadc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a807bdcd6ebd920c7c0a43c11980b7e51c3f3bf0e69a129b0331b142979d9c081654906548b03e35;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff6d65dfa3dbd1aee4f63de313a8a932f115b847937d4f0b2437fabf371a8fc45403a152eaff9465a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h824952a0124c0b719f4bc1a977a7e87e35ac126b1da2cd68d858b59b7528d702aee859b7cdb0d3f6c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd420fdc0a874de09849a99105ee439cfdda93bc9a0879af2bfc857eaeaaf51936e67284a5e139c39c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e9f6081b2c1f5c13f18436b87acaf45b51da6c3fe65b31abc4bd5c91234397bbdffcf921a35119b1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fb5ca0579c6e478d46662c073c30ea600f07f5753ac2dd0a4b26654866c8b051d6c897f153093b99;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c60fbdd8622f1b8762f6199f2e80fb3404b3a9d0ced99bb5a06f87a84a5cc26b5428decb0f5af37c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5357e36b70b10b7616cf43681c9be6f4ecba18908095133c6efbbc6a840b6882875d0ede4c8b661a0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha94ab41b9ae67081295acb1079ad8ee816d374fbef6cfe99c155cc65c9b90980026824856546750f9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf46be63aba92c0960eff15dc02dcd1f8e1eb632eafa7ad67e7c7be95397e2b8b28a4c3ed7a1e2ab4a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37576e3c55e6497efd56d5102254a2b7fc274334980aa2cf15018d215ae836e86b6c2113323afa03b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb95c69f7022057e052392b7b81e3bfe4058651ea32595c7ac95dc6255f8c3ef0aa19639e8b4db375;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd56d5300ff86f3fac4f3ab5a5c1eff69a00a5c10f61ce9670d8f61193c1f236ac16e31bee03e0422;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2eade6a435eace5758d2dafa35f6189620d9cda4d9435c9c37ed2562aa75460e63c4aa0a22bb1404;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h33bb5f2e2acc416cd9f0a76213e867515ef7361fa2bc0d48738c554581a4b2e7ca033ce6a7bfa57c0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbca24e3c88d14196eb66270851105be50bb7ef6068848e2bee92c5ac5763ff28a31cd29b8cafc6313;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8282989053256ac00e06dbdc16db68a9a546780750fc4e375705a0eb3f63ff553a46c7e6fa31c44f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1e3192ea47f678cdf58938c10b741df68181bf3d8a4ceec2e644ea58b79a04adaea83f7c35765241;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc72aafbec126b52973e93198caf3fdf1851f402ff357d7777a653c48d7515df8a7cb1f30a9f3176aa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed73f1788f5ec8846c736c28a074f30bc6dd44dbabba5fc6a13521656d142b783e7c3d0a61ec7bba8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec1cafaea11380507213bb00773f827cb9e525c23fe03bfb82d0eb66ab9a6ebaffd2078ae855a71fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2307ce202b254f7fb08e37e7ca04301f7e945225bf038840fb7b4de7ed9520a31ea245b8e8093a7ba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69138fe10a6321fed879fbb5a2acb6c4bba9cc065d3eb9c5d8aab2988c36a4d79c6063be13ff8cf2c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d4b392971c0df1f15b55b4a02b3d5b65a90c412941cc2742cd8be1de018a19101d39bbcebf3e02e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb9a981f51091c60789fccf6c7bbeed4b9a750f71ce7c9de89570d81156f6561c47c3e64a7caa1bb7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he99e9dad7d47d7ea400f8c18c887ac8eb466150eb7c50fd883b13544699d4198222070a1c3d3fd7a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4798032dd18052b277c1d0d12263a097baa5b1ea18162841b176e914e840f264d8665e475640689c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6b295af5ecfd20f69276df7ab24e8ec6012c21c303c22b9b78ac61283695e515922479241436bbeb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e1a099e2f90fdff05edd9d030347f0c824616db450a80ebcd7d030562b4fb08acc2e0b64c0590dd0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h637418e44bae4e85a9e0508d8fbf3d358d287e33e2eae2cfac36e036ee41a4d9b842926aa8926009f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf5321c0336fd6c43506aeb5b6a3c04dd91ac0a28f3808d0b579d166287e3e7e8f3d6f4eb7e99326f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9bbb342c4e8f7af07d5e9a3b0389e25ca8a6901c0ad9091e6bd94c191c3ee7b432291fdb3ecfb0fbd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6083043f58c41deca5f59e59911bcf6c8c59c71fbe664be232cf2cafa228b7abdd77173acd569851c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb16c6546787ec4ee86b30b2a147d2ccb80c3cfe9f66033f94502b0d3fd845167e97d3c6039bcee16b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7f1519caa1614890baf944fa915f0eb1d2190a89d53b3060451702418a406337855c5719b6a6b168;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2010ffae824c9c620e8cd5ad0f8b76055a9bae65e2ffea57d4bf86c9398af1a2d414fa95ca98e85f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h766d69efbe6c99305b7a4604ac83c74eadb8fe8e455e68065652f2605e56c93a438fcf8aae346400a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3b86d50a33a087b332aa192a1ecd86ce54fffe1c627894a572dbc3cae90ca86f31cacb64b9142f6d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8caada1b6ba87f092b5498839ea3d1c3b3d38a04bf749692830954ba93f0dc5729ad8f5778dd9992;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d4979c842fba715c6b1b8f37a9109e44578eee8cd7a3a8049fd43391b41a81976e49be812f0de06e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88a140d44bfdbcddeb9f3de9fb5c754f732b8a557fcab87045b1ce1f02de0153798e0e9d3e3301a37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e169b848377d4c14e71ac6eb8de4ffe84a9e6e4c1dc9ff69422baf7867dda61ac746cd8a121a7d23;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbf4e59881454173e1f1e56b48feb3795fb96b14641c26b33929522befc5a0debcf69745579ef869;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62d495825042bf41c8bb2a821df46f52c946057e3f4dc1e82d420ba6896b6564cdb72267dcf9bcc0a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1bd7647eae7ec653caddc2ac0fda888a6f924c4d145526eb3ff0b99ba3d568c7763b6eee2bbf1dc2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f3bf6245d88d173a6206802acc1d5e2686564ca1f6b3fde2bb7350ee60df4bcf470dc728c1d94525;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c91db6015388582d1300cb3e3ae3a4787f1931605be3587da8f910ed9ad25f87706e6bf1a685c80d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69e07bee9c2ee4ad89b21fe8003e2b3a614106d831f64f969ebf40d1e9d0e9b5ee62ea8cdf37d3b43;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h551bb6f97fbb1bee5f180450fd98089c15de16146d8009f56c0e325d8c2f3fff3b2edbcd29c3b6641;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h834ef1967af8783a9659eeff831eecb7f7146e2714df0a2637ff50b6bea198a6b93caab950478157e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61343a3dadd3aaac1a85efdb3a16672ed5a47aa0f72cd548545584533bd312aaff11729ae22060d22;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ae0de3cd86870d5a7868d5b0c53646f93ceb3d531616d8be361fed8305f97c7412a0e304df3f20b0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h642af25f0af2c7eb083cec04be8605edd54fce282bc9674cba7ae40ca23a3808ed9feea8bf888af36;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h297ca2c46ef0022d12ff5003a61bcd5c56dce9eef0929daa9cb3489a4fd6c01c71db4e5cf134eee8b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48eb24fd038dbd70bb49d2ff69fb23ce532fb1289a6879b49e01000f8c85dc9f837e68a5703330c6f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h589c0cbb8cac838344469599c0df9458600e533b8fbf4c4400b7ed9d5c7636d49b981ad6a72e2687b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd09031ac9d1ef517d5448d308c0d4be2315257fa92956982049d82e9b0211b5ec18d3416733ef640;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18369a077ae2e719c7ba8f758640dc4f28eb8f78e88ec776830ae279d3ef277de671a4f6353ddb2b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21ace79f69060ec5beb643557d38110a0845aa95920fb1d1c89d05cac34b35926d3b35fcf5586d263;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3223a46cf991d9382399cd1bef58e645d2ae0e0cd2b9005d8f5d6b0dbf167549d2f4ab44d7a338c7d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fbb4fe423ae19d198ffec6c5fcfad02f05b7ec784bc47a9ae7c8b67b2f1efbdb6a4a95e623774c11;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac224d6dda1ef3686c43aed718869c351526ca97efa91fc9566b70a45b8bc72bddff1582af3f744df;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he41b7e626bd2ac2b54c3f4a2fdc31f6bba58885f1646f064e3518bc812a10331b9f54a5b2f5fdbf4e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9bbf890e978961c6ee3cba3b57a20e35a90148011b8af3ffb804d3ec54bd343deb26a641fa087bb2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e68fccff97f0ddce143a85b339efbf27b9c7413308cdb9d6b261fc69148e58819fa3b98758c7b835;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5461dcd7f37a736a9d3c2d3c26d7be083fc44c0f22f8331af4f393471ea3f7f052a7731861a4114d9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6575adb1e74030cc9d1cd06aff900a69fb01d097515c26d0f0113b005c66bac2850a6d1d91c1c0d72;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e5e8d9b4eb34e91ca4be04b464080658ed065f9571d7f5e542830c7892ff5c398e6e6463bf7a0130;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7225a4df9314883f98a8cfe71e78cd14db488d3c65eb80dd661ee289d4f6e64b2e7d3a77fc027b00;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he49690b80e297c7067e3f9a3970d5539140f69d7c886f9158016d227e42e8c47ebd2ce6b7b57ef63b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2522e64c06c894acec4759aa46f8b4c77eee967090c789b839694a47e1c8f8a77415278dc25a1748e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd65f08b50c77b992f6b9c37a35ab74c0dc775fb530b676dd67f8298c31e5be7b4d2cf20d310e7eaf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3683f2183d81a72644047e3d642b58ea6fecea7e4fafc6a58003161c7eb224a29f1ea951faa02575;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90690b2dbe1772b904946b03102ab62b2cbbeba63c371834f11a4c2595ffbc215053612bf5e7c9f0c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d7aa2e4fba61b1e085378a7a945f170786095cf87b39711c4f1c6e067382662d9db18392e98209c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea75bf07c2bd7edbc9acfd32d359b3339f7e53abcc4d5a072ca6f081ba922ca8d6cf3ea57c18e1e78;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda6182773bd4f349a539d859213dc25cfd22b18ac4e293406d40508f30496f5e1b2c4f81ce4df255b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf6294edb199ca170987c78cfa61ca54147b74e7b825e057a9999a102c856a8a2de959462f75e270f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h716b57257f9b5fdcc6f1ca066ee210b0963ad3a38275cfd91eb35bf1f58885bb39439f4f66ea7ee28;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5cff4b7276dacdce64b66e195e967bcf98646d8ee8fd8966b4f4ba566300204d4fd4c18dfce9ba3fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf964df9f5bc183075974fb68e3cc4da241f4bbfc10035084d2f16e168d8f404c0dc3c1ed9817f61a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3fe9764c2e69dce258eca8bcdf37789d81745a17f3472411db38da79b53cb36791254148490237369;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63e2958722ddaaedf6f2768d763120e38ceb383c0f9829cb65ef3217357b29789f9891d44d1ad2235;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd36866decea08476a303092d1bd8d7963842a3bcb9df62aedca6cf1b8726cd17433211f6d59cfe56e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4150e10e300a3de2a4ab43db3d5cd2c02ecb3c36a538309c104cfc28b826819dca8c7863692f8a61;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47e03cfc88ba25b47f6b92d0756cdc1d1bcb2800c20af132d9bdc9cce622c1d629ad2cc282c43e6ea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8de7bcb11a7867fa69709f97030c92fc798d8960b6838a99e8d5b3d9cd8d7ceeb4b998669d8ea7ec1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38b28076f71324c2ecd85e320a342db45c756df4f866ffd92103d1569b91fca69143bbf8f9cbb197;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he714613cdec73a6f18cd8364540c8549fbf6b3853199f4e00c9e041de97507211d4efb7563656850d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5b9a8f7e7238a33225b79274ded100176dc1451afd8d0a3725367efc4cf839e461ad48772ba604d9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h544a8dee3895fd010c9635c39fa58e061157f285c2660612b9180675283c09d969dba5194ebab042b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he13fd0439655d67092bb757fd13b3516a141a807c8eafe06d10281b0cad790a3becc45d3469f14a7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4241bc16664eebdbc760f0df2fbf8e0d6771433d6d0884e2c7743fb8a67b416356e0184c61f792105;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf05948ba9f1ef8e675b78a9934b5b1d9e73e48bf620b64c076a0f2cc26fe14a032977e48aad0d75a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53aa33b2f842e1d1e4613ff8148ea3ff7d7b74625389e61cd8ad7fcf6e801b7f2237257eee650b566;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42fc6fe8406c1e92751b43a492067f710ec393907986541be98efd2829cc09362e48ad5856aa34ef3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4824f5477d8e3160a849e13ab5dde8c977599c8b3a8735711c5fcee0f3d4a954875f9632b493b6c2e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h644e2fa6a95d9e15cd31778fd4eec7480f9e9f2d09776368fe269d8dc312c48a549da4c6831919271;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ef4e5ad17b03a188ecc8f842044590dbeae0893c38af01d70f3fd4f95f030616a6874a06b4639aa9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5e83269d338e56590447d2acf900b933eac4379027946b7df4dc8e3398827f89852896f36f7b994a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h261925216692267339813341b74a998db1210a45f57f9530cde0c72ed18c5e02df80c9330b46aac3a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h432c1b4cde0e9484e5908b7cbcde2945b91d47fc941daa41b97859a47dbdae567876ce303cba6f3c0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha86bbcb206482e6224928de31ed58a77591eb9cbae02eba3be5c9f13842151e86915db5c2723185bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f6b0d9687c27a620d68671da8414236ce001fcb164ab28d04b8f609f142b9dcb61fb0ef00ffd2455;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2942f168a668d7ba602255a5726c37a4795736df7504626029d65e4e92f1dfae98f45d4689e7fd34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haeca44d4c95cdae90f1e19610de0831d919b723952da0a8beb73c800cc5cc007cf77a1ae97560d936;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74e79c95b3a3ee6ce98752f3ed43f783edecddd439938fd845af4e60fdc742395aeb2934c1eec47ad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7def4e36f884dda57aed452ff07ff11f765e39b622dc1139297b26d50391ee0a27a88f9ab1c418ac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb55e202fcd0f7fa123aaae897b88569ea1d78986ccf6662b9fb1819bc2852bfe59a98929abbc397db;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5bb7fa4baed529ff89e47f9e847fd3c7c016b426b0a31e786fdf4cc4996650795e34fc653b166ae7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e49905ef7a319a79c04669b4e6a8699d03946cb7f7cf0b73a780070e463c1dacb4f4bee89708262e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4191dc432088a91ab93855c7f2bcddc5d39f81d9430a046936254a89fc1a18740ee37798fc9c4c828;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ac40e1f3aaee5a7726c6b976bbd87fc2920138602b9a13917ef2dbd35e9532342b6d04b3aea00318;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f72d1407ffed4fc7e3cd2b4cbeae9d5f9f27b3664a461a275b67851948772dc50917878ad86770;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc235412cfac5e675d59e11a566eb4922106a440af1b968bda5565231b3ac0502a2be992a531cd6f4d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40ed2c291b7b37b1b8e7932b268f0b9772c3b1fe7260fa52deb9558ea36a9a91365468e229440e92b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b1589acf43e4a8e1fd0b0a531d7656f02e7174e334a7966ad1202a4001f0d9f1164b9e45e72d7283;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4867ea3f0934dd4e162cd983288850caa3e7512aecb2811d00c651eaf5abcd43e6cc7058e6edc14a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf56aabe18ca5603d52d6d0123c40e2296dac79d6e2a63a15ab3d379f1916d3bc70faf3da725676016;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc58b2ff0893f2e0858153f4a4067e50a749317d98a4f762a7298dba8bba953cc494c71eb8f48e05fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ed60b208138df0479b8f8c273a87c6be69c7f1bb9fed68eb6044d783f2e232d180282776a37ab9c9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3e0da63073de6171db5d79b82d5fa9737fa98a005104bbb5f645a8ecc426501320bdd1239397cb32;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a52d2533a9bf4e594445bb32eabcd6dd04748676445dce71cac6a4c9b4a583210276293a6aef3e4d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64d2154e1bf87e0c567938fe9516acec8e751506b8c664043630116f2270c29480776b8f0a066cc79;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5016775cab8fd1d70353469f1b05237e24d98ec98593fbf65f77747eb6be6c7c9d3e838e08a2b632c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c1fa79b9e38d90ef9bdeae6a867300fc764bf0c6c8c1858dc8e01fc12b843c2adbd340052b4e9d0e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h938a74ac49232dfcc1674f174402ae19412a807e39842a2b938a7b6b9aef62cf2bf1cdb33819d2fa4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ce61b466f33691e7c44220f21a66885fdf9cfbaaf5f7b0a40d5a18c911e5ddf8a7224d72b6d07c3e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a4160849cdf9fdc50ec1956538ab91d90355d073e6017dfbf41713663cf50cabd3c108548abf3251;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7da8d272291f932925f3e9d61c1332a1544989388091aca2dee8f1e36057f6ba32b23e020c3f3c8c9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h880832eff1ddf70baa1c75165da88c524c57d2b3a18184f580bbbc10da1da91a844a8ce22b1090c2a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73561cdc6d9d06e3005224a3812e88da98ada35bb86ea413d37a8f6084dd80ef5bc2807c382b0b374;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c111df43e5288d611d2f1594e1e6fe2eff1e6f7138513f3b6a49add5200a669d8f70f2461167f347;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4d7784b01e2ec5ee3d1323c534d98977e827810dbc9d46a6121a0a2a3e15f5acfb8c869986fa0e42;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85a2b98a01911ba869a2a56a97319c5f349da70e0d04c700d21ebcb5d1706c449cf5d84b9724aab89;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h236f2a282dbbe6f6c346b79b9fc7518047f8f7270bbb95c6d6f5e78a77c26cc77a9ed68eeeb7e1e65;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48741c41f5fd926a64ce439560d9ea8bfde83bf56e3d842041e920758c554ce1845cc32ae6dddffc6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd663b5da362c33bbb4fd9467cb50e96ea830ede5cbc44a5463248ed74e8186899da3959b03edcc6e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ce6353c55f471f2e1fe2b4a56854bc84b19fdc14e205d229c9cea8185919e8f1677f81ac35d495b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4aefb2abfba5f7b25cab1587f13517d23caf3870eb241665389ff5ef7665968b8437893c5b84e7745;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1fb02ed349c29d6871479df83635b24c75c55574394fb51b21f1ef0596e37b63f3d96d842ebf271d0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4c9a9185d612443d8dca91a849341fc6fdd7494805fb0aba4ac4151e3f28a8cbf4f43c003adf5bc5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1dce7bed3669e51fb9fdb33e2f487a48c339d0062379771c3d8365d51ea18bc51bf700ee725de87d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc48e4d6ac4541da0bd12a6369846f17d07c6372acb0919d52a32517d2838e4c5e6244c057ed0be2a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa930c6b5152e1cb166912d3099a3df6936eb7603afe998793a91c5ca6d77d71c6cdf918829ab3f2c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd84c9fa6398d6e3a152490f73d7c7826722799ef97782d98a79d3f3eba9df41e4f123d1f471c51eda;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1b84a25b36828b6381cf17941e2d32c281ed093820925e213a896002ad98129a4ac844bdb2b98c18;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a9d95f1abeee0ae99b3546eba063d2ba3eaa37ca4fc699a7da96d33722b7a83c578aacab8e83e748;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57fa070001530caf6e9af8cdb172d71124485b573a5a8bbf23024df328022823308827ea86b18ad0e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3fb6901956867d3232bccfa9eacf7aa5ff1ae8a13fd1e555a398f9bd853e9985eff6e5658c6e418ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f065e0e08981356c78d1bdfca24f202992095b0f1380a1da0052274d5456914ccc469cd454117481;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c513aeaa093106046a9f8feba000f8b94a2b147de0777456e6ea60a2ed77f97ca2e1ff662a10014f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58bd086005e4aeb80be6cd15c3f34774ab3cfda7b24bd8ee3e967b4623ee6c308c40bb33fdfc28687;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e7429c9ada76e32c4c49e456fe51047b420b742da3572d27cf2df251b5cfa8094009d95f9d38089;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c0d4ebeb6b40610599d141fb719e68b3c7b5ef2178fb9618538de45c84d15e8d67b1c479b5887379;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec62f72c1eeb858881de232bc797ab0108b099768def0f6c3a70caaf69ed47894d8d49a69c51a2feb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb917826355271d04fc55220d03c3046fd0b98bf9abb070845b32a933bb525c8fb1bedde4caeedf80f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e90a829167c5c0c1342ffd586f248d1b1ae1c531e9b8dea916c50d178499f28417fa67ca6be2a801;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a6e04a43cf599dd3efb581abaec2aeab358c929fe25c890de4374fe8ee623c5c9e60ead02e4a454a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h207ef2a4107741056eda276b6650f03f85fd92bf5186bc63f2cb48dc47d95e555e8b5795d77a71c3a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf92bde548bcc59ec36a1cd91b819dc13e82819da30c28850aee8faf0e7cad62d63d95859d274fbbee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbeb7286b08286f0df181f4278ba07cd9eead87e2098829e7d8b9d0e3fbcd3022c1c4fd3dd77eddd37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5420267ef4ebdfad3f445356e594aa3c1f31414df6c6afa5d635d3a3febef6f648d7ec621a2ab4b7d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8583e3611363787184c7b7655bf94d930b0d2ad439114cc5101bf1ff9771a365e0a2d5b16b43a981;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7e77d82d5d7e394a2bc74073f5065571ae41125769c751e57efabfdc19424fedc7edd803f1ff6cdd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18ac00b6abf58c03d3f028e709c3af8fc7597f8523b044236d81984ccd202fa78b1e4b144df816132;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd434370313a5a3217f8bb1c9951397a5275c49a74b03571613f1632af7989d5d27c24b3c54107eb91;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84c8030ba4aa0faad58ba21dd82bae33554ba0900f384390a20805ee7b0dfdda49c30653cd2be55b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57b972ef84c52a869826f66553d00ea3a2a7ce096a07980137589b8b275a368d244314dedcbbf698c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd851991050c2a32cc14dc7b59356b1c49792d6b2cf896f476fa29625be4ba31acd4041223bbcc16e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48843d18fa5200babefff42391e536e16b72d3750864ae4299ea719a2e3b494f199aca1e6e1d31177;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb33124a3bbbef35cb5a831ef278028aaa7df7b0f5b8914c38fad6da0eb559f1335222c69f3b7b08f2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h384ebb8d6b2c866c6a6cd31a511def4853c7b8b8f10dcfaa8c9a01001632982ffff7f6c404c90e0f8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc70f2f077ad94e4dc2db49a4bff0571a6cb56e7727648f0f7f478aa9dae328e99bb5f39b2b5032dd9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc56cb35b5f2deef4f3b9cdda411e45695dcc962d18acc6557a74752837c3ce53047f3a52e75e67a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5df729d929c098109b891fd66afc3f70622b2a718ec44b120f2da80da14484ac58d8f374bfef78515;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d28f1240c0a11a677d0659023aaa0435a6089e20765d4fdf1b5a967ad30040956e7351e78679e862;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13f74ae6f0b4672d4bde97b24aa25e241e25c1eecc2278676e21f1aa86c7973d9efec82fae88d5a62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd7c095e6dee70edf41cfd6c5ff3bb465f6f53b5f1c7e2f02d0accb764a64f77bc83c097f1d7dfff9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4daad524140d6b8bf6011013b6286e96e903e90ccd826e7bf43fbb948d44cdc2d26578dd298355a0c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a8ccda1e6050729c9184f2c639c47feb0b9afaf7aac74b886aba3e67e9407816e3a2039c9f62c641;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2e21074e78a0114882c521a08d2cd12d451ee7d1561325792da87ddfbea03790bd147090c604a8b1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60dd2594172adb43f100a234e0dc331ef13cb12b5b6419eb323e69385c281180d42ce4a53529c4d4b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf50332ccb07abc8001d6c5e1d091a3acca0cfb9bbc156c58b24ab99a232eb330fae626bc1cfa6eefd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf5baea99985507d4801fe6bb0454330717435733c871712158097b9b0e3c2666b4e091da29eb53a8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6df775acbcd877e678f7c0da8d71d62b8bd62631ea8c5567f2731a926adc9283fc17f36d0b265c609;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f7e79b20f895afb9a78e317959ef15ccbfb9f2622547903f3f1c937ab67d07aa2a4dfc3648c01ea3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h763827b7b1ce19eadf70a0b74bc2eabe0b7954c301f175835115b08a327db426f4709a1ab3aa3358e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf7f9e25ad2e1f5beacd537b8f486bc443056fbc0a11efd24c8add4197a8d6075bf30ae1c9555d5ce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58b9567738ef4353d2b9b2879812a431edd32b5420de246e02f309d8ea33bec40913a6a32be4cb408;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7abf009d087ba2429b8a4baa5e380c09216b89a56e10456211a7b5e5ba1aaeabe1718e68165c3cdae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he62423c814151c2c4008ad3b59c889f8037a8b408575e3582134ffc53aaffcba07cafa3af7d79c151;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcdd711a7dd944f177f14161e6e06b9c108f62d3b3224f8a3abae83cb316b2c367b43b084b79011138;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a420b9ecaa2ff8ba1926d5333deb33ecdce60ecb261c26473984ced3dbf743eac265c337553a172a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d79bc5b627459ad00b4c5ec030c3a3fd9c112430bf5a53291893c9ca8428aecc8379b78db74a74af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1710496deae4ab43f9691283ba093bb8e1ae820b682e7d4d47e2a341d763534198b1c920ccfcc211;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78c82f11a702ff389c0721aa0fb8d38ef56116277a0265c8adca6b6ac20d51f2a454a916fcfd32afc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b3422e3ec058b9b94f2dcf9633e5c34f7980e1e6f8d9aa76299392977a1c2944310c2068b45d35c2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha272f121f09cd9438b617fb315d812b704422d7f709203e9cf070ad0e9ac253af337922c734f04940;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc596d3e552d2e646cfa636d54448a87581c1c0357897f66e8b2f71ae05f4941a58b053243e2a3bfb2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8cbd243300942e54263b8cee8b81640bba793b18295ec757f7b96439f8aa19683164fba92e21215e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20e2e9d078ced9bada88f031f37ef202d02395da6a5e72c228344e5592bd35cfbc0ee878062bfee4c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ecdcf163c062ab00b3d307f5e9ed71f7ce14bf1703e9a19cc94de83d4b0fd62aaeacd5d968f71a5f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee70920bed8e3d7ccca7f03028af68547d607011be944df02af3e6653e09553b3dd4a6679f436df80;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h313b835b75063b44ef3e677100a7aad84d8ab39b0aeaecde254f4e0b10253e867b45b71ecef9a9a9d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6893567b719e38ab7976625d861ca160db10ee8fd6cc0ef2f1f11d3474ec84aa878a17b0f1b0a77f9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8d227e321fa2215f95f1f30c74976b575136716d371e6f483fb9cd6c306360d01dad91b9cc480267;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h743137d81e1475df03a67d3e8de38d9b975810ac54be4785a24904c0293707ae77402e925c7aeea1a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5082977327fb97fc2d52d0ab98e482c42ef6343b40cae0faf1591f969a8ba9323006edcb6d7461cbc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h227cfc4cf8022ec81487747a2ebf1a0e036327eba0518bebef9ecadf6cd277fbb45ade330b82e2a44;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59f5bb5b64057d5b72d84469db5d1a143702d4580d42c7e6e59a6fa7d8ca0f0e285dab09de987228f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a6b33428dccb90d6ff45ffa9a92714c8ec3da019967d76e701351822a8494e5e34207006a41ff1d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94bf09fc8589d5ac53402be201e7c849d78af9628c3fe38c2190b47d912f4317afc8c0622c0cd5932;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42dbdb88ae8271841ac0d3c259f926b1e187328645a6c5005b5e71a202b8c4d7afa4cec5464a5993f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68bfb278fdf6528ce80946d67b241e0ff852bd3390310b5036ff78b55ecd32001325d380e3836720f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3d2d7c87862d5536c76c8303d6201cc5c195e82532646d4438351479c4c00c5cd9d0876f3716115c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc79c119d8079bbdd949558f4a29a0bfedb34ef642f470e305a56db4a378175a035724aa0525598303;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5aeb53db8fc121cff6881b2289229ecde906ec0d1c16c930b26d4a87c32be56bacabe80517a768393;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb5c19e7057da3b5965cafe3a49edd0a081e561eb437a506e35803c634dbbdd8e9e6ebabbde92f1b2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf3cddba039d014648ed705ec57199a7eeb453a463b270640c39c1805b5ca35c6f49df6efc1988554;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8290f40c6b408fb61333fa79dab87e784711ac4b8642c5ef5ba891aa6bd0056c5a8934f8fa71812a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e44e2d9c55bf52f2962af35b49adca14452aca5103e3a6766bf66de3b573f40771ad6e9e6faa76fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6bc03f7e2e8849dea7eef996b2faa999dd1136f3a36da7dfe427ad6f83fc12907dc47444cced195c9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h642e5d37e87449a1883c78d4d25d2a6d24ea58c78df5f0d7f7d7f725a85af49b8a6d9893ce162002d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h613b2dd92db0debcf2854c8e6c85df68bdf0d8db5a57abeac29657582123481b98f98d4bb75b68c59;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb14d4940c05e930a0236673e2de5c9e42816ec736eb2876e2f0639276b706fb4308dabe17350195dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2225e6e22c1bbf5eab41d0d5229c4fc76bbdd81783260de8d1f723138f8c343bd8767e9f684dafe3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf486cbe7ab2c7dff59c1de416f75e41cc9f96270e61a107a9c4d63c1a025d36650fe5b806dbf1c4b8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50e0c2cbdc76137e845f90b6db35bdba2783f194fa5627d7968b838e5a3bfd9acb58afa65a2894807;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h382995470a5f2d0c474d83b4133f395116105dd17369973d3234a847036a2e5b83ccb8469d5c5ad7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10d129a119017415ab7e6d559d9442325972899759b78a9ca661ad449fa44f67f51e78f5c1a7b4ce0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31ffecf47ed5f2554dfb25d156e791e605763fa0a8e9950466eb84f5331ed121949c85910c42df5a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea8cb8ee0c0efa6424644a0a7a5639a3fc16c843d9b59ad8599b8f84ec1ca243459e8b539d1bd800f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6293f54825c9f7003969f6524af7764dfec870ca16a382aa84c2c7a5e676283f06661621fc011575;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha742c8de0028cdbb55390770713a40973e6926a01b038234ce0e634f826dd20757fe84b6c2a8b5fb8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3d922e6c38e7996bd40325a3bb93ba2293d48bcd20fad8e1144f10f7941ade7556f094ca260eb27b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96ab15d846eb77179c16f37f116999f50af18000f9f9dac2d30f41ee952fcccb6715f709332ac5ee3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f16e41f7acd199214b6d0aa1bdf2b834542850f71bf156eb472c23e79e1b09e5449bb889d4ccb8a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec2aac582c643cda378d4ecf40f39907ee1abb10b3d84d5eaf932be30bb8bce1503ee9cd605d792b5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11f90837f87e5723fec7c191ca6c05e9569be9a41183700022803df11ec2dd0a79dd4c0bb8ee1d63b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae0911f28b8530f7b3ad2e72ec493e9310dc0f591a2dd7810ba66db40dc69e7218a45a6a268447669;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d54ebf7f4bbccd6c214ebdba3d999dcb6a45ae742606b3b453cad52d1ba0dad8a91683d3b37bd978;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1b766774de7245d536ad806530dd16857c1cb04f24cb01bab4e58d9fe3a25fc73fc95f5597ae52af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4db502340b759ea1789eb0398acd587fddf2246844bbd05e3fe6549923236686d22e6b43e16ab47b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31bcaf5cb19e536b96cdeafc89a7b813eabf451c209b62aa4fcd222d13d7d1947eda301c5b0b9bd69;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16627098ed381a2222957c53708f0a713f4ee36da0db9772d6ea5eaeed4ac8f39d886d9a1ec8cbcb1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fe297f8b5b1ddab72f0871f237558a2560ebba138b75ffbc6d63bad79b5b99cf256c73608cbbc81e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafeb5711e2f052ceb1c54772a1102bbd35a49972542788e4ee67fa77bb9686aa3621be04cc94811d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4697da9818c9e33ddfb0513a7258bb82dccf34e39dd3ea76fe3052028fbafa51add6d76239c4a58b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a89a3493924a5379d32d1e9890483cf80342393529e20b6059fa28f1c90cb28557661a8e185cfb16;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61c452a93184b828c87aff29b581af31adddd4fb51762cc4e2c1abcb39dbc5d718ccbe4c10c63c7f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he68ea454719faf04c650f9ff9c39cafc970abba57a0041ba5589c280f000f4f6517456319783a0391;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0c00995b553f50729d15b6be0670a5953f20396f0ba0ab952758891c5f1f38311b3f2c4418b6790c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0337fed8e79454107629440308f96521dd656fdbe7b14a27179171870d87edd2fe0c04fc46113393;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h320d030d5f1081e5b63a1c25824561945cc6a0e14139b9490f64689d39c99fffcef14e4d9dd3c84fd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddd2c0542b991c60259e3bacffe0eecfd0c630bf5f49c603acf6362ef90901d4a29d625456fc4e5b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he47545c02e586ba298319e46d7b9b296abe0190c23f734e40673385bc9a4319d053a3c5e4645eca8d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0be92ff2673c518a73443400e8deff4b51f75b718a87b50a2a2ed644c8f2758c4b3cb33cb9578f84;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6320c9d9a6932a1b24802d0f78fed1f27f49683b55beacddcec5a3564c6b08a9ea340bffb22e1069b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac1c8e43dc0b54fa2333f2f5201afbaca83a6b08ad6da186c8d40004e3926717c72a1c02d68f3cc4b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ee045263927881bb574468ab979ae5b1ead2cf9523b6ff6cd76af4dc8653c9855c7bbe16dd7e8322;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8ed0c323f75413434cddf92902102ee47d396446733895c2e93366aea626d1793fbfbe4c232ae4c6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6233443e84f17b96cd5881ababf715da91161d9bad7af3f939dff31785c5a46d5358ad4a1adb99501;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5ab008a15ec0a946f1cf9b7bf398f04a17c8dda03fdf07de675133e29e59e7bce6d96804430eb477;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46707b5fcab53b1c40b27549a9d1134a3d5c2ca9a9b94ad87b0ea9f7161de1c17a79414e40e9aa583;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e4355fae299b42a7bd6c6823018908940737c47979c10f66b47ba3bcf6f79c1b0da1bb16bc4e460e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f31aecf4ccbe9d243c50f8d0b89b38c96d29c6e772ac65d94e909ef652d24f0442b6ef8e55eb8963;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4418fcdabac9ef0a5e998acbe7c4b4f74270dbdaccbbe7423c136f7c2237a6356323ddecc816dae3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0f0326b0a244b54b2649b3cf7ec5b6351afe6202bc6b6048136f7e9740a8abe8223399c8d3a50557;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1cf463ec5cbaa9e6e0f37e416fcc66b11015377b660f64d58cfaedba77c3d299bdfc26140ed532b0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h607ed78e5ede03d73811d1bf86650aabd6c4cc59917babb6ca63ee02cb66791e09ea683cc84f1d1f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27969105521df4a87efbc9a9b667113cb96e09a72d49c51afba44e6391c818b85aaf4bb484bc3050a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8413bd611e832ca9f9f8a78e38bbdb9ed6845756111f7b700f8161bb0367e82010ad1dfd01f93d78a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69bdb9385ff91845a75160c93a847b6873a61a6b7499631b418db5e42cb5c0dd63d22536488573300;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a79860d8c740a70c02c118bbeec31534a0669006f4279758e2b66ddc1627279d7ce85ea3e713299;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf076acb70fc5815ba745b7c58f963cc4e0b12862f02f8d9115af64c90445fdc5a48bd8f7d15ef1a06;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbb7b5bbe797f69d20f1de4e4cc1c1569c57684fec7a7159707aacd55469fde93c42a01eaad99ea74;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9b037a51929977c4fcc20f2a5d2916a186302016e7db80efd3968318fa00fde5fa92e07c0ed474c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea664ac07717aa67af193dad4a977b372baa7ab70570cf784e5f81724e94fab49be65dcb6096ba1ae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd09b9c57182f6c0c05eb5751c32ab6f668e691c1cb275e66ae41348e901a98577ba187729433eb3e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc647c9cdd3ca14968b87b58be6a1ca334c3d7d2c43984be0df68a0a0f6af61dcf15766ad0be006cb6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fc45a3f4a73a67a6e4af71a4ea9891919e302db9338b1b4d85c1f05a9cb3bb8aeab9be4cbfae54a7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4014c9bc99c3f09042d1d503b59bf3f0f8a03e532fc883c48106dc5eded31001bb5008ba2113ea605;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedd6ecb7f879e673b32b7caedd275484e19e9442667d244694518eb5c3014fc7fc5e3d1f6748c6bd8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6fdf5c42c1dfa780730e267b55c16825b678960b34724bf681826076049e3ca6847d19726539a6e02;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h427d481712a7a4f6c7ac211001b9aa6cfde7e7b69b9dfb5b659ca7b1fd611d7351cbcd44887982624;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb2c4b35be9133dccd0acc3d3baefa97fe2477d2110cbf61300e5477053c51fe0844799b02e69ff4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hecf5748edc3ff06a5f1999f23fe670b419281aac88215a6ce9d0f01c12aca9914dc7e4f5c0f63863b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53d6575d77ffab446d9e2d87dfa976f108be9fc8380c4b15b14a93714cdb5aa1b4c1b336722085de1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf3bccfdf0e8f1abacfb0a4ec691df7b487de04f737ebac38176a83f5d28957687fced50fdcac5788;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71406e31d1e0fb5f45901daffaa283ec33e4112fb484fcbc67d861ae3b62fc3032d102217de9918bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1f95f7e736eb2fe3f96f58b09a4f528e75d609211197503b4209c9120d0187a0afa7727813c0e159;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha59b536dc1a5198281bb641f0bef56c65f5aef523252e65c10a2f55fefac2e657cf982d139a89a607;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53e9d918af656d1da6d8ea0c396fdf050d33bb407024f8a90e4e6d4d6693e813da2cd238666942a37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5fa946b4cf64ab625776726baddff0f48865534f2973c4e72a523dcd5b80248cb543c2f8b629316f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87dd996fcb1332b60dd19d5f3d97d597beb51f58fc9816ff66956855b807cfb9ed91393620c0ba4b8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h370148df05b8b8b59db22a8c4d0025525b78f2ef1f2e334928f2e6d7ad04ca67dbbbf0a476aaaac71;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae8a6fddfbb20d07f02baac40228f8335714a57f8f4f958ff72ca2be1aae80ce84a089381afaadc97;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82077609ae313e25e9d50ea8f36dec8de49b48704676ab157a2fa5df2d4a6800ddd714d2c073df7db;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4efd904e97bec22c01d46283208ef3a69db153cfae92f00978cc6b167a70df5e49e2d9807a1e4f67a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85e7140d810796407bdd51fa2942b008a19d9d77e955d5ef4fe47a3fa6bead8b12c76f0d6118c01d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ae2205e1df3a9c00227600fe3fd08df95dbacd54392282537a87928c977dab9f9dc92010df9fec3d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8beaf2458ebc04005e1b69aa095caf77c7e38670e03971f590c7de84d48dd2fa91cac4772d9e577e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80d61fba636fb20840bbb2864f0d52dd639038ac3954023ad840de08a9e136209b4ef1789038c304;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1b02afc61cfb12467efa551e877cdc97c536d83eabf81ce5dc2bc224628af0f400fc50e7709ddb63;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96a8907dca0b0b81e27dc1bb1b4ce0251e97a99ca9dcb09e999b72b31e3dd9c82dfc0e9ba6a08539e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb237efbf6019cd383fb10ffbd9f5499f12be57cda4d4865216bca49e212a886c53fa11cfe8cdd7a0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6b8d47f9d7808704cd50e3bfd76a2c4d9daaa52f3d758791662e0cd3c52170599012f6662c85e320;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcacd5feb5fc75f450be45cdc7896de81ea69cd26545ddb659a0880001f32feb5f370f568e483edb2f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27c8724d54dbe835bb13f4ba3c2b11c32085eee0d85320bba9cd565394a9dbf11a90bdf2da41289dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72194ae93174e2fdfabbe08e765917a95dcc5588344c24232ef301716d1f05e243a78a2c0c5855127;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc323a6ac6f07dcc9435f1d2d4a0cb1484ba750ecba5848a5f7936ddbaed6fb47266a7a9c6920b34af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65330a34b87a2d81841dba7a8f65625994a6960524bde2f8c06b47d48b93eb36d9d70358ebe2529cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec7f69ec1cb55a6281314049330956ea572a8676683859eee2d255cd7c72a4bfc2dc393b983112f62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91f7a657e394c0537476c5fe43163c658532f7b0404a06eb0f9804b938aac12ef82fc051d3c56a92e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b8053ce3aef52074a379dafc019c24800e120988070809cbfc64d514193410cfb0b2072b4fb34404;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3169d185ac7f85fb55a5c14e2511afa88056541b797b711f8506cf8bf33e0b24ba93ec55d701c72e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c71a18edfbe0f026e07b403fe596fe434630446ffc4c9e5220e4f53a82d955d08da51eaf91a763d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf340a01593d80f192c097490ac4e000cf99f78812bf93edcc53896d0d59410f42a1e751ea20fa8b36;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c0ed62878f8151d30581747f0fd4a31741ff7c77de5eacba24d7c0b0f41ecd73379209e092668130;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6eac1a198fe32d3a9f633974b7ace9e16b7c8a8d571f9fe282d50f4fb3dc75e78f600689f17f0ca25;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd528cde7faf55831845907eb9275c41cc93333d148b77c00eeb606b9296ead81f285a940668a67fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbee27e38ca97f1843f95f579c6256c2723c6f221af69c53862c95978f8acf77b8ff6d0e7ad1cb2cf3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hecc3518c3fa22842485d87a2fdcef0b1fe7e973ac43bd5ceb442e00ae6ed38a1d6582269a843534ae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6013426b224102792b85395f34e48bd4a5f8b5e884f021593db4903543f250b3744bdbac76ec79536;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h800c53516469f06e20bab13e2f220953c1067d9e0c4c498f8c4d93f2d1cac50566ac91545a949808e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a83bc4f66a10afac1f3ea19088c250f96533416b40f0147440ea9401a13b11fae7692a1db9eb4470;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77042d8e312c8570f6a5ee6bb02c27c83a8ef5a06210208c49999bbd983cb95cb0ff60bf803051cc5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3a7f0c95d118e1edcf62d70b1dead4df303a89f60a7d098475b58493494d22ac925ed0444fa507a8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb0a8ce32d2f812122291b90e58ef4a502257c8ddba51329b63fd86930e8e47c7a886df973a0549f9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he248afe4aa6b5b3946fb1da34379335f43913e26284bfabc14f193a03f9d6e7c78bf2cd4906dcf25c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4df55887ac94fcc8cdeebe6d5c2cc40b1f77d5266a6422ae8cf2693430fa1c40ff21f662d0eb8984d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h285d3d7e713ef33fc0450c899427b69df06b884cc58b37a534f4782880cc884c90641f1abf416d79b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51e314bad1d60ef02276c23871e90a53fab4541f173eeca1748f92f2be5f375c7a4aff4f67da25c1f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3f7417c992fe18d0d8cb06d0b984c394220fd13026208af6aca9e2cd33693d48506fe49e48a63769;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5bed5fecd701e1ce183a47135bdea1a6ba808b2ae82ab858a82a1d51a6adf5a53203b6983ce0347d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27dba5c1e68ceee236b3d18dcee685c5b08afdf7713b6977ae7fe2da994b5304d98a4434ad36f08fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b8cb2164703d610d3e81e6dcde3ec1e71590725f7afdc13e8a40295dc487a71e050b74293479dd3b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50f0dd3dabdff83504e7cb013368c9538cb517a61d82645037fe5ecfb34cde21d8d55d167e09c0326;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf618bddc8b79d1f05c8f7136ae0579a2e5409d44a9818a94197741b815c1956520ac1669a0546b29f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15846458ecf4bbb7240828f61272cfa08f2776f436047ae4432eeb9154416298240946e9c764c64b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1789e578d84281a018433e56f893054273ed6e243b38db4ad6d7ecf2c98665a006464b9d94a0e66aa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b39a7dc16ce32e14e07437c6163de94f1e20b139ae5190e3c87da5b92fea7a7d237ec1af3d55876a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1176276205109716a480370e7738f07c54cc5fff31f18104d9429863e2a17b6985517117fd64cc434;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb536376438c7b5cd900982c8358f087b4a864787130d44b546be4a757d5842b6c7651f71a0a87c95;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0148fc468d9c581882c2e71fda1bdf838ca4c8064a81115a3eeb6f688be9bd975b8bacdd2e38481c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a4d61b3898eed1e84c62d0dedc4dd8fb83d819cb1a7707e1bc1782c187acb569eb119fc277dbe782;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a1b6ce8b475d792bc0292e3b599dd824ecb27f3b6e33e144254c39a4e35de30a5435c8c0d395057c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45e18b471374ab2adade88feaade23ea9e0a915e2b008030841eb0d76c286724e39fdd56c761b3055;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93109a430a0962dc50d886dc9a8126c5f9ce3bd2d007a8f0f765139aa9a5571a4e83fff88d9307fe1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3ae69794e6fb3a94c994bdbf95b4a8da4b5e43b57b9eb4f3e69047e955b313c9928768fd5ca5a8d1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a0d70eec3f40bcf81b2e535231b17e3d1eb5bd2f0a88f54efc8cc43a59a7951f5f917ddde72d3ab2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h631c21f5bc37757a212afe25379fd28024f43252008a0293e1f5c8e01984b43b09227eb1013cadbd3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6c828e5658eaaeb3f5e093c924e1ac748240de23e94ee7af2bc01562965c968f4c674f9a95bcfa8c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52fb71950ca7d2f34a8ee3eddcb93df831168b9da6b299c6befe171793e9eef1081f29971efb137cd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82c41064c1b030ce1b36fe7735f64115172869e3ffd8ed29b76a0fd0041b40dd91301e41e5796bc5c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d804e749c7a4635440bb3c1f1afb3cf9d29228a4fc5e9d7d8fbda5d87c25586818010cdb26ad729d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h246b0c2bdca1c662a8b7ffecee880a78345bc2d00030ef7b48b9db5cbb8ba641990b24cde777d239c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b940fcc2169bde22e5b919f61ffeac12ad3b6d7110d4da7373326522e6489181b1cca2893bc91b46;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8be261fac3230b17107305086780858c080468ff39a2d54a0d889349cef2ba1a9f80a115cad9e33ad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65bfd526049f6413604b08d4580384b0428ec0f3c6f66ba3e4e8e93960ad2938fc4b49d3c6dc9c5f2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha52ec93682e4e43f726f31665be967f71eb3c41bbd47564ba5fe7af5165ed59c5de3bb1db6ebb7316;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h870c5a435391e2591e3c9dfe2e004bcbad7f350541e2c7ed06fb4b2b78f3bb99145722f6963204c1a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec91d02049f6278712d2af28ca7374a9d9f446cd7dc201f6a1874f530281be485004dd36572fa192a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hccbb64431ef363e28835f0bc968eaf4749f258a9724d4aa3e5b8d4f4117ee0d0c4d0e088f9d9fdbbb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51a34abe583c4093d46f7bb0e33f546ad0f4d7a160d61c4c84c88a3d0996ea9d70f8109c629ffcbf0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdbcbc07060f182812f5674d950abc1e36d78b9f8f5fd74993195cdf4f8f3b3c928a95c83ae93eff33;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h469a866a95b99478f42a9b284c889c8c035b41aa1d2bce00ae749e2e5d64c245f2340c350aac0ed12;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h826a52db14b152a5599a4f45a0e8d6e62cd977637f6c369d29fef58e713eff8dcc7867af9629ecfff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66bbdddfd0c3bc38e1e90141c636dd1acc5ed79e5ece2b4538aa8e607dc533a92a3a7d53db3186ca3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7a88c70299408d11c842a94d91ec03ce5e1a2c26c4a9d0925b37180079c6335967b77f104ad385c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h102d81cfee0ee0686eca6c572441ef85fd40dae089cdb864d4fcf22406db2fd565c6658387def472a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h113be11b85d231dc80de66db415080fcece0e510dd38044b4557f9b9cdde2d632c15098e24db7cc9d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h666aa4f87fbdb876fe31ce1df856ee32c4f983c568307bde0133eecffe91bc2b082b8494a6619a1c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha926577907b29ed69e61148bf1a9d743e09897df557416c388287894119bb0d7854fb8d7adbbce68;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9407bf075da2bbfcf37979bf9664bb7aad545c3395a8d42eb769f74dd0ce34605d721da66a56efb84;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34c015cad31636aa352d2dea46e84294763188e138a31c24251485266fc1c06959595ccb183fc4b1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab3828d37a14c2383a5054008256e337b687ebbee805a6d4008dfccd8fbb27adcc11adce060594a25;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f457b3f68ee60ea5e6aea83de3bae60637d30b862939e27665deb49cfe636a7b6cb613f140c433fd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98a036da248bfe4265826eef217ceac74a1878c380ca5b31ed63c1629b5d0a55bd69155311fc48b0d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc18050d7e8a37c583f2ea9da23f5cd3a717c9c826ff99ab4a93e12cbec0af1ef6f08c1383b02da0c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18d18a70a2c33fe18eea05758750ba2669b0a54370c43a5021c6ed17f9b65fe8d4e7e6fc2b0fe7f10;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c01264671fe877b3cf4fff06c1f9e2fbfc2c3648a512ea997beda55c3d38e61af2224d8cec4aab05;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e905b4dd2bb4d6647ab37307301070782eaea4fdf5acea9ad18e7e0160d9c04ae1b34ae174802347;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8109e9680592706fd9797d08fabf76d1e80b50eabeab6f8a67562b4aa75b5419d255fd7c2dc5a0f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed096cc3f9ef511721cb4f873ba554bb776bb02e12b75985cf68155e443ef8582b17d1bb470a11b5a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4d2a789694d23a27315b51af54c02d4c2998328c7914b4164a119b991dd67a15f0c0edafd478b264;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87a88709bc3cf88b866ffbf9b74b6056587b0c1308bfd674bb0559b60973d23bd32345bdea7bb4860;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had5649f0dbcc989181fe01b95e804827854a2f12457acb6d8eb661849a0334b3fe9eb2691a67c1e9b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ff584614976107f6437c3b777ba1c842266e6e9b7b4e17b7ae6991c8fd493a1cce9f8e5f2a0511ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he560f353849c7893f7395846a0a6eb6bc70f0ec265b8bd350d00df86713cf86ec0aff4e46a6e47690;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe1c1f9b7ba8f20c8f9c0cb79539cc99e5f5b3e1de0e32fe5b811efb2a5f61e5097d548b576d70790;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27a5a9424f892ec974d015cc7a96a83d3f470414a60c300aa4397b5e5fde2a311231447deb716c9f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d04a2173f4fba04a50043b38623f74babc496de7a214baeab4f4dfbb0ec4a6ca599e3ec83693d7a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f8a0700ead893bed1d374a24efc9d7bb8dc04d6627498755b99541ab25b65fa66facf28d265bfcef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb5540e345dec51e23feed7ad75b3fa4207490b1c452023d8bfff27cb138b23abbc8d4311ae48f82f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38f1e3f695bc59083ec9a4103fb8d46fe76efc5c4b83eb69d7531e88fedd344ae83060b618dc8ebc5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heddb1b2b1e68026bbd4074961503459ac710543e27a4593d9559c6f5e15fb346d9b8505d2742db2b3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e4db3de3183302bfbc4e52949731aa5cd6762922dd7a5a7ef10f397593cd58cdf9e301a1680c52fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1cd7c7209fe42b2ffc76bd93f572fd9038ed5e077bb97212cfe9efff4f28b5919782082c83d96b730;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb1b7cd584b760716daf39f9a760bf2dc02331c0fb28da45989ad2873449128b2e3311dda216a29a7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75228f101733617787bb966059702b659a423490330c76027b237d8d7f5fff258f01e6a1c4e9d76c2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcd3a3fb9a505a1e082dee32c1e594be476ee58a0f15672a4b06732fcdf44f31ab29d8e9ea0e1d4e6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h954f9ef6fe0d66929ef016521a151e73f7ec3ef65a93e5a8517bab2c7988dff4894f70177b9cc341a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0e99309c376f618b37f119ea3a0e81b5ad9e9726c6577da62e1318d3eed9949bd207945604b8cf17;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a856ace55921e3cff77eb53f38e8e91674fa24349421335c66c08917863cb2de03bb598bfbeac538;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h736049d308c854b08b48e1620cea05f58c2b37f24f56104a09ee457e490341fcbbfd7d3b05a648ccb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e9a0fa45e0e5a30c0f3e8a848e883505f71ac926caf24ce7e4e812efc35bdfeff1a1cf829ad05015;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfdf99b055156b99b31a69fca8da7d2462fa24591a0ad7a6e3bd3b7872e0b483fbf82ab6cbe98f8093;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1565aa88e25a4730992ff1d82bd9694adb14b8fbe24b5e496503fe2c8384a644257160ec75f3c87c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha04bda72ce04dc9983e4d7477dd5a332e4003c1d2d83d492e8aae21e81b63a3704c09231a7c000bf8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac7e45334a2d8ebde1ca4b897415d3b4eabad4978386cd598a27238f6dd7c0c46470fc956e034ba5e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6be1657b4fcd00894f0e7cd75caa9384e78a2a1be777a720cf05f8ebdc473d509b103b9b9792061a5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haaa4a1d7bc082002ff1280dce3b0581ca1260eb29b70bf555e1c4a96172c5eb2c7228953aa7136fef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5370175f0833f80e3f26a17aa6ffb1e35ea782d352b8fbbee5697d9651117815a8ca4f615038d81c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb42d4a3988a6590ca87dc0dee7e1a0ce44e46d59d99de1303ad12b22aa13588794520f00f7a913e22;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6664a35e8c6c04a6242e5a567b1cf7d0ce2bf6c17a859015e816ea19dcb79eed27042593a4c5ad438;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7a1d44947b57cb89b08a7c8f389d485699b53c0046217828676889f422269c76ff61af16e1b77529;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h902867793ac7a934733463d32b5f9d466df8693a6307028dcdcfea4b0da6032c3fa5d0e52adb15ed0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3207300ee455ec9d4e035d61f789465308fe838955b45a944575c39c71fc04af6fb9cf29477b4f9c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b17ae865c73246c8d0aa0e93b8f41e4dd8ff417babc4a30251e62edf3491c49d6c144199fef8c0a8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc926493d232fb653b50db187be10ef0cf3686839f9a3e28a875545eba04fae11a5d7618a29a157f8a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c37389dcbfd29175ec69fa5b1c4203416f8a98097f7da1f8c1fe1fc745f808b7751d905ae39591b4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fa42f36c3da08891e8940699c06bf0b8c48a0145da9a3049b97c50ef27e81d56e15e3b515130a074;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9f37eacff5c2e900644c309651b66311f62c0f092809d05e774a9ca9b3d3789cead6d16134d13771;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61dadb97b3e119313ab2263d5cacdd9510ad7ad725276f4da757fa790d54baeabb662e1a14f4cb2db;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a03c6354c5c2910aaa385c96e8d5a441c6668a935190a2a1e7662febacd43b5e9361e35d730cf9dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h854fdcf978b65d7cf52d9da234f5df10f2d224f5e333345d235bdff6f01cb55b3d1909bf36c3aca0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba92123f85bc05a24dac5270b7615228bc1c5a1dd5f34327b96e57910b04f8cf5cd321cc77d1171de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc04fd58269b69c0f835daa015c60a0a010d0ac21695ab9eac99b73d00b87b2d826e3ddc0959852c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb30583c15fa0da1e0aa3813990fd280e9749493770261c664ba4ac72b073e8e095170cff536c77256;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97c24e6cbf4f011b426dd0b5f43e8119449972bb6020dcd9b20fccc60b67e3c36f6c472754c5043ce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b069dc688277e8b118c3a40acea49b977b2bc1d6e37a45b8b614921e6f1f26efd5ed16ddfdbd598f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6fa69e0ba7f41c20a916f599e553caf63708fd5f8cea3922bc35bc68008e7cfc80c185256f5b6b178;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c5624387c70975a23b355b1c34f60d2bb7f299c85b64e180473d9fc060af214b3c7639009883c0d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f0340ac5ce7a6892f94ed71c3df55cca9761fb95b0994fff9a27efbbf7403d5d0812764546aad62f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8de700b5ff178dcf461ba7c827b9b6c64a21b3d50e1c3bb87c20dbf0ed84ca2b2af971389d4dc95a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he13c52d9ee4b8178f60c283567a79fb825b570f147b9f55e0ef1050f90e134a45c9c2fbdfa8deb943;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95986c7137c049e98f27d00c1871dd4cdee30c30475c26f5789861138a74e14daef612a4d39ac0284;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf992ff748095e56970532098993439c2910779e2064304cda8e2a477b721ed46891c435a681a1124;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd38ef56486a8e277575efedc9343e73e948b456c5a455c3b79122562621f163edfa552f4efd09ad18;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h197b0d9b53756b107adf7ac053e5f8114ef7bb90816679fd1981f1a290ba7eb364e4a60da80d708d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e26b09557607abd5d56a7b0c08b1d16a852bd40fdd871f39990e39a92230f7e694b473208367af89;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5cde061688defd008ea33b316d29e4b7dd6c80fa77a7308f6dc0aa5beb57c4b5350f1c069dab049f7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h499f661b8a50ce1b8828fd155c6336d288b14457c52dff8d4329b4f1700c8ecd8dd59666b1d810f3d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h516aa5821d2b7551bca8f48a0dc8a7b9a1848d9dfca513811b8c75605739fbbeef8ade533972cd522;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45d3100bb2c8e5b0dd1e588a515443371b80ab6306d5fb10aa61bdc11ca830312ed96896aff57eca5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7039f30e776f9ccf4a3f23b280532c2bcac108abf65361c62301519a0e8ac6347a65ecff503c5924b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0ac2d51b08f143c8342d7e468a06e3886c110a64b4d2c3da243e2f3eeec36f213173cbddae79559;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e63a32c2d2fdab836fa25f89cf2c730fb8951d7f09151507987b051b0c6995cb2f9781b8f86c606c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99bbd648a735b8b112bb069eed0c3ecbc037c49446c7cb1ff307a47992a0cd81e8a6b55ee755aceaa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac1588bcf744b420d4fa23a35183bddde6a83fbb40e839f4dba6ac959802cb0e1f04b88b5c59c5373;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c9c1105457ff35395e17e8b96d03192cba8b7a7e59754e7c317c61b4fd35321dd751cc9f7ba375f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h574c4e111e527b26a92b2b831b5689950cef621c45764aceae34ecf331878287daf900185404671e2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e96c742eae2f34812be4bc2a76b174e262284427333cb6d85fe316a4a60425a107520eb7f33f4944;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4150da1973b2a2d81924d8a431d70cc6d778257c5cc8cee0abacd5af3dac9abec14c334cebd626be2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5328837756b413cab4a04ccdcab83f67b4754166503798ade19d4ab04c28d364adf58b77dc375abb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha07409c44c66226e43fa313bd28eacaaed821a72ae8827737dd3935b858a9a2fb5564f785753f3e19;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ad1b8511ea23af7b0d9c699b09ab22cb1ff87324eca0b70813ca57466b4bf079b08959396fdd4049;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he099dbd2e85e8eb828c865c43a18f46855607f8be2361cd496fdbef2577d099dac998c838d4bc4489;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ba20ddfc98597c75a2073a8edaa6b1009c39d2417b7059dd15a55638a48bc9230717845d55f2d987;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd958a8c489af0918b8de1ccf12f0277c526f9b3b3c455482e5d39b0623cd6926d39989b638ab8214;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9cacfda2c8b0d2586df8991752af1ad4f6e06fcd728b8d0c7498268d8b03ccaad73ba2fb58650e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h154ebf18d14d9fc67845122a1223b1ad4761b6df0a5a3e485ece71a12d917e64975dd7f4d42035d32;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90c36f12a14ea337ccdb43a8a52878223474b1b01f943c28974dda2d37519d6d49f6457303865685;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32190aabcc1d46f72329386a57d0babd1bdd4f56d63d0ea155b847854cded550aa56012c9d75d5b3c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd385d55936aab91342b5fa839c444db0d1eaf6407b72787e14636483a713a6944aaaa8f734f6c5e34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hebf25755baedab6ae1cfced84c3470bb7e09fc58d2744f72e70f9220a3c5caf53420a216b4911edaa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3c73fe6e14ee27b966527f7591d44eef5ddcc5f8c2882368b71c7037493aca4c442727e1f3300879;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7852784907fb4308694baffdb628fdf1a7441be4ac96150ee49536bec04ad11a72a0d39ea3570395b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5a706023cec539e3746afb30fb99339ca13d3b8bc896172d6c6deeea7f14c0e560ef77ab10642dd5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30156338db6428fbf739ccc1a26290e2e8b186ac8bb5d87d9a00a94b6a5320c5d239abb4c952240d5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h25c19904bf0a86b4626d67aa24299e6bc612c5e083b5408681c66b558a0e661603cb0f203eb36971;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h976fc282ef2a2b16a7d1fa57d139248726276fedb5e24b71e42f1fd6d487a3a2d7f0aa3ccab0bf0e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haeebe1febaf9b36b25442fb82a8b705affd4f9d3edfff0ff569a85a38666b66bc67130ba2f37bbf7b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6c10a74ddba9c53dee704f910b421eb7f99d00a91c043b6da492f2d7b8671739b9c8db5aeafd253e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20c8af800c8f0255268bc09d2b27812e8bd66d43c9b9cf71a976b3d402be724bb8c89e5694be22565;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30d8603da6a4a95838aaf3898495f52aefeb7b25cd2d45f654ad64d988a4689e4e5d63a0a2c9af1e3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h309bbd72ffc93a0dada8ad8dc2dd5a266953dd4ab68248cad413929688acbdb03f5f39664d52b2442;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfba2414baab82a2dfa6d5e10d165ca63ca440d4602398d8211b5e810baaab57bbc90ad735a28eed5d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcdfc970021f7b02366146025ea707be2c1c1e911a456a44c67a4d60f44795a676e739ff62017a9cf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87c8d5272c89f4bec4b39d4c35ae49da92a98e1d1a7d92eeebe6b5be8592b09a6f4ff6d0dc81672c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9dd13ed6bcce6fc1db5bfbb67630ebcbbdfda41c4bc8d281190d4a982a8c2c0eaed1e1d61bf095fae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b115cf886ec85748379d746db0325c3d7686100e4f62559b61703c350f79129a973628c6992289a7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4ddd1fb64b786c4b824f9080d7cfb671554b3ba13d5588723177c5b98b8f6a4e87e5e05d606b6f0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d118f0f3a457d73956e31f2f556f40bb8d57cd1de8ca724c31a78af637f607a90b79c8fe732cf45e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ebff648c6ac20691c21ae6bd2ec04033ff6a6178507c71f12f917797933fa0b8a50d196057e9b2cf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17b917c27720297ad1ca4e8761502cf23a97e7e996a9581fea0ba89ab225cb812ef825bda42a7b295;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ffeb950f0919e417e25aa2ee261d13e0b7fe601126e7ed9227c35fdd12c4d93212647ebebb32ea6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h133431adff6300f971be2869fac0420dbc6739f11fffdc03aa1fdc4c925050f083cc04cae5b850387;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h396f826626333563e3fe6b5cc41699ee34b449e85a159192f269516d68ef1fc2ba696967038095e23;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e0776bc20674aac50c89a134d7f3b239972cd5365f3b854be92db59079d727a0700acf8bfe58525b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7aa8bb49ea8a07eaba3fe28a5b4ebc148802fea76eca102f0e2d2fd802cf9c2188e9412598672d817;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98aca101a233ccfc7faae368df8904ceb4c5640fdd6fee24f2f669713947b8ba66d527ff7500de639;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h204669f2619dc8ce377e7731b561447925b4f0399caf2ec6613395c2a7adaed3a0c2a206693f3ab86;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39ccf1a8c6d315d52f4548d3aa8f7afff0eec4ec74594e5c543cb63f8c40fa0d092d25ca92c3721cc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36fbee8a62a1b0cda1d04d2108b82929eedad1468eb4d1733dd141f0783d3aff3bb4acdbe36dfc475;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h171e3bb0899f509b6f3597cb43132116d734b9dc78b2e384f91f665fef81ffb10ba4e57fe225ec148;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b475cf4005d6d57cee6c71fc817a2187bd7f83cf4b95ea6792c2b2b45501da09d331be42f04514fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e3edff254e1a8bdad972a7f418d9d7e2968e76aa99d985e7858c35fcb7bfed9f8fb7c24ac4d7b86e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1cf1bbac774810a4e6c7a93a41cc636d3caf7866756daf03bd0ff1c791fa75ca65c3a3df4f0ff933d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae93f4fc1cf3e552b0a73b1afa5188104220335a0517e6f500e94da9ec233b9b31a0d96eb4ea5ee60;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c9cabdb9da66e9888c106a9569ace6577b90483dc7b60150aff72012c8f8fcaa0b736d06dc1702a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ad93eadbd9d885e118c4d73016f1ed0d2b28a7477644b117b15d1f708ec03d57616114f02053eed3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77c62b6650c20452a01250a728b3d152eb483ad08720807a41977dbeb07c9e897ffcd98c7f89c5c87;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4cac82b87caed2f3b23b5cef65cf3419445bc1c01d86104964086846d4611e7125103d4b30701d02;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46a401197afd573fd2d5594f4829ef54197eedfdcbc2feaf6d59bf14cbd95ab129ec22c76b6acedbe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb834a1918499acc8c7fe4b02785a7512f66c2740828b2e8f5c7df9084e78c55e066f13b0f14c7e637;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haadc865f5a92f1d1b30b17e607828d6d1124b79caba01c7e97f0e9444c2ee6d61f1d1fb230f919d36;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82023e0b9937d349002c792405d69c1c59641b73263d864e3726ed3a012983fc4620d4238eb2970b1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b1cb8ad6a21e457f51143a16f2e82fd57a366db86918ad89a139bef5e0151d35439118519c1ee3d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f1ed698400de5b27a44562d3a23b14a351911991dd5ae39290148960bd051ebb1ae6643247b1b22f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h828268058a8d473cef62301efc04063e265ee5ad51c760ea14c1b52ccc0adf8cf70756eaa0052852f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67a55dcb41d3d6769c253701eeaf9c7f4977fca43e17cdb99efaef05f66ac6852cea178d45178b103;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h378e18a655a44f04779b27a3aa6692dade4683ea9822dd759a8e0a69029f086572910512b745da06c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde2855082ab52df66084c8599bbf862b5e21a441dedd21389cca983403fa79a9920477f14123cc6e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had9c7ce04d67ba9804378ea29d67de18262d8bc1f02c9b967d15f48fe482e9aede5facdc156a508e0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h845f339def3659b5b3549937fb074e18e30b2abff91bf25802a65a611b37c1f7305c361bc3da0e494;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed0d2b88413eae095bd818385c8c1e13cdb44998759abfa8a7f886c87d4b6de95a096e4c1b02d8f9c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he67e26a65e1c5991a9bcf26e7bb33c956f4fa8181b61b524996509c744e41447c77e573272e5adb85;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d781fd68946336a86caa447c1bb222edfa10a7e0cb6dbb7d271b774b6890470835d3a2a9d9479d59;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57b825dd290505e011ea8ecf0d3fbd1f66083de08565dea92557504fd8281e031f4304300de10e699;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d9bcff61bbca7ff8775bff3cec2e0a8558e189e7ed9fccb27af39eba02a1921fd05e746a874a4fd5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2623179fc1b05d3ff8dd33637fec32304393b610d2baeb25985353c62619eb8e66d4b893e5d7cba6c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0e4a98adaf8efae7bebb8385ac59f7f853b237272c2258dd6a3c246126b9d41b8f982b3981055937;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7031ed30ce338c7c5314491bea39d07eb2986a8b76d8e826cb99a292a5054c95993cfc7f2c6b7ac3e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdf7c9652937a0d6ad83cff7a5a3778acb695930b4d5fd18ca6949df2729434ac9bc03c1e2cc6e2933;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc9c813cb66dc3d3cac7a4dbafa22e153fc781c55b8094b23a1c0e6cbb2f6290df432a7518d16bc04;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f9c4537936eba33a6912f1ccd3b7e0dcbb26d8b24ada51933cb54083390c4bb660c4bf41fd2a0f91;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4f6f618d72f15e4caf17b676dc9e57169afdbd2a20e832d4622001ac1fbf72b4efb8ab94e4ddc0c9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2c799f64c274ebd5f20513b93f79941e294d3e680504774ff608575ea41df5f8b466fa5e0451b589;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha61e4c12c6d7da426152866667ec7642d71c6df60fe5155e105a4039ec6f1828d9a18e16cf1b23987;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52fa9e1c9ac35f42b2af44ba3b231c09f869be527c3b231b09da82d051c9fed13c2f87431a12ee279;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52b2d8ebdd1dd3cda5e4f1cde4756b9e3c56ec36304a8d73bac0047ca43e233ca1f004072a6df690c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ed49f8adc601166820af3b7ba0b249ad23ae4f182c1e1191429aadc33416b455d280b14fc0840467;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h972205145857f5d546ad7fa3ecb89e70c3930e5375fc84f628a14eec2b06407f73b7e9b35c14d7775;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2a2658cd10d5916147f8ed7545b16f8ed41bb01dd0bace9824aa104ec020f5aea0c25a68bc2966a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h803e9b12f14f0e32a35414f56e3924f2eae38e6538b0f2510126ade14374771315aff9695dd38704e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99559bdd13914c8e7ccff2db9b83973775f05214406c41e5fecb21941b69c617ca952343a3ef30ccc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5799a28849b4917abbc8dcfa1afe1aa5509cbf3a916df7e9893f2a6a418775db227a7aa50308ae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c9a6ca843a574cc2af00ebbfeccbcaa0fa721c49fd57942179d3e5711bf588471e94c7abb311d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8890333e9fc71910e9c348efc8b81ec644dcc23014d8760950a97ad429140fa5fe4d06e2c7610575;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha126cf1eb062bbdcfd2dc3af4380173e706884283399b2c7f7473ff348d48187369dbda03c858e453;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h182848c9a9eef21678590ff6f2409f52875119c8ed8f69fe5d53b5e053b5b5877f970f01e6d62a669;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf8e4866cb57dfdd1bc6998570441cc0c271a0dc442b67bb70d4f850906419b434439ce0030660c34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9786268c458a79a594e438d83695daf13baf568ca2d07559a331b90f6a8a29b8416e80ffcb2d15fa8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f2cd2f95ba109d6b60e65d8d2ed6e043b34a90b8d113b1b7d57b81ea862822d5cfdb4a6cb6096805;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8772aeea42954b905221dc639145d8b965be622be325d316e8eea80fb20d52105dc3b9017f29240f5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d48d1a196344d6cd300ab8683b2398cc77e548bc68fad01d621668fb331d5c7b90f433532bd698ae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h816d95d4308635a918a1ee6311ba1ae04e39d661420c47b6a0da67a7981cc07e64bec67ebc1eb2b33;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h240047e06e2dbed98cc42df29023dbae690f80d04871941b095078a5935771cd852d408f69a57cd52;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c65b647629de3679e936e1f0a90947ce2106626c6ee92992e64733600b874cacea302d0155c55f85;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9257b85a1f683abe33be16978d1ada8840d94fec7603881f095faad804ef949452b8b1e841dd10492;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3f8c3af84d60896f533d7bc1731380924a09101cf5517000de165d69aaf6e0ff46d56cc7a668cd42;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc61ac8464b5aeda459e3256516f45a574a12e38647f4c4aebb8dbabb08653500d12dd50df6cfefe58;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1dcbcb2efe6c7269d985c59819d6a01e7b33d2990bd5a1f5a33531b9385b703ebb09dc416eaf14f5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92f265fc64dfdea17347900940ce2bc2c25a81c5e613de21c6342fe9451a2cde480da964caac5e298;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9df19f9d02d31dbfb1ba079594a3eebcc0dbb32ee72ec0bf972f5b1a26b1939be2a7e6ff81825628a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbaa8dfba7e0ee70dcc07ea94f1f0dbddc46ede121e754b721c886f24a186ce033d714b75f6a861ddf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h507f3e1b4ac26deccc139f8f40fe70a6d4adf403986471eecd8bf0100b772cd299b2969ada4daa8f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca2fb30188aa2dfc2ae643c40c9ea04c1b5a98cbf5a6cd99e4488f995d7c88427e0f09d660bb25e24;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d2d5ad60c3afb6b825539b47c0332f06d86fb33fd0951ff647ae651b1ddf7d522648b561aa980c53;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef2048b4b1b2636b5d08ccc00bc19545da19c985e17a8ab0533754795670786c0100d9e93d760f1d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0970c85165d3fdd84a9d19e2146009a7543082f8f882ef9bc0197ac44701cba826f7025eb30cbc96;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36cf896b6a67a53b096f8ca951805a5658117f7393ee6a56f25276b8a23f44101dcf9b0efb702d449;
        #1
        $finish();
    end
endmodule
