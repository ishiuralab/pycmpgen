module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8a9888e091713a3abbcbec2433058820c328c18d7eff0c3a2f93886dc2b773c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6ba36a93a041e3c6d7eb3a7b9f9892ac64dbb83803f66f4ec81520aba35b71f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0c4763f7f4694c42085209654f8a6fd9879ecbafbcf453b04390c6c52d79de8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h79f6a3b1c0545ae569ba72d4ed85ed35987d140ffa197ec731db3fe4eb9ccd70;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h271e4d74acc397a2a23f34fb03743f78475450ee3861edca30ce16ab22babf7a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab4f503ce9ff37f07c7a88f178d94dae91745c37d0116108cc75ee48cadc96ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h990ed42372d7bcc6cb4361d707c463d4fe3acda5af80c9c08e2655ff9500a6a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8899b9a243a42f8a50b831ec060c758977e378063151b2220ccf031a6fa47ef6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b653bedde350507dfd6c093a2b1826fc3e61ba5f22e033a9f1fa96dabc9e15a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h82c778b42e053e6df5b10d6ee2154e8b47aa020b66636569a3a4e4325e374fc5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4f7b79c117001a4ff37312273f2c7d54b45c27badd663df8cf7319c72d8876a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24a227473f4373c534020ea7a86c9429bb271d56b779a399e63ca1c4d743a4bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ba50857e449e9f9e7b9f2441b19ddfb9ed6bf710a09b94892c6db5b2f6af048;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c6aa121b75eeef1853007e5364d5ca1fe04d7649d8e8d0565978161e82df50f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46bb119f80749d59e1e3825ab95c8e7b878d13277cb10e3e2cb2ee87a509e87b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12b4137188b6fe579f5d1140a62d3d1bfc40b40e3bfd8779e14661cc1487f5d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h27461e71e2f0902f71c92568ba6cd6314c3ace32cb0cf3cda029a17ac8d1f388;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he21ac0efc6190dfc134e4cf2bcc8b77a7ac6ff06a1f316d1644be8ed302d1c13;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb94b7930cb4ca80c282424d62dbb3d7930da51362bb73f0634cbdf79491671e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa54d27afd88f373e38f8f4d99de50ce965ffa01847ae17b77809b1bb1f93159;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31030c6641efc122c5d1203629266e35e4932457ce1e0bf7d0860d9ecc77a682;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h305082c14c06dee53b344af14196a9374bb0f66e7200142261eedd7ea231255;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc184b9bb787ba81124482f7fdaf746e57394392ee29faa8ee3e7d0ede91e40a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h90d09d3e7ac011f76bb5ecfe8c04045ab99fdf720f53ce94d474d290379a254b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc04911f340299213e2222fbde94b5d24a4bab026ee5de489ae1a08d50045e304;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5ac18bf286de41c179f36998c65610aacd27e741c6f32a4c9424a9ed69a5502;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec6acf9f42728ca3f08e95a2a23945f3884202e961cc2dbe6673532f5268955c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h348cc656822af7ab4fec387ae81a7186bbb46c2ce01dad3b85be3250a396a50b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc267f6bf985a801c7e3cd7cdc45d6c2b6b07a43396944e859a8202896de88402;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b2c2783523a8744af7dd8935ed9358059f3f1e605a7d5a2f345729a6eb4ea51;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbfdf8b2faef771e5f79ad6ae12279f54c571c67337a0351400acde85130d9f46;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h245011593db7586cc928a9e840c3d6a89007e77268f89641cc553a981dd974f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a721a1985860cf77ae37b7711df555dd859b42ac898a6ebc1c4d2fc99c07f22;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6b4527c3a0c7fa69d5124bf3e0fe5f0ad65dfec14c6117c76e9dd6a39bafd96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd250f6a6843cc62f7377e67b3e5f99e7316891fa23ec1109660af7a45c42ea9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f2246bc84699f28d2aef6282e60b4a1e20d3ff48660ba53dd4e0b625861a0b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd084c0f8bdb965175210bf2fdcdab41b501a11546cfb2f9c53207c8762758206;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfcf4ecb32ba7322d6aa7a70f5680a14872481c8b9feba56b7fc9add23b870a79;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h446c0a68e3277e19770dc9214d35f53783ee13b75900057af978ecdc23f89d9d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73e67d3beed24e9b1620a1edec3c77d232b560a5d86f5b649d347690bce6eff6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb84e6ab3e3d39d666ef87b1b2971fca36b1779b3e0c8e2bf26fbbe9f77558860;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h91e63e347f42f3dd9e5f069827acf72a4bc99f0db5185333535d5ff5e2c7c9c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hebbda55cdd9dcdd41247fc0e769ec068ae6a7bfd646b0b302ef8e74fc971b596;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5aa507b41c7059dfca495bef221df1f85536b58f4c41c7fd816cc5ad6fc2e2bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9288f41be3b2c2fb3699f82366138bb301873203e420fd16038714be50674a08;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7dad73b33e46d9e1427b934353d61e5b1200e2d802a82bb4499fe51af35337ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7bd1fb5a5ac7a9f203ec7b02733726b681d6b6d33618c81e5644334c5f7896aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h985015e45f8a3b36d20d2e9a924401089dd756bb53130285dce880c7c8b1d85f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ac0541dc5f4e8c315f31b87fd3431f38dfdfb42cfc4d7583252be483ac3073a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7178b77526d9123f1ce84116f5800bdf1369626c73d469ca50a6e682019de09;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a472255be31f9a4633cbab2c706e57e9da2eee9b702c210e97e7f8aeca04c32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb660ceefdcb9a4af58f0b0164f267ee8fe6ec281de4ed3b01e563ec9e7b0fc9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h71af108435d66a93abdbef6d4aff20823cd59046f69d251aead79c3e33045366;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha19a551aee722b654c9c977d4035eb64645b38bda6f4657ea3a749bdb27f543c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59d3e3cb3d7fd4a3447057f6647533069dbd27fa3aac516b173c5e630a31774d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hddf84f8b45bcee0411255953e332dffb3bb6714d6dbf04920b645d8fbf501608;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d5533b625edb796b17d77c892a1adbd8d6e7cbd21575481fb66aeb55aecaee6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e9631f03518209719e3d3d9683dfc1c1d91605e460571490cee2fd097f08a1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc3de6ad55170165bd74ff7ae3958dac8fffa4c92e004271f927b9ad1b25c7bf5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75acc298b563c60a0c2d734c2940fa53fcc3da65e24263f13824cfa447da00a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfadb59af51f199a0da8377474fdb7425ddc3c25960f1aae43a06c7264bbed2a1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8dd3b8091fdc9fb842887473c7cc8bc919f67815ec47a00819e6a429fd5089cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h381ae3e4b8f7709625dc923cd316c408799fe85b0e01eaf829511633d54b9c85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ccf1ca68437162c7eff35c7fcc5783895308f84227a6c3838beba5a577eab97;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1179f7f839f9487ec37b1cff384736e967cdaabfdaf00ab43741114352122b9a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h30364a49bcffd904c589e743f86e42010f87335decd5222979a9b2c917ac90e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h85839d8edcbc2c8edd80930d0976122b24f80e7f4c597faf35d12cfab68cf072;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1c07085c920bfd8338ba2137a9615e9426f65327b4de3787f1953ecad20bb1b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c45b2842b02a20182795f1456097aabdd37894bf277242fc5dae2ce1ef7a903;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9063b1eb49cdf5f2c50ad20e563c542f666eb70fba1e6a1c45ca4d26ad1a2fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8994e25a9eb54c017f14c952e9879b90cb271d31274193d77d421b5e273be9d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h177449efd772443d33d081bde0a7ea6af267fc9fd018dd07e96db23f194233de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb021eb78aa72740ba2309f344d51eea381f5c81b981ad416e48cb554dd4244cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd02a5e067a455435b634408e458afa60a4add85dc3c41d5f9d1766b56cb259a5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4095aa3cb60c6a8cfaa707e1562b96654c71659271c5a8a7eea059b395ed21b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45e388609df776edc2ca4911f578f8b90eecedc85d841efef39c036eae768e6b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3927b786f66805d403158aafea6ce7b7121544e2ae05ffce6e6e4d5fd455952b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd581c54d44aeb2c49b21540830e99d258505cc39ac2f4d91687285fb993cc5d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7bcaea18a50571e8a67030796ea13dcfe884fa9a507b6e1f992ab1bc2d9df0dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0de254471fd26a18764d5c15a288cae8c9005a87b02d092c0ce2a2a123259ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4ea3078bab726458e01da8651b6c8a207000863a7e16f69b55c1e0c7d90278d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4f4a60399b4a7a58161cf8f8a6cd730da95e542579d2eac7128d06d4bcbf12a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7264e96061ba249437b172cfe25cbe4370f6b150529d14a65671790fe7889c25;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9c057bae24f7fea32c690d2d74906e76ee16faf22690fecfb9746452f409a29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h374f89123b9a361b2f767953e007aa0a6d4dc42048a019fff98016d579d2341e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf705f28a53963ba3ccadfadb047e94cb1785689e6a01da3f0d5cd8fe1ae3ee0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f3f9f933cda8e39b488bd96aec97b8946e0aad337b7895ffe7df8cde96a0777;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b9a7cb0628bb9c1951f4e3e28f05c439f215c9789566d03270b647fdc0a6d54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h404ea53d598f005de3642f6edbeae542838b0c0d555509cce6999a5e2c48f05c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31e896b11a8e3676c7ce5fb19ab40e1473ff07675dea48c19765457886ecb94e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e735254304aef055a3c79cd6e5857914f84d6f09c4ab11e92f367eac2d49f60;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb1f26b7c433fb184b01ecf68a2d301614da031926a08b2d26013e1ab1bf40d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haff865247876fcdeefa656ffacc7e0b20c6dbb44684b96b6999fb55ecc1c833;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc23de843ff08b82f6099e745ac71acb7e767e34176095a8ba2819a9844393ad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he411f0fb74e4b90fd7fcc12c2a974d6b50e0487e42f879238831d30eac3bb13e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ee651d188abdc7ab25f9b7546d1ad5b5f9c85259cabd4b23616d19f723de206;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5108061c4d8da8ea1ed686e234ffc28900ced428c38c98cc8d5af9edb1ee9133;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5d2e995e72a4849b1d589414ca116518eed2c8dd6e8f270e4603ebff351774a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h432098a731455ad40bbcca046ff14dd1d9947a7388e5ea025ebd9954a3794c7e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb991d2694bfb1a5212188d8d37591decf6405e0202ece20e3aacaccf6614a932;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd5819c0bd548c23c494ecbcacaec81a9436aebdde46685dc32f0d9f8bf5779b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe570ad362171210a5974de19e7208b7e9fedb2946bd44dc6e10c4b6264ad0ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4c3b4a0e1d0f3425bf23f1569251911de25b5654fe86b7845b618527671608e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haeaecfba501fa28d56b076c07fb055842343856d9b11b03cc3167df0edc53030;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae83e44d5c71d54feee8e3c9cf81dfbf3fdb488be0d2e0affb91f3b0ce6355af;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h665fe094ba572c37134b90f413798c642c7c5879944d97673f7b0a3580941001;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2b1b6526c2c92dbb44c23b557b1cfd658fad35bac365bd08233f4970094f0d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h691a4e0953f5a4ba1dc1a1788b85c5b99a8b278ad16db1955b1a6fcb99923933;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h502fba30a2cb6f1e915bc5be6bd844f0b0aa789073aad2cce93bb0c5c10a68b3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8dadaa93a98d4f50f4045f44b1a3872b5f8971afa9c006453187a8bd19a258c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee4044f755eef8f7188f453edd736451701885ee3825895da7d3ba748b56d6e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86834a3e62a6aba874c993139055bba8069dd8380fde1b044dc5dd2ac6e3de06;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1d8d313574c5f44f426e3cacad6a0ed3ae68734471d4b523e73c92d59bd55da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd781961ad7a8bdd9e7ac39aaba78a43b94db59c0cf9b1ac7ab3315d5067b4d18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h879f9b9f6b806cb7c7ad7b871633a21ab182cebd9ea6bc20bbdfcfd2afb0840;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'head57b55338965a2711e65829c647b2e944407415b63c104221d3152e9e3d7e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57777ef18c04b8926803cabd47729ed69baa012a6158b2aa0e84c1e55c9765dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4e0a83b8cc8cf7d27b59d1f398cc93d34e4d9c22cdc883c34e829e83511422c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a3a675502f9246c43bd9922e666175c120f6b79e3479fafecc1cbb774e0a834;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6a2a1b4369f54608bd9f73881f501c459d21b8fbe406d4d5a568151251803b19;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1effb5c61949cb25041fd449f44367166d52f0e568ba971f9bcfe9582654be2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf1ac985ef5dcefad79ab716f68f6c2cdd5532d9ef4db134339c6210cd125715;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2b7172b257e23588d3bd1ee5275d5d5321fc9cbca8ca26625f49892c317a0cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7f2331344684db20f3914c25812de1a888588677c73095d7b1b50624ee48987a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2dcb53fd43ead87a2ea31095ab8e689d1ae84b089c1759a304caab3897e62f0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92ee99b294b9a111978c03075dbeb0600a2dba22902fef56c98d35384939c2d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he0a711df99a4a2fb65d40a7f2f67e85715ead1c890d97380d563e8ef10f32211;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6849e91c4b5bc50659857fb548bdaeeb0b06f321bbe77851647e18363cda279a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc6d500062734469659be8eb07d9c0b79fb543ff299e3127ecb14af57fdb4121;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h922860a426101a94d91f449ab50606957064cfe36442b234192c1aa980ad73d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d36d4512d9949397b7c059a3b5bc7372091a73953e6373b200400c4d4b22617;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23ddbbd72ab741fdaf50d5f82f8dc8eaa00326d66260cdac813ab9ac34f7a479;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46154af7f90dbddd99754d1782bd3974e93e73af4e1cef6c2986fdbf776ffaf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h296d2bda11ac9253955c8c73b00bee6043fec1cc07894ffee16cb2e17e37c182;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f6194573508d07837f0c6756d1abe10ae012b75cb81a6800e1cd8bf022825f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93f1db808ed6db6048e9856cb5475df5d4523c98a09962d2e75b44e6d40d574c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e57211d604b27d7c258ddae6f707a04a125b747eec9fbb8ba0affa41dfacec9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb12be119f2a20c691bf52db4135d831e31d9ed953bd2b4f9c3659f528daa9bc5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd97cd40423ff61f42f8baed1679de07147d00713ed807c02b295bfdf4162aed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbcea1becfe7abe56dff9146684cf8927e3cdd2413f3f6d83f256ecbab84fdfcf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8eb1632f27a12a1a4da1f0dd2fc360978ff5f5a5ea6898c821de042e025d52d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7029ffe2e6904a9160be8d2b10decd12493e9508bcdd900575cda9f66913733;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11e48ba0054b945b2bd08e4725989208fe2c7fed80cdba1d1e9b42da35dce6bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61b81f825f55e3e1a80d1fa9f971beef873ee3bb8474a3087efe610fde346b1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8062465f231b3dd4a7fc9e1e3ff2f49f9b6a197f15f07b0660f326b403595c52;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h991ac142c98c3c113af324dc545e8e54bef81620dc8a6b8bb2db0765650cec90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haeb3042472c0d4db217b64065dde99b3c044f413d806c24bfaeed87f85a2a461;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb80b816b83fd45312f33126b0166fd22346ada669b2982aea03da63aa725bf98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd560b7bd43e896f253a85a67c88f90037efd408a45cae23d891ad1d73ab6e182;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8522a36aeb1f22ff939ba117bd0391274fdc1ef5f140ab3f0b1bdbaee56e0b4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5cbfbdd86eacb05f8c5bb31ce94d3c5fdcdfc6040d71ba8978c68682ff5c761b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d39b7b5c0afb31e06d5d46ed251b53fcfcfdb79e22caa4577e5c5e9704c3de8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0533aace09b352db7ccf8fc6ee48d21b69f607300f65050ecd930c90a4c7bd3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf6f5cb4a4c16e3b3e48f20113221c9f96ba6ecf21fe58f18c43063001de8693;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h29e80a52a474b726dd747e1b1f2944c32c56fdd3e242e3b1fcf67b6f04e9e3a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hede3982258537b516514046015b9fc4a73703c4fbd93b3efed05929112e2122f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h211373ac704ace9e4bb5f330239c58543edac7aa07dfe6d753029d3249b7dcf7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5227914ecee45f45f5203ab738333f165779c1ebcd77a0d8bb00353db23461f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9bf5b4ea558b360b539f45b8faa51ad050557043899de11a93aabf191136ac94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f5bf54a3fdf158250e1c219ee910f2e9238889fc0ed4ae7162cca5dd5f109fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ad015166907b39e9b9e68ea9a8532f0aaab85f0046fec91305753ab2596872;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8eea123f3da9b8178a14a965fa5f17d9557d243113fc8bc7b36516acf1bfe88a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed34491b500e72d5a9da010c0068cfcce844dd3a494f0d1277709f7b7dd966;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33f6b971d67b92c9c2efc153513c02734a506f82b1464414269d3e858598b1d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6a8bd078d95a0011d79b0963e23547cec69ce86c70645a47888fe34a184c2595;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a3ac7ee0938153276ba9ee32d4536902a4f6731107fe4af31af4d2e907b17b3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ef3feb44580692a7a06dc5cbd01b0603b970cd6a317db30bd5d5e39384dd7f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec3ead8e676bea45ff4978eb5a03dd6ee529b5e65c76e6956acbd1eedee40f7d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5d2ed58f338679c606bcfa3b92999fcc2508c90b4e74dca6499f4d41ae1f212;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9d72adf4cbe200da4d4acb0983ad6d3e34aa8c6168329f72ac38f6d3f0d9f99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h647be11c5bd2e5295f26c7f38a103370b5ea67e89c08a1b761b748df5f55d80c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h299d5096563877459cc82c26cb02bc087808518ff856f69f72980562f0da6457;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb207bcb55edacd0599027391352a4d69caee06428916ab7879e9ab3bcfbb262;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d4c43b4123b5deef12eb7e26071bab2b51c5344b1c9a7651844fbbde475d896;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd8c4bba961b649294ad034187b69b3cfcefe96625f5334b60f37439545867be9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h231d9929a1619c6425148a149815641d6f61c5d721187f97f7abb21e80e47bb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h65bb1108be77e40d8953b8bc79163003581f4eeee63f741246286bf770d69987;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h423703c9a307bdca88f8b22c1a68723ece5d3d130a12616cd375721e9ab5031;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd9812efd6b75e66208085613837204fb0177bea6c301d2c26b2d1e58c317aac3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc2ce1b8af9e03d866df80c6a7c37b4a543dc61aafbc5a5726076235fdc6edbd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2447b75d642e73dfba22fb818da30acc50f7790ba05492203e7a3bc33608f605;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9908d415ce8ebfebfd278dc48525f2e1ba67920a86340c03692cedfc61f0c34;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he52db4fbe134bcd1873ce49e4b491ddbc0bb08d9b095377316d91e9a3e5d7aee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9874b078b841dbf1369fe7fd167e0722e2e1858d1a6767bd79dcd3767f511346;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h773b4b357441e3d0d783852d4ea9186f981d2b1ff0dfeeed279f536fe4131eda;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70abc59cdf1f877e8e0a7b11f5fd7e1fde94eff9d9f65c4fd6fb59cffa808484;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h780c7dfd38ca9e2b8a65940a33f751dd8dd0de34902a48c0288f2d72579f713a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd06c61f2450de3005512b90a59a0e371592e7d4f5049ede0726ac30f317a002;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6bc1b7c06debbc99c554bbda66334cb526adec482e5f16e97e7369f4312a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b5c388dfabb84e1533a10d9a946da1af4c85e2d79679f9c0ada7fc522d4d8ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfcff24c13c0044e9eadf85ed3c1b82b7f7a2334e00261cb875337ae6ea444ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he6d02433a5186b933b56a91b6f10b5dd502dc215301632ea5494565669aac703;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h732c89f2d4c8b61c75b6b5c4b041aa48db616120f49fba4d9aa8b44a8b5ffd93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2c933ed599a18c3c37350c7229425ae058f32c73db9e23b66ed9e7aa1e29f50;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e23f26ef17fd7bc233f4f22249f1f89d7ce3abc960aec42afff4c7865b96f6b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9fd8df895b3235f39b4f31fa0ef378675a3195bf4d6147937623c6d3f5633f8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4205a03209918a8d78c003ff96f2c2e06b71d1ba3ba2a68364b0dc8ff758f269;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2fd280857adbdd86e1ebc03396d76a1ec2c3231ff46521358f9a280f86196217;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3c24f7a8c1a5fa47e6d3153dca45225be7e357e7cd1bb50ddb8bbe954644ae59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b4fb3fcdbebdc7fc4073cfc70c07926c54ad82478ad4ca7a23f26cdb06e2d60;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfac5e1368ee749502e47c5f095be576a774064bf7a7e295f63b9f67a2a1c195b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3fcf2c403540fec02f0a7c089418c3db52f32d59e40da747cd52549393ccc92f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf458ff0e751974c265a37e0b1179a7511a10bcd014f6124046b2a7c3b72ee22;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3efaa78492e90b6dc08641013310c45b75ed5ef0248303bd018fb14455443aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc60d21aa100314ac5df5c4c170b95d215a81b074f9729914798b47e1f5fe5d04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4bbcd2d348e57691f28d5c90849ebbcc22e4585dbc2da87bc957ee1dd6459b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9699023feceebae4961c3c06d85c820479bf6fe01c31ddf7145e6a6986d559bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4726fc952ad6caafce0ec17bca1d0fa3e67d8d277da9869ced35f000380af31d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdcde90bd740b6972f92c2a8a79424cdc77628e4643d04e6528d2c0d5de0ff292;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ce3e964d76994356a6a0288d641349710aaeac033ab316facc42ad9b656e0d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1f5637599401309f00cbb307c1d44ad29b374b42ed96db871b4d588c8f604bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b92de491c734d16a2ca22d00ab01843ae6749570749b5b4d6a8402f9717e42b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2bc8e0f4fd913c54e85553a478f4021e591e9af787fc6ea2271437ab2030656;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h722a1fa672420d182551e65f667a1d9397eb82153fa9771e225e658ae6f154a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7addafb413fb167b86ff9983ed2c0a02fd6ef66e7378d124827cae253f9e4e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19db7b8cf2d0be49d4a09aa3635f2a713da34f3a12ccdde5c514c46625479e7f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10e9c982f94a84cbd79e59c3575cf0787c108c172a5cf6b124e58c2ec2a0a194;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h650a5a8887e66fade9bf94bee60042f37a1a9672b3c983b6495c6b1ff86b9ed4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb08bf56426b364970e1a09bfef31562424debf5fdb1bbba94f7a27affc98b56f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb0edc243b443e28b2f63f2087ffe153d8c6b47c1b251fa7372a6c8aa21a597e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f5b11816814f2f52d12686e7a063de26cb2c786fd1af92b17abe26e60f08818;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h16394d8a9d21f6d050f2dac0deb37131df528cdc690ba2c796d06a458d2bfeac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6bad24bf447e0f318d70c27e55a5d90c1d1c6db88029d1d8c5f5affa416aa893;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf27c27efd6b9d4c6aa0a0b3162eb9ba9f61ec37fbabf4e9983fea5eda2b0565d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9f5760b9c1e3482f33a86e978c7fc6851de1aafcf632ddd085c19c58cef2972;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53818a176caf0d1cec898fa73953854f56eac463ca43195cccf42e9f7b140ac7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf763e1a363a469b30424a52c831e6a0920165418e0e18d4e1871659b26406417;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce17d7383a8f58a1afc4f138fc8bc4b2c4c1f02a951970814ea7e236e8c7d37d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd956435cefcd3149060787cc41656b69a51524af61986cd2808c0e2c8e46d92e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1e59d1fd4eb6b5de7ecf13d98ac6ddfaf43ff46541c36d196c91e4770d4d35d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62dae0d0b58b4c5acae115307d045f0277317190d46dcd6ef4bb03dcb97fb7e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb292ebe5010b0f242bea51e09c391cf1e7056dadcf4b10ecade2be86a0c8f0c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e157c2a3c78f43f529fc49e4f9d0b4be0adf4a309300fdb10266ecf71551eb8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1610c9c38d9cb2e25e36b75e0e617666a526aa8b0157904c2e7c218e41a7e780;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d621345ed723895480c2e317c57427b751aa732347651f7568ed8085aaba4fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f89a4847a5b0c76fbd760c101361a21b6c6062e48e87b69e571518085177611;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75fd9a4c74a7abfca54f13fa97a6870341667888780b40061c5ff56eda1540c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e4c90b30b21b408371877ea34079c61697e4fbf1f884d3a35c7dfeac2a4417e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc32ceba7cf0f3d95e9612da53d5aabfa951dfb37885c54964538989d2a025542;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2bc534080945f406541c28fc78edd6d36bfc386534d40b8195ad14dc55d135dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25a425438cf0f2fc862207942c6546d97ce2af4d17946042b08241beb776aa59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94c4b9c81227d74aac76291b210f92aa84bb71914e174efcedd99a1943c126e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h609ea314b7ede325af2997aef301fa301f380d0e43b64d0ce93691c6d13b8ed6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4cd8fa39a7fb908a435dde92327bc9d743b4eea66cf75ad03f52dc53fc770c2c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h811fe008c7d59b42a3dcb3948efd0aa2aa9369a5798212205b95cc527efa3085;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he62246aaf3e000372718709ed9b78541630baf5278ecb17adb68a20f2d2b4c02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda482e18692794b0c1c23524949ecef9cb7257fd1fc727d336866c3b3d15425e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40a331abdff3ab6cf2c006231b244cd991eb92530176fe378df4e7f62349ee8c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h102bd7bdbb018fd15161d2327e8892d8aeb3ea70225da0b9e0a94305f13873e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h507e86817aaed45875087b3b40f8ede0e65a13eb4ff0b0e66b04c892ec9d021e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93723b8d859db25cfa16d44476e29fa40c1b2e94753e046e0b9a67e5bace06aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h786995e4ca413285a8c3ecb7088182dd610ea6ba2cc5e6d8ee8dffaaaa70cd6c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h832e5e4ee4469f2d974d76a17bd91e113c7501aebc482d8e82d0095b10c0d5b0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b73192eb11ccd0684e85365f8eecfac652db862b46114d6aaa94e1ab1628303;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb547b951ed46570f10654e7fa02bde6bbfd975a0c91c392b43f867134dff963b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h285b86f0a1084d408ae5c9a7430a0a0d8863745f82d6a6c45cbf176bab640a98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49a9540d7f300e746d3851b89e72ea52edd6cf50751b62ed40aa5f7c8f60e62d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h495999584c83fc12766c96a1a6453d1fddc031f064b5fc38cb9453229f3560eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72ee8b5ea329331eb398703053cbf6f0c01ce80bef16b67aec293605f72930cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd76dbfda34a546a843854f839e6b31a49818b79ae093aeec51659b4e7a42cfaa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcad1333a44091879343a87587b0d2a8c1e276d438141d18a66e39480a696bd7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a6aabf304134a051fc721eb2f980989cf01d297fbbc2e74d9e447b6f17a4da7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc3719fb08b334c474f1583d247edc9ddf16b774f52931a5ef0150bb3bd9944b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b96eacd87a3de72f5058f0b2f50ef5b806a403df5f88e79fd7b8aee89187a57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc8ad12d06fd4f58b7c8c92c09932024998edb4a54b6d3596e66000b02c45bdf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc960ed2a43b75a300dd4790b9e1557a28d7391cdf6e412db329c50c6bf613736;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75ed173ab4a9a755837c246805349650681f2287ab4b67b89d2f72c97cc52468;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h48efffb5af3e13ca92788a6ba4ec7a7aee02c955f0de8288926023eaaeca718d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73a2ccdf3c15a8bd593e0115755b5c97f81cf9fb0ac8f8398e9164148e3efb9c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e925b063d0fbce56d5419fee8100c1c41d4608930d145b35cc51ad7ea52260;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58448f502d5615ea496e21bb174b433efc5a9e9d693ea4259c180b9800d43cae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf4c984d35e6c82b2871d886ab90b210f0b94669cab65a773831a91891e09e2f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9524ab8ce14cd79262c7b4ce4908859d0f9440ac830a9fd770f2d1e86b7e3b79;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2c51134fce0419140bf17f1ad8d2771e5d7f641a16c38982764a78c6f8a7274;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd074ba92cd30837440c9c0a69585f5b8d9674ac05a1291886df57f355cd3d6c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h351bfd987f8e2d27aa62cb79a4b301afcd4015e119ee46fdf864ec43a32f0ce2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h108b50a071a0a33b8f38d1f8baa1dc5dfc83b7165d19b4f6711a1db6d89b6b5f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he523cf54ebf68891479759bc7440a0adf0c4389719cb049224280312e1a84303;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h856f559b4c409e77b52722ab92dd5a4cc011bfd6b1928687f74dcfb464fbe0a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7bd74eb63429b415d42fe9b07ebd4d3bf7d22d9cc4f13df08f3c168660d98c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1ed5cc241d4eeedf9fc483ce0f3f71ea4f91aeb1b2a97ab9f75aa72610f43c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb883f7be2c35310bfc23e839cb8a5bb2f2bcd3c5b2fd0e579f85f6177b462b46;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6bc798aa1fc88f6b1c36c767a85d5919a7b3ac199821f6c95cd86d0a5800fbb5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59ebe4000dc82e9128a526f729a748d52296da516afc2524915ced81d3e96aeb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h741cefed2082dc2e6eedea6551af58ff1f32edefab8098773cb9a0af18871038;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd46871fe9aa61b99d9d0fd4f4b7b8c7c7eb30c468ec0dab83c477516f306edcc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h51782656090b023f6a20bc6e0547dd12e90f684d9f8951b6ddaaab7acfc27fff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50e118b986baad21685caad1544375027696d2d93d69095b8e6f10f31d9b9476;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5323f6ea8307a1c5cc0056a1ff20851bddb57d0cde8108e0949509586dc16c98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa6769980f2a5d72d81e0fe0203d52ab38f22c40c75fa04aa1ba3a642397ed6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce571d6332ed0eec4679f1c4732adff4d3d2d6ea050816838d79d9225ef098c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had5036bdf8a8e1f50796498a432ea64acc748ac1a652b19a4536785048989d45;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4682094b91173b2b32f3509c852843956f93b9d76d9070763bcc44d5e39027da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7a63e00efe6c7b9185685e6ded32a5340ed5ad7cd36b019567a32cd86d0fc8c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3cf082507e4da067d96df2f435e7c54f35a68dbda2bbcd2503408249be84ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a2aa6ef1cdad1575089e9953530581156d0ceaed54efe5f6386bb127db23cd4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h85c8884e6aef26a92c6f5c0a1f18b430128347ea22e8fc0da640183132d213d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7591894292fbe002cea6ea1757bb42dfaf133414ee5c755f3e53b7c8bd9f8f10;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2244e8f37bc67bc48919140a50965bd4da1e97d00785310459c1aaa7460dcad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4ea813ecb4e2eced54166e25c041002c6b4ab087a4b6132085903b8279076d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ed9966d29cf90eb39c90852d165c9738e87205cef670dd610a621b6b658bda0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19ab1f32cce92d040c58292bca67ec35a6f62dc78ec3a68481b433ec2c807638;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8dad213e7858f1777be8cb0c13f2ce6d8ed5c0d861a5429cd0d32d33542c5bd4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6dadfca6ff1a1522021d7b6a5e7b46e7405aed95c75700037761577a88737dfb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h785a665ba6b8853df3f51481978d577eba20eb88f0a6dc7f1cf9c24ccdcd05c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6e76f0cc60eb0a8fc58dd11fe4df37489811cb0d4cb1c3b44b3dc5dfbaf9cf9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24404970129d29434c72d44e5735d25e4873dbcf962b65864858fb86be8a66d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h336bc738e0d501e95e04b48cf799eca883c4430f44efff5cd0b5fc7d3d03c88c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c84df4b3a1cac9c10ec1fca811e3f992e87affea9f6c7f146a74d7ab72a5be8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2caa3e44604ab371ba573a3413a595b304196028b3b4a2267573fb38fa894a1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf0995b8e1643494ba6d3cffc4deb1234d991e123071958fb4c99faecf9d433b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc3411438639621fad1cd6fa9451db1cc75e106303910022fdcf03076dff6f03e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4bb9216c1a8712326e0548539d1f30dc6b8bac87dee22cd0e8716a5d4bb49460;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0ffd3e6a44195f29a9cef0bf4790ad2da77bbe695c0da5bc8fe19b2df3acba2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17b95b48912a1edc67cf015b24cce496bd1295743c4ba0f6a54fe87cc90ea73e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd86e69d3be26fc24ada711e9a3c9b842a332038deed201fa8abd97089abaae9b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcebb949f8855575cb9b7dc41235f10e30b8bc0caf7fd25405191ba190e0b48db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8cb7121f63e32edfb355674d984e42bd1f67cf50d7e9c341fab269dd66848a9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h985f1307036cc61aaf3fbcf1271663b2d53048689018f116ce11e77ce0ccc0fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5ffd177413f316049f0c3edf61bcf8e2b39e7a43311840cacd1243cfa127dee3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9547eeef4d8cdb080e9a127e4593255a1964cbf212184a357cb1bad7d3b92e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19578ba78a659c80f758b4056fa633269c3e7c4799849dcc7309685f2f0a8427;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d7c937c7436ee2ed2641e4a0e0925367c5cee66154e5881aedc256663111a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2dfce47a54b6ed1e0f05a42e7e4171d5554c79bffe4955002cc03f5d8736986;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3ac3e0f41d462413f42c9779653ee5c98392534bfb91cfe432021d147e6a938;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb86d47e456a6d55df0a6b4b83ef5afa8efdf8f60d2720943f4f859220653a78;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d99904e4d7df96c32bfd0385d59a2f1e5b227fccc4efd005898d3d5da433a0b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe4a2948d14b198a0f55cd52585919a16659701c2ab21ee6a88493f2f79440c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he91a00623bc8017f093ec3d5525a7166a83430ec0634d46dd1e24e813a391c53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9bb9cd26fc1a3217780c739f7742d58f59a2daae44911fd85caae47d6b48927;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h588dc539c33e10f536709df804b947ca43a3388ed2a0296d55a4402afbe4d98b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb546f3fa2fe0e936f21d23514db4727bb99ce2c3d9502b670722b58d87d06b65;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17a3d243e969ceaecb3fa280ec20126aa545bffdafee398fdcffb0971e6c7c4c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdfa537046e5d8f56f11e458ff22ae28c699e058a8198185e1b0f484126205624;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hccf5f15e6c3fef1829044c95ce7e1039944bf3c69952277999332135e3c7f51e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h837221b4adbc973b7c1ce487d5ba920336551592c109f9cf9075ea1493eef1fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he344bcdb06d7037f6e2b7bbbb799e3fa4b3028f19b9ae60377b706bed7249bd6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda44a527d7fc6f04bab78f277d23c14af825fdb0006995665cfc5a1a8f442123;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ac18f86bdd673bdafc756a040e605b417378e07170d65a57aa2d4409069e8db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4bd2b9f17b764f62021e624147cfe4c935b5e424639e26029855c88c6e10501;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8fbe39521affcd99f9e810280a3aff68ade139a3b8e96de33807ae092f233f00;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7635a83f5346c81b8b2f14af94f8fa56e0eb346c4e80659d33c9ac7e927dd63c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdaff41cf51109c8a55b5e161c043a2a2e14d5ffc135fe57850320e07795f772c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb54193fc378dd880cfd649ec4f6f151bcd7b7b3a0edac0aaa164ad504c0bfb3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3738d51e353046334203626f7e2aaf551ce3041f96d5b48f15e1919374ba57b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6029ffb3a1e48b6af99411ba12758ea6f310353a55c7091c8b1972a3464e0efb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had276991ba5f3709ea7ca24cf71487599276b4928163e7cf3359ca799b5169a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa6991f9e6ba46785f7c991e1145e6999a8854e846dcdf6130bfc95139ddf12e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd891553573c0e1e5f8e3e8c03218056cd14f4690182a1003488bb98a15a456c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef3e089f8a1f1d2a5b8918b23517b0c13f0f6e4555ec71a0d9f970f1eb8f8034;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9419abcc9ba9daa2921c446f346122f70e1a95a40f6a0941d834ac014c404cd6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa74078a6db2064173aea78ccb99e786449ac887e4b40cd44366f50d42a8aa37;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f40d153e0a54a52a5d475bc5a621084831c394a550da2080700a1b16592ba9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c452e426354ae5b02ab55a6896f1612a14e5ab2bd3710ed132b1bf15985d3be;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2f5666eab0297cab1d44647adea5b213e0492ce3c7c121299a1e4a2b29d87e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h972dd4b1a43935aaa13ac23d6893ea99e40370c575caa8c856526c2eb568feba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha01ddfa57935a0c1e0e22b4ea80cfde82364f9677e523404bf36345e60ea31c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h419bce356af5694eda315f0f468302e0a72e2eb7a592863eaea3698d3f417908;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc5545a8f877b6658e16bf773ffe2f171b91ba96f4fb5b4cfd8e49fe52f091af;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h450c235bae10a6468b808a2b072d82033f63cf54355973c275884c040cb337ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb84143d1026d2f9c91ec00aea294acaf2b150e6889851f4cbc66089aaa79de1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba639e9bab3f8e5dfdef66799a827ef6f6afc6ecd21249505b17497188413f16;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b55ea58f665ce3d97f95ff3b925a965d3f151633c402e13a1d818937eafdfbc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca200d947f7b85855c17965ecc588c046c6371e4a0b968c3e9b70a93405b7c82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9248dee1c29626054f48bf7843165683fcf9bdf828f2f944d10110be04eac09;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h467ff7f9ef6d3387834644ce00b1d363fdf2b2e63ffe233ea91453d4d424ebb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbdaa3beaacf9624e29415b89ff28517dff334f3b0335a8881b25a3d8a9336ccc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25177197a4b7b1c83a9cf3aa3f2a6cdb2c7ca44f8d75adf1c4ffc56ac477de41;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed2df367eb24484b35458a1cd5ed515adaffacc9c804d06f11b510bbc6585afb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b4eb26f4b020642abfbeef4c770a4e47093e7ba839bf2c74816dab7976e575b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80f69a259171200fa22f89fdd14c1d2b750b3b8bdc71eb17c9b3a4ef3e9b3a33;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ce4c98011fa949321453e4735b2e456713bd1df2ba1a3feb3139fa2ebf3e124;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42ea7d7ed7f886b3049a35d508d94629ef6be5304e9c95e81790e27002a121fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb745fef69e877722edfe769e75d20bde0b73b2d9db4d881af906f71a231cf2ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6708ec57c6d6c3ec1a628fc70c4c44a49b0a58964de1bdb7f6b08e4c53126a49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4157ba6e6c7ff28c0ee7e1988c5f65668c418f11f6fecfde2bcd073ef70e7d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a1dc21814bd53005fa2127b2c0fc136b2082eccfd2612ecd007b1050748da50;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8da4eb3ba847e8f7e518491bbb11798f5e89ab8e8bc3c3efad3dd3053a59fa18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd7f1131880d1b5aa2ee0e53e09e6fffc268f44689317f801f9644b7806d5335;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd60fc2861bfd4a090af2a42c34fcbd3aa314a6b863aabf6508bee3052f459a92;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d35abae763918e5f935efb8d173451e9d4f88b40ea008ce8fcdcc6fff450abf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e33d799ec7c5296351c51ffefc77fc8f01d75462d13cfea8b782487c730851a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd88c0b919ade4a4ea583a9324b4f235ea695b45b941a01f38ff76acc866ab39a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7903ed44e17a00654341109daf3f7b367810bd6b8809ed18f0dd4705635432db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb6cab2b3702b89e5079f2623f2b1842d83971535e7ee5cbf7c88bb7a65ed3aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he87775dc73cbb045cc13ff6099ec34d328996c1f625a95c501c9ae3b3238b5ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ac75423e8c9c1efa19af2864a81670b9282b4fa5f362b7ae380e7d542d33295;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hde4fa74f0d81dbfdce96c0319c1e9843aca07b3c84c050174ce1c6ca12f124d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc1469d7d17b0f0eba042a79d8997ca16e0868c2b96ded67d4f27a31e271b2d04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h947c69929911171ad7476e9411651e8cc5483804849492bc9de7e161d8f26fab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h34c87ca560972d5370f867a85e43c547321cab01c4f3bf0b74c61c41256541ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb163ecff936f89546792cb728949d0f2f088a6abc7c51fc06661638adc6a6fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4af2f7762cb334635026656bd2ada61f2f26239b97817d90bbb34414031173f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb15a2005c76ede8a26bc40ae5ccfef5d096003f7df53f68a9c1707c7e1928a83;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9962d91e10de9b1f80e94a2b757f9dd3c2fce3d29cfc64c42f3c3942e1db519;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15b16d57551d6f4c0d157f7f576a382153b73902112c8e831d5833e502959af6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c03692b84b4012114eb5934bd72d6cd6861ac3a0593f08104f39af8cedc3b8c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b8b2bfb91ea2dd6720b94fb06c8dd225e2b099ed2abb297b287850667bdd85b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc44b4b995fcbd54cc579dca03400efc32ea72faa08b5a8a01da109dcf4189fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a68dabea29d84ff35cc073ab091b8324cfeaf1f6abd76f5ea4bc2d3719ec775;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2cf33b1a71633cd251077f1f99a7621bae35fe7e38ce2b51308e63872ca7436;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca5438e8152afe205385dfdf16d8bc08fce44ba6d5350073c68cf53ae5f4fcc1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33f6b666e2a50d7b80b2527ee6b038ca64b318a506dc3159b1f622817b8e369c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8f8c3d74964b3be369112ada3047103c8a1119e40aed278f5d04423b6c60f5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc325684ed8d94b509642a879d228899867821099e9bf1f501bb2c11393472721;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hade0949e1078f83157249b121ffd20c624e050d007173b597b01d1f56374a2d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88d94416d1ce28d4556b9b5b080e43760b96de9e50c9fa8e013596cc2331b12f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4cb579bee4acd429f95d0b68c0e74f40beb6b15ebefbf421df5a7e075e8ded53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb877230f2e15671f8c307950469b18fec529ce9d7480c2068a3f4665fcacf82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf8402cdd7360ce756924712b28c240890d0a93ddd6e14a7941345b74d80f862;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha36bf5cb6c44f11cc30f9d7b0f8d454b26a391f7c1b0eea96c94de6bb93dd44f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b2ffbd61ff8e486d5763cdc24ab3fc0b8b2bef43ca9f9a15852eea73c2922fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h739f0cb6b8ea7ad6515bd993dcfed8d1a1886230eb63d762aec8e4560baa23a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3720e9671fdb6dbb81b66592327185b1b2d5a942eeb8649cf5b039c41f5e3b5f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h564280a352fc22f8e361a659d80494d5783f5ff2860be9540dbb035b0eef47df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdfa01e90a607863051cf4da601c372646c4916d23dca3c7823bcb53bfb6eff15;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h76908a92e1c4110927697764492f0abb6724236918d834718b0ca50d033bc6d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c775ac5c15dc2317c74f2132a611bad3a0642b87d2f4e1d9be0ea115613238b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had28c339370696ffed38bb3f2be8467381c0d0c205b285922906c5cee2f0312;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b777e7319de92f69943e203caae90891e6891dbb410e8a55533d5cd165f6c7e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h955a6dda45aaa342e47e5ad6121a7376d867be91d109f7f576b2f22a0f9e7977;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5ad85dabe7f00d04798e848db88ce0038f6145ffe651fb4fdd665feddbfcb3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5691836b1f3f7feac925a9b197ad424dc7499efed92a495d36d4cb00a0f4b43e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hacbedef0752c34469ceda6e89c55cb2c8b43af1c8f5ae3807711585f7c1d619;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a1cba3290ce39c8e5252fb62088234a6c27d63770538409cca8743f1f75ec2d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heec4b30b5512c14c1c7c4bd9d4c8bf9c99369aac3f412c0f5bad8b0cde3bbe19;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd20c4a5441e3d7a01de308b6f36ae61aba8c454685a4580d4b6965452694575a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h84b713f852c8a1465703fe139e2ef232e815ad926f1d1408850ad2f22d71df35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ea0e5be84b756124ae18b6715f1c05f82862f6a095757ed2e4556bc96b3abbc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb840a876c335b393a903695670821f30a25efa83fa42145282fd663346bf007f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd88787611b5c9d811552ea2466a6d235d72015a3efb15029e05b6e7f1ebda6ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4dd21a58586c954f1fe414fd9a1de1dd6f2af691270ff4d95f9f2ace9199ab59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5d796a5953bb99038c746f098ed9e5fec5c4bdadaacfae87fa0c6dd9420db72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h76c29844a81fdca645980212fa3cc9182455f63b26e0f9e42115c6372c515a94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0b036d1fc86d220c44ae61f2b43871f8d89e15dc5ee0d2356711890e5e007e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f0fed6d4a0191301fd1421ed9f59e755586b5d8a203bb5dda4c4f77699dba9e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e3feb5475b937119673010ce7a74a4d97736c5c15993457d81eadcad03b4ff6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8a9e3c2a9f9508669bd226f9a4faab884b01bbe837ef2cfb6db8ff1c11a6634;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf85db7bf4037bf0a8b01b8ab92f0b92ab9cd68074c9002261f774755ebfadb7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc482e680b8f1763e1d32b6da5397a3c2f6d427b468bb2a500c5b76154ac04c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2694342d6bc75054353fc9b7e5073b09942b8f55fcc6a3a7a5b9229a0b7204c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7abc4092ba12a55871fa8661533b068106be3e387d9cea2b44f80272b3115e3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ca261d0494922273ca06951c84bc830a8bc9ddf18d2b8ede86b006f1c6a4c1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha79858eb84cb31d8d4a222e7fdf1195b9c9c1a2ed055f7ba4f97e405981bb4d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he31062f212c71fcee63b1fc83d4ff477373b1f49112d138d69f2ff21c33fed2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f43767c9bd7b374088edba77ee5df17ea685fd4a48ea00bc83330f0ea5f01d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5fd62fb252fb8ad14704162b40b2b9dac6866aa38b36beb082690b2d403dbc1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96a6817fdb171a6cd7582e185500aa0835e508b0348ae80d966a1996d2278171;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfad6a3a6cde1f9c625367093260a71b65e0ea7e3c1ef4c517e061a614a230e5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb3ff162a0c61d38f5b36fc065e9e322a8933a4b5111f4fb38403f1f993def383;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h678f66ad3ec3dad483b07c474bfef45046c22c5d85aea62c269a59e1ffcea2ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f07e0c19bc71bf9d212f3a849bc11944c0cc957356b3553d0901baad2514564;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h639ad0943e1d643b85ee84be76165733cb13874d34ecc930c0a8051a81c639f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h549e4d4ebdd54a2e1442f001cc6042020c54fd35bb7a1e3c106bab6348d95adb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ff2b48459851b12c751a4ad36cc4757c7509100dfb811203fade35c38547acf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ae69af1a6d5039635a4f451bd7fca181b7c487d84e24c47c2e5a7337263a824;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73b7501b3b84453f51ba50998184ffbdaaf9d9f2898cbc28a1c1aa4e524ce34d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4b2e382445d8997d4ef76124279838bb5f68f50134e56b5ca55154c11eec191;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h161f8d7587d40bcb6310075fe75f175f30b90f1f31a2f68c22c50e4285cc2fb7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haeba888ceacf8e25cfaa3fee5e8478151d05e6e2d57abec0578bacd64c349efc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e587d1aef6d2e32a4ed7e787fcfc47d91f0775b5dc3493392523fd40509a040;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17026db826cdc60775e7e6a137dcde94fcd3869b92c8a47d7cca39bb340dc5c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h243a083e6293b19a570d691db46572d5528a387519f9450b29a62a217b4291db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3db36f80060828d0f5356ccbfc90cb98fa3b2dcf584b62a4b07873d3b27d0c18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8b57a7890ef7cfa06d5fcdec044d1698ed89fcfb90d47705005e46ab644da49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52ac402f19b4d9974e6fcaadd8740952c4cd1d5977d60db2971fe2242740e55e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6caa80c4177e20dcc5867abb83a42e97fa1af028c6677fe1c39e305507895832;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6f873cf28de0861717bc3e4813447cdbb04f9c9914ca2d4148529f0a25e1213e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a662ecf9e5ce722c16612e1a9bfca7d331bf2ee4a347016a86d416c2700e131;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h55abc7609d8b95ea3c91436560449cf0a07d3cc88be7549242bc4640f6303a3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbbf8466fd6a5a672a3a17779bf324c41f1f088d1451fa9140080101c9fdc9e60;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h666dfebbe60cbbdc8f4aa9942c9ef350ff6943a05b8aa07c2c66e2e36b5948d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3c99349390ae5f82c31f452029eaca22a320da5a33d90ff4bb027614c046bb5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h416731f4460416e60e94e6167e4403f09950906656cf1144c8369345aadd48df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8164ae33f0331b2697c0e10c930c858b297cea819736d4b0e310ca959f6047ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hddadfa280dcf921850bd91af4ffa635db8ffb0bb5b75e1b97926ae9f5c04e3ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h27dd460295bc81d5c20578648d6fe17fe364e0f64f4ccd23c11007b1d8230f54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b558535e42c67143e9654616a8a0675a49383eccc087b20bba98cc02a8733c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4138e4823200c51d3e6d23fc88b3c073528b6505e2807d8d2f53a0efc24be819;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b1a163cb6bce7d9d9ce038040fd6572dcceaa31b77f90669761b4b51b46c7b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'habfb3544b011f9b801766400c2a46ab8247a10101948262f535f28f4ef5bee26;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hddefda25e40e65e67b25da145ce12eb2e837f42edf0263c604500d8c0ff4a206;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbcde25d2c39663ec859b88cc185b9b39c86abf5c1792371aa13bba57ef0884bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b1994452b669f6d8fb97bdc14ee12c13ce31d0349336d33a134e6a220db102d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36b06d1ca77e5727e0ecdbd0a3227d75beb183cbfe555ff2bcfc43b1cdf0983b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd81617f88da9f45e7038c279e5bd57fbe409d3646c18411e7504e1739ba238c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcfda813e0e1ceb58fd4c4b28ec0f668a2af309f05e493d292af33f58e372d2c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd84a634d2faa440d804d491d70e7c03445a3441c74189c9d954deca2baf60a44;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d3bc5cc460fdcb9817f8e4ea04081cd3016e5598215b0f65e78197d9a378f0a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h672fdb2bbdfef11ecd8772996cb8c08932d03473f651bf36664b63f0e4e9a290;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h100b7b4753cc64f0132a6ad1bbdfd577432fe1050de611112946ff14f8fa29f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf0ed6dd49d1b85b1263c6e93a13fa52127f3369d09e6526d7814b4ea140e22a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h815aa359fd27833ff973c634b1456646bc7790a29700ea4e1f3b3972f7283ae2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h220f06bee6813df77972cabf1c64c6c610a02a4e1abe1f147172d1f0d72a7e54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8adcd299d61f7d05c14ceda0f726decc16a1a56fa2e21d3fffd92f5b60919bff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6827a34a3396b67c816cc4d1d8653f4e2d91e3602646dd76f9ac4d1ae907c85d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd8506736446019c34fddbd21075ac5a3992df342eb463b6c488e8a2fd97c8288;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'habec77963fac244c5a83f32eb9203f4cd6b2d8b8bc7b8a4def6393bef40ebd36;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a861bce8e6bd968b315bc77474198d2f9c53bc767dd16d463430f8493b670dc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7215cccbf3571d7aab15371c4d02774f5428a07563675bec4bd056b59f698d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7097e60534dc0fd6f57df8715cb535e693491f9b0f4d32847d1d2f27fad168b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e47f372894642d881f4960f166bbedb841ce05491953d41df51eece4b9ddd4c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd77764172effbe1ec751380811491cd954792dd752c99d348d07b3fe7903edf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8813c3faac2639730b6a5d3c32f29f4e01aade311f933d09b8bea7b7bdb76946;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee43e21e3e441f1657311adcee8edce6d2192ee41bbd522d8427e895c36d5945;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9941657bf8ebf6698280ef93b7ba815f05477cf022fb47679e61804f9bf903f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h557cd06b7c66a187c1dfad953c6ef51857dd3679df218d9197cc0313d98eed7d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60da5f5ec22123e50466d24f13bd6adc3d225d1558733ae6cef273df9d22c0f0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59029f10b18e8e9d6943182a2e659598a6bbe437aef3d5a91f7bd6ddee107446;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74b8d9b17f94a242352792304f95332ced61035634d216c616749f11c0e6ddec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda89022a23da4a06f4f82aa35db89930048b818dce9e567b995ac90015e628d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdeb7af1dc5fea9b1efef552b793d1882976d3f48b4fb35a7918b20bf551eaddf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7e2ce6ee8b0a7133713e2e79fb7ef5bf022a7f4334c165c7529f50c1b3dc3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7260399a561c65209a99e9f467a49251a9d042982dd6dcafcf1446e7875909c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5bf2c94f3f819764f7be45b2487cbd047251829afab1e0e37c4454e1b439365c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h34e538acb403304773425318ed9cb653276fe7c2e692faa35cfd57d527ff6ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62badc8267caab5f77f494e4812583e93bc1a1c614efc334ca392ec63aa6c9ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h206e33d4c8e68852707d0aea2154b1e7f4cde7533402238ace6232a39a837b00;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb05d93a00b7e30c4a2ffab051ba92e8d60aa3880beaad5e3f2267f8f757b6e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haba91049f4e551df2e5ac87376449964109a924ab5409af42cc34bdcd6e15808;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49c65b9d4be43c37627b9a48e13a895724029698be8aebf46dcb789fc2dcb938;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3eb472b0e6c777f5ecac7d96901ff8e32289079d3e5538e2c150e17186cde70a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h269222c203d6decf5c2cedf8c21de11adc36f0719dc544f6d4e1aab35691d61b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6d48c4f706844edcc7d574017c9f543c4ce982553b4355cd66009f2b50b68ba9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1434bc61a7eda0ed18ccf6c0764a3007d75012a1aa4afa6bb22dc9dc496a67b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ef1fb0374125e51f7403a16d65e3a16eaeb1ca99f7c858dc87db62545e5ea4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h99149dc365c748d80ba2bd70e94bf8196f22c6ac084483dff32d08e2b2d966fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha44fd713aaf91ac2aa6847073deaf12f902631862b8e2feb98ccc46b47445211;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2adab40dcc2dcfd13de8ffc17b7e400755429157efca66558772ab99f986de4d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h985116a65a91ccb6a08edcb08807b6468554a6d36beab85875192b0a28112e3d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h307ac73f3d5ef6f6db4cbb8b6358fa5b82d8f70c66a8543bd036a3653f4502ad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc97fe9e028c3bc1af55df9c4f90a3a79938d2b08e76032c4a1deec6bf578a313;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha1a2d76a74b357b0dac68eb63d0071740f94c82b0717d668abad2745050c9ced;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b7a02f82522c0f8e5f767c5e8dceebae215f36578dfede4ccf91cefde18cc6a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5ead47d72e6e00d43e584051847c59c0a0c478da2083ca9f32bb8442330d9c2a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec86a2eaaa5773809da11053366387739a3f9274b33e12367518c4ee190c209c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d9d3af625d2bf382ed3e5e63c1aa04b9b94db4394e09a406b606053f020c22c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9d69b6f8b46e02d2ceb2cc2f7985e52ec4d89fbd4db08b9ab635fc5f3957d53f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c95224b2eda0fd82053dd14174d7b8520b84920d6a63dd0010aa4f8e12c6ad5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68703514f1628b2b00117d24d5eb3eed96b7318bd8b4e57528edc8bb9952a32b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3571eb357210a6b844ceb820a61ba3fd8a2232addfd84adfc8e2934ea8e00781;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h911d9c330c6b4925510598219983b76b7012ec959fe4d15009fa498a5f497c41;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae2b4c26183d9730ab16f1c886b5f087c2f3b95ac54874ca1bfdcd6ccafd5cf1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b52220c2a10f7d5de41244f52f8f80092237948ba7db0f3a6ebc7a50849e9d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hccd77cee24b40c84044a7e2d076be01a6df82adda1387578a0e52c8ef09dab49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd3b7e48dde9d63ab0b93187d8cef7b359ff54677fba361130339d304794007c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9f6ea6c0c0c751fde104e4958a46d8f6172bdb1791e3b3a7344751c50475866;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e7daf1bf29c978c1d28f457f2c4fd84a8fb6e8e6d2f50412230b3aa0c883129;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5aaa1b7717decc2b8e55291e005fe3f5fd92768f94ef0ab75975706cda7ea45e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1702867f98c46f157698da51aff42efd249b99d3bf75df4719b834fb5a316a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h153a9595dd5bb6b215534344aa05cb0b652542bf319b8688fc96e4cdc21b9ca5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c903f2d34ecbc7221b3dc9ca8ad42bb7177d9098d7990d2c63cb7e9185169c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hece543b2f83d4681168ddefed854b717b0395a055d6479cd79bff3a0e73c8bb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4329c5741eeb6c1eb9fbd52e6cf0133b2617ebd7ba38dd79e3a9573134ca3df9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf967bc56465757efe41ffc7bb3ba49e1e4fff22cfb8019ac913fa0d88a731e4d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e7f675a3680e0e4d42594376eadd89b7a40671a07a9fbae2a3042c085a03e4c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haee3ec6f7901c803e05848b6eaa7da32624219f834ba22ac3bd869c7e00d331c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3751aef7e2b4156e1bb929a013fc15bb745ea4c39772a844f75edd9887aa8833;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1db2694bff0b6161e70530dec0f54b46c2fe11e6991e663e4c75a089d0d8ac58;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6372d3047f1766a67fcf60bce63cb576c6ad4788d391270ec1263c16a3ae86ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4845d2cc330a366322c8467e6c9810a24cfd1a5e9498bc02a93d27debafe2237;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12e10f56eac0137229fd29561416b01ada230e32114a69371bcd92208192e087;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h894faf1b46b42ee02f31e0372c401de4feed11dcea338c043629d59fe257ee32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9c686683dfb9f99aa2c407e129860a6aac5d7c17e3a95cd77deb910866479b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h285fa1d68e0f553a54b3a17f871ae4011edbe0eb4259d6a1486891f2068d82fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f96468fe6825f33f3029b6774f28c93059d2bd2e9acdee1df91bb8820126e04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h693c25e8c31f6d3514008ea5dbcf5f502cedbd9c4e1197bc5be588a239886021;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74cf8e3a1611c3f9c7cb27c988e40e07d01a6eb27bb1b6a859239ddc89bf6071;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h865753c97835bbc3c8006f62762a184eac474646a53e1a575e7babf82094d233;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42e5bcc81bc7ec6e80aabea431f5f7b7bf0eff7e81a8a9994a50cc11af181ccd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a348092116481feadd9083ae9671199570c98fadad1781ed4992c28da517041;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b0b6c144d04c29165fb5920bfdb57f3adbb336e9cbc66c73904a30a5f0a2e96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52218707c98a87901090ee6b54e10691e493dfee32fdb88083580968b8245250;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h355c4ae7c81059454ce09d5a0d931730e5c1418b9ff3417cb749d38df491f9e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa112af51348609e0fa27ba95079f7e2241de067cd5684b8cb1609f95700b5d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3919f5fc6c213ea0209f3fd88915cf76e233d2fe9cfcfe1ba46610ebbe9cd72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha98c6934a5a3a1052c0e57862046c5a91464939f71797448f64c500895d61d48;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5599d4b6d3b74267257e5867685d0da8f53e9120eda2a93dde09ede19c7fc61a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3ebd66725e4911b1856f6926c267bb7d324eb5a1160765d00063a427b092d78;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe547de62b244520cef59f0b6da9425be1be9c4f32902ac9975579342cf60de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0cabedcddea9f51833704ff67c5eee4a8d4662845887f7e8b6ade26d7f8a0fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23526e5795a6e0a9f8c0e8d3908f0073f053cc92410aeb81b918019b33c41e07;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e99942442878697a19d86479b40623645902d3ae6e09541a4466863f3860bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89f1b23b6e3b91693ff39b466051796c06cbb2b57b7d2961c4ea6ad84770c778;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6f23eccad6077021a85b300ed1ee30c1faf5ba46705e28d90e0c59a82902c5b5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h730e3aa2f5c492e896a92be8e1250b0d06c1ba93b16355e1c731bc183faca895;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3b3fd370a3cf3fb831791b9c3e7529e98b2143f812a9577882944f1561344d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc94503c9a8d11d8834cd767c6f3112691d5a7d6b147984ae6883668fc466c128;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5120548e234df034e2bd5abcb44fa24e32f6a7185c1cd7eef1c8af6c599d879d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3268670b2b4ca14811e06c5327cd3b629bd51b04c8129533452e4985f08534b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff73b37d61ec745d6613fc834615c53d8cbbb1520cbd08d3e777b8ffca91299a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7287b09a12ff10183d72b31f8d7403654ffd305d835137967a8baea90140089;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a3465c4212175fc46d8dcce3bf8094e72dd63018f40691465a84b0781c683e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e493f2a68f5ee909383da370c2226606b158ff66a0bf16a377faefe2d719084;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47e74cda0e642c0cef26ed0416caf2763ba0f04299bcee53498fd9a064ca14b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ec43c1cc41f3d7d31b2734582f2cb46d16be887cd3f098d0052fc6052898aaa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf48b846f2ded2ba804ad58d515207d62ba662e4a6d37cda57a55de0d1f3b2d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf66ff6f250507b8bf418a6cccd639e9b002566062e6297e9db9d21696e5669c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36907ebe8e41f48ae22fd79df909891653c31c691deeee422c5300bab7e81ad5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h640dd94d20741239f286cd4c7c2a65886adf37091be817ce2c768a8385404ac1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a16dd18240e114f0b830a8898040bb2017d762e5ff1c02c8cc945b2a657e339;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e06daa886664e822be82e07e60f72960b3754f6866f64ffc07f3c03dfe9df09;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15a5d7b5efaba657af8aec9757058116376bb8d7267c7f75e2fa119070000a76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1dc0b82baec360b1c4a0fba25aece9f199d6bee5de97a026605c8f4b3b2c852;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e368ca62355805a5bb08213293343c1c8d0b039894ea1d5fffc052b7899dccf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9756d2373c5d8a196cd572ccc8ee8e392844bd5b26d941bc8db159da9956f49d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec266a04cfd780e8f9f421c82d187ac16217ba1ca597feb517e0cf49a1f3f96b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47f18bf8fd3920b0de66f4d4335da9fbe3cea9ab2f98e2ff17828d026a4b640a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf00523ceae0b8873bcabaabe51d6a30afdaae57b241c0bec76d6c7eeaa6b4c14;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1869b762e0953f7aa6b0570d27d8ab47c6e1d5a758e79afef0f28fa0a73b55c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haaa355263418a536846e6c061777fe65c12cced72d159ebaf85dd506c51936d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1065b926d24bed32a69dc7ba47a6f17beb9024f49612f5bdd6e814a95120e483;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2d5d538e31bcebab27c78d8275dcf1c5ced13725a6add0865fa54c59b1a1a04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h593bd0a06477ec9c52b488072e0167d4d506a8f8cbeb14915bfef989229a4026;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52fa2bd4f19f9437dacc88f04e20653125e930fe1d4150d0f9f52e586ade4f47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h670af343586557b5fe465055e8511d19b829716c6199f9a3a85f6f1d15faca80;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h621ff9d0df8bbf222df7878fc0a2d0e87d0af0771f2475169b2183c9f8aa344c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8849558a63af9aa5ef339211c4d441e715d4026cb520aa71bd39561872fd8b61;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53cc6a6b67c1f3bc0eeb73275e2047388b6e10ef7575ad31f745863e992bfed8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53d3e33cb696e36b18933fe1c405ee8d0963d43957c13b876581a8a5a7052bcd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6292f3a94550d7fc53c8718487f7c3a0559614440348c265e620ff0f6e8e290;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee76db68e2e5aa66a7ed9545da07556c19fd791c9adf1b8c82d904e2aa7e340d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7755c80fa8b8787629ada27439837aa8b675b825848c93ad4b3601c155e26d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf901159c6371252c6cb59c0f0546129033e7d9bf4a9cba7fc664b05eeae949f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h257ba876586712c32b96a0d2470ca5fcc73664c7b1fd47dff44913920a0b7b17;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5dcc8960649aedcdecac5f57843dc7232fc37c3d9447158485460e7040d292fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0a8115476871c79cdd1f54336c8bdc81569813ff97cc963e013084c573f85f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7c3f350f5984227defe7e38368ad337e1328a62db0a6b1454f79252657f3189;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h34538114661c66d33ed5c2fc70af6eb1a69c31226dfe20ad9a2a7701a10020be;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54432340de2045b91f54bec2521a68df660288473587a790efaf73e6fd42872d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he03e03738da4ebe14e12841223eacb6ea990789c2a2cccfc66ea2be5d57f8c98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2dfe25aa108080c0dba0feacffdf3eb966fd31c47c162e9320540c2da8fab37;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h669abad8c02543d8b94471817a773bc42b5f112fcf72bfbc091a2b0701d1b907;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9de4a3657e2ec4fbc36c0281a16a6407e0845ffce9de5632bfa6853a24c3c13;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31dc67fbe1993c57d552dd969f68bb6cce2fdaa4ba3199101d3a553bdd4861a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7cc071214f251071bb41039fa5acaafde217ea7a74fc057e7b8cd29f8db5fe71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0536c05822627ed8d095616c01b8a53e0baa4022746c827958f23da70076416;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c60bd1d16f0ccc25ff2464d93a7f0b9375d8bbb6e3a97ed3f9162c0a60dc4b0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc626fd946fe8dd4d676d84c22de00a8908307aec364c89a21fb856e3306e2922;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h95e580ba5d31beaae428c05d0786135c5afe7a91f5fb6caeb48deae8d148ef77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f195e0203a34015a3317b8e33cf6aad8c807273d338ea72c4c3ee53e5611908;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h766466753d506078700cee9d9584d4a03d01f2135f6b716466d2876f47e7dae3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46d9ad86304fea433d2eacbec3951d7cec0fa139952490da569331136e133520;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b2669b6a4b827bc6b43753f7288c93ad20b98e2ac5d8e1a78a1f1c59473a79b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbddc6c0456b3b1810f54720a218631caaaa8f1de4971e7ef545c79651c8a73c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd43f7168c1bb54c4229b8367bba089074caaf572f824e70ae082c4a414adf32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha817d3709435ee09bc5b07abe82954a24f54838a020c7b589c93bd0cd42fa64f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe1888ea02e27b603382c9745e4c3f76c4a588b397fac5e985d324d5a77196af;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5468acf7c18a8d7b28055550722d388c0f094f220cb9084aa34a2c4ad8f99631;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h678869f4930bcc0ae7652247ca737344db3dfaf0c9c01654d42b5a1454aac12d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b010c9ad49c0d05dbd945f7d3b97044bda4574faaa57ba040ecebf2fd106573;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab1675093bbaab070b6c996c7e9a1e52f39e7c3f83696f01a601b861b024daea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6dfc8c72e7640bdd48a759cac7fe27aac0630a6f3f59e806579fa2f0c1365532;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h87a505ac135f97169bf5c0d7e6426b07eb6ad75fedc0a8b7530af15b0bf4a8f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77465570c4a6719b7ceefc0c315c06eb84c0944e391600f400393692a7365d9d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2040cee6d5f8a1abe6e514f1f3f418ce98e08f9e94e087f91549034b160da1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56b14858b68bf1115f700d32255bd73056c75e9bd88eb54927935e05459b0f5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9725919cff18d28e059c6ee0f12d3bd901d75a346b6567ff40b939c7f22d31c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72844ee72cb5329cd61e579e31ac6e78acd3d685ed78709776a636d7f3a437b5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hafe675967fc8b3706f8ada4c069ed8bbcb6b3921978398f085f87bafb144007c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h27486f8b3e5ce54a594abee2a5109322acbb2192fa4c4b6f871f0abc87a132b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h90b05eb24cbe105105dfd06c03d603458ceeaabdcf736291a72f6c24dccc61c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb6af562888c0517743bdbcb9de08c770cdd12b91a7f937b72d6c83077aa635b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9690a31bb0f2c0f6903ff2ed70c899f4807ef77e7ab89fddc0761d09c879e513;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c19e41f326ccc87e29980a338b97bc1c8380b05bd9903ea9d587923398c4f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92110c68c74490f420e356233a9e7f28106505d9315afa37f6393b64cd1d4017;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb62e8f7859fe941e92fff0d66732035cb5fcea3ce948cb47c94b88bfd6833235;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce5cf83e9c2cd4e7ce07f6e4609b0f65f73a13bd92bd0e113cc26f287bf17e72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f32d28f4b93d8c53becc0fbbba7cc5647853bf4134c772e84589dd4fd18719c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb88daf5cbaae20dc1a810b78aee3b6a76bfac8e9d76790c581c5dc6705f0388;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74861a9ef1a1a4b91a24b492b90b452d5b543cafd079476bec438e0ff43f77cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hadd93b8081b45767639384d8b30ba0c23d079f69d4afde44ee067b509b14b983;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha62687608d82696bbca2ed23bab6616c82dd40d452bafff479a25adf32dffae0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c30dad92f46034913a37e2eaf9d8e4896c0542bc08a41e1c54eb7f778205401;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdbfb091a7a4dc67ac846aabfb7e4fa4387cab74fa98105b0bcf16bd6c59d1c91;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h417d4bfa9c27e6f70d51448eb6ba7aa987f396cb6e2e728037d475eb22161f85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h55cf309c1604714f211b15b34b84b250ef1189b0c3efc03b2b9009c8495c0e61;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc26210c85404b36c11e4a0c826bafb40091bd1ae6c52f2ac9e02200eb89777b5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1086c0732d464392642d534c0d56403eceee38e0dbb2e445e5ab7248e8c93e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcae1ebee456ce229dd578551da9b3d1dfb8a50f76ad711e642b63b8efefd2168;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89cc51767ed42f6f718de76fdecfd6e91a11bdc84607dcad4bdeea768776404f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h29167bff1618b996604cd99768548c1241ccde84f99cffe037c7d504c784ce6b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44e72667cfb7c7ed6f5151b358bef65312f31ed3f4074c6be56d653b9a2cf03f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf7d3db2422eb29c07ee302610176eaf68ac53b524fa75e3fa5aa6114a92c43a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ff74765960e43de0058922153693264769db7616e6e276867f7cf9b55578977;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5418ab4b56552b5af5e2589c5d060ee6f9f2b83e33927073ecbb6b5d84400c6d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc894d856c2dc411c4ba407387d1a73f4c30f1f761c166b642bf2404e2e092465;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h115f9c9a166171ff5d1fd60fcfea79fd808131cfc41b64b4397b665432f18302;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h99dca282d2e21e15085846dd1f3bf64f594739bc079a02383d8d8502b8f88065;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd897b40e2420500c6f7d85e21cc5b46eef5ae70d9b9a9654a7e97051f6ea2e4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8cb86621bbe42aa405aa3f97e8fdcab22573fd62a44227d7070d46a75fb4b9d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h304d9f064c9f800fb35fd0506a5d45fb929582d99f2409f131e86de94215e32f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc3ea94cb78299484ee3a410058f79f4ee06ce1f7cee37e0572116e9de7bc5f4d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3de063ed452816b7052e67e2349f8b5e579e246f96dff29cbcf69a25ff189077;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h13206ffdcf84a2aa7d5d4c4ee62f8375c938b76d79dbcb39406e82643bbe7839;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6e725486ec14d2260aa69aa76a355a39d1a6547773c9c632893e870887c9677;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6c192d69ce702c6967881706689d9681902489e9dd47f087a5ddc173c8e8094;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f3ecf1995b347476e62c9f46380f4398c5637105de4f03f8d02c6e2495d43ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56e969d151afdef5be579fc5534da287cdef10fc8b4f9010b175ba64ff6aa08;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf7ad721ebf4ac6e55c660ffc39958bb43b9ad5c969208f73b2100d39e91341a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8236427db33222452fd2ca10a531524ef1eed6c4e6b2ff43039ea651cf5213fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5ec1297b89dd92367534e27d02909b726a76a1d45e3f26b4df132257c96c189;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1fe21f189f95792cdb95ac84defef314ff0da4d555e60185bd98b2fdde9de08;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f61e41b95be197b9dd6df836e4aa416b249afd98e2cda0f365aa8d02fed0f04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3c02140379b874961b075d25a05cb03159db1c2ae1ad1325404749da661998a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb7f2b34631072f18fd137a9af41f899b53218a2ef474ecb31fe1cd6faaf5f8a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h604ac8abc3afaf20efb7ec26a74619d600b2402ccd419a4032442c3288e1a0b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha050769bcc0f44cdc4d58c749951a9336a34957d254f5d8e2c5a9c14eba6713f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10f9ecebff8a3d13bbbe6b4e5ad9e0710ae5f097c06f8051d4c2c8e852ae169e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h480902dd4af884d2dff5a30b8125914e746dc5f8eafbd88fb58ae57102910c98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b8dc7752573b0025278108ab62653c3d6b058ab6c9e4911acd9aea42dd33478;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6d1f0a20829def6e2a3c48c20e106441f13d49e27a2b6df7c84b929626edfeb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfefececa7f47cbd56d329d6fd01c05a458b81b66269b5b258d4057c2c364a3bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d21acf3c64a11dbf8d6aa6db14cc8d7a23f312d97bdfdf5822aa8bff4f7018d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50183eeed9c09a1d1f8f3f73c7343cfb808c17641e1f931ce6560a4065d08891;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he07c6e2eb37a7ba058160f0ade74f58dcc8de3407016ddeca4e8dd944294a991;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4bc532ed770d8cb720c5a03edb85a39be77d1236eb6d40ba34133baea11c82bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he0921d8f523ff595b4941a8c3181a2980c7698120d7b435d2aba09703387154;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h76b99c092391596b6702bbb2cfdb7382ac73c54920e6cc85fc4928bf316050c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41c28428e56356497108de5e8a7f566cb974380bf8f82c541a8e76b8c41da713;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f81fee540783753b7c40ee83811ad5e42a559f4551e686419f49323ce235288;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0683142ff7360b0c8362333489a4ac3ae86e2646277c81a3c80ff413df65a95;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60b4ad6acfec13ad3c6357f09b2bafeb72e59fea0ba5e31542459d2896f5fa15;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6a5a978528ed499fb2193fc28465c7b3c2b14045bb71440a118732f013841ea5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h472099579f56ae61d39dedfac47b029ad8b1f61c74d6ef1dbc48cae0221ad06a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e4697bfe7d7914478b9b6635141d1fabf19e003b5ecafa7d3dac4c5e268ed79;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h125c98a45a6ae7e89a802b95243307a436b4a4f28eeb813603016afd4c8a759f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h142f84b215fa9702bc9b83d25740b44bea0744d211e57e79ffd74f8d2242dfbc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e5beaa48ebb612e4b95f11d39c78c8e25d8d795dc821dadec683c741750ff93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3c6f6ad839457bd49906f2b07a69ff9c0cd9416341b96134a4d467a6a1bb4d55;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfebbc930ff4df9f1239fd24b413d614bfd9e7fc66048f92f74d502c67b526612;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbaa3abe010ef286042b47c7323228b4f12b8ed45f013d3fde6ed09a17fd4ad97;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ae9caf925cd43193f0d2982e6e9987cf5fc59dcc15886dc0787d92d4355a1d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2a84d1f4b3163646117ef9f284f84f712a1308e5740aaee9ca599742730b705;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he516022a4d933aa4ca66db15022f9e8d605b30a809b83a7ee4adafc4170b0338;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37eb040ffc63eaf4a4c15097963acde702e53661fc29c2c3804ae12620e3667;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdaa27bed7e4db65339b65564e6e7dcbbf644b175c52bbfc6fa3505b28a33b2fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd461745305cd273f6ea0b4727ca560d24a7bb45a0f83a370658ae56a348aeb1f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he98fded4fe65fb5341267c5986c05f54b322c6388be53af932ea288f09cbfcd7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3655bcecfb60ecaecf653e2ac4ca2713ea33813dce87997d3434ad54fca8946;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h91a0cc166f3d9a13e53b1d6bbc43e80888b2f307589f86fa0645bef6fea25b57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3170a5ad51a9b88c8ba639e07fd2cf539dfe9cbdf7b697eda1f55a67306eff79;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3939706c802da4837b8e42db093cced4b32f2efae253060a37e1c635dffb02f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h383b9789841ac425d0e82c00a1f69733905a98416f8637aa992500edd2f90920;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59b36e6a9505c149de6dd9e638e76557600e945e4be9b84f4ca984c5bd2bcd11;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h132931a3d1bb8e7cb2334a36e7d5bdf4dbb70d2027a7fade81b8415c259bf728;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he49dbf2cd25b14199101381317fee45d4538fe4d9878f61251bc1fd346bfb64b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h84cde5f2a278f7ac8b4430a81a34ddeba961b8faaff2375550c1a5f7c4216bb3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9bb7f116ef508190c271f977a99555148e30de4ebab57c89e28f29106fdcf282;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h55c248982ba5c015f8f86165f7dde11a9bd52071d869d77ddca80bf0a1851c7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9978bb146bedabf5e53d28b75d00b5923cd56ecd736d5b01b58452e8c8b2f4e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe3d117428a664041a0e7f3fb6fe9d680a8627e9d37c1b80f3bea2260bcb9a6d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd9199ab4b793a4ec96285ddffaf26d68751e66b1b1ebe25a85e5265af6b4e4e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8d5a3b434dae8f33c0614e877a58f22d7e89af6549e19eb60f60f19fdab3266;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c9071c02b1ebaf06d22963d570550cba549465f5f9da6ea38766000e4aede70;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf98feef495063271e523b1d901238068bf52c8322fb455a2e35e75c68a199ceb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc43abadb48143344107da9f85de84830c2aa71a45ad8d20d9a52bf4f7f5369b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38608a9ce20a680a888bc7b93cb62c70ea4b5df9ec0d58807065a9b660ec0b05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b87036edb4a83a869df73a6b002613f5b20962744e898df2ed57f019d5a635f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h239de48f57a3a353b7e4fafb423bf2674179a10c973823360e7069cb183cba75;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b4008dad7fb44b9e1906adec0c3395cb55cbdada13c36764a22a99e3ad75674;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62f56eca3068a48c52094dc23651d5c1bdd55736a50abdf3793b153e0e5b7ed3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40cb740622642f666680a9b6672808413b84bb0ed73b038a1c08c3b57e6bac91;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c20ec73c902481d6ff939ee7e8237b90cc6fbdb3f45980e09b120272b0669bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa2c13e392d5dbb1f310f25b6ea38d3f81c1adcf72539745fdd5a7c73505a1d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9d6725767815684d340b20d3fe38a45541c86303090214c5652dfd0b6356bb3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b357ac58f7bb0077e27d235c91b9f6c18f2e43d4493edec86c032957b72c4c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc10945b81dccc660fdd4af31d1a321f22e7a8dd0eb0fb2e4b59f2ad56087c02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54afa66c852f9cbde0fe5d26a6bd78a5e34def4bd79db5208c7267ba150b276e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93454cc2ccedfc64ab4926348976e73e5d772d9911550476224c889b70bc8dc0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97ce11405882e16c777f754e75097ddfad9ebf927e98989b583940b1bc5fccb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h51c1e3d54bc868b85649158cb674acaca9aecb99f82ee95163847543d3e27326;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e21df5a8f61677e6ae33a3a4f5c00638c532cf6d72f9265a0bd42b840bff42f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff9392632985bedca05f80e8dfe9a3c1bed18839c987aec2ff44882fae89d4ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd503bd01645ba8cf673efe4550c67b42b7ef1f03b20533febb5d6734aad9c67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d42fa36fb277490ce499bf03cb32a438490c43d248ae99a6d196b972c6d35a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f7758cb6513eb9ebe01b8f0e9223da71fba016c5178318df5340dbbc67e3611;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca9b93d9896993e972913f222da59cce4b52a13b71b2a7b50f115be17986839f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3c7a5a51574a2bef690f1c88cf370c225812aba4018b144eeb09f25ab33b0b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2eb9a6c475bcf9dbfc2a16fa6da1e214af12c8c2848edd9d4835ea1a1241605;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15ab08750d361945913dc24719af8dee6e5d426152e7d960cdb65b87bf5f910e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9952b2f40ccf4a669c1e04a7f00f86be5db7931cbe45237636c95b5eb7778d3d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9c6c44e947253ce099be14a085db400502b0f73345ce890fc9ee4a84503a3a59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38234482d0a65758cd41cb4dee8fadeb190c17f8eb4b46e24e8366f4600574fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb6825a076895261b7921fc0a625014954aaf6fdee0df98ee72fff27a9c12e43;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he622f36953b317c92a19b2c4f41527a910fb8f292b6c669a02ffcb959240da0e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h130ec0087e90685b7e9159f3b2f90b39f8448c897e018a40bc30f79513f4c51b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h659c957d4450424fc3a4caad10a465c17ecc7cf7f880787f7688334caab84241;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8cf8811e1eb1662739d991df7c72cb3222811dacfd0ece23a9f0bc95428aeedf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h307af40efa7c49127e40c4039deabf04314b209b99ba134090ccc673d12a43ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a14380778e96607a2a1bf8780af1499380237dc1b1f3da1a7e421c96c6c5760;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69beedf993299531e3b918bbb978e393c793526a171f4d96505de778a57de2f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he44aa2cc20ebf7bd23913ca7e4d1c018bf35d3cd261bd1bce0720a7361395e21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e90b855d8467fc9c2be2cffaebae1cef24ed02d01a1cf865787e6ae4817f894;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2808d6409a1ff7552e645971fc4ba1c973c7118beb05d632a9d59f1611e5df57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h184fc51b58c1e7d22b6ed71d353a1c1bba86ef17fa5a9c32e331f62ebb5baf41;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a5a895105b36e1f056104f801517fecb56c168f27edf8d5ccb1141382787f39;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h22e5df53158aa0174da020e524f14fac81e7740f9672a8ab388524470fdb9165;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf363ca5d7a6f2424121d28dea17216752c09e4c675157aaecdd22e7155ea441;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha699f6d3655b1216f2465c0b5a16ae8bd8bc50488ce9e9db8236a10007353b32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a53ff13c5503cae661b37910702237f03d0f9f4c2c53238370d1fcab8bb6fec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5bc1ab33405628351cfa5dc511d0ba5f4618a1a15397dedd67c8331be775d09;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h345e018505fb7d123eb8837ee2f4cf36d4df6358689cb7620d60716551669d1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8d21261f0011593a74325d439f9e6d7aa92ea108867944183801a45a6eb6355;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8073c462aab33116529cb655d88c10513aea5d29a6481176b591cc8e36aa0968;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1887e05306c223e74e622cd028484c9ae2b87c4990d06ee7b1c3c099a1b37b7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h81f16a93d223e334510c0ee648e5f2b969c47c53276ad34612fd9acceb257961;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53031e0e45a883be6db301726390671e625bafe848940b3ba3d3074e8694bb1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1362e23fcbc63912ba0783ddbbc792a8d752d7998468695322058edaef5a4ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2404c0640b4f695ffc20a7e4742e113082faf151a03ba7ef1072c0db9a2697a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17e5e7d0fad8c4b7e48b1e6042dc935a8f63f3796a0233aeb01bd61b24fef515;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38861a584bb2e564b270aae574ccac4f7acef62ee6fbc347bae18039afc3f412;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h438ed8b60854faf9e535f41cc01966bfc7618b812ca67bca144a3262e0dab974;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he83a4e7de30bcc1ca4b166e0d554f9ec6bb92203cf840663813d32588f75602a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff867b2a86fdf9ad190c8055d69538aec656c248ba86f7cbf9109abb9f3afbc1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b72b21f2c348ca05e41e0ee2e87270f04bdf8eb00d895a6e052f981a667d0bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he51172925776c70cbf458c76c7fc451cfe7fed4a8fb3b87fcfc262a2b69c285a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h51c65ac0c25e30c867367c0ef268feb542622ac206a7cd76a5f558878ec17fca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h215c2ef8db68152e4ffc75b42ef0a6d8273829f78b485bebb65dadc6f700629c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h675ad152373206abede82a9d7312770ae4885b733483e101f5eec6d0b572ebe2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b3f835b67f95cb482ff479dae21ef1b8fc0205d13344fa92cdece6e0fcc63a1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3c69e98aa3c7dbdd301305159ba329c344a0877bba24c0a986291a8b4a8196;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c2ca13793fac129b43c601cb62b68a5d2b038a9b70686192fbe5e5e1727f328;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb56f04d8d3271442fa26acae92fbfee8b37233dbbf5cb932b6c10dec9c81acd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4240ef7eaa080012afbf9de92bb4ea18278b4a165b83e150668dd910e2d32c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hefda027ffcad14cc34c5e432a630276aa2d3d752760024e5b36c906b386c6d0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77d4c7b47f32800d9cbdc96fd6040c47a8fe7c803b966344960f6f8b6a2ec681;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1825aa220877119336b8028744179a9d0fcab7221cfba6e61e9fefd9f2b9efa1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a65b44772cfa7e251155fb7b19972f944b5b8ea47a3c336453da6d1270e31d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h353b87e091e60125a0787cef2ca7c3ad7e03fabbc27fa258852e1a4d70096f2b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h84a237400c5799d7578730d69841cf417c121f22d4e4c7705da5ffba90a44816;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7de3337c4bd7e75701d33151f28998f65004c9602650d312d9ddbed204d1ec99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h522a21b7257074be47615bb3b4f128e24c1cb20d22c30fe33774204cab083a85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8cdc01e5e4fedd9288ac1f7c3c7986e683a2a89d45c1c6097c5bd036bbb0ee57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15d62164c1b6c119f92bc606109c4ef78f601eed960eec58048b112bc6e09b44;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97d05b7938bed9c00239f88f423bc110f319590b7f30d1d3b442c6e92ef395c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd27ecbbbbccbd5064f62905abb50b6e8ca7de71abc0dfece202bd43c80c662a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4cf28c87428eea12a6864f85d4cb1dedcec5295e1faacff88ff2e338ca359022;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbae5ce64d727365ccad41804aa1d449afc9f0d21996e69f92d13779ab2e7bda3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b96c15ccf9ef1639b873652d254b08d8c58cbbcffa39ce56228cdd0f19d5552;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c0651ffa17f8f8e1ed236375a1f398ad4f77a28431b5f8cfd95c8650108633c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h866f55d33a6afd496824089c4d0c1dc588bf59fbed978c070a857e4d38cf6179;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17ec8cb14709d9e3e1aaac3903968fe835d6f8aab2854a73e24b353ed6aaea7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0ad9f4072661fe4b194d72b77335a532a10520b6e6198eec90d461993f8c897;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5148e1b9d1b4c24c152659924c94f9ddde53ee975af1381bec900764ac70a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf0c082f75a84ba34e241fc420c202baf294655e7d99ed35c77764b0ae41d3f12;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a614d4efbb988cb6d49f924e0a4c17f3eecabf7b1ac84d6e93ac89fa6ed3f0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb4a5f445a3d4dcd4ae1eedfc9681a2b11f26b9d3598cc586042bc69e97bb75c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1525a57e27cc289dbc7f0009c03fad1d965c0cd0860afbdfd77334fb0ea43f59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h81a518bcf185c6efae9761701ee55b116375a3e6c67af967f4430f7f85af7c47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8de84fc337f26a52040ea37dc85a6d3ec3672c67d9bc0a379218b4011ac4f27;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89b71c8687104355160670f476bd17591ce3c48ec9b0aab9d0759704e05448c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h976f896c3b027f905e71febd959c742980edf5a89b00b65c0078105d47b6f95c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f75d3494d16d8ddad7859831d8c8a2e62c7f3efd12ca467cd7c605b08273213;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h71361d1bd9c3d869689cce1667d119ea3e59bfd0268d7c07f078d2975e136081;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4bb7ab38167102c528a3c4cf784ef71e1bae3938db4186c68da68687b8898ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f98b9cc2081a3ace1e72ab438a3a5b8fb65c6d995d2e2ba4f312cf721454b9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31256ba055df7c003cc02a4f927b7240e9c906cb92825ab771fffd1668fbfcdf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7cfebba669d0d66ff647022d37bdfddf878da8d8fb1f732e8a8f81244dc103b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3de065c1dba70af9b283bb1853e444b9c4de87c833c09c99f2dfda1184626e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1bcaf43f32e0d5fa4f3d093e64257133b5815d739e8204ca723f98890e476530;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h65adc722906ba3b40ee4f9bdcbf2ccb4bca6aa56cd747a8f6d71c4d1ce74187c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77633f0c720907a9d56e61dd6429164af7ada5a1c4a962f05677598db39daa9a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfedfcc144b929fa6d471b5af83b33ea839861825cc3abfd1fffb9121fbe5cc4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf792a689739c536aaa9b88e5ce810ea92ebd82e90ab78ad5381abe98795a728;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe74613bff9fe7b3edf7e4f4b250c602f24b521945c4a3f271d6ff4b5c6fe666;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a9c31c366c5555af52811db5da644436a802e26a0b2af2b1d7ec3eedbcd7484;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd85a1f8403438c04d8ceb807a5bb44dde27588f04d894cd6bcb18b849285855;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e7e9d893cce5cf59ab6bcf3084dbe9ca8ee46af8ef205a01f78f469d9ac3db4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc53ee004a78b548111959231d9e8a84b7aa759ca7948c5218cf3914e63bf81f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e603cc279da34396ad521630a376252e46c822293fe12ba4d63b053204bf5d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4c9407e2dc1dd9286a250fc3e93f806da22dc1dce4e9476c3b749ecdf4c3352a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50f6b0f2905a5408ca4a5ae70ef16b340b9c70ae828c1fe819ab20ed3d8a2375;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h51128a2ce1bcc3105578ecd1b67d6b7a785fa43cc8868d5ac4e7596cbfcdfd7e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0ed486c5bdb714c80a778577c8d1c488420236ca9dad66cf06f105120de19e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b4edfa51fbdf71ba3cd117ed0ea65385d17c3738e311bbdb039ef6c496b2f1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0016e0e6eedbd4d53ffbc9fa30f423d52ed2141300c77dec3ed864585b6ca8d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2d33f0aa7df06af2080980212379c4bcf7768f56d62ab3596fe32e9f3f3622a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab51b5539696c13fd625187920e71ad066b5abd314a91fe230e69f8b743f6611;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50847f56ed0d1b543bfe5fbb4a87843684c9ac0f099506eb63c487720b60041a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62e036b219bf646ec6fcc9abec6465f6b712c46cc4a40835bfa83264cce2bd8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h843aa9ea817861e093a527cd674312d33eed92709ef3aa6205770a1a84c0828f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdea82e34006685ab9e1bded7926c5d801c881f884994f115f5767ac98123c9ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he128114f18dead53b8d5663a3ac25ba2577fd97d24fa866ee852076eddfbbf01;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d19626dd97c7c96e8666ebe731b5fad01d1923742eb2b7f231a8a7998d9f09d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3695fe6d75ccbc946e327c8cbce01eb92e9f9231e8ad8c444ab51e6435bf3bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2455208822a83eaf6e3e1f3160b70ec02af430b09ee99a708a2d5b9f42950d67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe222e6fca1a48cacd9d4a434fd057e9e8032eabb50491c3f03b1a74fb2e4687;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe43273e4632afa84e0ad04ad7450276f2008c0810deca7fdd53dfec819d83ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h366ba6b6811a76cf3413389b7ba15a4b2335b521594ba6598f73a4b9616a7a16;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa49af05a75edb28f030ec015ccc112e4aca5dea3f1ba6a1ef22c6a878109e59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50a7b7cc9e3753e8baa1d2dafb8c450aa7086c1321c2e9591f2fb0f91c3aeb5c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h14fbadb76b4177f629dc91a3f69e37a32859229d51ce2d7c744a9a8a7e66e498;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd186dc9323f80899a7706ff402f1008acb1306aaa4d6ff48c971c17027c3d2a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88544fb165cf9fd803651847eafc8167e7c299600bd28676f1fe7f30905a6669;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8438a22710a41acee9ed7013f4ae0e91d8c046a2a61233fd4806f697b5c5a094;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h409efee677e1d217432e10cd4c287fb4bb22d17436dc0d35ec6b20b39832182b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42794cbfb344e79e000587b56ff5894eba841f2af2afe01cb644eed2a55b143f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbcf8c98b25473ea59b13eaf38b9dee8e600f4a5cf91a5ee71cdb62e00f795c35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9920d57e26e71e1932f799a5b96fd947edb98382f3f25c7eda59f7e5986459f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e5a0055ad548c39bcada413587a8c27ce8e54752a8fd7a8b1045e7759604f00;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3cd045f3bcf434a3a1290612ca69cfc786f0fe35b60b480c08076de73eb8ba18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h95bcfd89ccc46578ce3096638377a501c87c7899115aced9c62bf78444550836;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe94384a411aacc7af62358f15caba23ea25755780693dbed6a475fda907be8d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98fc87f2a326cda7b1c8eb6e855fd7d8cdb48d96e77a07362855e7835c45f486;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9ac5d337431a624f1c03f937149a255cf5734c65076361057fe7776ce3facb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f0e471d1ee8d8d38a211ae34e64e4bc625e76520235eeeeef91b67feb8a269b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53f702cffffbea7d5e1ef90ff7a5c7a1bd34498751486a35a690fc5a2da2f683;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h105f2a24bd79e9ebe0d380c2449076193a22bc735ca24f3c24fd4dec51ec5bc6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98bf3e80a6ff6b8b20cb0735a2cfd477fbe645bab8b531a0a5ac2d025b5ff74a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb878077ac1b1c1a0f13d6daeec1cd65690d684581acb327a1327d03e5419b61;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h84413702cf7fff6e057ed26bcc39f9042ed2f723a7def691d86d59b1f90f2b4f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f12a2a67e5bb5ea158a5ec14b2b53a77b9928728e9c4392c668624085dbdc60;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h99508564a4e3fa537a851b31d1391c40613e0a4d54012d6dd22a26b4bbbf9f32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he95aca12e7b8e57ff6b2e2e4e42655b47e3bd3c673ca0a256d2e203124d07571;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4c6153bb1c160dbd4340c1a8e70a68914e3bfac36e023581bb7e35902979cec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8953909173f7bbf84b679abe6dcbab8c1f62b34f814d0623dbec0413851fb89;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b4819257406f4d23d5d3b85aa0202b79ae712cd309da9ea69305d755030ce0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd329b8cf263bcd3583d158984e261e52adbc069bc79dee6119d69711f6f304d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb65deba8afe4e26bf2d567b46fd050a2318d90fc87edc3b8886a806d18d4fed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h34c52b2b0f49c992cf08cb2d8e793bdf626fec4f78102ab9e3563bfd27ef40b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6837849764dcbcae7ddef565e251dd54795733b6ff17cc296a26fb9b0c79685e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b9027e4b7cbe975551b2f0346cd0e259705c13e1649a29dc85f38e74e677a3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbbe600d4a8e860851a3eb71b89597ebd1f696bf01897fb512dcd91b9c9d07f10;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92ab77626e76a37d1d6a5cebdfcc537cf7b737e1b693b6cc47a4e5117be4034a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75e74a9830c5acfa5e54af1bda20ed9f414146414575dcfca151e8b00375e525;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40a9bc487aeed1dbb82614dfd3fdb27f78df89da9f869d6b8ee8515c4358b04a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd118f0cfd8af936a4c057be4466a528e01023c9775f348c61f63991b13acb774;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf0fa9ca1e81f85ca9f61a5e635289f59109b5a59e360790b4be5f66c8cf3278b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1912550bf8c6b8d28a9448409d87a36c316b1dc0f7bb6fd207cc2b305d12bc54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf73e71b45ef9cf3568672d3b08ffd6c8533bd93d6468c72fac6881cd837581d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd1a922ed54da0ca5712a0f5e885265136fcc5712648163a1528e2f4b885e35f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb0937f76c1f40a9ec7d7dd6871fb3cc9b8470c54f51307a8ae2acd92d2c43167;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57f9db9fd750440d563ded84a50e4b8c124c836fa26aa826c016bce155937bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h454c8cc1ab1ea88916e77b6c4673c7d4db43b2308eef6266b47bbd1590ba235;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc213109c27f7108a34538412fd2ba1a7dc5a9af0c2c3660c84a3d80b8b9b3cc9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28550383e2706242bd54fa5337e07038a7c06478d189c5d4bdda0a3f912e9a65;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe874ec0ef2da4d23ecac99c6589f711100f929fe4f6af32d948a3a648bdf1b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4865f15a34d99e71bbf2710cdac84d198047aed1d17fcd2c020cbce5d65e17d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7312e12e2ed01b7bccb85f815b8673789d72614974b5dc5ab6b595c87d7ec47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h349f98b181d3db449e187a740ca3a96ee4653ee63462b39d54c39b6ead9c50d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e7d56fbc5cff5b0843c391419a0f122ef141599f2401a2e4724c5e4cf63cb44;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h686e45c7adb6d94a2dc4e0d2afd7ffbf38e67df3177112894911760ccd8aeec0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5edfec2240a067e6ce6ac21fdb5dec4e0ba03168007993cfefb975092e0389c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ecbaf82aa559593240394db44847f07b0226c7d123fe64bc93d3c6aeef31527;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9cf597e4d2b45a39b4219e93fdafa75df14d050ca26ff483b4f8b6f82f651ec5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96425cf40c6e41d92c17a93225dc4a86eddc720f4cee5006818963c154c4f003;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4beb15973a43db825c0222d68322675e7ace442f629d863e32a8572b317b0cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47c8daa05ab892398d1876685a3f2e653022ecbbdc43b8bbe6d48f4e6aa6050d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h207e03a96e94f3f31df9bccf7ff1ffbc7beb7c7fdc133b11ddde73166d5b1425;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1edab72345d7ee740bb8a3fa26e88194898d2f3cfedd49d75f384f63f8274c58;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a34565cbe12b7b8327c69da868908c2b952620d4a26863576cc711ce1721b8a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a9ad72bb71e1d4f8acf4f930723094181f84334ab2fa202627f571bd9e85c8a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60b5ae2eaee33bad55c0d8209768e1d49d66f20f5eaaee9bc4a621c7bd404b85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d261ad703ca091bc1c03cb3e93210bf64a5c1214223b0219d511ef1b09875f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb3d2c095cba3de062e99c7772d11150987938e76202fb7b15a5f890f68fb9964;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3d3c6a7a2eab084cdc23dbcc8a5a5aece6c054d42d7efe7e88213db77385e35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h567c6ce81cf11eaf4b40fdd5ab77fd26d8ca8ff9311c8091705b06f6d6c1ac1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h81e946f1ec8da821ea572277a82a423535175ecdadf5f3351b9869ea320320cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haaf97d20ae3306dd64fa26d007c99e75dec387949ac628eec4ffe07c52828e3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf6518382e8f86c8e6ea02cf5f7d1f32260942b6e8d7a4e87bed39a07665a88e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89d60f3e7f1cb17aa6851b7703695716853ac71d1f7d11e711b42b47edfbe11a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6ba8b111ae479228e8843bf57c228c67d9a628bf10c4d91036c59d6ed662392;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f2dc9c71c8a3d8838f768532e3838b5894d95ff129a2efdf69d413fc17828f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he843c4bbe3e803c9b954fd24d87e705434d6339a732f1c1239fab33171ed6218;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef396cf3e6643f940fc8d733da36187bdc787a7641b6189b2e31faabdd996565;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3b6ae47c7486a9a9e1fee72be2670c5fa6435a542bcc007a1d7816b03a6e9c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h852ee993c7b36f79b771b64101e7fefc71d45a614dc3db0b96555fa934391efd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe1451efe41b73fe555da5d4fa0bab2872d0fab9815cb8dfd2d1f358dd5f4f3a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb411af274fc3f4693e856d1f1c840d04d6726fae285b79b3666baacd75eac4bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb20e0e60ed97ada71df6a26cdba27babee6e8ad57b52a3cb8854b7eb1abe4bda;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h22d3f171b901699c061ca8bee62fda5d4b356af9d26f7929ece6d3588c681dd4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3832b75394d7cfa768e58834ec08606db90d6dfaae3c9171883b3f87693654ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4c23ae9ba3af646397aff1ad222e6d796b1dab43bd7e4f241f0cbb1ababfc15;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36be60dc7e9029143f1011e94a70a19450b49cfb29730629b6c3d3a4c4efdf20;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3869b6d286340fbdc210b340bd07520ba7049b9b9f547fdd3e84c1bda2d79be;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfbba28dde39ba3261fc0c7673e429f93b16a11eb4b7204e18194113e35ace34c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2324b4425969f84c0e8200d8dd63d19af5eb25c10c794e4e0ee6d6f1dfecd8f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he32ae16adcdc0bd8405561f9037155aa03e363e8c3e1dd67ac1ecabaf6ec1ae0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4f840238a0babe046fc21432b5c92ec5523618fe314520c565f3dfce4014e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha587f48e4db772fba22ac651407d48058367d904de0f02400164e9b03ee88841;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0551ed78217833a03602fd682401ee13f602a44114ca0bc083046aac983b786;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he528ca40849366ce793972442d2060358487b4d6e6f7c2f054fef1bf6022ae9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40058eb69d25a9b4777aef528ba7b9321c329fe4968b91a979937892e32087ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9e75e187232bb28c9d22179ffeb459e8a7bed1910367f60a41b198909f0600bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h578aef1ff1ce9295a02979ab4341de90bf1e16816205d25d4478236a82fc5d88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcaf9178eccf4d990674821c733479dfce497aabae439bbdb9f733bf9ff1f8ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41b3b8112acaac269543c494ab6f08504941bda7a6f30d4b7c3773f30a583866;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc240021d1b70abe734de260745ffde7a210deb280fdd71f4bc9d7f1f8136cc2c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8cf7e1d8025ac5edfd2abfb7d7e9393aef8fc730ad554ba7b9311d6f4dc9f642;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7003c19c68b0b906e143a7372e089fca96d2a81ac869cc742f1bcf8aef8561e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e595446c18e3bb2599e40d08483dce43c7145d11dad083cfba3234aba48f156;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb593aa3b63502235961c9d163691afc8af2cd97aaef37cf08d3c5987c3fe7266;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89ec7df8102e895af3b7b412b6415d5880d444a24a9bd07af84f466157e17c26;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73f81130bdd5cb32c3e9df6d74d987e8e93b621374149210f7b5084e70d89bfd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a959fe6f20187c05450ed73a76794eb6c10fa5f51fd829c70c0a2bb57326ca4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20ddc74f4c001c681afc776d73a787790c0f4e84111f414142d546eab9672f5d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h196347ea69000f98116d98e83aa05d05f20cc2145efec0d53b0bf8fa6f41f22c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd728fdf96a2b161079520bf49cfa5b98fb4253930306ad35361be0381a7c76ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa36ce9cd655ab0b67b3542f6d41fa35782b25c4c5cf25bb91322abdcf09a3a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1829f15b2b19697837fc695e027aa38418cfe04b6c9dbf6a3e0f940dbe5582cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h55abbc12e88851642c05f898bc1e955506c41debc8809ab952933d615c6d9c86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a07d7e87a18421ca8336f02de98d0a17d8fcb7a14c751ccc3ef6ffa415465f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc77988c8f768bf45d11e634e3c7bb5566c8bbb21fcf21517bed7f2bc2f0b68d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d7ab12318dfcb8b41a0a07e70915642437607023a4f5c4ec51a577672949d14;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h251fc7e87374f78e55592863ae3453685abf9f5b64ea3ba8309898550138a1ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb72e593eb6ef2a61ccb620261cbfb0baf123d1bd1d78e1f2b011696d822f4251;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68502e3bb28a0f50d438e529f9793686b4ec1d91641cf238f4d9ed47fae4db34;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61b47124a9becd7fc6735d903c83d9a3636ba22bed3dadbfa0595a3b22b0b935;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba435e22d1efb4b95cab16296ba3abab9d9a5ed8809374fd19cfd2d01da69246;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b72c915fb5a5cfd3b8f95e287c75b7cb0cab6216f108fb495832a7247921c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf24774348a5412b9053861a17e3771903b28a8b5ea1b0018e17ca76c87b78366;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9e01b8e76fb7729bea49e05348dc910fce2e91199f1ce22651623d3da9ded9da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31f79f42cdf93a4839e535ed4e4973d62e387b855cb5b6fd2c6934c7f904db93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88e96441ebe755a5456d9f03e03366cc62ba3f51b8f289cf98a2182cdf90903a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h911f62d21b849e57261e2b5c53662f1db43c11c62a9623db9d24a3f3cfad1f9e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h51798b4ddeb0eaa3b6857a4e05706d67a88c93642ac391f5a98fcb292dc249e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h114981704d37b2fba034c73d14efed7b37582ef977f08cec2cd24a31d8cd04bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9e4db3420e2168db9e1e1912f42b2cfa3e557b0ed6c7a8730883b08928bb9d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4eb9eeff613bbd6ffd82fb1f3da42f89612c0baa30ce85bda2e72d0b6e1f11e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69288601e027f018a13df5aeb3744fb8ca0d6ac991c23b946417fa3ccf6d8e83;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a4476d6361dcba46b380bc051bf3918e3127d3da02312a0a8ad0529d75be74a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6daa9ab32531df2cd5679eb2a9a7c42de0778603f7dc01eb80fedf7ff7972625;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b846d2faa0caa13069e0926a3b4cf5fef82f142ddcdfcc2c5758fbda3da2ea8;
        #1
        $finish();
    end
endmodule
